// SPDX-FileCopyrightText: 2022 SH CONSULTING K.K.
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

module j202_soc_core_wrapper ( wb_clk_i, wb_rst_i, wbs_stb_i, wbs_cyc_i, 
        wbs_we_i, wbs_sel_i, wbs_dat_i, wbs_adr_i, wbs_ack_o, wbs_dat_o, 
        la_data_in, la_data_out, la_oenb, io_in, io_out, io_oeb, analog_io, 
        user_clock2, user_irq );
  input [3:0] wbs_sel_i;
  input [31:0] wbs_dat_i;
  input [31:0] wbs_adr_i;
  output [31:0] wbs_dat_o;
  input [127:0] la_data_in;
  output [127:0] la_data_out;
  input [127:0] la_oenb;
  input [37:0] io_in;
  output [37:0] io_out;
  output [37:0] io_oeb;
  inout [28:0] analog_io;
  output [2:0] user_irq;
  input wb_clk_i, wb_rst_i, wbs_stb_i, wbs_cyc_i, wbs_we_i, user_clock2;
  output wbs_ack_o;
  wire   n3, n4, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n220, n230, n240, n250, n260, n270, n280, n290, n300, n310, n320,
         n330, n340, n350, n360, n370, n380, n390, n400, n410, n420, n430,
         n440, n450, n460, n470, j202_soc_core_qspi_wb_we,
         j202_soc_core_qspi_wb_cyc, j202_soc_core_qspi_wb_ack,
         j202_soc_core_aquc_STB_, j202_soc_core_aquc_ADR__0_,
         j202_soc_core_aquc_ADR__1_, j202_soc_core_aquc_ADR__2_,
         j202_soc_core_aquc_ADR__3_, j202_soc_core_aquc_ADR__4_,
         j202_soc_core_aquc_ADR__5_, j202_soc_core_aquc_ADR__6_,
         j202_soc_core_aquc_ADR__7_, j202_soc_core_aquc_SEL__0_,
         j202_soc_core_aquc_SEL__2_, j202_soc_core_aquc_SEL__3_,
         j202_soc_core_aquc_WE_, j202_soc_core_aquc_CE__0_,
         j202_soc_core_aquc_CE__1_, j202_soc_core_bldc_int,
         j202_soc_core_qspi_int, j202_soc_core_intr_vec__0_,
         j202_soc_core_intr_vec__1_, j202_soc_core_intr_vec__2_,
         j202_soc_core_intr_vec__3_, j202_soc_core_intr_vec__4_,
         j202_soc_core_intr_vec__6_, j202_soc_core_intr_level__0_,
         j202_soc_core_intr_level__1_, j202_soc_core_intr_level__2_,
         j202_soc_core_intr_level__3_, j202_soc_core_intr_level__4_,
         j202_soc_core_intr_req_, j202_soc_core_rst, j202_soc_core_rst1,
         j202_soc_core_rst0, j202_soc_core_j22_cpu_regop_M_Wm__0_,
         j202_soc_core_j22_cpu_regop_M_Wm__1_,
         j202_soc_core_j22_cpu_regop_M_Wm__2_,
         j202_soc_core_j22_cpu_regop_M_Wm__3_,
         j202_soc_core_j22_cpu_regop_M_Rn__0_,
         j202_soc_core_j22_cpu_regop_M_Rn__1_,
         j202_soc_core_j22_cpu_regop_M_Rn__2_,
         j202_soc_core_j22_cpu_regop_M_Rn__3_,
         j202_soc_core_j22_cpu_regop_Wm__0_,
         j202_soc_core_j22_cpu_regop_Wm__1_,
         j202_soc_core_j22_cpu_regop_Wm__2_,
         j202_soc_core_j22_cpu_regop_Wm__3_,
         j202_soc_core_j22_cpu_regop_We__0_,
         j202_soc_core_j22_cpu_regop_We__2_,
         j202_soc_core_j22_cpu_regop_We__3_,
         j202_soc_core_j22_cpu_regop_Rs__0_,
         j202_soc_core_j22_cpu_regop_Rs__1_,
         j202_soc_core_j22_cpu_regop_Rb__1_,
         j202_soc_core_j22_cpu_regop_Ra__0_,
         j202_soc_core_j22_cpu_regop_Ra__1_,
         j202_soc_core_j22_cpu_regop_other__0_,
         j202_soc_core_j22_cpu_regop_other__1_,
         j202_soc_core_j22_cpu_regop_other__2_,
         j202_soc_core_j22_cpu_regop_imm__0_,
         j202_soc_core_j22_cpu_regop_imm__1_,
         j202_soc_core_j22_cpu_regop_imm__2_,
         j202_soc_core_j22_cpu_regop_imm__3_,
         j202_soc_core_j22_cpu_regop_imm__4_,
         j202_soc_core_j22_cpu_regop_imm__5_,
         j202_soc_core_j22_cpu_regop_imm__6_,
         j202_soc_core_j22_cpu_regop_imm__7_,
         j202_soc_core_j22_cpu_regop_imm__8_,
         j202_soc_core_j22_cpu_regop_imm__9_,
         j202_soc_core_j22_cpu_regop_imm__10_,
         j202_soc_core_j22_cpu_regop_imm__11_,
         j202_soc_core_j22_cpu_regop_imm__12_,
         j202_soc_core_j22_cpu_regop_Rm__0_,
         j202_soc_core_j22_cpu_regop_Rm__1_,
         j202_soc_core_j22_cpu_regop_Rm__2_,
         j202_soc_core_j22_cpu_regop_Rm__3_, j202_soc_core_j22_cpu_ifetch,
         j202_soc_core_j22_cpu_memop_Ma__0_,
         j202_soc_core_j22_cpu_memop_Ma__1_,
         j202_soc_core_j22_cpu_memop_MEM__0_,
         j202_soc_core_j22_cpu_memop_MEM__1_,
         j202_soc_core_j22_cpu_memop_MEM__3_, j202_soc_core_j22_cpu_pc_hold,
         j202_soc_core_j22_cpu_istall, j202_soc_core_j22_cpu_intack,
         j202_soc_core_j22_cpu_rte4, j202_soc_core_j22_cpu_rfuo_sr__t_,
         j202_soc_core_j22_cpu_rfuo_sr__s_,
         j202_soc_core_j22_cpu_rfuo_sr__i__0_,
         j202_soc_core_j22_cpu_rfuo_sr__i__1_,
         j202_soc_core_j22_cpu_rfuo_sr__i__2_,
         j202_soc_core_j22_cpu_rfuo_sr__i__3_,
         j202_soc_core_j22_cpu_rfuo_sr__q_, j202_soc_core_j22_cpu_rfuo_sr__m_,
         j202_soc_core_j22_cpu_ifetchl, j202_soc_core_j22_cpu_id_opn_v_,
         j202_soc_core_j22_cpu_id_opn_inst__0_,
         j202_soc_core_j22_cpu_id_opn_inst__1_,
         j202_soc_core_j22_cpu_id_opn_inst__2_,
         j202_soc_core_j22_cpu_id_opn_inst__3_,
         j202_soc_core_j22_cpu_id_opn_inst__4_,
         j202_soc_core_j22_cpu_id_opn_inst__5_,
         j202_soc_core_j22_cpu_id_opn_inst__6_,
         j202_soc_core_j22_cpu_id_opn_inst__7_,
         j202_soc_core_j22_cpu_id_opn_inst__8_,
         j202_soc_core_j22_cpu_id_opn_inst__9_,
         j202_soc_core_j22_cpu_id_opn_inst__10_,
         j202_soc_core_j22_cpu_id_opn_inst__11_,
         j202_soc_core_j22_cpu_id_opn_inst__12_,
         j202_soc_core_j22_cpu_id_opn_inst__13_,
         j202_soc_core_j22_cpu_id_opn_inst__14_,
         j202_soc_core_j22_cpu_id_opn_inst__15_,
         j202_soc_core_j22_cpu_id_op2_v_,
         j202_soc_core_j22_cpu_id_op2_inst__0_,
         j202_soc_core_j22_cpu_id_op2_inst__1_,
         j202_soc_core_j22_cpu_id_op2_inst__2_,
         j202_soc_core_j22_cpu_id_op2_inst__3_,
         j202_soc_core_j22_cpu_id_op2_inst__4_,
         j202_soc_core_j22_cpu_id_op2_inst__5_,
         j202_soc_core_j22_cpu_id_op2_inst__6_,
         j202_soc_core_j22_cpu_id_op2_inst__7_,
         j202_soc_core_j22_cpu_id_op2_inst__8_,
         j202_soc_core_j22_cpu_id_op2_inst__9_,
         j202_soc_core_j22_cpu_id_op2_inst__10_,
         j202_soc_core_j22_cpu_id_op2_inst__11_,
         j202_soc_core_j22_cpu_id_op2_inst__12_,
         j202_soc_core_j22_cpu_id_op2_inst__13_,
         j202_soc_core_j22_cpu_id_op2_inst__14_,
         j202_soc_core_j22_cpu_id_op2_inst__15_,
         j202_soc_core_j22_cpu_id_idec_N959,
         j202_soc_core_j22_cpu_id_idec_N958,
         j202_soc_core_j22_cpu_id_idec_N957,
         j202_soc_core_j22_cpu_id_idec_N956,
         j202_soc_core_j22_cpu_id_idec_N937,
         j202_soc_core_j22_cpu_id_idec_N917,
         j202_soc_core_j22_cpu_id_idec_N900,
         j202_soc_core_j22_cpu_id_idec_N894,
         j202_soc_core_j22_cpu_id_idec_N822, j202_soc_core_j22_cpu_rf_N3392,
         j202_soc_core_j22_cpu_rf_N3391, j202_soc_core_j22_cpu_rf_N3390,
         j202_soc_core_j22_cpu_rf_N3388, j202_soc_core_j22_cpu_rf_N3386,
         j202_soc_core_j22_cpu_rf_N3379, j202_soc_core_j22_cpu_rf_N3378,
         j202_soc_core_j22_cpu_rf_N3377, j202_soc_core_j22_cpu_rf_N3376,
         j202_soc_core_j22_cpu_rf_N3375, j202_soc_core_j22_cpu_rf_N3374,
         j202_soc_core_j22_cpu_rf_N3373, j202_soc_core_j22_cpu_rf_N3372,
         j202_soc_core_j22_cpu_rf_N3371, j202_soc_core_j22_cpu_rf_N3370,
         j202_soc_core_j22_cpu_rf_N3369, j202_soc_core_j22_cpu_rf_N3368,
         j202_soc_core_j22_cpu_rf_N3367, j202_soc_core_j22_cpu_rf_N3366,
         j202_soc_core_j22_cpu_rf_N3365, j202_soc_core_j22_cpu_rf_N3364,
         j202_soc_core_j22_cpu_rf_N3363, j202_soc_core_j22_cpu_rf_N3361,
         j202_soc_core_j22_cpu_rf_N3360, j202_soc_core_j22_cpu_rf_N3359,
         j202_soc_core_j22_cpu_rf_N3358, j202_soc_core_j22_cpu_rf_N3357,
         j202_soc_core_j22_cpu_rf_N3356, j202_soc_core_j22_cpu_rf_N3355,
         j202_soc_core_j22_cpu_rf_N3354, j202_soc_core_j22_cpu_rf_N3352,
         j202_soc_core_j22_cpu_rf_N3351, j202_soc_core_j22_cpu_rf_N3350,
         j202_soc_core_j22_cpu_rf_N3349, j202_soc_core_j22_cpu_rf_N3348,
         j202_soc_core_j22_cpu_rf_N3347, j202_soc_core_j22_cpu_rf_N3346,
         j202_soc_core_j22_cpu_rf_N3345, j202_soc_core_j22_cpu_rf_N3343,
         j202_soc_core_j22_cpu_rf_N3342, j202_soc_core_j22_cpu_rf_N3341,
         j202_soc_core_j22_cpu_rf_N3340, j202_soc_core_j22_cpu_rf_N3339,
         j202_soc_core_j22_cpu_rf_N3338, j202_soc_core_j22_cpu_rf_N3337,
         j202_soc_core_j22_cpu_rf_N3336, j202_soc_core_j22_cpu_rf_N3335,
         j202_soc_core_j22_cpu_rf_N3334, j202_soc_core_j22_cpu_rf_N3333,
         j202_soc_core_j22_cpu_rf_N3331, j202_soc_core_j22_cpu_rf_N3330,
         j202_soc_core_j22_cpu_rf_N3329, j202_soc_core_j22_cpu_rf_N3328,
         j202_soc_core_j22_cpu_rf_N3327, j202_soc_core_j22_cpu_rf_N3326,
         j202_soc_core_j22_cpu_rf_N3325, j202_soc_core_j22_cpu_rf_N3324,
         j202_soc_core_j22_cpu_rf_N3323, j202_soc_core_j22_cpu_rf_N3322,
         j202_soc_core_j22_cpu_rf_N3321, j202_soc_core_j22_cpu_rf_N3319,
         j202_soc_core_j22_cpu_rf_N3318, j202_soc_core_j22_cpu_rf_N3317,
         j202_soc_core_j22_cpu_rf_N3316, j202_soc_core_j22_cpu_rf_N3315,
         j202_soc_core_j22_cpu_rf_N3314, j202_soc_core_j22_cpu_rf_N3313,
         j202_soc_core_j22_cpu_rf_N3311, j202_soc_core_j22_cpu_rf_N3309,
         j202_soc_core_j22_cpu_rf_N3307, j202_soc_core_j22_cpu_rf_N3305,
         j202_soc_core_j22_cpu_rf_N3304, j202_soc_core_j22_cpu_rf_N3303,
         j202_soc_core_j22_cpu_rf_N3302, j202_soc_core_j22_cpu_rf_N3301,
         j202_soc_core_j22_cpu_rf_N3300, j202_soc_core_j22_cpu_rf_N3299,
         j202_soc_core_j22_cpu_rf_N3298, j202_soc_core_j22_cpu_rf_N3297,
         j202_soc_core_j22_cpu_rf_N3296, j202_soc_core_j22_cpu_rf_N3295,
         j202_soc_core_j22_cpu_rf_N3294, j202_soc_core_j22_cpu_rf_N3292,
         j202_soc_core_j22_cpu_rf_N3291, j202_soc_core_j22_cpu_rf_N3290,
         j202_soc_core_j22_cpu_rf_N3289, j202_soc_core_j22_cpu_rf_N3288,
         j202_soc_core_j22_cpu_rf_N3287, j202_soc_core_j22_cpu_rf_N3286,
         j202_soc_core_j22_cpu_rf_N3284, j202_soc_core_j22_cpu_rf_N3283,
         j202_soc_core_j22_cpu_rf_N3282, j202_soc_core_j22_cpu_rf_N3281,
         j202_soc_core_j22_cpu_rf_N3280, j202_soc_core_j22_cpu_rf_N3279,
         j202_soc_core_j22_cpu_rf_N3278, j202_soc_core_j22_cpu_rf_N3276,
         j202_soc_core_j22_cpu_rf_N3275, j202_soc_core_j22_cpu_rf_N3274,
         j202_soc_core_j22_cpu_rf_N3273, j202_soc_core_j22_cpu_rf_N3272,
         j202_soc_core_j22_cpu_rf_N3271, j202_soc_core_j22_cpu_rf_N3270,
         j202_soc_core_j22_cpu_rf_N3268, j202_soc_core_j22_cpu_rf_N3267,
         j202_soc_core_j22_cpu_rf_N3266, j202_soc_core_j22_cpu_rf_N3265,
         j202_soc_core_j22_cpu_rf_N3263, j202_soc_core_j22_cpu_rf_N3262,
         j202_soc_core_j22_cpu_rf_N3261, j202_soc_core_j22_cpu_rf_N3260,
         j202_soc_core_j22_cpu_rf_N3259, j202_soc_core_j22_cpu_rf_N3258,
         j202_soc_core_j22_cpu_rf_N3257, j202_soc_core_j22_cpu_rf_N3255,
         j202_soc_core_j22_cpu_rf_N3254, j202_soc_core_j22_cpu_rf_N3253,
         j202_soc_core_j22_cpu_rf_N3252, j202_soc_core_j22_cpu_rf_N3251,
         j202_soc_core_j22_cpu_rf_N3250, j202_soc_core_j22_cpu_rf_N3249,
         j202_soc_core_j22_cpu_rf_N3247, j202_soc_core_j22_cpu_rf_N3246,
         j202_soc_core_j22_cpu_rf_N3245, j202_soc_core_j22_cpu_rf_N3244,
         j202_soc_core_j22_cpu_rf_N3243, j202_soc_core_j22_cpu_rf_N3242,
         j202_soc_core_j22_cpu_rf_N3241, j202_soc_core_j22_cpu_rf_N3239,
         j202_soc_core_j22_cpu_rf_N3238, j202_soc_core_j22_cpu_rf_N3237,
         j202_soc_core_j22_cpu_rf_N3236, j202_soc_core_j22_cpu_rf_N3235,
         j202_soc_core_j22_cpu_rf_N3234, j202_soc_core_j22_cpu_rf_N3233,
         j202_soc_core_j22_cpu_rf_N3231, j202_soc_core_j22_cpu_rf_N3230,
         j202_soc_core_j22_cpu_rf_N3229, j202_soc_core_j22_cpu_rf_N3228,
         j202_soc_core_j22_cpu_rf_N3227, j202_soc_core_j22_cpu_rf_N3226,
         j202_soc_core_j22_cpu_rf_N3225, j202_soc_core_j22_cpu_rf_N3224,
         j202_soc_core_j22_cpu_rf_N3223, j202_soc_core_j22_cpu_rf_N3222,
         j202_soc_core_j22_cpu_rf_N3221, j202_soc_core_j22_cpu_rf_N3220,
         j202_soc_core_j22_cpu_rf_N3218, j202_soc_core_j22_cpu_rf_N3217,
         j202_soc_core_j22_cpu_rf_N3216, j202_soc_core_j22_cpu_rf_N3215,
         j202_soc_core_j22_cpu_rf_N3214, j202_soc_core_j22_cpu_rf_N3213,
         j202_soc_core_j22_cpu_rf_N3212, j202_soc_core_j22_cpu_rf_N3210,
         j202_soc_core_j22_cpu_rf_N3209, j202_soc_core_j22_cpu_rf_N3208,
         j202_soc_core_j22_cpu_rf_N3207, j202_soc_core_j22_cpu_rf_N3206,
         j202_soc_core_j22_cpu_rf_N3205, j202_soc_core_j22_cpu_rf_N3204,
         j202_soc_core_j22_cpu_rf_N3202, j202_soc_core_j22_cpu_rf_N3201,
         j202_soc_core_j22_cpu_rf_N3200, j202_soc_core_j22_cpu_rf_N3199,
         j202_soc_core_j22_cpu_rf_N3198, j202_soc_core_j22_cpu_rf_N3197,
         j202_soc_core_j22_cpu_rf_N3196, j202_soc_core_j22_cpu_rf_N3194,
         j202_soc_core_j22_cpu_rf_N3193, j202_soc_core_j22_cpu_rf_N3192,
         j202_soc_core_j22_cpu_rf_N3191, j202_soc_core_j22_cpu_rf_N3190,
         j202_soc_core_j22_cpu_rf_N3189, j202_soc_core_j22_cpu_rf_N3188,
         j202_soc_core_j22_cpu_rf_N3187, j202_soc_core_j22_cpu_rf_N3186,
         j202_soc_core_j22_cpu_rf_N3185, j202_soc_core_j22_cpu_rf_N3184,
         j202_soc_core_j22_cpu_rf_N3183, j202_soc_core_j22_cpu_rf_N3181,
         j202_soc_core_j22_cpu_rf_N3180, j202_soc_core_j22_cpu_rf_N3179,
         j202_soc_core_j22_cpu_rf_N3178, j202_soc_core_j22_cpu_rf_N3177,
         j202_soc_core_j22_cpu_rf_N3176, j202_soc_core_j22_cpu_rf_N3175,
         j202_soc_core_j22_cpu_rf_N3173, j202_soc_core_j22_cpu_rf_N3172,
         j202_soc_core_j22_cpu_rf_N3171, j202_soc_core_j22_cpu_rf_N3170,
         j202_soc_core_j22_cpu_rf_N3169, j202_soc_core_j22_cpu_rf_N3168,
         j202_soc_core_j22_cpu_rf_N3167, j202_soc_core_j22_cpu_rf_N3165,
         j202_soc_core_j22_cpu_rf_N3164, j202_soc_core_j22_cpu_rf_N3163,
         j202_soc_core_j22_cpu_rf_N3162, j202_soc_core_j22_cpu_rf_N3161,
         j202_soc_core_j22_cpu_rf_N3160, j202_soc_core_j22_cpu_rf_N3159,
         j202_soc_core_j22_cpu_rf_N3157, j202_soc_core_j22_cpu_rf_N3156,
         j202_soc_core_j22_cpu_rf_N3155, j202_soc_core_j22_cpu_rf_N3154,
         j202_soc_core_j22_cpu_rf_N3153, j202_soc_core_j22_cpu_rf_N3152,
         j202_soc_core_j22_cpu_rf_N3151, j202_soc_core_j22_cpu_rf_N3150,
         j202_soc_core_j22_cpu_rf_N3149, j202_soc_core_j22_cpu_rf_N3148,
         j202_soc_core_j22_cpu_rf_N3147, j202_soc_core_j22_cpu_rf_N3146,
         j202_soc_core_j22_cpu_rf_N3144, j202_soc_core_j22_cpu_rf_N3143,
         j202_soc_core_j22_cpu_rf_N3142, j202_soc_core_j22_cpu_rf_N3141,
         j202_soc_core_j22_cpu_rf_N3140, j202_soc_core_j22_cpu_rf_N3139,
         j202_soc_core_j22_cpu_rf_N3138, j202_soc_core_j22_cpu_rf_N3136,
         j202_soc_core_j22_cpu_rf_N3135, j202_soc_core_j22_cpu_rf_N3134,
         j202_soc_core_j22_cpu_rf_N3133, j202_soc_core_j22_cpu_rf_N3132,
         j202_soc_core_j22_cpu_rf_N3131, j202_soc_core_j22_cpu_rf_N3130,
         j202_soc_core_j22_cpu_rf_N3128, j202_soc_core_j22_cpu_rf_N3127,
         j202_soc_core_j22_cpu_rf_N3126, j202_soc_core_j22_cpu_rf_N3125,
         j202_soc_core_j22_cpu_rf_N3124, j202_soc_core_j22_cpu_rf_N3123,
         j202_soc_core_j22_cpu_rf_N3122, j202_soc_core_j22_cpu_rf_N3120,
         j202_soc_core_j22_cpu_rf_N3119, j202_soc_core_j22_cpu_rf_N3118,
         j202_soc_core_j22_cpu_rf_N3117, j202_soc_core_j22_cpu_rf_N3116,
         j202_soc_core_j22_cpu_rf_N3115, j202_soc_core_j22_cpu_rf_N3114,
         j202_soc_core_j22_cpu_rf_N3113, j202_soc_core_j22_cpu_rf_N3112,
         j202_soc_core_j22_cpu_rf_N3111, j202_soc_core_j22_cpu_rf_N3110,
         j202_soc_core_j22_cpu_rf_N3109, j202_soc_core_j22_cpu_rf_N3107,
         j202_soc_core_j22_cpu_rf_N3106, j202_soc_core_j22_cpu_rf_N3105,
         j202_soc_core_j22_cpu_rf_N3104, j202_soc_core_j22_cpu_rf_N3103,
         j202_soc_core_j22_cpu_rf_N3102, j202_soc_core_j22_cpu_rf_N3101,
         j202_soc_core_j22_cpu_rf_N3099, j202_soc_core_j22_cpu_rf_N3098,
         j202_soc_core_j22_cpu_rf_N3097, j202_soc_core_j22_cpu_rf_N3096,
         j202_soc_core_j22_cpu_rf_N3095, j202_soc_core_j22_cpu_rf_N3094,
         j202_soc_core_j22_cpu_rf_N3093, j202_soc_core_j22_cpu_rf_N3091,
         j202_soc_core_j22_cpu_rf_N3090, j202_soc_core_j22_cpu_rf_N3089,
         j202_soc_core_j22_cpu_rf_N3088, j202_soc_core_j22_cpu_rf_N3087,
         j202_soc_core_j22_cpu_rf_N3086, j202_soc_core_j22_cpu_rf_N3085,
         j202_soc_core_j22_cpu_rf_N3083, j202_soc_core_j22_cpu_rf_N3082,
         j202_soc_core_j22_cpu_rf_N3081, j202_soc_core_j22_cpu_rf_N3080,
         j202_soc_core_j22_cpu_rf_N3079, j202_soc_core_j22_cpu_rf_N3078,
         j202_soc_core_j22_cpu_rf_N3077, j202_soc_core_j22_cpu_rf_N3076,
         j202_soc_core_j22_cpu_rf_N3075, j202_soc_core_j22_cpu_rf_N3074,
         j202_soc_core_j22_cpu_rf_N3073, j202_soc_core_j22_cpu_rf_N3072,
         j202_soc_core_j22_cpu_rf_N3070, j202_soc_core_j22_cpu_rf_N3069,
         j202_soc_core_j22_cpu_rf_N3068, j202_soc_core_j22_cpu_rf_N3067,
         j202_soc_core_j22_cpu_rf_N3066, j202_soc_core_j22_cpu_rf_N3065,
         j202_soc_core_j22_cpu_rf_N3064, j202_soc_core_j22_cpu_rf_N3062,
         j202_soc_core_j22_cpu_rf_N3061, j202_soc_core_j22_cpu_rf_N3060,
         j202_soc_core_j22_cpu_rf_N3059, j202_soc_core_j22_cpu_rf_N3058,
         j202_soc_core_j22_cpu_rf_N3057, j202_soc_core_j22_cpu_rf_N3056,
         j202_soc_core_j22_cpu_rf_N3054, j202_soc_core_j22_cpu_rf_N3053,
         j202_soc_core_j22_cpu_rf_N3052, j202_soc_core_j22_cpu_rf_N3051,
         j202_soc_core_j22_cpu_rf_N3050, j202_soc_core_j22_cpu_rf_N3049,
         j202_soc_core_j22_cpu_rf_N3048, j202_soc_core_j22_cpu_rf_N3046,
         j202_soc_core_j22_cpu_rf_N3045, j202_soc_core_j22_cpu_rf_N3044,
         j202_soc_core_j22_cpu_rf_N3043, j202_soc_core_j22_cpu_rf_N3042,
         j202_soc_core_j22_cpu_rf_N3041, j202_soc_core_j22_cpu_rf_N3040,
         j202_soc_core_j22_cpu_rf_N3039, j202_soc_core_j22_cpu_rf_N3038,
         j202_soc_core_j22_cpu_rf_N3037, j202_soc_core_j22_cpu_rf_N3036,
         j202_soc_core_j22_cpu_rf_N3035, j202_soc_core_j22_cpu_rf_N3033,
         j202_soc_core_j22_cpu_rf_N3032, j202_soc_core_j22_cpu_rf_N3031,
         j202_soc_core_j22_cpu_rf_N3030, j202_soc_core_j22_cpu_rf_N3029,
         j202_soc_core_j22_cpu_rf_N3028, j202_soc_core_j22_cpu_rf_N3027,
         j202_soc_core_j22_cpu_rf_N3025, j202_soc_core_j22_cpu_rf_N3024,
         j202_soc_core_j22_cpu_rf_N3023, j202_soc_core_j22_cpu_rf_N3022,
         j202_soc_core_j22_cpu_rf_N3021, j202_soc_core_j22_cpu_rf_N3020,
         j202_soc_core_j22_cpu_rf_N3019, j202_soc_core_j22_cpu_rf_N3017,
         j202_soc_core_j22_cpu_rf_N3016, j202_soc_core_j22_cpu_rf_N3015,
         j202_soc_core_j22_cpu_rf_N3014, j202_soc_core_j22_cpu_rf_N3013,
         j202_soc_core_j22_cpu_rf_N3012, j202_soc_core_j22_cpu_rf_N3011,
         j202_soc_core_j22_cpu_rf_N3009, j202_soc_core_j22_cpu_rf_N3008,
         j202_soc_core_j22_cpu_rf_N3007, j202_soc_core_j22_cpu_rf_N3006,
         j202_soc_core_j22_cpu_rf_N3005, j202_soc_core_j22_cpu_rf_N3004,
         j202_soc_core_j22_cpu_rf_N3003, j202_soc_core_j22_cpu_rf_N3002,
         j202_soc_core_j22_cpu_rf_N3001, j202_soc_core_j22_cpu_rf_N3000,
         j202_soc_core_j22_cpu_rf_N2999, j202_soc_core_j22_cpu_rf_N2998,
         j202_soc_core_j22_cpu_rf_N2996, j202_soc_core_j22_cpu_rf_N2995,
         j202_soc_core_j22_cpu_rf_N2994, j202_soc_core_j22_cpu_rf_N2993,
         j202_soc_core_j22_cpu_rf_N2992, j202_soc_core_j22_cpu_rf_N2991,
         j202_soc_core_j22_cpu_rf_N2990, j202_soc_core_j22_cpu_rf_N2988,
         j202_soc_core_j22_cpu_rf_N2987, j202_soc_core_j22_cpu_rf_N2986,
         j202_soc_core_j22_cpu_rf_N2985, j202_soc_core_j22_cpu_rf_N2984,
         j202_soc_core_j22_cpu_rf_N2983, j202_soc_core_j22_cpu_rf_N2982,
         j202_soc_core_j22_cpu_rf_N2980, j202_soc_core_j22_cpu_rf_N2979,
         j202_soc_core_j22_cpu_rf_N2978, j202_soc_core_j22_cpu_rf_N2977,
         j202_soc_core_j22_cpu_rf_N2976, j202_soc_core_j22_cpu_rf_N2975,
         j202_soc_core_j22_cpu_rf_N2974, j202_soc_core_j22_cpu_rf_N2972,
         j202_soc_core_j22_cpu_rf_N2971, j202_soc_core_j22_cpu_rf_N2970,
         j202_soc_core_j22_cpu_rf_N2969, j202_soc_core_j22_cpu_rf_N2968,
         j202_soc_core_j22_cpu_rf_N2967, j202_soc_core_j22_cpu_rf_N2966,
         j202_soc_core_j22_cpu_rf_N2965, j202_soc_core_j22_cpu_rf_N2964,
         j202_soc_core_j22_cpu_rf_N2963, j202_soc_core_j22_cpu_rf_N2962,
         j202_soc_core_j22_cpu_rf_N2961, j202_soc_core_j22_cpu_rf_N2959,
         j202_soc_core_j22_cpu_rf_N2958, j202_soc_core_j22_cpu_rf_N2957,
         j202_soc_core_j22_cpu_rf_N2956, j202_soc_core_j22_cpu_rf_N2955,
         j202_soc_core_j22_cpu_rf_N2954, j202_soc_core_j22_cpu_rf_N2953,
         j202_soc_core_j22_cpu_rf_N2951, j202_soc_core_j22_cpu_rf_N2950,
         j202_soc_core_j22_cpu_rf_N2949, j202_soc_core_j22_cpu_rf_N2948,
         j202_soc_core_j22_cpu_rf_N2947, j202_soc_core_j22_cpu_rf_N2946,
         j202_soc_core_j22_cpu_rf_N2945, j202_soc_core_j22_cpu_rf_N2943,
         j202_soc_core_j22_cpu_rf_N2942, j202_soc_core_j22_cpu_rf_N2941,
         j202_soc_core_j22_cpu_rf_N2940, j202_soc_core_j22_cpu_rf_N2939,
         j202_soc_core_j22_cpu_rf_N2938, j202_soc_core_j22_cpu_rf_N2937,
         j202_soc_core_j22_cpu_rf_N2935, j202_soc_core_j22_cpu_rf_N2934,
         j202_soc_core_j22_cpu_rf_N2933, j202_soc_core_j22_cpu_rf_N2932,
         j202_soc_core_j22_cpu_rf_N2931, j202_soc_core_j22_cpu_rf_N2930,
         j202_soc_core_j22_cpu_rf_N2929, j202_soc_core_j22_cpu_rf_N2928,
         j202_soc_core_j22_cpu_rf_N2927, j202_soc_core_j22_cpu_rf_N2926,
         j202_soc_core_j22_cpu_rf_N2925, j202_soc_core_j22_cpu_rf_N2924,
         j202_soc_core_j22_cpu_rf_N2922, j202_soc_core_j22_cpu_rf_N2921,
         j202_soc_core_j22_cpu_rf_N2920, j202_soc_core_j22_cpu_rf_N2919,
         j202_soc_core_j22_cpu_rf_N2918, j202_soc_core_j22_cpu_rf_N2917,
         j202_soc_core_j22_cpu_rf_N2916, j202_soc_core_j22_cpu_rf_N2914,
         j202_soc_core_j22_cpu_rf_N2913, j202_soc_core_j22_cpu_rf_N2912,
         j202_soc_core_j22_cpu_rf_N2911, j202_soc_core_j22_cpu_rf_N2910,
         j202_soc_core_j22_cpu_rf_N2909, j202_soc_core_j22_cpu_rf_N2908,
         j202_soc_core_j22_cpu_rf_N2906, j202_soc_core_j22_cpu_rf_N2905,
         j202_soc_core_j22_cpu_rf_N2904, j202_soc_core_j22_cpu_rf_N2903,
         j202_soc_core_j22_cpu_rf_N2902, j202_soc_core_j22_cpu_rf_N2901,
         j202_soc_core_j22_cpu_rf_N2900, j202_soc_core_j22_cpu_rf_N2898,
         j202_soc_core_j22_cpu_rf_N2897, j202_soc_core_j22_cpu_rf_N2896,
         j202_soc_core_j22_cpu_rf_N2895, j202_soc_core_j22_cpu_rf_N2894,
         j202_soc_core_j22_cpu_rf_N2893, j202_soc_core_j22_cpu_rf_N2892,
         j202_soc_core_j22_cpu_rf_N2891, j202_soc_core_j22_cpu_rf_N2890,
         j202_soc_core_j22_cpu_rf_N2889, j202_soc_core_j22_cpu_rf_N2888,
         j202_soc_core_j22_cpu_rf_N2887, j202_soc_core_j22_cpu_rf_N2885,
         j202_soc_core_j22_cpu_rf_N2884, j202_soc_core_j22_cpu_rf_N2883,
         j202_soc_core_j22_cpu_rf_N2882, j202_soc_core_j22_cpu_rf_N2881,
         j202_soc_core_j22_cpu_rf_N2880, j202_soc_core_j22_cpu_rf_N2879,
         j202_soc_core_j22_cpu_rf_N2877, j202_soc_core_j22_cpu_rf_N2876,
         j202_soc_core_j22_cpu_rf_N2875, j202_soc_core_j22_cpu_rf_N2874,
         j202_soc_core_j22_cpu_rf_N2873, j202_soc_core_j22_cpu_rf_N2872,
         j202_soc_core_j22_cpu_rf_N2871, j202_soc_core_j22_cpu_rf_N2869,
         j202_soc_core_j22_cpu_rf_N2868, j202_soc_core_j22_cpu_rf_N2867,
         j202_soc_core_j22_cpu_rf_N2866, j202_soc_core_j22_cpu_rf_N2865,
         j202_soc_core_j22_cpu_rf_N2864, j202_soc_core_j22_cpu_rf_N2863,
         j202_soc_core_j22_cpu_rf_N2861, j202_soc_core_j22_cpu_rf_N2860,
         j202_soc_core_j22_cpu_rf_N2859, j202_soc_core_j22_cpu_rf_N2858,
         j202_soc_core_j22_cpu_rf_N2857, j202_soc_core_j22_cpu_rf_N2856,
         j202_soc_core_j22_cpu_rf_N2855, j202_soc_core_j22_cpu_rf_N2854,
         j202_soc_core_j22_cpu_rf_N2853, j202_soc_core_j22_cpu_rf_N2852,
         j202_soc_core_j22_cpu_rf_N2851, j202_soc_core_j22_cpu_rf_N2850,
         j202_soc_core_j22_cpu_rf_N2848, j202_soc_core_j22_cpu_rf_N2847,
         j202_soc_core_j22_cpu_rf_N2846, j202_soc_core_j22_cpu_rf_N2845,
         j202_soc_core_j22_cpu_rf_N2844, j202_soc_core_j22_cpu_rf_N2843,
         j202_soc_core_j22_cpu_rf_N2842, j202_soc_core_j22_cpu_rf_N2840,
         j202_soc_core_j22_cpu_rf_N2839, j202_soc_core_j22_cpu_rf_N2838,
         j202_soc_core_j22_cpu_rf_N2837, j202_soc_core_j22_cpu_rf_N2836,
         j202_soc_core_j22_cpu_rf_N2835, j202_soc_core_j22_cpu_rf_N2834,
         j202_soc_core_j22_cpu_rf_N2832, j202_soc_core_j22_cpu_rf_N2831,
         j202_soc_core_j22_cpu_rf_N2830, j202_soc_core_j22_cpu_rf_N2829,
         j202_soc_core_j22_cpu_rf_N2828, j202_soc_core_j22_cpu_rf_N2827,
         j202_soc_core_j22_cpu_rf_N2826, j202_soc_core_j22_cpu_rf_N2824,
         j202_soc_core_j22_cpu_rf_N2823, j202_soc_core_j22_cpu_rf_N2822,
         j202_soc_core_j22_cpu_rf_N2821, j202_soc_core_j22_cpu_rf_N2820,
         j202_soc_core_j22_cpu_rf_N2819, j202_soc_core_j22_cpu_rf_N2818,
         j202_soc_core_j22_cpu_rf_N2817, j202_soc_core_j22_cpu_rf_N2816,
         j202_soc_core_j22_cpu_rf_N2815, j202_soc_core_j22_cpu_rf_N2814,
         j202_soc_core_j22_cpu_rf_N2813, j202_soc_core_j22_cpu_rf_N2811,
         j202_soc_core_j22_cpu_rf_N2810, j202_soc_core_j22_cpu_rf_N2809,
         j202_soc_core_j22_cpu_rf_N2808, j202_soc_core_j22_cpu_rf_N2807,
         j202_soc_core_j22_cpu_rf_N2806, j202_soc_core_j22_cpu_rf_N2805,
         j202_soc_core_j22_cpu_rf_N2803, j202_soc_core_j22_cpu_rf_N2802,
         j202_soc_core_j22_cpu_rf_N2801, j202_soc_core_j22_cpu_rf_N2800,
         j202_soc_core_j22_cpu_rf_N2799, j202_soc_core_j22_cpu_rf_N2798,
         j202_soc_core_j22_cpu_rf_N2797, j202_soc_core_j22_cpu_rf_N2795,
         j202_soc_core_j22_cpu_rf_N2794, j202_soc_core_j22_cpu_rf_N2793,
         j202_soc_core_j22_cpu_rf_N2792, j202_soc_core_j22_cpu_rf_N2791,
         j202_soc_core_j22_cpu_rf_N2790, j202_soc_core_j22_cpu_rf_N2789,
         j202_soc_core_j22_cpu_rf_N2787, j202_soc_core_j22_cpu_rf_N2786,
         j202_soc_core_j22_cpu_rf_N2785, j202_soc_core_j22_cpu_rf_N2784,
         j202_soc_core_j22_cpu_rf_N2783, j202_soc_core_j22_cpu_rf_N2782,
         j202_soc_core_j22_cpu_rf_N2781, j202_soc_core_j22_cpu_rf_N2780,
         j202_soc_core_j22_cpu_rf_N2779, j202_soc_core_j22_cpu_rf_N2778,
         j202_soc_core_j22_cpu_rf_N2777, j202_soc_core_j22_cpu_rf_N2776,
         j202_soc_core_j22_cpu_rf_N2774, j202_soc_core_j22_cpu_rf_N2773,
         j202_soc_core_j22_cpu_rf_N2772, j202_soc_core_j22_cpu_rf_N2771,
         j202_soc_core_j22_cpu_rf_N2770, j202_soc_core_j22_cpu_rf_N2769,
         j202_soc_core_j22_cpu_rf_N2768, j202_soc_core_j22_cpu_rf_N2766,
         j202_soc_core_j22_cpu_rf_N2765, j202_soc_core_j22_cpu_rf_N2764,
         j202_soc_core_j22_cpu_rf_N2763, j202_soc_core_j22_cpu_rf_N2762,
         j202_soc_core_j22_cpu_rf_N2761, j202_soc_core_j22_cpu_rf_N2760,
         j202_soc_core_j22_cpu_rf_N2758, j202_soc_core_j22_cpu_rf_N2757,
         j202_soc_core_j22_cpu_rf_N2756, j202_soc_core_j22_cpu_rf_N2755,
         j202_soc_core_j22_cpu_rf_N2754, j202_soc_core_j22_cpu_rf_N2753,
         j202_soc_core_j22_cpu_rf_N2752, j202_soc_core_j22_cpu_rf_N2750,
         j202_soc_core_j22_cpu_rf_N2749, j202_soc_core_j22_cpu_rf_N2748,
         j202_soc_core_j22_cpu_rf_N2747, j202_soc_core_j22_cpu_rf_N2746,
         j202_soc_core_j22_cpu_rf_N2745, j202_soc_core_j22_cpu_rf_N2744,
         j202_soc_core_j22_cpu_rf_N2743, j202_soc_core_j22_cpu_rf_N2742,
         j202_soc_core_j22_cpu_rf_N2741, j202_soc_core_j22_cpu_rf_N2740,
         j202_soc_core_j22_cpu_rf_N2739, j202_soc_core_j22_cpu_rf_N2737,
         j202_soc_core_j22_cpu_rf_N2736, j202_soc_core_j22_cpu_rf_N2735,
         j202_soc_core_j22_cpu_rf_N2734, j202_soc_core_j22_cpu_rf_N2733,
         j202_soc_core_j22_cpu_rf_N2732, j202_soc_core_j22_cpu_rf_N2731,
         j202_soc_core_j22_cpu_rf_N2729, j202_soc_core_j22_cpu_rf_N2728,
         j202_soc_core_j22_cpu_rf_N2727, j202_soc_core_j22_cpu_rf_N2726,
         j202_soc_core_j22_cpu_rf_N2725, j202_soc_core_j22_cpu_rf_N2724,
         j202_soc_core_j22_cpu_rf_N2723, j202_soc_core_j22_cpu_rf_N2721,
         j202_soc_core_j22_cpu_rf_N2720, j202_soc_core_j22_cpu_rf_N2719,
         j202_soc_core_j22_cpu_rf_N2718, j202_soc_core_j22_cpu_rf_N2717,
         j202_soc_core_j22_cpu_rf_N2716, j202_soc_core_j22_cpu_rf_N2715,
         j202_soc_core_j22_cpu_rf_N2713, j202_soc_core_j22_cpu_rf_N2712,
         j202_soc_core_j22_cpu_rf_N2711, j202_soc_core_j22_cpu_rf_N2710,
         j202_soc_core_j22_cpu_rf_N2709, j202_soc_core_j22_cpu_rf_N2708,
         j202_soc_core_j22_cpu_rf_N2707, j202_soc_core_j22_cpu_rf_N2706,
         j202_soc_core_j22_cpu_rf_N2705, j202_soc_core_j22_cpu_rf_N2704,
         j202_soc_core_j22_cpu_rf_N2703, j202_soc_core_j22_cpu_rf_N2702,
         j202_soc_core_j22_cpu_rf_N2700, j202_soc_core_j22_cpu_rf_N2699,
         j202_soc_core_j22_cpu_rf_N2698, j202_soc_core_j22_cpu_rf_N2697,
         j202_soc_core_j22_cpu_rf_N2696, j202_soc_core_j22_cpu_rf_N2695,
         j202_soc_core_j22_cpu_rf_N2694, j202_soc_core_j22_cpu_rf_N2692,
         j202_soc_core_j22_cpu_rf_N2691, j202_soc_core_j22_cpu_rf_N2690,
         j202_soc_core_j22_cpu_rf_N2689, j202_soc_core_j22_cpu_rf_N2688,
         j202_soc_core_j22_cpu_rf_N2687, j202_soc_core_j22_cpu_rf_N2686,
         j202_soc_core_j22_cpu_rf_N2684, j202_soc_core_j22_cpu_rf_N2683,
         j202_soc_core_j22_cpu_rf_N2682, j202_soc_core_j22_cpu_rf_N2681,
         j202_soc_core_j22_cpu_rf_N2680, j202_soc_core_j22_cpu_rf_N2679,
         j202_soc_core_j22_cpu_rf_N2678, j202_soc_core_j22_cpu_rf_N2676,
         j202_soc_core_j22_cpu_rf_N2670, j202_soc_core_j22_cpu_rf_N2668,
         j202_soc_core_j22_cpu_rf_N2658, j202_soc_core_j22_cpu_rf_N2657,
         j202_soc_core_j22_cpu_rf_N2656, j202_soc_core_j22_cpu_rf_N2655,
         j202_soc_core_j22_cpu_rf_N2654, j202_soc_core_j22_cpu_rf_N2653,
         j202_soc_core_j22_cpu_rf_N2652, j202_soc_core_j22_cpu_rf_N2651,
         j202_soc_core_j22_cpu_rf_N2649, j202_soc_core_j22_cpu_rf_N2648,
         j202_soc_core_j22_cpu_rf_N2647, j202_soc_core_j22_cpu_rf_N2646,
         j202_soc_core_j22_cpu_rf_N2645, j202_soc_core_j22_cpu_rf_N2644,
         j202_soc_core_j22_cpu_rf_N2643, j202_soc_core_j22_cpu_rf_N2642,
         j202_soc_core_j22_cpu_rf_N2640, j202_soc_core_j22_cpu_rf_N2639,
         j202_soc_core_j22_cpu_rf_N2638, j202_soc_core_j22_cpu_rf_N2637,
         j202_soc_core_j22_cpu_rf_N2628, j202_soc_core_j22_cpu_rf_N2627,
         j202_soc_core_j22_cpu_rf_N2626, j202_soc_core_j22_cpu_rf_N2625,
         j202_soc_core_j22_cpu_rf_N328, j202_soc_core_j22_cpu_rf_N327,
         j202_soc_core_j22_cpu_rf_N326, j202_soc_core_j22_cpu_rf_N325,
         j202_soc_core_j22_cpu_rf_N324, j202_soc_core_j22_cpu_rf_N323,
         j202_soc_core_j22_cpu_rf_N322, j202_soc_core_j22_cpu_rf_N321,
         j202_soc_core_j22_cpu_rf_N320, j202_soc_core_j22_cpu_rf_N319,
         j202_soc_core_j22_cpu_rf_N318, j202_soc_core_j22_cpu_rf_N317,
         j202_soc_core_j22_cpu_rf_N316, j202_soc_core_j22_cpu_rf_N315,
         j202_soc_core_j22_cpu_rf_N314, j202_soc_core_j22_cpu_rf_N313,
         j202_soc_core_j22_cpu_rf_N312, j202_soc_core_j22_cpu_rf_N311,
         j202_soc_core_j22_cpu_rf_N310, j202_soc_core_j22_cpu_rf_N309,
         j202_soc_core_j22_cpu_rf_N308, j202_soc_core_j22_cpu_rf_N307,
         j202_soc_core_j22_cpu_rf_N306, j202_soc_core_j22_cpu_rf_N305,
         j202_soc_core_j22_cpu_rf_N304, j202_soc_core_j22_cpu_rf_N303,
         j202_soc_core_j22_cpu_rf_N302, j202_soc_core_j22_cpu_rf_N301,
         j202_soc_core_j22_cpu_rf_N300, j202_soc_core_j22_cpu_rf_N299,
         j202_soc_core_j22_cpu_rf_N298, j202_soc_core_j22_cpu_ma_N56,
         j202_soc_core_j22_cpu_ma_N55, j202_soc_core_j22_cpu_ma_N54,
         j202_soc_core_j22_cpu_ma_N53, j202_soc_core_j22_cpu_ml_N429,
         j202_soc_core_j22_cpu_ml_N428, j202_soc_core_j22_cpu_ml_N427,
         j202_soc_core_j22_cpu_ml_N426, j202_soc_core_j22_cpu_ml_N425,
         j202_soc_core_j22_cpu_ml_N424, j202_soc_core_j22_cpu_ml_N423,
         j202_soc_core_j22_cpu_ml_N422, j202_soc_core_j22_cpu_ml_N421,
         j202_soc_core_j22_cpu_ml_N420, j202_soc_core_j22_cpu_ml_N419,
         j202_soc_core_j22_cpu_ml_N418, j202_soc_core_j22_cpu_ml_N417,
         j202_soc_core_j22_cpu_ml_N416, j202_soc_core_j22_cpu_ml_N415,
         j202_soc_core_j22_cpu_ml_N414, j202_soc_core_j22_cpu_ml_N413,
         j202_soc_core_j22_cpu_ml_N412, j202_soc_core_j22_cpu_ml_N370,
         j202_soc_core_j22_cpu_ml_N369, j202_soc_core_j22_cpu_ml_N368,
         j202_soc_core_j22_cpu_ml_N367, j202_soc_core_j22_cpu_ml_N366,
         j202_soc_core_j22_cpu_ml_N365, j202_soc_core_j22_cpu_ml_N364,
         j202_soc_core_j22_cpu_ml_N363, j202_soc_core_j22_cpu_ml_N362,
         j202_soc_core_j22_cpu_ml_N361, j202_soc_core_j22_cpu_ml_N360,
         j202_soc_core_j22_cpu_ml_N359, j202_soc_core_j22_cpu_ml_N357,
         j202_soc_core_j22_cpu_ml_N356, j202_soc_core_j22_cpu_ml_N355,
         j202_soc_core_j22_cpu_ml_N354, j202_soc_core_j22_cpu_ml_N336,
         j202_soc_core_j22_cpu_ml_N335, j202_soc_core_j22_cpu_ml_N334,
         j202_soc_core_j22_cpu_ml_N333, j202_soc_core_j22_cpu_ml_N332,
         j202_soc_core_j22_cpu_ml_N331, j202_soc_core_j22_cpu_ml_N330,
         j202_soc_core_j22_cpu_ml_N329, j202_soc_core_j22_cpu_ml_N328,
         j202_soc_core_j22_cpu_ml_N327, j202_soc_core_j22_cpu_ml_N326,
         j202_soc_core_j22_cpu_ml_N325, j202_soc_core_j22_cpu_ml_N324,
         j202_soc_core_j22_cpu_ml_N322, j202_soc_core_j22_cpu_ml_N321,
         j202_soc_core_j22_cpu_ml_N320, j202_soc_core_j22_cpu_ml_N319,
         j202_soc_core_j22_cpu_ml_N318, j202_soc_core_j22_cpu_ml_N317,
         j202_soc_core_j22_cpu_ml_N316, j202_soc_core_j22_cpu_ml_N315,
         j202_soc_core_j22_cpu_ml_N314, j202_soc_core_j22_cpu_ml_N313,
         j202_soc_core_j22_cpu_ml_N312, j202_soc_core_j22_cpu_ml_N311,
         j202_soc_core_j22_cpu_ml_N310, j202_soc_core_j22_cpu_ml_N309,
         j202_soc_core_j22_cpu_ml_N308, j202_soc_core_j22_cpu_ml_N307,
         j202_soc_core_j22_cpu_ml_N306, j202_soc_core_j22_cpu_ml_N305,
         j202_soc_core_j22_cpu_ml_N304, j202_soc_core_j22_cpu_ml_N303,
         j202_soc_core_j22_cpu_ml_N195, j202_soc_core_j22_cpu_ml_N194,
         j202_soc_core_j22_cpu_ml_N193, j202_soc_core_j22_cpu_ml_N192,
         j202_soc_core_j22_cpu_ml_N191, j202_soc_core_j22_cpu_ml_N156,
         j202_soc_core_j22_cpu_ml_N155, j202_soc_core_j22_cpu_ml_N154,
         j202_soc_core_j22_cpu_ml_N153, j202_soc_core_j22_cpu_ml_N152,
         j202_soc_core_ahb2apb_00_N143, j202_soc_core_ahb2apb_00_N142,
         j202_soc_core_ahb2apb_00_N141, j202_soc_core_ahb2apb_00_N140,
         j202_soc_core_ahb2apb_00_N139, j202_soc_core_ahb2apb_00_N138,
         j202_soc_core_ahb2apb_00_N137, j202_soc_core_ahb2apb_00_N136,
         j202_soc_core_ahb2apb_00_N135, j202_soc_core_ahb2apb_00_N134,
         j202_soc_core_ahb2apb_00_N133, j202_soc_core_ahb2apb_00_N132,
         j202_soc_core_ahb2apb_00_N131, j202_soc_core_ahb2apb_00_N130,
         j202_soc_core_ahb2apb_00_N129, j202_soc_core_ahb2apb_00_N128,
         j202_soc_core_ahb2apb_00_N127, j202_soc_core_cmt_core_00_cmf1,
         j202_soc_core_cmt_core_00_cmf0, j202_soc_core_cmt_core_00_str1,
         j202_soc_core_cmt_core_00_str0,
         j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_2,
         j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_1,
         j202_soc_core_cmt_core_00_cmt_apb_00_nxt_state_0_,
         j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen,
         j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_nxt_latch_status_0_,
         j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_0_,
         j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_nxt_latch_status_0_,
         j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_0_,
         j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt1_to1,
         j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt0_to1,
         j202_soc_core_ahb2apb_01_N159, j202_soc_core_ahb2apb_01_N158,
         j202_soc_core_ahb2apb_01_N157, j202_soc_core_ahb2apb_01_N156,
         j202_soc_core_ahb2apb_01_N155, j202_soc_core_ahb2apb_01_N154,
         j202_soc_core_ahb2apb_01_N153, j202_soc_core_ahb2apb_01_N152,
         j202_soc_core_ahb2apb_01_N151, j202_soc_core_ahb2apb_01_N150,
         j202_soc_core_ahb2apb_01_N149, j202_soc_core_ahb2apb_01_N148,
         j202_soc_core_ahb2apb_01_N147, j202_soc_core_ahb2apb_01_N146,
         j202_soc_core_ahb2apb_01_N145, j202_soc_core_ahb2apb_01_N144,
         j202_soc_core_ahb2apb_01_N143, j202_soc_core_ahb2apb_01_N142,
         j202_soc_core_ahb2apb_01_N141, j202_soc_core_ahb2apb_01_N140,
         j202_soc_core_ahb2apb_01_N139, j202_soc_core_ahb2apb_01_N138,
         j202_soc_core_ahb2apb_01_N137, j202_soc_core_ahb2apb_01_N136,
         j202_soc_core_ahb2apb_01_N135, j202_soc_core_ahb2apb_01_N134,
         j202_soc_core_ahb2apb_01_N133, j202_soc_core_ahb2apb_01_N132,
         j202_soc_core_ahb2apb_01_N131, j202_soc_core_ahb2apb_01_N130,
         j202_soc_core_ahb2apb_01_N129, j202_soc_core_ahb2apb_01_N128,
         j202_soc_core_ahb2apb_01_N123, j202_soc_core_ahb2apb_01_N91,
         j202_soc_core_ahb2apb_01_N90, j202_soc_core_ahb2apb_01_N89,
         j202_soc_core_ahb2apb_01_N57, j202_soc_core_ahb2apb_01_N56,
         j202_soc_core_ahb2apb_01_N55, j202_soc_core_ahb2apb_01_N34,
         j202_soc_core_ahb2apb_01_N33, j202_soc_core_ahb2apb_01_N32,
         j202_soc_core_ahb2apb_01_N31, j202_soc_core_ahb2apb_01_N30,
         j202_soc_core_ahb2apb_01_N29, j202_soc_core_ahb2apb_01_N28,
         j202_soc_core_ahb2apb_01_N27, j202_soc_core_ahb2apb_01_N26,
         j202_soc_core_ahb2apb_01_N25, j202_soc_core_ahb2apb_01_N24,
         j202_soc_core_ahb2apb_01_N23,
         j202_soc_core_intc_core_00_cp_intack_all_0_,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_0__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_1__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_2__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_3__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_4__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_5__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_6__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_7__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_8__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_9__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_10__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_11__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_12__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_13__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_14__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_15__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N23,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N22,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N21,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N20,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N19,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N18,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N17,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N16,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N15,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N14,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N13,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N12,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N11,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N10,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N9,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N8,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N7,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N6,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N5,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N4,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N23,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N22,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N21,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N20,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N18,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N17,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N16,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N15,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N14,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N13,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N12,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N11,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N10,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N9,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N8,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N7,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N6,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N5,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N4,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N3,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_req_N3,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N6,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N5,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N4,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N3,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N6,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N5,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N4,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N3,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N9,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N7,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N6,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N5,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N4,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N3,
         j202_soc_core_ahb2apb_02_N159, j202_soc_core_ahb2apb_02_N158,
         j202_soc_core_ahb2apb_02_N157, j202_soc_core_ahb2apb_02_N156,
         j202_soc_core_ahb2apb_02_N155, j202_soc_core_ahb2apb_02_N154,
         j202_soc_core_ahb2apb_02_N153, j202_soc_core_ahb2apb_02_N152,
         j202_soc_core_ahb2apb_02_N151, j202_soc_core_ahb2apb_02_N150,
         j202_soc_core_ahb2apb_02_N149, j202_soc_core_ahb2apb_02_N148,
         j202_soc_core_ahb2apb_02_N147, j202_soc_core_ahb2apb_02_N146,
         j202_soc_core_ahb2apb_02_N145, j202_soc_core_ahb2apb_02_N144,
         j202_soc_core_ahb2apb_02_N143, j202_soc_core_ahb2apb_02_N142,
         j202_soc_core_ahb2apb_02_N141, j202_soc_core_ahb2apb_02_N140,
         j202_soc_core_ahb2apb_02_N139, j202_soc_core_ahb2apb_02_N138,
         j202_soc_core_ahb2apb_02_N137, j202_soc_core_ahb2apb_02_N136,
         j202_soc_core_ahb2apb_02_N135, j202_soc_core_ahb2apb_02_N134,
         j202_soc_core_ahb2apb_02_N133, j202_soc_core_ahb2apb_02_N132,
         j202_soc_core_ahb2apb_02_N131, j202_soc_core_ahb2apb_02_N130,
         j202_soc_core_ahb2apb_02_N129, j202_soc_core_ahb2apb_02_N128,
         j202_soc_core_ahb2apb_02_N127, j202_soc_core_ahb2apb_02_N123,
         j202_soc_core_ahb2apb_02_N89, j202_soc_core_ahb2apb_02_N57,
         j202_soc_core_ahb2apb_02_N56, j202_soc_core_ahb2apb_02_N55,
         j202_soc_core_ahb2apb_02_N30, j202_soc_core_ahb2apb_02_N29,
         j202_soc_core_ahb2apb_02_N28, j202_soc_core_ahb2apb_02_N27,
         j202_soc_core_ahb2apb_02_N26, j202_soc_core_ahb2apb_02_N25,
         j202_soc_core_ahb2apb_02_N24, j202_soc_core_ahb2apb_02_N23,
         j202_soc_core_ahb2apb_02_N22,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N34,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N33,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N32,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N31,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N30,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N29,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N28,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N27,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N26,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N25,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N24,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N23,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N22,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N21,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N20,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N19,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N18,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N17,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N16,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N15,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N14,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N13,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N12,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N11,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N10,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N9,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N8,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N7,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N6,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N5,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N4,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N3,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N71,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N70,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N69,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N68,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N67,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N66,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N65,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N64,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N63,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N62,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N61,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N60,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N59,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N58,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N57,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N56,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N55,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N54,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N53,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N52,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N51,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N50,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N49,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N48,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N47,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N46,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N45,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N44,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N43,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N42,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N41,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N40,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N34,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N33,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N32,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N28,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N26,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N24,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N23,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N22,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N20,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N19,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N15,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N14,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N13,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N12,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N11,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N7,
         j202_soc_core_ahb2aqu_00_N164, j202_soc_core_ahb2aqu_00_N163,
         j202_soc_core_ahb2aqu_00_N161, j202_soc_core_ahb2aqu_00_N128,
         j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N98,
         j202_soc_core_ahb2aqu_00_N97, j202_soc_core_ahb2aqu_00_N95,
         j202_soc_core_ahb2aqu_00_N93, j202_soc_core_ahb2aqu_00_aqu_st_0_,
         j202_soc_core_uart_sio_ce_x4, j202_soc_core_uart_sio_ce,
         j202_soc_core_uart_RDRXD1, j202_soc_core_uart_WRTXD1,
         j202_soc_core_uart_TOP_N137, j202_soc_core_uart_TOP_N128,
         j202_soc_core_uart_TOP_N123, j202_soc_core_uart_TOP_N118,
         j202_soc_core_uart_TOP_rx_sio_ce_r2,
         j202_soc_core_uart_TOP_rx_sio_ce_r1, j202_soc_core_uart_TOP_N102,
         j202_soc_core_uart_TOP_N101, j202_soc_core_uart_TOP_change,
         j202_soc_core_uart_TOP_N95, j202_soc_core_uart_TOP_rx_valid_r,
         j202_soc_core_uart_TOP_rx_valid, j202_soc_core_uart_TOP_N89,
         j202_soc_core_uart_TOP_N88, j202_soc_core_uart_TOP_N87,
         j202_soc_core_uart_TOP_N85, j202_soc_core_uart_TOP_rx_sio_ce,
         j202_soc_core_uart_TOP_rx_go, j202_soc_core_uart_TOP_rxd_r,
         j202_soc_core_uart_TOP_rxd_s, j202_soc_core_uart_TOP_N61,
         j202_soc_core_uart_TOP_N58, j202_soc_core_uart_TOP_N57,
         j202_soc_core_uart_TOP_N43, j202_soc_core_uart_TOP_shift_en_r,
         j202_soc_core_uart_TOP_N33, j202_soc_core_uart_TOP_N32,
         j202_soc_core_uart_TOP_N31, j202_soc_core_uart_TOP_N30,
         j202_soc_core_uart_TOP_N29, j202_soc_core_uart_TOP_N28,
         j202_soc_core_uart_TOP_N27, j202_soc_core_uart_TOP_N26,
         j202_soc_core_uart_TOP_N25, j202_soc_core_uart_TOP_N24,
         j202_soc_core_uart_TOP_load, j202_soc_core_uart_TOP_shift_en,
         j202_soc_core_uart_TOP_N16, j202_soc_core_uart_TOP_txf_empty_r,
         j202_soc_core_uart_TOP_tx_fifo_N42,
         j202_soc_core_uart_TOP_tx_fifo_N41, j202_soc_core_uart_TOP_tx_fifo_gb,
         j202_soc_core_uart_TOP_rx_fifo_N42,
         j202_soc_core_uart_TOP_rx_fifo_N41, j202_soc_core_uart_TOP_rx_fifo_gb,
         j202_soc_core_uart_BRG_N59, j202_soc_core_uart_BRG_sio_ce_r,
         j202_soc_core_uart_BRG_N57, j202_soc_core_uart_BRG_N55,
         j202_soc_core_uart_BRG_sio_ce_x4_t,
         j202_soc_core_uart_BRG_sio_ce_x4_r, j202_soc_core_uart_BRG_N47,
         j202_soc_core_uart_BRG_N42, j202_soc_core_uart_BRG_N41,
         j202_soc_core_uart_BRG_N40, j202_soc_core_uart_BRG_N39,
         j202_soc_core_uart_BRG_N38, j202_soc_core_uart_BRG_N37,
         j202_soc_core_uart_BRG_N36, j202_soc_core_uart_BRG_N35,
         j202_soc_core_uart_BRG_br_clr, j202_soc_core_uart_BRG_N21,
         j202_soc_core_uart_BRG_N19, j202_soc_core_uart_BRG_N18,
         j202_soc_core_uart_BRG_N17, j202_soc_core_uart_BRG_N16,
         j202_soc_core_uart_BRG_N15, j202_soc_core_uart_BRG_N14,
         j202_soc_core_uart_BRG_N13, j202_soc_core_uart_BRG_N12,
         j202_soc_core_uart_BRG_ps_clr, j202_soc_core_bldc_core_00_adc_en,
         j202_soc_core_bldc_core_00_pwm_en,
         j202_soc_core_bldc_core_00_bldc_wb_slave_00_nxt_state_1_,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_nxt_bldc_int,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_0_,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_wen,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_nxt_latch_status_0_,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_0_,
         j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_2,
         j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1,
         j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posc,
         j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_negb,
         j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posb,
         j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posa,
         j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld,
         j202_soc_core_ahb2wbqspi_00_stb_o, j202_soc_core_wbqspiflash_00_N750,
         j202_soc_core_wbqspiflash_00_N749, j202_soc_core_wbqspiflash_00_N747,
         j202_soc_core_wbqspiflash_00_N746, j202_soc_core_wbqspiflash_00_N745,
         j202_soc_core_wbqspiflash_00_N744, j202_soc_core_wbqspiflash_00_N743,
         j202_soc_core_wbqspiflash_00_N742, j202_soc_core_wbqspiflash_00_N741,
         j202_soc_core_wbqspiflash_00_N740, j202_soc_core_wbqspiflash_00_N739,
         j202_soc_core_wbqspiflash_00_N738, j202_soc_core_wbqspiflash_00_N737,
         j202_soc_core_wbqspiflash_00_N736, j202_soc_core_wbqspiflash_00_N735,
         j202_soc_core_wbqspiflash_00_N734, j202_soc_core_wbqspiflash_00_N733,
         j202_soc_core_wbqspiflash_00_N730, j202_soc_core_wbqspiflash_00_N729,
         j202_soc_core_wbqspiflash_00_N728, j202_soc_core_wbqspiflash_00_N727,
         j202_soc_core_wbqspiflash_00_N726, j202_soc_core_wbqspiflash_00_N725,
         j202_soc_core_wbqspiflash_00_N724, j202_soc_core_wbqspiflash_00_N723,
         j202_soc_core_wbqspiflash_00_N722, j202_soc_core_wbqspiflash_00_N721,
         j202_soc_core_wbqspiflash_00_N720, j202_soc_core_wbqspiflash_00_N719,
         j202_soc_core_wbqspiflash_00_N718, j202_soc_core_wbqspiflash_00_N717,
         j202_soc_core_wbqspiflash_00_N716, j202_soc_core_wbqspiflash_00_N715,
         j202_soc_core_wbqspiflash_00_N714, j202_soc_core_wbqspiflash_00_N713,
         j202_soc_core_wbqspiflash_00_N712, j202_soc_core_wbqspiflash_00_N711,
         j202_soc_core_wbqspiflash_00_N710, j202_soc_core_wbqspiflash_00_N709,
         j202_soc_core_wbqspiflash_00_N708, j202_soc_core_wbqspiflash_00_N698,
         j202_soc_core_wbqspiflash_00_N697, j202_soc_core_wbqspiflash_00_N696,
         j202_soc_core_wbqspiflash_00_N695, j202_soc_core_wbqspiflash_00_N694,
         j202_soc_core_wbqspiflash_00_N688, j202_soc_core_wbqspiflash_00_N687,
         j202_soc_core_wbqspiflash_00_N686, j202_soc_core_wbqspiflash_00_N685,
         j202_soc_core_wbqspiflash_00_N684, j202_soc_core_wbqspiflash_00_N683,
         j202_soc_core_wbqspiflash_00_N682, j202_soc_core_wbqspiflash_00_N681,
         j202_soc_core_wbqspiflash_00_N674, j202_soc_core_wbqspiflash_00_N673,
         j202_soc_core_wbqspiflash_00_N672, j202_soc_core_wbqspiflash_00_N671,
         j202_soc_core_wbqspiflash_00_N670, j202_soc_core_wbqspiflash_00_N669,
         j202_soc_core_wbqspiflash_00_N668, j202_soc_core_wbqspiflash_00_N667,
         j202_soc_core_wbqspiflash_00_N663, j202_soc_core_wbqspiflash_00_N629,
         j202_soc_core_wbqspiflash_00_N628, j202_soc_core_wbqspiflash_00_N623,
         j202_soc_core_wbqspiflash_00_N622, j202_soc_core_wbqspiflash_00_N621,
         j202_soc_core_wbqspiflash_00_N620, j202_soc_core_wbqspiflash_00_N619,
         j202_soc_core_wbqspiflash_00_N618, j202_soc_core_wbqspiflash_00_N617,
         j202_soc_core_wbqspiflash_00_N616, j202_soc_core_wbqspiflash_00_N615,
         j202_soc_core_wbqspiflash_00_N614, j202_soc_core_wbqspiflash_00_N613,
         j202_soc_core_wbqspiflash_00_N612, j202_soc_core_wbqspiflash_00_N611,
         j202_soc_core_wbqspiflash_00_N609, j202_soc_core_wbqspiflash_00_N608,
         j202_soc_core_wbqspiflash_00_N607, j202_soc_core_wbqspiflash_00_N606,
         j202_soc_core_wbqspiflash_00_N605, j202_soc_core_wbqspiflash_00_N594,
         j202_soc_core_wbqspiflash_00_N592, j202_soc_core_wbqspiflash_00_N590,
         j202_soc_core_wbqspiflash_00_spif_cmd,
         j202_soc_core_wbqspiflash_00_spif_req,
         j202_soc_core_wbqspiflash_00_N86,
         j202_soc_core_wbqspiflash_00_alt_ctrl,
         j202_soc_core_wbqspiflash_00_N85,
         j202_soc_core_wbqspiflash_00_alt_cmd,
         j202_soc_core_wbqspiflash_00_spif_ctrl,
         j202_soc_core_wbqspiflash_00_spif_override,
         j202_soc_core_wbqspiflash_00_quad_mode_enabled,
         j202_soc_core_wbqspiflash_00_write_protect,
         j202_soc_core_wbqspiflash_00_dirty_sector,
         j202_soc_core_wbqspiflash_00_write_in_progress,
         j202_soc_core_wbqspiflash_00_w_qspi_cs_n,
         j202_soc_core_wbqspiflash_00_w_qspi_sck,
         j202_soc_core_wbqspiflash_00_spi_busy,
         j202_soc_core_wbqspiflash_00_spi_valid,
         j202_soc_core_wbqspiflash_00_spi_dir,
         j202_soc_core_wbqspiflash_00_spi_spd,
         j202_soc_core_wbqspiflash_00_spi_hold,
         j202_soc_core_wbqspiflash_00_spi_wr,
         j202_soc_core_wbqspiflash_00_lldriver_N430,
         j202_soc_core_wbqspiflash_00_lldriver_N429,
         j202_soc_core_wbqspiflash_00_lldriver_N428,
         j202_soc_core_wbqspiflash_00_lldriver_N427,
         j202_soc_core_wbqspiflash_00_lldriver_N426,
         j202_soc_core_wbqspiflash_00_lldriver_N425,
         j202_soc_core_wbqspiflash_00_lldriver_N424,
         j202_soc_core_wbqspiflash_00_lldriver_N423,
         j202_soc_core_wbqspiflash_00_lldriver_N422,
         j202_soc_core_wbqspiflash_00_lldriver_N421,
         j202_soc_core_wbqspiflash_00_lldriver_N420,
         j202_soc_core_wbqspiflash_00_lldriver_N419,
         j202_soc_core_wbqspiflash_00_lldriver_N418,
         j202_soc_core_wbqspiflash_00_lldriver_N417,
         j202_soc_core_wbqspiflash_00_lldriver_N416,
         j202_soc_core_wbqspiflash_00_lldriver_N415,
         j202_soc_core_wbqspiflash_00_lldriver_N414,
         j202_soc_core_wbqspiflash_00_lldriver_N413,
         j202_soc_core_wbqspiflash_00_lldriver_N412,
         j202_soc_core_wbqspiflash_00_lldriver_N411,
         j202_soc_core_wbqspiflash_00_lldriver_N410,
         j202_soc_core_wbqspiflash_00_lldriver_N409,
         j202_soc_core_wbqspiflash_00_lldriver_N408,
         j202_soc_core_wbqspiflash_00_lldriver_N407,
         j202_soc_core_wbqspiflash_00_lldriver_N406,
         j202_soc_core_wbqspiflash_00_lldriver_N405,
         j202_soc_core_wbqspiflash_00_lldriver_N404,
         j202_soc_core_wbqspiflash_00_lldriver_N403,
         j202_soc_core_wbqspiflash_00_lldriver_N402,
         j202_soc_core_wbqspiflash_00_lldriver_N401,
         j202_soc_core_wbqspiflash_00_lldriver_N400,
         j202_soc_core_wbqspiflash_00_lldriver_N399,
         j202_soc_core_wbqspiflash_00_lldriver_N398,
         j202_soc_core_wbqspiflash_00_lldriver_N397,
         j202_soc_core_wbqspiflash_00_lldriver_N396,
         j202_soc_core_wbqspiflash_00_lldriver_N395,
         j202_soc_core_wbqspiflash_00_lldriver_N394,
         j202_soc_core_wbqspiflash_00_lldriver_N393,
         j202_soc_core_wbqspiflash_00_lldriver_N392,
         j202_soc_core_wbqspiflash_00_lldriver_N391,
         j202_soc_core_wbqspiflash_00_lldriver_N390,
         j202_soc_core_wbqspiflash_00_lldriver_N389,
         j202_soc_core_wbqspiflash_00_lldriver_N361,
         j202_soc_core_wbqspiflash_00_lldriver_N360,
         j202_soc_core_wbqspiflash_00_lldriver_N359,
         j202_soc_core_wbqspiflash_00_lldriver_N358,
         j202_soc_core_wbqspiflash_00_lldriver_N356,
         j202_soc_core_wbqspiflash_00_lldriver_N355,
         j202_soc_core_wbqspiflash_00_lldriver_N354,
         j202_soc_core_wbqspiflash_00_lldriver_N353,
         j202_soc_core_wbqspiflash_00_lldriver_N352,
         j202_soc_core_wbqspiflash_00_lldriver_N351,
         j202_soc_core_wbqspiflash_00_lldriver_N350,
         j202_soc_core_wbqspiflash_00_lldriver_N349,
         j202_soc_core_wbqspiflash_00_lldriver_N348,
         j202_soc_core_wbqspiflash_00_lldriver_N347,
         j202_soc_core_wbqspiflash_00_lldriver_N346,
         j202_soc_core_wbqspiflash_00_lldriver_N345,
         j202_soc_core_wbqspiflash_00_lldriver_N344,
         j202_soc_core_wbqspiflash_00_lldriver_N343,
         j202_soc_core_wbqspiflash_00_lldriver_N342,
         j202_soc_core_wbqspiflash_00_lldriver_N341,
         j202_soc_core_wbqspiflash_00_lldriver_N340,
         j202_soc_core_wbqspiflash_00_lldriver_N339,
         j202_soc_core_wbqspiflash_00_lldriver_N338,
         j202_soc_core_wbqspiflash_00_lldriver_N337,
         j202_soc_core_wbqspiflash_00_lldriver_N336,
         j202_soc_core_wbqspiflash_00_lldriver_N335,
         j202_soc_core_wbqspiflash_00_lldriver_N334,
         j202_soc_core_wbqspiflash_00_lldriver_N333,
         j202_soc_core_wbqspiflash_00_lldriver_N332,
         j202_soc_core_wbqspiflash_00_lldriver_N331,
         j202_soc_core_wbqspiflash_00_lldriver_N330,
         j202_soc_core_wbqspiflash_00_lldriver_N329,
         j202_soc_core_wbqspiflash_00_lldriver_N328,
         j202_soc_core_wbqspiflash_00_lldriver_N327,
         j202_soc_core_wbqspiflash_00_lldriver_N326,
         j202_soc_core_wbqspiflash_00_lldriver_N325,
         j202_soc_core_wbqspiflash_00_lldriver_N324,
         j202_soc_core_wbqspiflash_00_lldriver_N323,
         j202_soc_core_wbqspiflash_00_lldriver_N321,
         j202_soc_core_wbqspiflash_00_lldriver_N319,
         j202_soc_core_wbqspiflash_00_lldriver_N318,
         j202_soc_core_wbqspiflash_00_lldriver_N317,
         j202_soc_core_wbqspiflash_00_lldriver_N316,
         j202_soc_core_wbqspiflash_00_lldriver_N315,
         j202_soc_core_wbqspiflash_00_lldriver_N314,
         j202_soc_core_wbqspiflash_00_lldriver_N313,
         j202_soc_core_wbqspiflash_00_lldriver_N312,
         j202_soc_core_wbqspiflash_00_lldriver_N311,
         j202_soc_core_wbqspiflash_00_lldriver_N309,
         j202_soc_core_wbqspiflash_00_lldriver_N308,
         j202_soc_core_wbqspiflash_00_lldriver_N307,
         j202_soc_core_wbqspiflash_00_lldriver_r_dir,
         j202_soc_core_wbqspiflash_00_lldriver_r_spd,
         j202_soc_core_bootrom_00_sel_w, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10577, n10578,
         n10579, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10599, n10600, n10601, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10624, n10625, n10626, n10627, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10643, n10644, n10645, n10646, n10651, n10655, n10711,
         n10712, n10714, n10716, n10717, n10783, n10784, n10785, n10786,
         n10942, n10943, n10944, n10945, n10949, DP_OP_1508J1_126_2326_n3,
         DP_OP_1508J1_126_2326_n4, DP_OP_1508J1_126_2326_n6,
         U7_RSOP_1495_C3_DATA3_2, n10957, n10958, n10959, n10960, n10962,
         n10965, n10966, n10967, n10968, n10969, n10971, n10972, n10975,
         n10976, n10977, n10978, n10979, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10998, n11000, n11001, n11002, n11005, n11006,
         n11007, n11008, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11036, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11118,
         n11119, n11120, n11121, n11123, n11124, n11125, n11127, n11129,
         n11130, n11131, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11207, n11208, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11375, n11377, n11378, n11379, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11394, n11395, n11396, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11497, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11522, n11523, n11524, n11525, n11528, n11529, n11530,
         n11531, n11532, n11533, n11535, n11536, n11537, n11538, n11540,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11586, n11587, n11588, n11589, n11590, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11641, n11642,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11721, n11722, n11723, n11724, n11725, n11726, n11728,
         n11729, n11730, n11731, n11732, n11733, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11894, n11895, n11896, n11900, n11901,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11978, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12063, n12064, n12065, n12066, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12295, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12321, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12461,
         n12462, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12574, n12575, n12576, n12577,
         n12578, n12579, n12581, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12778, n12779, n12780, n12781, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12853, n12854, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18504, n18505, n18506,
         n18507, n18508, n18509, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
         n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
         n20945, n20946, n20947, n20948, n20949, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
         n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
         n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
         n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
         n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
         n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
         n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
         n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372,
         n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
         n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
         n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396,
         n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404,
         n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
         n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
         n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428,
         n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
         n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444,
         n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
         n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
         n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468,
         n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
         n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
         n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492,
         n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500,
         n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508,
         n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516,
         n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524,
         n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
         n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540,
         n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548,
         n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
         n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564,
         n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
         n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580,
         n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588,
         n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
         n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
         n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
         n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
         n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
         n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
         n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660,
         n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
         n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
         n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684,
         n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
         n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700,
         n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708,
         n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716,
         n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724,
         n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732,
         n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
         n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
         n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756,
         n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764,
         n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772,
         n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780,
         n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788,
         n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796,
         n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804,
         n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
         n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
         n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828,
         n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836,
         n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844,
         n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852,
         n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
         n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868,
         n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876,
         n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884,
         n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
         n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900,
         n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908,
         n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
         n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924,
         n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932,
         n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940,
         n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948,
         n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956,
         n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
         n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972,
         n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980,
         n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
         n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996,
         n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
         n22005, n22007, n22008, n22009, n22010, n22011, n22012, n22013,
         n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021,
         n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029,
         n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037,
         n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045,
         n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053,
         n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061,
         n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069,
         n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077,
         n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085,
         n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093,
         n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101,
         n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109,
         n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117,
         n22118, n22120, n22121, n22122, n22123, n22124, n22125, n22126,
         n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134,
         n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142,
         n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150,
         n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158,
         n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166,
         n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174,
         n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182,
         n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190,
         n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198,
         n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206,
         n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214,
         n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222,
         n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230,
         n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238,
         n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246,
         n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254,
         n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262,
         n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270,
         n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278,
         n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286,
         n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294,
         n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302,
         n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310,
         n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318,
         n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326,
         n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334,
         n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342,
         n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350,
         n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358,
         n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366,
         n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374,
         n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382,
         n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390,
         n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398,
         n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406,
         n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414,
         n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422,
         n22423, n22424, n22425, n22427, n22428, n22429, n22430, n22431,
         n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439,
         n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
         n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455,
         n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463,
         n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
         n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479,
         n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487,
         n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495,
         n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503,
         n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511,
         n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519,
         n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527,
         n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535,
         n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543,
         n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551,
         n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559,
         n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567,
         n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575,
         n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583,
         n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591,
         n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599,
         n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607,
         n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615,
         n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623,
         n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631,
         n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639,
         n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647,
         n22648, n22649, n22650, n22651, n22653, n22654, n22655, n22656,
         n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664,
         n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672,
         n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680,
         n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688,
         n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696,
         n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704,
         n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712,
         n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720,
         n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728,
         n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736,
         n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744,
         n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752,
         n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760,
         n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768,
         n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776,
         n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784,
         n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792,
         n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800,
         n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808,
         n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816,
         n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824,
         n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832,
         n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840,
         n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848,
         n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856,
         n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864,
         n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872,
         n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880,
         n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888,
         n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896,
         n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904,
         n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912,
         n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920,
         n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928,
         n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936,
         n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944,
         n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952,
         n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960,
         n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968,
         n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976,
         n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984,
         n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992,
         n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000,
         n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008,
         n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016,
         n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024,
         n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032,
         n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040,
         n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048,
         n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056,
         n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064,
         n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072,
         n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080,
         n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088,
         n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096,
         n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104,
         n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112,
         n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120,
         n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128,
         n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136,
         n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144,
         n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152,
         n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160,
         n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168,
         n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176,
         n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184,
         n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192,
         n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200,
         n23201, n23202, n23203, n23204, n23205, n23208, n23209, n23210,
         n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218,
         n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226,
         n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234,
         n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242,
         n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250,
         n23251, n23252, n23254, n23255, n23256, n23257, n23258, n23259,
         n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
         n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
         n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283,
         n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
         n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299,
         n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
         n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315,
         n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
         n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
         n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339,
         n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
         n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23356,
         n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364,
         n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372,
         n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380,
         n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388,
         n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396,
         n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404,
         n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412,
         n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420,
         n23421, n23422, n23424, n23425, n23426, n23427, n23428, n23429,
         n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437,
         n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445,
         n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453,
         n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461,
         n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469,
         n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477,
         n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485,
         n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493,
         n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501,
         n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509,
         n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517,
         n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525,
         n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533,
         n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541,
         n23542, n23543, n23544, n23545, n23547, n23548, n23549, n23550,
         n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558,
         n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566,
         n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574,
         n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582,
         n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590,
         n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598,
         n23599, n23600, n23602, n23603, n23604, n23605, n23606, n23607,
         n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615,
         n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623,
         n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631,
         n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639,
         n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647,
         n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655,
         n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663,
         n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671,
         n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679,
         n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687,
         n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695,
         n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703,
         n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711,
         n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719,
         n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727,
         n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735,
         n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743,
         n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751,
         n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759,
         n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767,
         n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775,
         n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783,
         n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791,
         n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799,
         n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807,
         n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815,
         n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823,
         n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831,
         n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839,
         n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847,
         n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855,
         n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863,
         n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871,
         n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879,
         n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887,
         n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895,
         n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903,
         n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911,
         n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919,
         n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927,
         n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935,
         n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943,
         n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951,
         n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959,
         n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967,
         n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975,
         n23976, n23977, n23978, n23979, n23980, n23982, n23983, n23984,
         n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992,
         n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000,
         n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008,
         n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016,
         n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024,
         n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032,
         n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040,
         n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048,
         n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056,
         n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064,
         n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072,
         n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080,
         n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088,
         n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096,
         n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104,
         n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112,
         n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120,
         n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128,
         n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136,
         n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144,
         n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152,
         n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160,
         n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168,
         n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176,
         n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184,
         n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192,
         n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200,
         n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208,
         n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216,
         n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224,
         n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232,
         n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240,
         n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248,
         n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256,
         n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264,
         n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272,
         n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280,
         n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288,
         n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296,
         n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304,
         n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312,
         n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320,
         n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328,
         n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336,
         n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344,
         n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352,
         n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360,
         n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368,
         n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376,
         n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384,
         n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392,
         n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400,
         n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408,
         n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416,
         n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424,
         n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432,
         n24433, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24450,
         n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458,
         n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466,
         n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474,
         n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484,
         n24489, n24490, n24491, n24492, n24493, n24494, n24496, n24497,
         n24498, n24499, n24500, n24501, n24503, n24504, n24505, n24506,
         n24507, n24508, n24513, n24514, n24515, n24516, n24517, n24518,
         n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526,
         n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534,
         n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542,
         n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550,
         n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558,
         n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566,
         n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574,
         n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582,
         n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590,
         n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598,
         n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606,
         n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614,
         n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622,
         n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630,
         n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638,
         n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646,
         n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654,
         n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662,
         n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670,
         n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678,
         n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686,
         n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694,
         n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702,
         n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710,
         n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718,
         n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726,
         n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734,
         n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742,
         n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750,
         n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758,
         n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766,
         n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774,
         n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782,
         n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790,
         n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798,
         n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806,
         n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814,
         n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822,
         n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830,
         n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838,
         n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846,
         n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854,
         n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862,
         n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870,
         n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878,
         n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886,
         n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894,
         n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902,
         n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910,
         n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918,
         n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926,
         n24927, n24928, n24929, n24930, n24931, n24933, n24934, n24935,
         n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943,
         n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951,
         n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959,
         n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967,
         n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975,
         n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983,
         n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991,
         n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999,
         n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007,
         n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015,
         n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023,
         n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031,
         n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040,
         n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048,
         n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056,
         n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064,
         n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072,
         n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080,
         n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088,
         n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096,
         n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104,
         n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112,
         n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120,
         n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128,
         n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136,
         n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144,
         n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152,
         n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160,
         n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168,
         n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176,
         n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184,
         n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192,
         n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200,
         n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208,
         n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216,
         n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224,
         n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232,
         n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240,
         n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248,
         n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256,
         n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264,
         n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272,
         n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280,
         n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288,
         n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296,
         n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304,
         n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312,
         n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320,
         n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328,
         n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336,
         n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344,
         n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352,
         n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360,
         n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368,
         n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376,
         n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384,
         n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392,
         n25393, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25594,
         n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602,
         n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610,
         n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618,
         n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626,
         n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634,
         n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642,
         n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650,
         n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658,
         n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666,
         n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674,
         n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682,
         n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690,
         n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698,
         n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706,
         n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714,
         n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722,
         n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730,
         n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738,
         n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746,
         n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754,
         n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762,
         n25763, n25765, n25766, n25767, n25768, n25769, n25770, n25771,
         n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779,
         n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787,
         n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
         n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803,
         n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
         n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819,
         n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827,
         n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835,
         n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843,
         n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851,
         n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
         n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867,
         n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875,
         n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
         n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891,
         n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899,
         n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907,
         n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915,
         n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923,
         n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
         n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939,
         n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947,
         n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955,
         n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963,
         n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971,
         n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979,
         n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987,
         n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995,
         n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003,
         n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
         n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019,
         n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027,
         n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035,
         n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043,
         n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051,
         n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059,
         n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067,
         n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075,
         n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083,
         n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091,
         n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099,
         n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107,
         n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115,
         n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123,
         n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131,
         n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139,
         n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147,
         n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155,
         n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163,
         n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171,
         n26172, n26173, n26174, n26175, n26176, n26177, n26179, n26180,
         n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188,
         n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196,
         n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204,
         n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212,
         n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220,
         n26221, n26222, n26223, n26224, n26225, n26226, n26227, n26228,
         n26229, n26230, n26231, n26232, n26233, n26234, n26235, n26236,
         n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244,
         n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252,
         n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260,
         n26261, n26262, n26263, n26264, n26265, n26266, n26267, n26268,
         n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276,
         n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284,
         n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292,
         n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300,
         n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308,
         n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316,
         n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324,
         n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332,
         n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340,
         n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348,
         n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356,
         n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364,
         n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372,
         n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380,
         n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388,
         n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396,
         n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404,
         n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412,
         n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420,
         n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428,
         n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436,
         n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444,
         n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452,
         n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460,
         n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468,
         n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476,
         n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484,
         n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26492,
         n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500,
         n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508,
         n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516,
         n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524,
         n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532,
         n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540,
         n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548,
         n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556,
         n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564,
         n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572,
         n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580,
         n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588,
         n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596,
         n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604,
         n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612,
         n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620,
         n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628,
         n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636,
         n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644,
         n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652,
         n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660,
         n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668,
         n26669, n26670, n26671, n26672, n26674, n26675, n26676, n26677,
         n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685,
         n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693,
         n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701,
         n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709,
         n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717,
         n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725,
         n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733,
         n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741,
         n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749,
         n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757,
         n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765,
         n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773,
         n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781,
         n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789,
         n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797,
         n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805,
         n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813,
         n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821,
         n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829,
         n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837,
         n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845,
         n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853,
         n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861,
         n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869,
         n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877,
         n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885,
         n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893,
         n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901,
         n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909,
         n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917,
         n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925,
         n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933,
         n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941,
         n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949,
         n26950, n26951, n26952, n26953, n26954, n26955, n26956, n26957,
         n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965,
         n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973,
         n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981,
         n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989,
         n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997,
         n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005,
         n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013,
         n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021,
         n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029,
         n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037,
         n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045,
         n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053,
         n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061,
         n27062, n27064, n27065, n27066, n27067, n27068, n27069, n27070,
         n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078,
         n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086,
         n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094,
         n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102,
         n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110,
         n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118,
         n27119, n27122, n27123, n27124, n27125, n27126, n27127, n27128,
         n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136,
         n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144,
         n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152,
         n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160,
         n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168,
         n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176,
         n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184,
         n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192,
         n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200,
         n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208,
         n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216,
         n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224,
         n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232,
         n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240,
         n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248,
         n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256,
         n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264,
         n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272,
         n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280,
         n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288,
         n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296,
         n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304,
         n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312,
         n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320,
         n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328,
         n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336,
         n27337, n27338, n27339, n27340, n27341, n27342, n27343, n27344,
         n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352,
         n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360,
         n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368,
         n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376,
         n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384,
         n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392,
         n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400,
         n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408,
         n27409, n27410, n27411, n27412, n27413, n27414, n27415, n27416,
         n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424,
         n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432,
         n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440,
         n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448,
         n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456,
         n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464,
         n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472,
         n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480,
         n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488,
         n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496,
         n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504,
         n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512,
         n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520,
         n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528,
         n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536,
         n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544,
         n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552,
         n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560,
         n27561, n27562, n27563, n27564, n27565, n27566, n27567, n27568,
         n27569, n27570, n27571, n27572, n27573, n27574, n27575, n27576,
         n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584,
         n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592,
         n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600,
         n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608,
         n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616,
         n27617, n27618, n27619, n27620, n27621, n27622, n27623, n27624,
         n27625, n27626, n27627, n27628, n27629, n27630, n27631, n27632,
         n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640,
         n27641, n27642, n27643, n27644, n27645, n27646, n27647, n27648,
         n27649, n27650, n27651, n27652, n27653, n27654, n27655, n27656,
         n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664,
         n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672,
         n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680,
         n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688,
         n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696,
         n27697, n27698, n27699, n27700, n27701, n27702, n27703, n27704,
         n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712,
         n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720,
         n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728,
         n27729, n27730, n27731, n27732, n27733, n27734, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27889, n27890,
         n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898,
         n27899, n27900, n27901, n27902, n27903, n27905, n27906, n27907,
         n27908, n27909, n27910, n27912, n27913, n27914, n27915, n27916,
         n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924,
         n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932,
         n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940,
         n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948,
         n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956,
         n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964,
         n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972,
         n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980,
         n27981, n27982, n27983, n27985, n27986, n27987, n27988, n27989,
         n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997,
         n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005,
         n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013,
         n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021,
         n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029,
         n28030, n28031, n28032, n28033, n28034, n28035, n28036, n28037,
         n28038, n28039, n28040, n28041, n28042, n28043, n28044, n28045,
         n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053,
         n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061,
         n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069,
         n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077,
         n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085,
         n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093,
         n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28101,
         n28102, n28103, n28104, n28105, n28106, n28107, n28108, n28109,
         n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28117,
         n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125,
         n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133,
         n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141,
         n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149,
         n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157,
         n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165,
         n28166, n28167, n28168, n28169, n28170, n28171, n28172, n28173,
         n28174, n28175, n28176, n28177, n28178, n28179, n28180, n28181,
         n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189,
         n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197,
         n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205,
         n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213,
         n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221,
         n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229,
         n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237,
         n28238, n28239, n28240, n28241, n28242, n28243, n28244, n28245,
         n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28253,
         n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261,
         n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269,
         n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277,
         n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285,
         n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293,
         n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301,
         n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309,
         n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317,
         n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325,
         n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333,
         n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341,
         n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349,
         n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357,
         n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365,
         n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373,
         n28374, n28375, n28376, n28377, n28378, n28379, n28380, n28381,
         n28382, n28383, n28384, n28385, n28386, n28387, n28388, n28389,
         n28390, n28391, n28392, n28393, n28394, n28395, n28396, n28397,
         n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405,
         n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413,
         n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421,
         n28422, n28423, n28424, n28425, n28427, n28428, n28429, n28430,
         n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438,
         n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446,
         n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454,
         n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462,
         n28463, n28464, n28466, n28467, n28468, n28469, n28470, n28471,
         n28472, n28473, n28474, n28475, n28476, n28477, n28478, n28479,
         n28480, n28481, n28482, n28483, n28484, n28485, n28486, n28487,
         n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495,
         n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503,
         n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511,
         n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519,
         n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527,
         n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535,
         n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543,
         n28544, n28545, n28546, n28547, n28548, n28549, n28550, n28551,
         n28552, n28553, n28554, n28555, n28556, n28557, n28558, n28559,
         n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567,
         n28568, n28569, n28570, n28571, n28572, n28573, n28574, n28575,
         n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583,
         n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591,
         n28592, n28593, n28594, n28595, n28596, n28597, n28598, n28599,
         n28600, n28601, n28602, n28603, n28604, n28605, n28606, n28607,
         n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615,
         n28616, n28617, n28618, n28619, n28620, n28621, n28622, n28623,
         n28624, n28625, n28626, n28627, n28628, n28629, n28630, n28631,
         n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639,
         n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647,
         n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655,
         n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663,
         n28664, n28665, n28666, n28667, n28668, n28669, n28670, n28671,
         n28672, n28673, n28674, n28675, n28676, n28677, n28678, n28679,
         n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687,
         n28688, n28689, n28690, n28691, n28692, n28693, n28694, n28695,
         n28696, n28697, n28698, n28699, n28700, n28701, n28702, n28703,
         n28704, n28705, n28706, n28707, n28708, n28709, n28710, n28711,
         n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719,
         n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727,
         n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735,
         n28736, n28737, n28738, n28739, n28740, n28741, n28742, n28743,
         n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751,
         n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759,
         n28760, n28761, n28762, n28763, n28764, n28765, n28766, n28767,
         n28768, n28769, n28770, n28771, n28772, n28773, n28774, n28775,
         n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783,
         n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791,
         n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799,
         n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807,
         n28808, n28809, n28810, n28811, n28812, n28813, n28814, n28815,
         n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823,
         n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831,
         n28832, n28833, n28834, n28835, n28836, n28837, n28838, n28839,
         n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847,
         n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855,
         n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863,
         n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871,
         n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879,
         n28880, n28881, n28882, n28883, n28884, n28885, n28886, n28887,
         n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895,
         n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903,
         n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911,
         n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919,
         n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927,
         n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935,
         n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943,
         n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951,
         n28952, n28953, n28954, n28955, n28956, n28957, n28958, n28959,
         n28960, n28961, n28962, n28963, n28964, n28965, n28966, n28967,
         n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975,
         n28976, n28977, n28978, n28979, n28980, n28981, n28982, n28983,
         n28984, n28985, n28986, n28987, n28988, n28989, n28990, n28991,
         n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999,
         n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007,
         n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015,
         n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29023,
         n29024, n29025, n29026, n29027, n29028, n29029, n29030, n29031,
         n29032, n29033, n29034, n29035, n29036, n29037, n29038, n29039,
         n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047,
         n29048, n29049, n29050, n29051, n29052, n29053, n29054, n29055,
         n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063,
         n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071,
         n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079,
         n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087,
         n29088, n29089, n29090, n29091, n29092, n29093, n29094, n29095,
         n29096, n29097, n29098, n29099, n29100, n29101, n29102, n29103,
         n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111,
         n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119,
         n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127,
         n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135,
         n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143,
         n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151,
         n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159,
         n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167,
         n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175,
         n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183,
         n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191,
         n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199,
         n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207,
         n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215,
         n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223,
         n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231,
         n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239,
         n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247,
         n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255,
         n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263,
         n29264, n29265, n29266, n29267, n29268, n29269, n29270, n29271,
         n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279,
         n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287,
         n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295,
         n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303,
         n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311,
         n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319,
         n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327,
         n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335,
         n29336, n29337, n29338, n29339, n29340, n29341, n29342, n29343,
         n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351,
         n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359,
         n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367,
         n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375,
         n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383,
         n29384, n29385, n29386, n29387, n29388, n29389, n29390, n29391,
         n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399,
         n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407,
         n29408, n29409, n29410, n29411, n29412, n29413, n29414, n29415,
         n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423,
         n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431,
         n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439,
         n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447,
         n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29455,
         n29456, n29457, n29458, n29459, n29460, n29461, n29462, n29463,
         n29464, n29465, n29466, n29467, n29468, n29469, n29470, n29471,
         n29472, n29473, n29474, n29475, n29477, n29478, n29479, n29480,
         n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488,
         n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496,
         n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504,
         n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512,
         n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520,
         n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528,
         n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536,
         n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544,
         n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552,
         n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560,
         n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568,
         n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576,
         n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584,
         n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592,
         n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600,
         n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608,
         n29609, n29610, n29630, n29631, n29632, n29633, n29634, n29635,
         n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643,
         n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651,
         n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659,
         n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667,
         n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675,
         n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683,
         n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691,
         n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699,
         n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707,
         n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715,
         n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723,
         n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731,
         n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739,
         n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747,
         n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755,
         n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763,
         n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771,
         n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779,
         n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787,
         n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795,
         n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803,
         n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811,
         n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29820,
         n29821, n29822, n29823, n29824, n29825, n29826, n29827, n29828,
         n29830, n29832, n29833, n29834, n29835, n29836, n29837, n29838,
         n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846,
         n29847, n29848, n29849, n29863, n29864, n29865, n29866, n29868,
         n29869, n29870, n29873, n29874, n29875, n29876, n29877, n29879,
         n29880, n29882, n29883, n29884, n29885, n30010, n30011, n30012,
         n30013, n30014, n30015, n30016, n30017, n30018, n30019, n30020,
         n30021, n30022, n30023, n30024, n30025, n30026, n30027, n30028,
         n30029, n30030, n30031, n30032, n30033, n30034, n30035, n30036,
         n30037, n30038, n30039, n30040, n30041, n30042, n30043, n30044,
         n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052,
         n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060,
         n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068,
         n30069, n30070, n30071, n30072, n30073, n30074, n30075, n30076,
         n30077, n30078, n30079, n30080, n30081, n30082, n30083, n30084,
         n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092,
         n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100,
         n30101, n30102, n30103, n30104, n30105, n30106, n30107, n30108,
         n30109, n30110, n30111, n30112, n30113, n30114, n30115, n30116,
         n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124,
         n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132,
         n30133, n30134, n30135, n30136, n30137, n30138, n30139, n30140,
         n30141, n30142, n30143, n30144, n30145, n30146, n30147, n30148,
         n30149, n30150, n30151, n30152, n30153, n30154, n30155, n30156,
         n30157, n30158, n30159, n30160, n30161, n30162, n30163, n30164,
         n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172,
         n30173, n30174, n30175, n30176, n30177, n30178, n30179, n30180,
         n30181, n30182, n30183, n30184, n30185, n30186, n30187, n30188,
         n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196,
         n30197, n30198, n30199, n30200, n30201, n30202, n30203,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412,
         SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414,
         SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416,
         SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418,
         SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420,
         SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422,
         SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424,
         SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426,
         SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428,
         SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430,
         SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432,
         SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434,
         SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436,
         SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438,
         SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440,
         SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442,
         SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444,
         SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446,
         SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448,
         SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450,
         SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452,
         SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454,
         SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456,
         SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458,
         SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460,
         SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_462,
         SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_464,
         SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_466,
         SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_468,
         SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_470,
         SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_472,
         SYNOPSYS_UNCONNECTED_473, SYNOPSYS_UNCONNECTED_474,
         SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_476,
         SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_478,
         SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_480,
         SYNOPSYS_UNCONNECTED_481, SYNOPSYS_UNCONNECTED_482,
         SYNOPSYS_UNCONNECTED_483, SYNOPSYS_UNCONNECTED_484,
         SYNOPSYS_UNCONNECTED_485, SYNOPSYS_UNCONNECTED_486,
         SYNOPSYS_UNCONNECTED_487, SYNOPSYS_UNCONNECTED_488,
         SYNOPSYS_UNCONNECTED_489, SYNOPSYS_UNCONNECTED_490,
         SYNOPSYS_UNCONNECTED_491, SYNOPSYS_UNCONNECTED_492,
         SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_494,
         SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_496,
         SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_498,
         SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_500,
         SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_502,
         SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_504,
         SYNOPSYS_UNCONNECTED_505, SYNOPSYS_UNCONNECTED_506,
         SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_508,
         SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_510,
         SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_512;
  wire   [31:0] gpio_en_o;
  wire   [1:0] start_n_reg;
  wire   [31:0] j202_soc_core_qspi_wb_wdat;
  wire   [24:2] j202_soc_core_qspi_wb_addr;
  wire   [15:0] j202_soc_core_prdata;
  wire   [7:0] j202_soc_core_paddr;
  wire   [7:0] j202_soc_core_pstrb;
  wire   [0:2] j202_soc_core_pwrite;
  wire   [5:0] j202_soc_core_j22_cpu_exuop_EXU_;
  wire   [4:0] j202_soc_core_j22_cpu_macop_MAC_;
  wire   [31:0] j202_soc_core_j22_cpu_pc;
  wire   [4:0] j202_soc_core_j22_cpu_opst;
  wire   [31:0] j202_soc_core_j22_cpu_rf_tmp;
  wire   [31:0] j202_soc_core_j22_cpu_rf_vbr;
  wire   [31:0] j202_soc_core_j22_cpu_rf_gbr;
  wire   [31:0] j202_soc_core_j22_cpu_rf_pr;
  wire   [510:0] j202_soc_core_j22_cpu_rf_gpr;
  wire   [1:0] j202_soc_core_j22_cpu_ma_M_address;
  wire   [1:0] j202_soc_core_j22_cpu_ma_M_area;
  wire   [3:0] j202_soc_core_j22_cpu_ma_M_MEM;
  wire   [31:0] j202_soc_core_j22_cpu_ml_maclj;
  wire   [23:0] j202_soc_core_j22_cpu_ml_machj;
  wire   [31:0] j202_soc_core_j22_cpu_ml_mach;
  wire   [31:0] j202_soc_core_j22_cpu_ml_macl;
  wire   [32:0] j202_soc_core_j22_cpu_ml_bufb;
  wire   [32:0] j202_soc_core_j22_cpu_ml_bufa;
  wire   [4:0] j202_soc_core_j22_cpu_ml_X_macop_MAC_;
  wire   [4:0] j202_soc_core_j22_cpu_ml_M_macop_MAC_;
  wire   [511:0] j202_soc_core_memory0_ram_dout0;
  wire   [15:0] j202_soc_core_memory0_ram_dout0_sel;
  wire   [111:0] j202_soc_core_ahblite_interconnect_s_hrdata;
  wire  
         [0:6] j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel
;
  wire   [2:0] j202_soc_core_ahb2apb_00_state;
  wire   [15:0] j202_soc_core_cmt_core_00_cnt1;
  wire   [15:0] j202_soc_core_cmt_core_00_cnt0;
  wire   [15:0] j202_soc_core_cmt_core_00_const1;
  wire   [15:0] j202_soc_core_cmt_core_00_const0;
  wire   [15:0] j202_soc_core_cmt_core_00_wdata_cnt0;
  wire   [1:0] j202_soc_core_cmt_core_00_cks1;
  wire   [1:0] j202_soc_core_cmt_core_00_cks0;
  wire   [7:0] j202_soc_core_cmt_core_00_reg_addr;
  wire   [1:0] j202_soc_core_cmt_core_00_cmt_apb_00_state;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata;
  wire   [6:2] j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1;
  wire   [6:2] j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1;
  wire   [9:0] j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1;
  wire   [9:0] j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0;
  wire   [9:0] j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0;
  wire   [9:0] j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0;
  wire   [2:0] j202_soc_core_ahb2apb_01_state;
  wire   [1:0] j202_soc_core_ahb2apb_01_hsize_buf;
  wire   [20:0] j202_soc_core_intc_core_00_in_intreq;
  wire   [127:0] j202_soc_core_intc_core_00_rg_ipr;
  wire   [127:0] j202_soc_core_intc_core_00_rg_itgt;
  wire   [20:0] j202_soc_core_intc_core_00_rg_irqc;
  wire   [31:0] j202_soc_core_intc_core_00_rg_ie;
  wire   [7:0] j202_soc_core_intc_core_00_rg_eimk;
  wire   [15:0] j202_soc_core_intc_core_00_rg_sint;
  wire   [11:0] j202_soc_core_intc_core_00_bs_addr;
  wire  
         [20:0] j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int
;
  wire  
         [6:0] j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch
;
  wire   [2:0] j202_soc_core_ahb2apb_02_state;
  wire   [1:0] j202_soc_core_ahb2apb_02_hsize_buf;
  wire   [7:0] j202_soc_core_gpio_core_00_reg_addr;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_dtr;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_isr;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_ier;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1;
  wire   [7:0] j202_soc_core_uart_din_i;
  wire   [7:0] j202_soc_core_uart_div1;
  wire   [7:0] j202_soc_core_uart_div0;
  wire   [1:0] j202_soc_core_uart_TOP_dpll_state;
  wire   [3:0] j202_soc_core_uart_TOP_rx_bit_cnt;
  wire   [3:0] j202_soc_core_uart_TOP_tx_bit_cnt;
  wire   [8:0] j202_soc_core_uart_TOP_hold_reg;
  wire   [9:2] j202_soc_core_uart_TOP_rxr;
  wire   [31:0] j202_soc_core_uart_TOP_tx_fifo_mem;
  wire   [1:0] j202_soc_core_uart_TOP_tx_fifo_rp;
  wire   [1:0] j202_soc_core_uart_TOP_tx_fifo_wp;
  wire   [31:0] j202_soc_core_uart_TOP_rx_fifo_mem;
  wire   [1:0] j202_soc_core_uart_TOP_rx_fifo_rp;
  wire   [1:0] j202_soc_core_uart_TOP_rx_fifo_wp;
  wire   [1:0] j202_soc_core_uart_BRG_cnt;
  wire   [7:0] j202_soc_core_uart_BRG_br_cnt;
  wire   [7:0] j202_soc_core_uart_BRG_ps;
  wire   [2:0] j202_soc_core_bldc_core_00_hall_value;
  wire   [2:0] j202_soc_core_bldc_core_00_comm;
  wire   [11:0] j202_soc_core_bldc_core_00_pwm_period;
  wire   [11:0] j202_soc_core_bldc_core_00_pwm_duty;
  wire   [23:0] j202_soc_core_bldc_core_00_wdata;
  wire   [7:0] j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1;
  wire   [1:0] j202_soc_core_bldc_core_00_bldc_wb_slave_00_state;
  wire  
         [2:0] j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status
;
  wire   [2:0] j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3;
  wire   [2:0] j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2;
  wire   [2:0] j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1;
  wire   [11:1] j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt;
  wire   [11:0] j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt;
  wire   [31:0] j202_soc_core_wbqspiflash_00_spif_data;
  wire   [7:0] j202_soc_core_wbqspiflash_00_last_status;
  wire   [9:0] j202_soc_core_wbqspiflash_00_reset_counter;
  wire   [4:0] j202_soc_core_wbqspiflash_00_state;
  wire   [7:0] j202_soc_core_wbqspiflash_00_erased_sector;
  wire   [23:2] j202_soc_core_wbqspiflash_00_w_spif_addr;
  wire   [3:0] j202_soc_core_wbqspiflash_00_w_qspi_dat;
  wire   [1:0] j202_soc_core_wbqspiflash_00_w_qspi_mod;
  wire   [31:0] j202_soc_core_wbqspiflash_00_spi_out;
  wire   [1:0] j202_soc_core_wbqspiflash_00_spi_len;
  wire   [31:0] j202_soc_core_wbqspiflash_00_spi_in;
  wire   [5:0] j202_soc_core_wbqspiflash_00_lldriver_spi_len;
  wire   [31:0] j202_soc_core_wbqspiflash_00_lldriver_r_word;
  wire   [30:0] j202_soc_core_wbqspiflash_00_lldriver_r_input;
  wire   [2:0] j202_soc_core_wbqspiflash_00_lldriver_state;
  wire   [17:2] j202_soc_core_bootrom_00_address_w;

  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_15__ram ( 
        .din0({n29805, n29803, n12242, n29799, n29797, n29795, n29793, n29791, 
        n29789, n29787, n29785, n29783, n29780, n29778, n29776, n29774, n12207, 
        n29770, n29768, n12319, n29766, n29764, n29817, n24516, n29815, n29813, 
        n29811, n29809, n29807, n29801, n29781, n29762}), .dout0(
        j202_soc_core_memory0_ram_dout0[511:480]), .addr0({n11090, n11076, 
        n11082, n11045, n11041, n11053, n11079, n11057, n11049}), .wmask0({
        n11031, n11065, n12313, n11121}), .dout1({SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_1}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10596), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_14__ram ( 
        .din0({n29806, n29804, n12243, n29800, n29798, n29796, n29794, n29792, 
        n29790, n29788, n29786, n29784, n12043, n29779, n29777, n29775, n29773, 
        n29770, n29768, n12231, n29767, n29765, n29818, n24516, n29816, n29814, 
        n29812, n29810, n29808, n29802, n29782, n29763}), .dout0(
        j202_soc_core_memory0_ram_dout0[479:448]), .addr0({n11090, n30100, 
        n12070, n12076, n12072, n12074, n11021, n12078, n12080}), .wmask0({
        n11069, n11071, n11120, n11121}), .dout1({SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_33}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10595), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_13__ram ( 
        .din0({n29805, n29803, n12242, n29799, n29797, n29795, n29793, n29791, 
        n29789, n29787, n29785, n29783, n12043, n29778, n29776, n29774, n29772, 
        n29770, n29768, n12319, n29766, n29764, n29817, n24516, n29815, n29813, 
        n29811, n29809, n29807, n29801, n29781, n29762}), .dout0(
        j202_soc_core_memory0_ram_dout0[447:416]), .addr0({n11089, n11026, 
        n12388, n12077, n12073, n12075, n11080, n12079, n12081}), .wmask0({
        n11074, n11028, n11127, n11162}), .dout1({SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_96, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_90, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_65}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10594), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_12__ram ( 
        .din0({n29806, n29804, n12243, n29800, n29798, n29796, n29794, n29792, 
        n29790, n29788, n29786, n29784, n12043, n29779, n29777, n29775, n29773, 
        n29770, n29768, n12231, n29767, n29765, n29818, n24516, n29816, n29814, 
        n29812, n29810, n29808, n29802, n29782, n29763}), .dout0(
        j202_soc_core_memory0_ram_dout0[415:384]), .addr0({n11016, n30093, 
        n12311, n12308, n12300, n12306, n11022, n12304, n12302}), .wmask0({
        n11068, n11070, n11120, n10988}), .dout1({SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_118, 
        SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_116, 
        SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_114, 
        SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_112, 
        SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_110, 
        SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_128, 
        SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_126, 
        SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_124, 
        SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_122, 
        SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_108, 
        SYNOPSYS_UNCONNECTED_97}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10593), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_11__ram ( 
        .din0({n29805, n29803, n12243, n29799, n29797, n29795, n29793, n29791, 
        n29789, n29787, n29785, n29783, n29780, n29778, n29776, n29774, n12207, 
        n29770, n29768, n12319, n29766, n29764, n29817, n24516, n29815, n29813, 
        n29811, n29809, n29807, n29801, n29781, n29762}), .dout0(
        j202_soc_core_memory0_ram_dout0[383:352]), .addr0({n11088, n30096, 
        n12311, n12308, n12300, n12306, n11080, n12304, n12302}), .wmask0({
        n11067, n11071, n12312, n11162}), .dout1({SYNOPSYS_UNCONNECTED_153, 
        SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_140, 
        SYNOPSYS_UNCONNECTED_129}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10592), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_10__ram ( 
        .din0({n29806, n29804, n12242, n29800, n29798, n29796, n29794, n29792, 
        n29790, n29788, n29786, n29784, n29780, n29779, n29777, n29775, n29773, 
        n29770, n29768, n12231, n29767, n29765, n29818, n24516, n29816, n29814, 
        n29812, n29810, n29808, n29802, n29782, n29763}), .dout0(
        j202_soc_core_memory0_ram_dout0[351:320]), .addr0({n11016, n30096, 
        n12289, n11044, n11040, n11052, n11086, n11056, n11048}), .wmask0({
        n11068, n11070, n12312, n10989}), .dout1({SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_178, 
        SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_176, 
        SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_174, 
        SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_171, 
        SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_169, 
        SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_167, 
        SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_165, 
        SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_163, 
        SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_192, 
        SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_190, 
        SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_188, 
        SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_186, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_172, 
        SYNOPSYS_UNCONNECTED_161}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10591), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_9__ram ( 
        .din0({n29805, n29803, n12243, n29799, n29797, n29795, n29793, n29791, 
        n29789, n29787, n29785, n29783, n29780, n29778, n29776, n29774, n29772, 
        n29770, n29768, n12231, n29766, n29764, n29817, n24516, n29815, n29813, 
        n29811, n29809, n29807, n29801, n29781, n29762}), .dout0(
        j202_soc_core_memory0_ram_dout0[319:288]), .addr0({n11017, n11033, 
        n12388, n11047, n11043, n11055, n11086, n11059, n11051}), .wmask0({
        n11073, n11029, n11155, n10989}), .dout1({SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_214, 
        SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_212, 
        SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_210, 
        SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_208, 
        SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_206, 
        SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_224, 
        SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_222, 
        SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_220, 
        SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_218, 
        SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_204, 
        SYNOPSYS_UNCONNECTED_193}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10590), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_8__ram ( 
        .din0({n29806, n29804, n12242, n29800, n29798, n29796, n29794, n29792, 
        n29790, n29788, n29786, n29784, n12043, n29779, n29777, n29775, n29773, 
        n29770, n29768, n12319, n29767, n29765, n29818, n24516, n29816, n29814, 
        n29812, n29810, n29808, n29802, n29782, n29763}), .dout0(
        j202_soc_core_memory0_ram_dout0[287:256]), .addr0({n11017, n11075, 
        n12290, n12077, n12073, n12075, n11063, n12079, n12081}), .wmask0({
        n11023, n11066, n12314, n29820}), .dout1({SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_246, 
        SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_244, 
        SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_242, 
        SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_240, 
        SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_238, 
        SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_256, 
        SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_254, 
        SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_252, 
        SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_250, 
        SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_236, 
        SYNOPSYS_UNCONNECTED_225}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10589), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_7__ram ( 
        .din0({n29805, n29803, n12242, n29799, n29797, n29795, n29793, n29791, 
        n29789, n29787, n29785, n29783, n29780, n29778, n29776, n29774, n12207, 
        n29771, n29769, n12231, n29766, n29764, n29817, n24516, n29815, n29813, 
        n29811, n29809, n29807, n29801, n29781, n29762}), .dout0(
        j202_soc_core_memory0_ram_dout0[255:224]), .addr0({n11034, n30091, 
        n12071, n12384, n12376, n12382, n11063, n12380, n12378}), .wmask0({
        n10987, n11039, n10984, n12315}), .dout1({SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_278, 
        SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_276, 
        SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_274, 
        SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_272, 
        SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_270, 
        SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_288, 
        SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_286, 
        SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_284, 
        SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_282, 
        SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_268, 
        SYNOPSYS_UNCONNECTED_257}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10588), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_6__ram ( 
        .din0({n29806, n29804, n12242, n29800, n29798, n29796, n29794, n29792, 
        n29790, n29788, n29786, n29784, n12043, n29779, n29777, n29775, n29773, 
        n29771, n29769, n12319, n29767, n29765, n29818, n24516, n29816, n29814, 
        n29812, n29810, n29808, n29802, n29782, n29763}), .dout0(
        j202_soc_core_memory0_ram_dout0[223:192]), .addr0({n30094, n11077, 
        n12387, n12385, n12377, n12383, n11021, n12381, n12379}), .wmask0({
        n11072, n11064, n12313, n10986}), .dout1({SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_299, 
        SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_297, 
        SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_295, 
        SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_293, 
        SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_291, 
        SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_320, 
        SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_318, 
        SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_316, 
        SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_314, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_289}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10587), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_5__ram ( 
        .din0({n29805, n29803, n12242, n29799, n29797, n29795, n29793, n29791, 
        n29789, n29787, n29785, n29783, n29780, n29778, n29776, n29774, n29772, 
        n29771, n29769, n12319, n29766, n29764, n29817, n24516, n29815, n29813, 
        n29811, n29809, n29807, n29801, n29781, n29762}), .dout0(
        j202_soc_core_memory0_ram_dout0[191:160]), .addr0({n11018, n11032, 
        n12071, n12384, n12376, n12382, n11022, n12380, n12378}), .wmask0({
        n11030, n11025, n11127, n10986}), .dout1({SYNOPSYS_UNCONNECTED_345, 
        SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_338, 
        SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_336, 
        SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_334, 
        SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_331, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_352, 
        SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_350, 
        SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_348, 
        SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_346, 
        SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_332, 
        SYNOPSYS_UNCONNECTED_321}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10586), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_4__ram ( 
        .din0({n29806, n29804, n12243, n29800, n29798, n29796, n29794, n29792, 
        n29790, n29788, n29786, n29784, n12043, n29779, n29777, n29775, n29773, 
        n29771, n29769, n12231, n29767, n29765, n29818, n24516, n29816, n29814, 
        n29812, n29810, n29808, n29802, n29782, n29763}), .dout0(
        j202_soc_core_memory0_ram_dout0[159:128]), .addr0({n11089, n11136, 
        n12310, n12309, n12301, n12307, n11020, n12305, n12303}), .wmask0({
        n11036, n11029, n10984, n10988}), .dout1({SYNOPSYS_UNCONNECTED_377, 
        SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_374, 
        SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_372, 
        SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_370, 
        SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_368, 
        SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_366, 
        SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_363, 
        SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_361, 
        SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_359, 
        SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_357, 
        SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_355, 
        SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_384, 
        SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_382, 
        SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_380, 
        SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_378, 
        SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_364, 
        SYNOPSYS_UNCONNECTED_353}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10585), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_3__ram ( 
        .din0({n29805, n29803, n12243, n29799, n29797, n29795, n29793, n29791, 
        n29789, n29787, n29785, n29783, n29780, n29778, n29776, n29774, n12207, 
        n29771, n29769, n12231, n29766, n29764, n29817, n24516, n29815, n29813, 
        n29811, n29809, n29807, n29801, n29781, n29762}), .dout0(
        j202_soc_core_memory0_ram_dout0[127:96]), .addr0({n11019, n11078, 
        n12387, n12385, n12377, n12383, n11020, n12381, n12379}), .wmask0({
        n11024, n11065, n12314, n29820}), .dout1({SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_406, 
        SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_404, 
        SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_402, 
        SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_400, 
        SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_398, 
        SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_389, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_416, 
        SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_414, 
        SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_412, 
        SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_410, 
        SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_396, 
        SYNOPSYS_UNCONNECTED_385}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10584), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_2__ram ( 
        .din0({n29806, n29804, n12243, n29800, n29798, n29796, n29794, n29792, 
        n29790, n29788, n29786, n29784, n12043, n29779, n29777, n29775, n29773, 
        n29771, n29769, n12319, n29767, n29765, n29818, n24516, n29816, n29814, 
        n29812, n29810, n29808, n29802, n29782, n29763}), .dout0(
        j202_soc_core_memory0_ram_dout0[95:64]), .addr0({n11018, n30100, 
        n12070, n12076, n12072, n12074, n11163, n12078, n12080}), .wmask0({
        n11038, n30097, n10983, n10985}), .dout1({SYNOPSYS_UNCONNECTED_441, 
        SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_438, 
        SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_436, 
        SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_434, 
        SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_432, 
        SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_430, 
        SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_427, 
        SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_425, 
        SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_423, 
        SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_421, 
        SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_419, 
        SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_448, 
        SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_446, 
        SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_444, 
        SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_442, 
        SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_428, 
        SYNOPSYS_UNCONNECTED_417}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10583), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_1__ram ( 
        .din0({n29805, n29803, n12243, n29799, n29797, n29795, n29793, n29791, 
        n29789, n29787, n29785, n29783, n29780, n29778, n29776, n29774, n29772, 
        n29771, n29769, n12319, n29766, n29764, n29817, n24516, n29815, n29813, 
        n29811, n29809, n29807, n29801, n29781, n29762}), .dout0(
        j202_soc_core_memory0_ram_dout0[63:32]), .addr0({n11088, n11027, 
        n11082, n11046, n11042, n11054, n11079, n11058, n11050}), .wmask0({
        n11073, n30098, n11155, n12315}), .dout1({SYNOPSYS_UNCONNECTED_473, 
        SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_470, 
        SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_468, 
        SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_466, 
        SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_464, 
        SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_462, 
        SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_459, 
        SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_457, 
        SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_455, 
        SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_453, 
        SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_451, 
        SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_480, 
        SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_478, 
        SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_476, 
        SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_474, 
        SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_460, 
        SYNOPSYS_UNCONNECTED_449}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10582), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_0__ram ( 
        .din0({n29806, n29804, n12242, n29800, n29798, n29796, n29794, n29792, 
        n29790, n29788, n29786, n29784, n12043, n29779, n29777, n29775, n29773, 
        n29771, n29769, n12231, n29767, n29765, n29818, n24516, n29816, n29814, 
        n29812, n29810, n29808, n29802, n29782, n29763}), .dout0(
        j202_soc_core_memory0_ram_dout0[31:0]), .addr0({n11019, n11136, n12310, 
        n12309, n12301, n12307, n11163, n12305, n12303}), .wmask0({n10987, 
        n11064, n10983, n10985}), .dout1({SYNOPSYS_UNCONNECTED_505, 
        SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_502, 
        SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_500, 
        SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_498, 
        SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_496, 
        SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_494, 
        SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_491, 
        SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_489, 
        SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_487, 
        SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_485, 
        SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_483, 
        SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_512, 
        SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_510, 
        SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_508, 
        SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_506, 
        SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_492, 
        SYNOPSYS_UNCONNECTED_481}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10581), .web0(n23989), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_fd_sc_hd__dfxtp_1 start_n_reg_reg_0_ ( .D(n3), .CLK(wb_clk_i), .Q(
        start_n_reg[0]) );
  sky130_fd_sc_hd__dfxtp_1 start_n_reg_reg_1_ ( .D(n4), .CLK(wb_clk_i), .Q(
        start_n_reg[1]) );
  sky130_fd_sc_hd__edfxtp_1 ready_reg ( .D(n29610), .DE(n470), .CLK(wb_clk_i), 
        .Q(wbs_ack_o) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_31_ ( .D(n460), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[31]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_30_ ( .D(n450), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[30]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_29_ ( .D(n440), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[29]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_28_ ( .D(n430), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[28]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_27_ ( .D(n420), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[27]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_26_ ( .D(n410), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[26]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_25_ ( .D(n400), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[25]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_24_ ( .D(n390), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[24]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_23_ ( .D(n370), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[23]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_22_ ( .D(n360), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[22]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_21_ ( .D(n350), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[21]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_20_ ( .D(n340), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[20]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_19_ ( .D(n330), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[19]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_18_ ( .D(n320), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[18]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_17_ ( .D(n310), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[17]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_16_ ( .D(n300), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[16]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_15_ ( .D(n280), .DE(n20), .CLK(
        wb_clk_i), .Q(wbs_dat_o[15]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_14_ ( .D(n270), .DE(n20), .CLK(
        wb_clk_i), .Q(wbs_dat_o[14]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_13_ ( .D(n260), .DE(n20), .CLK(
        wb_clk_i), .Q(wbs_dat_o[13]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_12_ ( .D(n250), .DE(n20), .CLK(
        wb_clk_i), .Q(wbs_dat_o[12]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_11_ ( .D(n240), .DE(n20), .CLK(
        wb_clk_i), .Q(wbs_dat_o[11]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_10_ ( .D(n230), .DE(n20), .CLK(
        wb_clk_i), .Q(wbs_dat_o[10]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_9_ ( .D(n220), .DE(n20), .CLK(wb_clk_i), .Q(wbs_dat_o[9]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_8_ ( .D(n21), .DE(n20), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[8]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_7_ ( .D(n19), .DE(n12), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[7]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_6_ ( .D(n18), .DE(n12), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[6]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_5_ ( .D(n17), .DE(n12), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[5]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_4_ ( .D(n16), .DE(n12), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[4]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_3_ ( .D(n15), .DE(n12), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[3]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_2_ ( .D(n14), .DE(n12), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[2]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_1_ ( .D(n13), .DE(n12), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[1]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_0_ ( .D(n11), .DE(n10), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_rst0_reg ( .D(n10525), .CLK(wb_clk_i), 
        .Q(j202_soc_core_rst0) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_rst1_reg ( .D(j202_soc_core_rst0), 
        .CLK(wb_clk_i), .Q(j202_soc_core_rst1) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_0_ ( 
        .D(n29682), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_1_ ( 
        .D(n29681), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_2_ ( 
        .D(n29680), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_3_ ( 
        .D(n29679), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_4_ ( 
        .D(n29678), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_5_ ( 
        .D(n29677), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_6_ ( 
        .D(n29676), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_7_ ( 
        .D(n29675), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_8_ ( 
        .D(n29674), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_9_ ( 
        .D(n29673), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_10_ ( 
        .D(n29672), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_11_ ( 
        .D(n29632), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_12_ ( 
        .D(n29671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_13_ ( 
        .D(n29670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_14_ ( 
        .D(n29669), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_15_ ( 
        .D(n29668), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_16_ ( 
        .D(n29667), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_17_ ( 
        .D(n29666), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_18_ ( 
        .D(n29665), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_19_ ( 
        .D(n29664), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_20_ ( 
        .D(n29663), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_21_ ( 
        .D(n29662), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_22_ ( 
        .D(n29661), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_23_ ( 
        .D(n29660), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_24_ ( 
        .D(n29659), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_25_ ( 
        .D(n29658), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_26_ ( 
        .D(n29657), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_27_ ( 
        .D(n29656), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_28_ ( 
        .D(n29655), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_29_ ( 
        .D(n29654), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_30_ ( 
        .D(n29653), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_31_ ( 
        .D(n29652), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_0_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N3), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_1_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N4), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_2_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N5), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_3_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N6), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_4_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N7), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_5_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N8), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_6_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N9), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_7_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N10), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_8_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N11), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_9_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N12), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_10_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N13), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[10])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_11_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N14), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[11])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_12_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N15), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[12])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_13_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N16), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_14_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N17), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_15_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N18), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_16_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N19), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_17_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N20), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[17])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_18_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N21), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[18])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_19_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N22), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[19])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_20_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N23), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[20])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_21_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[21])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_22_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N25), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[22])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_23_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N26), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[23])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_24_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N27), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[24])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_25_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N28), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[25])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_26_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N29), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[26])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_27_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N30), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[27])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_28_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N31), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[28])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_29_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N32), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[29])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_30_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N33), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[30])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_31_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N34), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[31])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_0_ ( 
        .D(n29598), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_1_ ( 
        .D(n29739), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_2_ ( 
        .D(n29736), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_3_ ( 
        .D(n29727), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_4_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N7), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_5_ ( 
        .D(n29728), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_6_ ( 
        .D(n29734), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_7_ ( 
        .D(n29737), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_8_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N11), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_9_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N12), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_10_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N13), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[10])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_11_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N14), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[11])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_12_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N15), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[12])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_13_ ( 
        .D(n29738), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_14_ ( 
        .D(n29729), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_15_ ( 
        .D(n29735), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_16_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N19), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[16])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_17_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N20), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[17])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_18_ ( 
        .D(n29604), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_19_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N22), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[19])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_20_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N23), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[20])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_21_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[21])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_22_ ( 
        .D(n29579), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_23_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N26), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[23])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_24_ ( 
        .D(n29605), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_25_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N28), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[25])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_26_ ( 
        .D(n29578), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_27_ ( 
        .D(n29577), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_28_ ( 
        .D(n29606), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_29_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N32), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[29])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_30_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N33), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[30])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_31_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N34), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[31])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rxd_s_reg ( .D(io_in[5]), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rxd_s) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rxd_r_reg ( .D(
        j202_soc_core_uart_TOP_rxd_s), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rxd_r) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1_reg_0_ ( 
        .D(io_in[22]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2_reg_0_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[0]), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3_reg_0_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[0]), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1_reg_1_ ( 
        .D(io_in[23]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2_reg_1_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[1]), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3_reg_1_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[1]), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1_reg_2_ ( 
        .D(io_in[24]), .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2_reg_2_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[2]), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3_reg_2_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[2]), .CLK(
        wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1_reg ( 
        .D(n29599), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_2_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1), .CLK(
        wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_2) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_o_reg_2_ ( 
        .D(n138), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_hall_value[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status_reg_2_ ( 
        .D(j202_soc_core_bldc_core_00_hall_value[2]), .CLK(wb_clk_i), 
        .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_o_reg_0_ ( 
        .D(n137), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_hall_value[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status_reg_0_ ( 
        .D(j202_soc_core_bldc_core_00_hall_value[0]), .CLK(wb_clk_i), 
        .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_o_reg_1_ ( 
        .D(n136), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_hall_value[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status_reg_1_ ( 
        .D(j202_soc_core_bldc_core_00_hall_value[1]), .CLK(wb_clk_i), 
        .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_0_ ( 
        .D(n29493), .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_1_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[1]), .CLK(
        wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_2_ ( 
        .D(n29694), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_3_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[3]), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_4_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[4]), .CLK(
        wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_5_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[5]), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_6_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[6]), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_7_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[7]), .CLK(
        wb_clk_i), .RESET_B(n12069), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_8_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[8]), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_9_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[9]), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_10_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[10]), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_11_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[11]), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_bootrom_00_sel_w_reg ( .D(n30030), 
        .CLK(wb_clk_i), .Q(j202_soc_core_bootrom_00_sel_w) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_other__2_ ( 
        .D(n10526), .DE(n10622), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_other__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_ifetchl_reg ( .D(
        j202_soc_core_j22_cpu_ifetch), .DE(n29746), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ifetchl) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_area_reg_0_ ( .D(n10579), .DE(n10600), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ma_M_area[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aqu_st_reg_0_ ( .D(
        j202_soc_core_ahb2aqu_00_N93), .DE(j202_soc_core_ahb2aqu_00_N95), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2aqu_00_aqu_st_0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_STB_ ( .D(
        j202_soc_core_ahb2aqu_00_N128), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_STB_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_area_reg_1_ ( .D(n10578), .DE(n10600), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ma_M_area[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_WE_ ( .D(n29496), .DE(j202_soc_core_ahb2aqu_00_N95), .CLK(wb_clk_i), .Q(j202_soc_core_aquc_WE_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_state_reg_0_ ( 
        .D(n29435), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_1_ ( .D(
        n10605), .DE(n10601), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_opst[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rb__1_ ( 
        .D(n10620), .DE(n10609), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rb__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__2_ ( .D(
        n12145), .DE(j202_soc_core_ahb2aqu_00_N127), .CLK(wb_clk_i), .Q(
        j202_soc_core_aquc_ADR__2_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_2_ ( 
        .D(j202_soc_core_aquc_ADR__2_), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_2_ ( .D(
        n29557), .DE(n10998), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_other__0_ ( 
        .D(n10528), .DE(n10622), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_other__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__15_ ( 
        .D(n29502), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_15_ ( 
        .D(j202_soc_core_qspi_wb_wdat[15]), .CLK(wb_clk_i), .RESET_B(n29827), 
        .Q(j202_soc_core_bldc_core_00_wdata[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_15_ ( 
        .D(j202_soc_core_qspi_wb_wdat[15]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_15_ ( 
        .D(n29446), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_15_ ( .D(
        j202_soc_core_ahb2apb_02_N143), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[47]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__7_ ( 
        .D(n10534), .DE(n12364), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__7_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__7_ ( .D(
        n12148), .DE(j202_soc_core_ahb2aqu_00_N127), .CLK(wb_clk_i), .Q(
        j202_soc_core_aquc_ADR__7_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_7_ ( 
        .D(j202_soc_core_aquc_ADR__7_), .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_7_ ( .D(
        n29556), .DE(n10998), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__10_ ( 
        .D(n29499), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_10_ ( 
        .D(j202_soc_core_qspi_wb_wdat[10]), .CLK(wb_clk_i), .RESET_B(n29745), 
        .Q(j202_soc_core_bldc_core_00_wdata[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_10_ ( 
        .D(j202_soc_core_qspi_wb_wdat[10]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_10_ ( 
        .D(n29448), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_10_ ( .D(
        j202_soc_core_ahb2apb_02_N138), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[42]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__0_ ( 
        .D(n10624), .DE(n10601), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__4_ ( .D(
        j202_soc_core_j22_cpu_ml_N195), .DE(n29746), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_4_ ( 
        .D(n29633), .DE(n10600), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_other__1_ ( 
        .D(n10527), .DE(n10622), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_other__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_20_ ( .D(
        j202_soc_core_j22_cpu_rf_N318), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_We__0_ ( 
        .D(n10616), .DE(n10645), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_We__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Wm__3_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N900), .DE(n10645), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_Wm__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_2_ ( .D(
        n10604), .DE(n10601), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_opst[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__4_ ( 
        .D(n29540), .DE(n10601), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__1_ ( 
        .D(n10540), .DE(n12364), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_address_reg_1_ ( .D(
        n29581), .DE(n29882), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_address[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__1_ ( .D(
        n13088), .DE(j202_soc_core_ahb2aqu_00_N127), .CLK(wb_clk_i), .Q(
        j202_soc_core_aquc_ADR__1_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_1_ ( 
        .D(j202_soc_core_aquc_ADR__1_), .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_SEL__3_ ( .D(
        j202_soc_core_ahb2aqu_00_N164), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_SEL__3_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_1_ ( .D(n135), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_uart_div0[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__3_ ( .D(
        n12144), .DE(j202_soc_core_ahb2aqu_00_N127), .CLK(wb_clk_i), .Q(
        j202_soc_core_aquc_ADR__3_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_3_ ( 
        .D(j202_soc_core_aquc_ADR__3_), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_3_ ( .D(
        n29553), .DE(n10998), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__0_ ( 
        .D(n10632), .DE(n10609), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_istall_reg ( .D(n10597), 
        .DE(n10646), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_istall) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_v_ ( .D(n29484), 
        .DE(n29746), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_id_op2_v_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__0_ ( .D(
        n12317), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__1_ ( .D(
        n12417), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__2_ ( .D(
        n11395), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__3_ ( .D(
        n29491), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__7_ ( .D(
        n12208), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__7_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__8_ ( .D(
        n29593), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__8_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__9_ ( .D(
        n12669), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__9_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__10_ ( .D(
        n29587), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__10_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__11_ ( .D(
        n11182), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__11_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__12_ ( .D(
        n29481), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__12_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__15_ ( .D(
        n11545), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__15_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_30_ ( .D(
        j202_soc_core_j22_cpu_rf_N328), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_5_ ( 
        .D(n29438), .DE(n10600), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_2_ ( .D(
        n29557), .DE(n13109), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_3_ ( .D(
        n29553), .DE(n13109), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_7_ ( .D(
        n29556), .DE(n30067), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_18_ ( 
        .D(n29436), .DE(n13109), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_20_ ( 
        .D(n12353), .DE(n13109), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_hwrite_temp_reg ( .D(
        n29496), .DE(n13109), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_we) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_req_reg ( .D(
        n10543), .DE(n29651), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_req) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_ack_reg ( .D(
        j202_soc_core_wbqspiflash_00_N730), .DE(
        j202_soc_core_wbqspiflash_00_N729), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_ack) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_stb_o_reg ( .D(n30068), 
        .DE(n10577), .CLK(wb_clk_i), .Q(j202_soc_core_ahb2wbqspi_00_stb_o) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_cyc_o_reg ( .D(n30067), 
        .DE(n10577), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_cyc) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_1_ ( .D(
        j202_soc_core_wbqspiflash_00_N725), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_hold_reg ( .D(
        j202_soc_core_wbqspiflash_00_N590), .DE(
        j202_soc_core_wbqspiflash_00_N745), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_hold) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_state_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N308), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N307), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_state[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_busy_reg ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N321), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_busy) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_write_in_progress_reg ( 
        .D(j202_soc_core_wbqspiflash_00_N709), .DE(
        j202_soc_core_wbqspiflash_00_N708), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_write_in_progress) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_31_ ( .D(
        n10544), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_2_ ( .D(
        j202_soc_core_wbqspiflash_00_N726), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_0_ ( .D(
        j202_soc_core_wbqspiflash_00_N724), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_len_reg_1_ ( .D(
        j202_soc_core_wbqspiflash_00_N737), .DE(
        j202_soc_core_wbqspiflash_00_N735), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_len[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N429), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_state_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N309), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N307), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_state_reg_2_ ( 
        .D(n29563), .DE(j202_soc_core_wbqspiflash_00_lldriver_N307), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_state[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_valid_reg ( 
        .D(n29603), .CLK(wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_valid)
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_sck_reg ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N312), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_sck) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_cs_n_reg ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N314), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N313), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_cs_n) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_write_protect_reg ( 
        .D(j202_soc_core_wbqspiflash_00_N722), .DE(
        j202_soc_core_wbqspiflash_00_N721), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_write_protect) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_28_ ( 
        .D(j202_soc_core_wbqspiflash_00_N695), .DE(n29754), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_0_ ( 
        .D(n10966), .DE(n10600), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_00_state_reg_0_ ( .D(n29645), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2apb_00_state[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_00_state_reg_2_ ( .D(n29741), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2apb_00_state[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_state_reg_1_ ( 
        .D(n29485), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_state_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_apb_00_nxt_state_0_), .CLK(wb_clk_i), 
        .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_apb_00_state[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_hwrite_buf_reg ( .D(
        n29644), .DE(n30055), .CLK(wb_clk_i), .Q(j202_soc_core_pwrite[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_1_reg ( 
        .D(j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen), .CLK(wb_clk_i), 
        .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_1)
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_2_reg ( 
        .D(j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_1), .CLK(wb_clk_i), 
        .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_2)
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_7_ ( .D(
        n29643), .DE(n30055), .CLK(wb_clk_i), .Q(j202_soc_core_paddr[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_7_ ( 
        .D(j202_soc_core_paddr[7]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_reg_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_3_ ( .D(
        n29642), .DE(n30056), .CLK(wb_clk_i), .Q(j202_soc_core_paddr[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_3_ ( 
        .D(j202_soc_core_paddr[3]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_reg_addr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_2_ ( .D(
        n29641), .DE(n12277), .CLK(wb_clk_i), .Q(j202_soc_core_paddr[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_2_ ( 
        .D(j202_soc_core_paddr[2]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_reg_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_1_ ( .D(
        n29640), .DE(n30056), .CLK(wb_clk_i), .Q(j202_soc_core_paddr[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_1_ ( 
        .D(j202_soc_core_paddr[1]), .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_cmt_core_00_reg_addr[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_6_ ( 
        .D(n134), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_16_ ( 
        .D(n29874), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[16])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_16_ ( 
        .D(n29722), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_in_intreq[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__0_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__3_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_4_ ( 
        .D(n29583), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__4_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_6_ ( 
        .D(n29480), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__6_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__2_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__1_ ( .D(
        n11102), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__2_ ( .D(
        n20255), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__3_ ( .D(
        n29848), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__7_ ( .D(
        n29439), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__7_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__8_ ( .D(
        n29486), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__8_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__10_ ( .D(
        n29845), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__10_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__11_ ( .D(
        n29846), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__11_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__12_ ( .D(
        n29487), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__12_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__15_ ( .D(
        n29495), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__15_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__0_ ( .D(
        n29444), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_v_ ( .D(n29747), 
        .DE(n10574), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_id_opn_v_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__6_ ( .D(
        n29559), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__6_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rs__1_ ( 
        .D(n10643), .DE(n10609), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rs__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__13_ ( .D(
        n29564), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__13_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__13_ ( .D(
        n29488), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__13_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Ra__0_ ( 
        .D(n10644), .DE(n10609), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Ra__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_21_ ( 
        .D(n12334), .DE(n13109), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_19_ ( 
        .D(j202_soc_core_qspi_wb_addr[21]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_dirty_sector_reg ( 
        .D(j202_soc_core_wbqspiflash_00_N720), .DE(
        j202_soc_core_wbqspiflash_00_N719), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_dirty_sector) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_30_ ( 
        .D(j202_soc_core_wbqspiflash_00_N697), .DE(n29876), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__14_ ( .D(
        n29595), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__14_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_21_ ( .D(
        j202_soc_core_j22_cpu_rf_N319), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__14_ ( .D(
        n29847), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__14_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_14_ ( 
        .D(n29547), .DE(n30068), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_0_ ( .D(
        n29532), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__11_ ( 
        .D(n29500), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_11_ ( 
        .D(j202_soc_core_qspi_wb_wdat[11]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_bldc_core_00_wdata[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_11_ ( 
        .D(j202_soc_core_qspi_wb_wdat[11]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_11_ ( 
        .D(n29447), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_11_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N51), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_18_ ( 
        .D(n29580), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[18])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_18_ ( .D(
        j202_soc_core_ahb2apb_01_N146), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[82]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__t_ ( .D(
        j202_soc_core_j22_cpu_rf_N2626), .DE(j202_soc_core_j22_cpu_rf_N2625), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__t_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_18_ ( .D(
        j202_soc_core_j22_cpu_rf_N316), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_16_ ( 
        .D(n29482), .DE(n30068), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_3_ ( 
        .D(n29551), .DE(n10600), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_CE__1_ ( .D(
        j202_soc_core_ahb2aqu_00_N98), .DE(j202_soc_core_ahb2aqu_00_N95), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_CE__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_17_ ( 
        .D(n29441), .DE(n30067), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_17_ ( .D(
        n29441), .DE(n30030), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__6_ ( .D(
        n11796), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__6_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_6_ ( .D(
        n29639), .DE(n30055), .CLK(wb_clk_i), .Q(j202_soc_core_paddr[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_6_ ( 
        .D(j202_soc_core_paddr[6]), .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_cmt_core_00_reg_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__6_ ( .D(
        n12149), .DE(j202_soc_core_ahb2aqu_00_N127), .CLK(wb_clk_i), .Q(
        j202_soc_core_aquc_ADR__6_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_6_ ( 
        .D(j202_soc_core_aquc_ADR__6_), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_6_ ( .D(
        n29555), .DE(n30068), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_6_ ( .D(
        n29555), .DE(n30030), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__9_ ( .D(
        n11185), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__9_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_9_ ( .D(
        n29546), .DE(n30067), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_9_ ( .D(
        n29546), .DE(n30030), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3204), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[454]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__14_ ( 
        .D(n10651), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_14_ ( 
        .D(j202_soc_core_qspi_wb_wdat[14]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_bldc_core_00_wdata[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_14_ ( 
        .D(j202_soc_core_qspi_wb_wdat[14]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__i__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3390), .DE(j202_soc_core_j22_cpu_rf_N3391), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__i__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_6_ ( .D(
        j202_soc_core_j22_cpu_rf_N304), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__4_ ( .D(
        n11520), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__4_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__0_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N917), .DE(n12364), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_imm__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__6_ ( 
        .D(n10535), .DE(n12364), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__6_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__13_ ( 
        .D(n10655), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_13_ ( 
        .D(j202_soc_core_qspi_wb_wdat[13]), .CLK(wb_clk_i), .RESET_B(n29828), 
        .Q(j202_soc_core_bldc_core_00_wdata[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_13_ ( 
        .D(j202_soc_core_qspi_wb_wdat[13]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__i__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3388), .DE(j202_soc_core_j22_cpu_rf_N3391), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__i__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_5_ ( .D(
        n29638), .DE(n30056), .CLK(wb_clk_i), .Q(j202_soc_core_paddr[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_5_ ( 
        .D(j202_soc_core_paddr[5]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_reg_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__5_ ( .D(
        n12147), .DE(j202_soc_core_ahb2aqu_00_N127), .CLK(wb_clk_i), .Q(
        j202_soc_core_aquc_ADR__5_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_5_ ( 
        .D(j202_soc_core_aquc_ADR__5_), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_5_ ( .D(
        n29554), .DE(n30067), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_5_ ( .D(
        n29554), .DE(n30030), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_27_ ( .D(
        j202_soc_core_j22_cpu_rf_N325), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_27_ ( .D(n13098), 
        .DE(j202_soc_core_j22_cpu_rf_N2668), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_29_ ( .D(n12135), 
        .DE(j202_soc_core_j22_cpu_rf_N2668), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_16_ ( .D(
        n29482), .DE(n10998), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_14_ ( .D(
        n29547), .DE(n30030), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_6_ ( 
        .D(n29634), .DE(n10600), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_23_ ( .D(
        j202_soc_core_j22_cpu_rf_N321), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_23_ ( .D(n12134), 
        .DE(j202_soc_core_j22_cpu_rf_N2668), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2676), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__8_ ( .D(
        n29526), .DE(n30189), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_8_ ( 
        .D(j202_soc_core_qspi_wb_wdat[8]), .CLK(wb_clk_i), .RESET_B(n29827), 
        .Q(j202_soc_core_bldc_core_00_wdata[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_8_ ( 
        .D(j202_soc_core_qspi_wb_wdat[8]), .CLK(wb_clk_i), .RESET_B(n29745), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__i__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3386), .DE(j202_soc_core_j22_cpu_rf_N3391), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__i__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_4_ ( .D(
        n29637), .DE(n12277), .CLK(wb_clk_i), .Q(j202_soc_core_paddr[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_4_ ( 
        .D(j202_soc_core_paddr[4]), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_cmt_core_00_reg_addr[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_14_ ( 
        .D(n133), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_const0[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_13_ ( 
        .D(n132), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_const0[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_11_ ( 
        .D(n131), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_const0[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_10_ ( 
        .D(n130), .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_cmt_core_00_const0[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_8_ ( 
        .D(n129), .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_cmt_core_00_const0[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_15_ ( 
        .D(n128), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_const0[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_14_ ( 
        .D(n127), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_const1[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_13_ ( 
        .D(n126), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_const1[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_11_ ( 
        .D(n125), .CLK(wb_clk_i), .RESET_B(n12069), .Q(
        j202_soc_core_cmt_core_00_const1[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_10_ ( 
        .D(n124), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_const1[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_8_ ( 
        .D(n123), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_const1[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_15_ ( 
        .D(n122), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_const1[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__4_ ( .D(
        n12146), .DE(j202_soc_core_ahb2aqu_00_N127), .CLK(wb_clk_i), .Q(
        j202_soc_core_aquc_ADR__4_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_4_ ( 
        .D(j202_soc_core_aquc_ADR__4_), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_4_ ( .D(
        n29545), .DE(n30068), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_4_ ( .D(
        n29545), .DE(n30030), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_26_ ( .D(
        j202_soc_core_j22_cpu_rf_N324), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_26_ ( .D(n13097), 
        .DE(j202_soc_core_j22_cpu_rf_N2668), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_28_ ( .D(n12133), 
        .DE(j202_soc_core_j22_cpu_rf_N2668), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_30_ ( .D(n13102), 
        .DE(j202_soc_core_j22_cpu_rf_N2668), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_22_ ( .D(n12132), 
        .DE(j202_soc_core_j22_cpu_rf_N2668), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_24_ ( .D(n29635), 
        .DE(j202_soc_core_j22_cpu_rf_N2668), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_24_ ( 
        .D(n29442), .DE(n30067), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_len_reg_0_ ( .D(
        j202_soc_core_wbqspiflash_00_N736), .DE(
        j202_soc_core_wbqspiflash_00_N735), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_len[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_N671), .DE(n29754), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__4_ ( .D(
        n29443), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__4_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__12_ ( 
        .D(n29501), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_12_ ( 
        .D(j202_soc_core_qspi_wb_wdat[12]), .CLK(wb_clk_i), .RESET_B(n29745), 
        .Q(j202_soc_core_bldc_core_00_wdata[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_12_ ( 
        .D(j202_soc_core_qspi_wb_wdat[12]), .CLK(wb_clk_i), .RESET_B(n29828), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_12_ ( 
        .D(n121), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_const1[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_12_ ( 
        .D(n120), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_cmt_core_00_const0[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[12]), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cnt1[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[12]), .CLK(wb_clk_i), .RESET_B(
        n29830), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmf1_o_reg ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt1_to1), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cmf1) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[5]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cnt1[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[5]), .CLK(wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[5]), .CLK(wb_clk_i), 
        .RESET_B(n29827), .Q(j202_soc_core_prdata[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_5_ ( .D(
        j202_soc_core_ahb2apb_00_N133), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[101])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__5_ ( .D(
        n29445), .DE(n29747), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__5_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__5_ ( .D(
        n29560), .DE(n29647), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__5_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__5_ ( 
        .D(n10536), .DE(n12364), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__5_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_5_ ( .D(
        j202_soc_core_j22_cpu_ml_N308), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_6_ ( .D(
        j202_soc_core_j22_cpu_ml_N309), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_0_ ( .D(
        j202_soc_core_j22_cpu_rf_N298), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_0_ ( .D(
        n29636), .DE(n12277), .CLK(wb_clk_i), .Q(j202_soc_core_paddr[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_0_ ( 
        .D(j202_soc_core_paddr[0]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_reg_addr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__0_ ( .D(
        n12142), .DE(j202_soc_core_ahb2aqu_00_N127), .CLK(wb_clk_i), .Q(
        j202_soc_core_aquc_ADR__0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_0_ ( 
        .D(j202_soc_core_aquc_ADR__0_), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_address_reg_0_ ( .D(
        n29565), .DE(n29882), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_address[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_29_ ( .D(
        j202_soc_core_j22_cpu_rf_N327), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2656), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2658), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2670), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__m_ ( .D(
        j202_soc_core_j22_cpu_rf_N2640), .DE(j202_soc_core_j22_cpu_rf_N2639), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__m_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__1_ ( .D(
        n29507), .DE(n30189), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_1_ ( 
        .D(j202_soc_core_qspi_wb_wdat[1]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_bldc_core_00_wdata[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_1_ ( 
        .D(j202_soc_core_qspi_wb_wdat[1]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_1_ ( 
        .D(n119), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_cmt_core_00_const1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_1_ ( 
        .D(n118), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_const0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_1_ ( 
        .D(n117), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_cks1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_1_ ( 
        .D(n116), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_cks0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmstr_reg_reg_o_reg_1_ ( 
        .D(n115), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_str1) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_3_ ( .D(
        j202_soc_core_j22_cpu_id_idec_N894), .DE(n10601), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_opst[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_MEM_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ma_N55), .DE(n10600), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_MEM[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__5_ ( 
        .D(n10637), .DE(n10609), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__1_ ( 
        .D(n10633), .DE(n10609), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_4_ ( .D(
        n10606), .DE(n10601), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_opst[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rs__0_ ( 
        .D(n29597), .DE(n10609), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rs__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Wm__1_ ( 
        .D(n10639), .DE(n10645), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Wm__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_0_ ( .D(
        n10608), .DE(n10601), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_opst[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_MEM__3_ ( 
        .D(n10631), .DE(n10601), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_memop_MEM__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_MEM_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ma_N56), .DE(n10600), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_MEM[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_intack_reg ( .D(
        j202_soc_core_j22_cpu_id_idec_N822), .DE(n10603), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_intack) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intack_all_dout_reg_0_ ( 
        .D(n29542), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_cp_intack_all_0_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N3), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N4), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N5), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N6), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N9), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rte4_reg ( .D(n29649), .DE(
        n10603), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rte4) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Wm__2_ ( 
        .D(n10640), .DE(n10645), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Wm__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Wm__0_ ( 
        .D(n10638), .DE(n10645), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Wm__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_MEM__0_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N937), .DE(n10601), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_memop_MEM__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_MEM_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ma_N53), .DE(n10600), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_MEM[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_pc_hold_reg ( .D(
        n10607), .DE(n10601), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_pc_hold) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rm__0_ ( 
        .D(n11520), .DE(n11112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rm__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rm__1_ ( 
        .D(n29560), .DE(n11112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rm__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rm__2_ ( 
        .D(n29559), .DE(n11112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rm__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rm__3_ ( 
        .D(n12208), .DE(n11112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rm__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_We__2_ ( 
        .D(n10617), .DE(n10645), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_We__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_Ma__0_ ( 
        .D(n10542), .DE(n10611), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_memop_Ma__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__4_ ( 
        .D(n10537), .DE(n12364), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__4_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__8_ ( 
        .D(n10533), .DE(n12364), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__8_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__10_ ( 
        .D(n10531), .DE(n12364), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__10_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__4_ ( 
        .D(n10636), .DE(n10609), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__3_ ( 
        .D(n10635), .DE(n10609), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__2_ ( 
        .D(n10634), .DE(n10609), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_We__3_ ( 
        .D(n10618), .DE(n10645), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_We__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2652), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2643), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2644), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2645), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2646), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2647), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2648), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2649), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2642), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__3_ ( 
        .D(n10627), .DE(n10601), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__2_ ( 
        .D(n10626), .DE(n10601), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__1_ ( 
        .D(n10625), .DE(n10601), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_MEM__1_ ( 
        .D(n10629), .DE(n10601), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_memop_MEM__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_MEM_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ma_N54), .DE(n10600), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_MEM[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Rn__0_ ( 
        .D(n12339), .DE(n29879), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_M_Rn__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Rn__3_ ( 
        .D(n12340), .DE(n29879), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_M_Rn__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Rn__2_ ( 
        .D(n12032), .DE(n29879), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_M_Rn__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Rn__1_ ( 
        .D(n12030), .DE(n29879), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_M_Rn__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Wm__0_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N956), .DE(n10599), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Wm__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Wm__3_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N959), .DE(n10599), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Wm__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Wm__2_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N958), .DE(n10599), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Wm__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Wm__1_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N957), .DE(n10599), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Wm__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3337), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3336), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3335), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3334), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3324), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3313), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3314), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3316), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3317), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3319), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3311), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3326), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3309), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3338), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3340), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3341), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3342), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3343), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3307), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3302), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3303), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3304), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3305), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3300), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3299), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3298), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3297), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3296), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3295), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3287), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3284), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3280), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3278), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3276), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3274), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3273), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3272), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3271), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3270), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__s_ ( .D(
        j202_soc_core_j22_cpu_rf_N2628), .DE(j202_soc_core_j22_cpu_rf_N2627), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__s_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__0_ ( .D(
        j202_soc_core_j22_cpu_ml_N191), .DE(n29746), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__2_ ( .D(
        j202_soc_core_j22_cpu_ml_N193), .DE(n29746), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__3_ ( .D(
        j202_soc_core_j22_cpu_ml_N194), .DE(n29746), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__1_ ( .D(
        j202_soc_core_j22_cpu_ml_N192), .DE(n29746), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_5_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[5]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_6_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[6]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_7_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[7]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_5_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[5]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_6_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[6]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ml_N304), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[1]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[1]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_7_ ( .D(
        j202_soc_core_j22_cpu_ml_N310), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_7_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[7]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_20_ ( .D(
        j202_soc_core_j22_cpu_ml_N359), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_4_ ( .D(
        j202_soc_core_j22_cpu_ml_N416), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_26_ ( .D(
        j202_soc_core_j22_cpu_ml_N365), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_30_ ( .D(
        j202_soc_core_j22_cpu_ml_N369), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_18_ ( .D(
        j202_soc_core_j22_cpu_ml_N356), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ml_N414), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3372), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3373), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3374), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3375), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3376), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3377), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3378), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3379), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3370), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3369), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3361), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3359), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3355), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3352), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3349), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3348), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3347), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3345), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2710), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2713), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2712), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2711), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2703), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2704), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2705), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2706), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2707), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2708), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2695), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2688), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2692), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2686), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2679), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2680), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2681), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2682), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2684), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2678), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2784), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[92]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2787), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[95]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2786), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[94]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2785), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[93]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2777), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[86]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2778), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[87]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2779), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[88]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2780), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[89]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2781), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[90]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2782), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[91]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2769), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[79]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2762), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[73]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2766), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[77]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2760), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[71]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2753), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[65]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2754), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[66]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2755), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[67]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2756), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[68]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2752), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[64]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2747), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[60]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2750), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[63]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2749), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[62]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2748), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[61]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2740), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[54]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2741), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[55]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2742), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[56]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2743), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[57]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2744), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[58]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2745), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[59]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2732), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[47]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2725), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[41]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2729), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[45]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2723), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[39]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2716), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[33]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2717), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[34]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2718), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[35]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2719), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[36]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2715), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[32]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2821), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[124]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2824), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[127]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2823), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[126]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2822), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[125]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2814), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[118]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2815), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[119]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2816), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[120]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2817), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[121]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2818), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[122]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2819), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[123]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2806), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[111]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2799), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[105]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2803), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[109]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2797), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[103]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2790), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[97]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2791), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[98]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2792), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[99]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2793), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[100]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2789), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[96]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2858), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[156]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2861), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[159]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2860), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[158]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2859), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[157]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2851), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[150]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2852), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[151]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2853), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[152]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2854), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[153]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2855), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[154]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2856), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[155]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2843), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[143]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2836), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[137]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2840), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[141]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2834), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[135]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2827), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[129]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2828), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[130]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2829), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[131]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2830), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[132]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2826), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[128]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2895), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[188]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2898), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[191]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2897), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[190]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2896), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[189]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2888), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[182]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2889), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[183]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2890), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[184]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2891), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[185]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2892), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[186]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2893), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[187]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2880), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[175]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2873), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[169]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2877), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[173]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2871), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[167]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2864), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[161]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2865), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[162]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2866), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[163]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2867), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[164]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2863), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[160]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2932), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[220]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2935), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[223]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2934), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[222]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2933), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[221]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2925), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[214]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2926), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[215]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2927), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[216]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2928), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[217]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2929), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[218]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2930), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[219]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2917), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[207]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2910), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[201]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2914), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[205]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2908), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[199]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2901), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[193]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2902), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[194]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2903), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[195]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2904), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[196]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2900), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[192]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2969), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[252]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2972), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[255]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2971), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[254]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2970), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[253]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2962), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[246]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2963), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[247]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2964), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[248]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2965), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[249]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2966), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[250]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2967), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[251]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2954), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[239]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2947), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[233]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2951), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[237]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2945), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[231]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2938), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[225]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2939), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[226]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2940), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[227]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2941), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[228]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2937), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[224]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3006), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[284]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3009), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[287]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3008), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[286]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3007), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[285]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2999), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[278]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3000), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[279]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3001), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[280]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3002), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[281]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3003), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[282]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3004), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[283]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2991), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[271]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2984), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[265]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2988), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[269]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2982), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[263]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2975), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[257]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2976), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[258]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2977), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[259]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2978), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[260]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2974), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[256]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3046), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[318]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3045), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[317]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3044), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[316]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3036), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[310]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3037), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[311]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3038), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[312]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3039), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[313]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3040), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[314]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3041), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[315]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3028), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[303]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3021), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[297]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3025), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[301]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3019), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[295]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3012), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[289]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3013), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[290]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3014), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[291]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3015), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[292]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3011), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[288]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3080), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[347]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3083), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[350]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3082), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[349]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3081), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[348]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3073), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[341]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3074), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[342]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3075), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[343]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3076), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[344]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3077), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[345]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3078), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[346]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3065), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[334]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3058), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[328]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3062), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[332]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3056), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[326]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3049), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[320]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3050), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[321]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3051), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[322]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3052), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[323]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3048), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[319]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3117), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[379]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3120), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[382]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3119), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[381]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3118), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[380]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3110), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[373]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3111), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[374]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3112), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[375]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3113), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[376]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3114), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[377]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3115), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[378]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3102), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[366]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3095), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[360]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3099), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[364]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3093), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[358]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3086), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[352]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3087), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[353]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3088), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[354]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3089), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[355]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3085), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[351]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3154), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[411]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3157), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[414]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3156), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[413]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3155), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[412]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3147), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[405]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3148), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[406]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3149), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[407]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3150), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[408]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3151), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[409]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3152), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[410]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3139), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[398]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3132), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[392]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3136), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[396]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3130), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[390]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3123), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[384]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3124), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[385]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3125), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[386]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3126), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[387]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3122), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[383]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3191), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[443]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3194), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[446]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3193), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[445]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3192), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[444]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3184), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[437]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3185), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[438]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3186), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[439]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3187), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[440]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3188), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[441]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3189), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[442]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3176), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[430]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3169), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[424]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3173), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[428]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3167), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[422]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3160), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[416]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3161), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[417]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3162), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[418]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3163), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[419]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3159), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[415]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3228), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[475]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3231), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[478]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3230), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[477]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3229), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[476]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3221), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[469]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3222), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[470]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3223), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[471]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3224), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[472]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3225), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[473]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3226), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[474]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3213), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[462]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3206), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[456]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3210), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[460]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3197), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[448]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3198), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[449]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3199), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[450]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3200), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[451]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3196), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[447]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3265), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[507]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3268), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[510]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3267), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[509]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3266), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[508]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3258), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[501]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3259), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[502]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3260), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[503]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3261), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[504]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3262), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[505]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3263), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[506]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3250), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[494]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3243), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[488]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3247), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[492]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3241), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[486]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3234), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[480]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3235), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[481]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3236), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[482]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3237), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[483]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3239), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[485]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3233), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[479]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__23_ ( 
        .D(n29511), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[23]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_23_ ( 
        .D(j202_soc_core_qspi_wb_wdat[23]), .CLK(wb_clk_i), .RESET_B(n29827), 
        .Q(j202_soc_core_bldc_core_00_wdata[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__22_ ( 
        .D(n29510), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[22]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_22_ ( 
        .D(j202_soc_core_qspi_wb_wdat[22]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_bldc_core_00_wdata[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__21_ ( 
        .D(n29509), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[21]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_21_ ( 
        .D(j202_soc_core_qspi_wb_wdat[21]), .CLK(wb_clk_i), .RESET_B(n29827), 
        .Q(j202_soc_core_bldc_core_00_wdata[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__20_ ( 
        .D(n29508), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[20]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_20_ ( 
        .D(j202_soc_core_qspi_wb_wdat[20]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_bldc_core_00_wdata[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__18_ ( 
        .D(n29505), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[18]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_18_ ( 
        .D(j202_soc_core_qspi_wb_wdat[18]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_bldc_core_00_wdata[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__7_ ( .D(
        n29525), .DE(n30189), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_7_ ( 
        .D(j202_soc_core_qspi_wb_wdat[7]), .CLK(wb_clk_i), .RESET_B(n29827), 
        .Q(j202_soc_core_bldc_core_00_wdata[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_7_ ( 
        .D(j202_soc_core_qspi_wb_wdat[7]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_7_ ( 
        .D(n114), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_const1[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_7_ ( 
        .D(n113), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_cmt_core_00_const0[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_nxt_latch_status_0_), 
        .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__6_ ( .D(
        n29524), .DE(n30189), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_6_ ( 
        .D(j202_soc_core_qspi_wb_wdat[6]), .CLK(wb_clk_i), .RESET_B(n29827), 
        .Q(j202_soc_core_bldc_core_00_wdata[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_6_ ( 
        .D(j202_soc_core_qspi_wb_wdat[6]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_6_ ( 
        .D(n112), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_const1[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_6_ ( 
        .D(n111), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_cmt_core_00_const0[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_6_ ( 
        .D(n110), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_17_ ( 
        .D(n29875), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[17])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__5_ ( .D(
        n29523), .DE(n30189), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_5_ ( 
        .D(j202_soc_core_qspi_wb_wdat[5]), .CLK(wb_clk_i), .RESET_B(n29827), 
        .Q(j202_soc_core_bldc_core_00_wdata[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_5_ ( 
        .D(j202_soc_core_qspi_wb_wdat[5]), .CLK(wb_clk_i), .RESET_B(n29827), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_5_ ( 
        .D(n109), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_const1[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_5_ ( 
        .D(n108), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_const0[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_5_ ( 
        .D(n107), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_5_ ( 
        .D(n106), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_SEL__0_ ( .D(
        j202_soc_core_ahb2aqu_00_N161), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_SEL__0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_RDRXD1_reg ( .D(n29541), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_uart_RDRXD1) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_rx_fifo_rp_reg_0_ ( .D(n105), 
        .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_uart_TOP_rx_fifo_rp[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_rx_fifo_rp_reg_1_ ( .D(n104), 
        .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_uart_TOP_rx_fifo_rp[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_1_ ( .D(n103), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_uart_din_i[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_5_ ( .D(n102), .CLK(
        wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_uart_din_i[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_6_ ( .D(n101), .CLK(
        wb_clk_i), .RESET_B(n29828), .Q(j202_soc_core_uart_din_i[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_7_ ( .D(n100), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_uart_din_i[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_WRTXD1_reg ( .D(n29483), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_uart_WRTXD1) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_tx_fifo_wp_reg_0_ ( .D(n99), 
        .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_uart_TOP_tx_fifo_wp[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_tx_fifo_wp_reg_1_ ( .D(n98), 
        .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_uart_TOP_tx_fifo_wp[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__7_ ( .D(
        j202_soc_core_uart_din_i[7]), .DE(n29864), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__6_ ( .D(
        j202_soc_core_uart_din_i[6]), .DE(n29864), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__5_ ( .D(
        j202_soc_core_uart_din_i[5]), .DE(n29864), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__1_ ( .D(
        j202_soc_core_uart_din_i[1]), .DE(n29864), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__7_ ( .D(
        j202_soc_core_uart_din_i[7]), .DE(n29863), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__6_ ( .D(
        j202_soc_core_uart_din_i[6]), .DE(n29863), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__5_ ( .D(
        j202_soc_core_uart_din_i[5]), .DE(n29863), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__1_ ( .D(
        j202_soc_core_uart_din_i[1]), .DE(n29863), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__7_ ( .D(
        j202_soc_core_uart_din_i[7]), .DE(n29880), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__6_ ( .D(
        j202_soc_core_uart_din_i[6]), .DE(n29880), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__5_ ( .D(
        j202_soc_core_uart_din_i[5]), .DE(n29880), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__1_ ( .D(
        j202_soc_core_uart_din_i[1]), .DE(n29880), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__7_ ( .D(
        j202_soc_core_uart_din_i[7]), .DE(n29865), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__6_ ( .D(
        j202_soc_core_uart_din_i[6]), .DE(n29865), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__5_ ( .D(
        j202_soc_core_uart_din_i[5]), .DE(n29865), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__1_ ( .D(
        j202_soc_core_uart_din_i[1]), .DE(n29865), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_SEL__2_ ( .D(
        j202_soc_core_ahb2aqu_00_N163), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_SEL__2_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_7_ ( .D(n97), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_uart_div1[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_6_ ( .D(n96), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_uart_div1[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_5_ ( .D(n95), .CLK(
        wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_uart_div1[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_4_ ( .D(n94), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_uart_div1[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_2_ ( .D(n93), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_uart_div1[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_2_ ( .D(
        j202_soc_core_j22_cpu_rf_N300), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N301), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N302), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_1_ ( .D(
        j202_soc_core_j22_cpu_rf_N299), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3346), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_28_ ( .D(
        j202_soc_core_j22_cpu_rf_N326), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_28_ ( .D(
        j202_soc_core_j22_cpu_ml_N367), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_31_ ( .D(n29646), 
        .DE(n29748), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_pc[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_31_ ( .D(
        j202_soc_core_j22_cpu_ml_N370), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_25_ ( .D(
        j202_soc_core_j22_cpu_rf_N323), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_25_ ( .D(
        j202_soc_core_j22_cpu_ml_N364), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_9_ ( .D(
        j202_soc_core_j22_cpu_ml_N421), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_24_ ( .D(
        j202_soc_core_j22_cpu_rf_N322), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_24_ ( .D(
        j202_soc_core_j22_cpu_ml_N363), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_22_ ( .D(
        j202_soc_core_j22_cpu_rf_N320), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_22_ ( .D(
        j202_soc_core_j22_cpu_ml_N361), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Ra__1_ ( 
        .D(n10621), .DE(n10609), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Ra__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_Ma__1_ ( 
        .D(n10541), .DE(n10611), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_memop_Ma__1_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_req_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_req_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intr_req_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ml_N303), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[0]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[0]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__0_ ( .D(
        n29498), .DE(n30189), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_0_ ( 
        .D(j202_soc_core_qspi_wb_wdat[0]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_bldc_core_00_wdata[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_0_ ( .D(n92), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_uart_din_i[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__0_ ( .D(
        j202_soc_core_uart_din_i[0]), .DE(n29865), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__0_ ( .D(
        j202_soc_core_uart_din_i[0]), .DE(n29880), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__0_ ( .D(
        j202_soc_core_uart_din_i[0]), .DE(n29863), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__0_ ( .D(
        j202_soc_core_uart_din_i[0]), .DE(n29864), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_0_ ( 
        .D(j202_soc_core_qspi_wb_wdat[0]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_0_ ( 
        .D(n91), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_const1[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_0_ ( 
        .D(n90), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_cmt_core_00_const0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_0_ ( 
        .D(n89), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_cmt_core_00_cks1[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[0]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[1]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cnt1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[1]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[1]), .CLK(wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[2]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[3]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[4]), .CLK(wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[5]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[6]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[7]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[8]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[9]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_0_ ( 
        .D(n88), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_cks0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmstr_reg_reg_o_reg_0_ ( 
        .D(n87), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_cmt_core_00_str0) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[9]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[0]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_1_ ( 
        .D(n29733), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_2_ ( 
        .D(n29725), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_3_ ( 
        .D(n29732), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_4_ ( 
        .D(n29724), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[5]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_6_ ( 
        .D(n29726), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[7]), .CLK(wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[8]), .CLK(wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[8]) );
  sky130_fd_sc_hd__dfstp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[0]), .CLK(wb_clk_i), .SET_B(n29827), .Q(j202_soc_core_cmt_core_00_cnt1[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[0]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ml_N305), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[2]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[2]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__2_ ( .D(
        n29518), .DE(n30189), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_2_ ( 
        .D(j202_soc_core_qspi_wb_wdat[2]), .CLK(wb_clk_i), .RESET_B(n29745), 
        .Q(j202_soc_core_bldc_core_00_wdata[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_2_ ( .D(n86), .CLK(
        wb_clk_i), .RESET_B(n29828), .Q(j202_soc_core_uart_din_i[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__2_ ( .D(
        j202_soc_core_uart_din_i[2]), .DE(n29865), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__2_ ( .D(
        j202_soc_core_uart_din_i[2]), .DE(n29880), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__2_ ( .D(
        j202_soc_core_uart_din_i[2]), .DE(n29863), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__2_ ( .D(
        j202_soc_core_uart_din_i[2]), .DE(n29864), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_2_ ( 
        .D(j202_soc_core_qspi_wb_wdat[2]), .CLK(wb_clk_i), .RESET_B(n29827), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_2_ ( 
        .D(n85), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_const1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_2_ ( 
        .D(n84), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_const0[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_2_ ( 
        .D(n83), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_2_ ( 
        .D(n82), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[2]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cnt1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[2]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ml_N306), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[3]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[3]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__3_ ( .D(
        n29521), .DE(n30189), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_3_ ( 
        .D(j202_soc_core_qspi_wb_wdat[3]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_bldc_core_00_wdata[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_3_ ( .D(n81), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_uart_din_i[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__3_ ( .D(
        j202_soc_core_uart_din_i[3]), .DE(n29865), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__3_ ( .D(
        j202_soc_core_uart_din_i[3]), .DE(n29880), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__3_ ( .D(
        j202_soc_core_uart_din_i[3]), .DE(n29863), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__3_ ( .D(
        j202_soc_core_uart_din_i[3]), .DE(n29864), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_3_ ( 
        .D(j202_soc_core_qspi_wb_wdat[3]), .CLK(wb_clk_i), .RESET_B(n29828), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_3_ ( 
        .D(n80), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_cmt_core_00_const1[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_3_ ( 
        .D(n79), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_const0[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_3_ ( 
        .D(n78), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_3_ ( 
        .D(n77), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[3]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cnt1[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[3]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_4_ ( .D(
        j202_soc_core_j22_cpu_ml_N307), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_4_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[4]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_4_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[4]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__4_ ( .D(
        n29522), .DE(n30189), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_4_ ( 
        .D(j202_soc_core_qspi_wb_wdat[4]), .CLK(wb_clk_i), .RESET_B(n29827), 
        .Q(j202_soc_core_bldc_core_00_wdata[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_4_ ( .D(n76), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_uart_din_i[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__4_ ( .D(
        j202_soc_core_uart_din_i[4]), .DE(n29865), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__4_ ( .D(
        j202_soc_core_uart_din_i[4]), .DE(n29880), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__4_ ( .D(
        j202_soc_core_uart_din_i[4]), .DE(n29863), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__4_ ( .D(
        j202_soc_core_uart_din_i[4]), .DE(n29864), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_4_ ( 
        .D(j202_soc_core_qspi_wb_wdat[4]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_4_ ( 
        .D(n75), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_const1[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_4_ ( 
        .D(n74), .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_cmt_core_00_const0[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_4_ ( 
        .D(n73), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_4_ ( 
        .D(n72), .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[4]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cnt1[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[4]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_9_ ( .D(
        j202_soc_core_j22_cpu_ml_N312), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_9_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[9]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_9_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[9]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_15_ ( .D(
        j202_soc_core_j22_cpu_ml_N318), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_15_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[15]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_15_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[15]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_18_ ( .D(
        j202_soc_core_j22_cpu_ml_N321), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_18_ ( .D(n29844), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_mach[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_18_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[18]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_20_ ( .D(
        j202_soc_core_j22_cpu_ml_N324), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_20_ ( .D(n29843), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_mach[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_20_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[20]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_22_ ( .D(
        j202_soc_core_j22_cpu_ml_N326), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_22_ ( .D(n29842), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_mach[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_22_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[22]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_23_ ( .D(
        j202_soc_core_j22_cpu_ml_N327), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_23_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[23]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_23_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[23]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_24_ ( .D(
        j202_soc_core_j22_cpu_ml_N328), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_24_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[24]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_24_ ( .D(n29841), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_mach[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_25_ ( .D(
        j202_soc_core_j22_cpu_ml_N329), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_25_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[25]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_25_ ( .D(n29840), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_mach[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_26_ ( .D(
        j202_soc_core_j22_cpu_ml_N330), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_26_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[26]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_26_ ( .D(n29839), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_mach[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_27_ ( .D(
        j202_soc_core_j22_cpu_ml_N331), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_27_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[27]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_27_ ( .D(n29838), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_mach[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_28_ ( .D(
        j202_soc_core_j22_cpu_ml_N332), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_28_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[28]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_28_ ( .D(n29837), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_mach[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_29_ ( .D(
        j202_soc_core_j22_cpu_ml_N333), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_29_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[29]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_29_ ( .D(n29836), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_mach[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_30_ ( .D(
        j202_soc_core_j22_cpu_ml_N334), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_30_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[30]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_30_ ( .D(n29835), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_mach[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_31_ ( .D(
        j202_soc_core_j22_cpu_ml_N335), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_31_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[31]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_31_ ( .D(n29834), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_mach[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__31_ ( 
        .D(n29520), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[31]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_7_ ( .D(n71), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_uart_div0[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_3_ ( .D(
        j202_soc_core_wbqspiflash_00_N727), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_9_ ( 
        .D(j202_soc_core_wbqspiflash_00_N623), .DE(n29631), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_N614), .DE(n29631), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_8_ ( 
        .D(j202_soc_core_wbqspiflash_00_N622), .DE(n29631), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_N621), .DE(n29631), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_N620), .DE(n29631), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_N619), .DE(n29631), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_N618), .DE(n29631), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_N617), .DE(n29631), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_N616), .DE(n29631), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_N615), .DE(n29631), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_alt_ctrl_reg ( .D(
        j202_soc_core_wbqspiflash_00_N86), .DE(n29745), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_alt_ctrl) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_alt_cmd_reg ( .D(
        j202_soc_core_wbqspiflash_00_N85), .DE(n29830), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_alt_cmd) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_ctrl_reg ( .D(
        j202_soc_core_wbqspiflash_00_N744), .DE(
        j202_soc_core_wbqspiflash_00_N743), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_ctrl) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_wr_reg ( .D(
        j202_soc_core_wbqspiflash_00_N734), .DE(
        j202_soc_core_wbqspiflash_00_N733), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_wr) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_0_ ( 
        .D(j202_soc_core_qspi_wb_addr[2]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_18_ ( 
        .D(j202_soc_core_qspi_wb_addr[20]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_16_ ( 
        .D(j202_soc_core_qspi_wb_addr[18]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_15_ ( 
        .D(j202_soc_core_qspi_wb_addr[17]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_14_ ( 
        .D(j202_soc_core_qspi_wb_addr[16]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_12_ ( 
        .D(j202_soc_core_qspi_wb_addr[14]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_7_ ( 
        .D(j202_soc_core_qspi_wb_addr[9]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_5_ ( 
        .D(j202_soc_core_qspi_wb_addr[7]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_4_ ( 
        .D(j202_soc_core_qspi_wb_addr[6]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_3_ ( 
        .D(j202_soc_core_qspi_wb_addr[5]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_2_ ( 
        .D(j202_soc_core_qspi_wb_addr[4]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_1_ ( 
        .D(j202_soc_core_qspi_wb_addr[3]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_4_ ( .D(
        j202_soc_core_wbqspiflash_00_N728), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_spd_reg ( .D(
        j202_soc_core_wbqspiflash_00_N592), .DE(
        j202_soc_core_wbqspiflash_00_N746), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_spd) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_spd_reg ( 
        .D(j202_soc_core_wbqspiflash_00_spi_spd), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N423), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_mod_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N356), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N354), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N358), .DE(n23851), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_interrupt_reg ( .D(
        j202_soc_core_wbqspiflash_00_N741), .DE(
        j202_soc_core_wbqspiflash_00_N740), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_int) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_20_ ( 
        .D(n29582), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[20])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N323), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N359), .DE(n23851), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N324), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N360), .DE(n23851), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N325), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N361), .DE(n23851), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N326), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_4_ ( 
        .D(n29702), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N327), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_5_ ( 
        .D(n29715), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N328), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_6_ ( 
        .D(n29719), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N329), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_7_ ( 
        .D(n29714), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N330), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_8_ ( 
        .D(n29705), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_8_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N331), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_9_ ( 
        .D(n29713), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_9_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N332), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_10_ ( 
        .D(n29701), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_10_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N333), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_11_ ( 
        .D(n29712), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_11_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N334), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_12_ ( 
        .D(n29721), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_12_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N335), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_13_ ( 
        .D(n29711), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_13_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N336), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_14_ ( 
        .D(n29718), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_14_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N337), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_15_ ( 
        .D(n29710), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_15_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N338), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_16_ ( 
        .D(n29720), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_16_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N339), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_17_ ( 
        .D(n29709), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_17_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N340), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_18_ ( 
        .D(n29717), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_18_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N341), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_19_ ( 
        .D(n29704), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_19_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N342), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_20_ ( 
        .D(n29700), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_20_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N343), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_21_ ( 
        .D(n29699), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_21_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N344), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_22_ ( 
        .D(n29698), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_22_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N345), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_23_ ( 
        .D(n29697), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_23_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N346), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_24_ ( 
        .D(n29696), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_24_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N347), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_25_ ( 
        .D(n29716), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_25_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N348), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_26_ ( 
        .D(n29703), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_26_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N349), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_27_ ( 
        .D(n29708), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_27_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N350), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_28_ ( 
        .D(n29695), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_28_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N351), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_29_ ( 
        .D(n29707), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_29_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N352), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_30_ ( 
        .D(n29706), .DE(n23851), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_30_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N353), .DE(n29753), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_31_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N389), .DE(n23851), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_dir_reg ( .D(
        j202_soc_core_wbqspiflash_00_N594), .DE(
        j202_soc_core_wbqspiflash_00_N747), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_dir) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_dir_reg ( 
        .D(j202_soc_core_wbqspiflash_00_spi_dir), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N423), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_dir) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_mod_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N355), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N354), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_cmd_reg ( .D(
        j202_soc_core_wbqspiflash_00_N663), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_cmd) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_31_ ( 
        .D(j202_soc_core_qspi_wb_wdat[31]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_23_ ( 
        .D(j202_soc_core_qspi_wb_wdat[23]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_22_ ( 
        .D(j202_soc_core_qspi_wb_wdat[22]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_21_ ( 
        .D(j202_soc_core_qspi_wb_wdat[21]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_N718), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_20_ ( 
        .D(j202_soc_core_qspi_wb_wdat[20]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_N717), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_18_ ( 
        .D(j202_soc_core_qspi_wb_wdat[18]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_N715), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_15_ ( 
        .D(j202_soc_core_qspi_wb_wdat[15]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_N712), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_14_ ( 
        .D(j202_soc_core_qspi_wb_wdat[14]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_N711), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_13_ ( 
        .D(j202_soc_core_qspi_wb_wdat[13]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_11_ ( 
        .D(j202_soc_core_qspi_wb_wdat[11]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_10_ ( 
        .D(j202_soc_core_qspi_wb_wdat[10]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_8_ ( 
        .D(j202_soc_core_qspi_wb_wdat[8]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_7_ ( 
        .D(j202_soc_core_qspi_wb_wdat[7]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_6_ ( 
        .D(j202_soc_core_qspi_wb_wdat[6]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_6_ ( .D(
        n10569), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_5_ ( 
        .D(j202_soc_core_qspi_wb_wdat[5]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_4_ ( 
        .D(j202_soc_core_qspi_wb_wdat[4]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_4_ ( .D(
        n10571), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_3_ ( 
        .D(j202_soc_core_qspi_wb_wdat[3]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_2_ ( 
        .D(j202_soc_core_qspi_wb_wdat[2]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_2_ ( .D(
        n10573), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_1_ ( 
        .D(j202_soc_core_qspi_wb_wdat[1]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_1_ ( .D(
        j202_soc_core_wbqspiflash_00_N629), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_0_ ( 
        .D(j202_soc_core_qspi_wb_wdat[0]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_0_ ( .D(
        j202_soc_core_wbqspiflash_00_N628), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_N611), .DE(
        j202_soc_core_wbqspiflash_00_N750), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_N612), .DE(
        j202_soc_core_wbqspiflash_00_N750), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_N605), .DE(
        j202_soc_core_wbqspiflash_00_N749), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_N606), .DE(
        j202_soc_core_wbqspiflash_00_N749), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_N607), .DE(
        j202_soc_core_wbqspiflash_00_N749), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_N608), .DE(
        j202_soc_core_wbqspiflash_00_N749), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_N609), .DE(
        j202_soc_core_wbqspiflash_00_N749), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_N613), .DE(
        j202_soc_core_wbqspiflash_00_N749), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_8_ ( 
        .D(n29693), .DE(n29876), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_9_ ( 
        .D(n29692), .DE(n29876), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_10_ ( 
        .D(n29691), .DE(n29876), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_11_ ( 
        .D(n29690), .DE(n29876), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_12_ ( 
        .D(n29689), .DE(n29754), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_13_ ( 
        .D(n29688), .DE(n29876), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_22_ ( 
        .D(n29687), .DE(n29754), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_23_ ( 
        .D(n29686), .DE(n29876), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_24_ ( 
        .D(n29685), .DE(n29876), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_25_ ( 
        .D(n29684), .DE(n29876), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_26_ ( 
        .D(n29683), .DE(n29754), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_quad_mode_enabled_reg ( 
        .D(j202_soc_core_wbqspiflash_00_N739), .DE(
        j202_soc_core_wbqspiflash_00_N738), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_N667), .DE(n29754), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_N672), .DE(n29876), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_N673), .DE(n29876), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_N674), .DE(n29754), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_3_ ( .D(
        n10572), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_14_ ( 
        .D(j202_soc_core_wbqspiflash_00_N681), .DE(n29754), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_15_ ( 
        .D(j202_soc_core_wbqspiflash_00_N682), .DE(n29754), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_18_ ( 
        .D(j202_soc_core_wbqspiflash_00_N685), .DE(n29876), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_20_ ( 
        .D(j202_soc_core_wbqspiflash_00_N687), .DE(n29754), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_21_ ( 
        .D(j202_soc_core_wbqspiflash_00_N688), .DE(n29754), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_27_ ( 
        .D(j202_soc_core_wbqspiflash_00_N694), .DE(n29754), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_29_ ( 
        .D(j202_soc_core_wbqspiflash_00_N696), .DE(n29876), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_31_ ( 
        .D(j202_soc_core_wbqspiflash_00_N698), .DE(n29754), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_32_ ( .D(
        j202_soc_core_j22_cpu_ml_N336), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[32]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_19_ ( .D(
        j202_soc_core_j22_cpu_ml_N322), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_19_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[19]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_19_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[19]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3364), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3328), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3289), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2697), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2734), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[49]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2771), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[81]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2808), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[113]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2845), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[145]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2882), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[177]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2919), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[209]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2956), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[241]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2993), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[273]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3030), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[305]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3067), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[336]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3104), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[368]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3141), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[400]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3178), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[432]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3215), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[464]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3252), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[496]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_17_ ( .D(n13092), 
        .DE(j202_soc_core_j22_cpu_rf_N2668), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3363), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3327), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3288), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2696), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2733), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[48]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2770), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[80]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2807), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[112]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2844), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[144]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2881), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[176]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2918), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[208]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2955), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[240]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2992), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[272]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3029), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[304]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3066), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[335]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3103), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[367]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3140), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[399]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3177), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[431]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3214), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[463]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3251), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[495]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_16_ ( .D(n12131), 
        .DE(j202_soc_core_j22_cpu_rf_N2668), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3354), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3318), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3279), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2687), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2724), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[40]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2761), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[72]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2798), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[104]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2835), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[136]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2872), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[168]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2909), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[200]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2946), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[232]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2983), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[264]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3020), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[296]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3057), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[327]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3094), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[359]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3131), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[391]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3168), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[423]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3205), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[455]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3242), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[487]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2651), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3356), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3321), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3281), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2689), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2726), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[42]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2763), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[74]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2800), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[106]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2837), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[138]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2874), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[170]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2911), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[202]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2948), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[234]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2985), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[266]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3022), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[298]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3059), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[329]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3096), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[361]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3133), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[393]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3170), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[425]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3207), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[457]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3244), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[489]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2653), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3358), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3283), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2691), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2728), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[44]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2765), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[76]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2802), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[108]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2839), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[140]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2876), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[172]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2913), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[204]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2950), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[236]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2987), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[268]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3024), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[300]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3061), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[331]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3098), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[363]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3135), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[395]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3172), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[427]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3209), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[459]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3246), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[491]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2655), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3357), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3322), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3282), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2690), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2727), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[43]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2764), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[75]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2801), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[107]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2838), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[139]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2875), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[171]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2912), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[203]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2949), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[235]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2986), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[267]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3023), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[299]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3060), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[330]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3097), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[362]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3134), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[394]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3171), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[426]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3208), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[458]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3245), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[490]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2654), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_11_ ( .D(
        j202_soc_core_j22_cpu_ml_N314), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_11_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[11]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_11_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[11]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_11_ ( .D(
        j202_soc_core_j22_cpu_rf_N309), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__27_ ( 
        .D(n29515), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[27]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_3_ ( .D(n70), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_uart_div0[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_27_ ( 
        .D(j202_soc_core_qspi_wb_wdat[27]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_11_ ( 
        .D(n29549), .DE(n30067), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_9_ ( 
        .D(j202_soc_core_qspi_wb_addr[11]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_11_ ( .D(
        n29549), .DE(n30030), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3360), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3325), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3286), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2694), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2731), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[46]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2768), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[78]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2805), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[110]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2842), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[142]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2879), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[174]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2916), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[206]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2953), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[238]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2990), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[270]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3027), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[302]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3064), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[333]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3101), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[365]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3138), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[397]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3175), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[429]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3212), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[461]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3249), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[493]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2657), .DE(j202_soc_core_j22_cpu_rf_N2668), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_14_ ( .D(
        j202_soc_core_j22_cpu_ml_N317), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_14_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[14]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_14_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[14]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_14_ ( .D(
        j202_soc_core_j22_cpu_ml_N426), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_14_ ( .D(
        j202_soc_core_j22_cpu_rf_N312), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__30_ ( 
        .D(n29519), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[30]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_6_ ( .D(n69), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_uart_div0[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_30_ ( 
        .D(j202_soc_core_qspi_wb_wdat[30]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_12_ ( .D(
        j202_soc_core_j22_cpu_ml_N315), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_12_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[12]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_12_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[12]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_12_ ( .D(
        j202_soc_core_j22_cpu_ml_N424), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_12_ ( .D(
        j202_soc_core_j22_cpu_rf_N310), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__28_ ( 
        .D(n29516), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[28]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_4_ ( .D(n68), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_uart_div0[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_28_ ( 
        .D(j202_soc_core_qspi_wb_wdat[28]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_1_ ( 
        .D(n29866), .DE(n10600), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_01_state_reg_0_ ( .D(
        j202_soc_core_ahb2apb_01_N89), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_01_state[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_01_state_reg_2_ ( .D(
        j202_soc_core_ahb2apb_01_N91), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_01_state[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_01_state_reg_1_ ( .D(
        j202_soc_core_ahb2apb_01_N90), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_01_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_01_N23), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_hsize_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_01_N57), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_01_hsize_buf[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_hsize_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_01_N56), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_01_hsize_buf[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_hwrite_buf_reg ( .D(
        j202_soc_core_ahb2apb_01_N55), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_pwrite[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_11_ ( .D(
        j202_soc_core_ahb2apb_01_N34), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_9_ ( .D(
        j202_soc_core_ahb2apb_01_N32), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_7_ ( .D(
        j202_soc_core_ahb2apb_01_N30), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_6_ ( .D(
        j202_soc_core_ahb2apb_01_N29), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_5_ ( .D(
        j202_soc_core_ahb2apb_01_N28), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_4_ ( .D(
        j202_soc_core_ahb2apb_01_N27), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_3_ ( .D(
        j202_soc_core_ahb2apb_01_N26), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_2_ ( .D(
        j202_soc_core_ahb2apb_01_N25), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_01_N24), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_12_ ( 
        .D(n29473), .DE(n30068), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_10_ ( 
        .D(j202_soc_core_qspi_wb_addr[12]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_12_ ( .D(
        n29473), .DE(n10998), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_10_ ( .D(
        j202_soc_core_j22_cpu_ml_N313), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_10_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[10]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_10_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[10]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_10_ ( .D(
        j202_soc_core_j22_cpu_ml_N422), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N308), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__26_ ( 
        .D(n29514), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[26]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_2_ ( .D(n67), .CLK(
        wb_clk_i), .RESET_B(n29828), .Q(j202_soc_core_uart_div0[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_26_ ( 
        .D(j202_soc_core_qspi_wb_wdat[26]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_10_ ( .D(
        j202_soc_core_ahb2apb_01_N33), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_10_ ( 
        .D(n29548), .DE(n30068), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_8_ ( 
        .D(j202_soc_core_qspi_wb_addr[10]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_10_ ( .D(
        n29548), .DE(n10998), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_8_ ( .D(
        j202_soc_core_j22_cpu_ml_N311), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_8_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[8]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_8_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[8]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__q_ ( .D(
        j202_soc_core_j22_cpu_rf_N2638), .DE(j202_soc_core_j22_cpu_rf_N2637), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__q_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_8_ ( .D(
        j202_soc_core_j22_cpu_ml_N420), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_8_ ( .D(
        j202_soc_core_j22_cpu_rf_N306), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__24_ ( 
        .D(n29512), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[24]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_0_ ( .D(n66), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_uart_div0[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_24_ ( 
        .D(j202_soc_core_qspi_wb_wdat[24]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_8_ ( .D(
        j202_soc_core_ahb2apb_01_N31), .DE(n12276), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_15__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_15__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_15_ ( 
        .D(n29567), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[15])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_14__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_14__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_14_ ( 
        .D(n29576), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[14])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_13__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_13__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_13_ ( 
        .D(n29566), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[13])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_12__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_12__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_12_ ( 
        .D(n29562), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[12])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_11__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_11__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_11_ ( 
        .D(n29590), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[11])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_10__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_10__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_10_ ( 
        .D(n29558), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[10])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_9__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_9__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_9_ ( 
        .D(n29574), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_8__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_8__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_8_ ( 
        .D(n29575), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_7__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_7__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_7_ ( 
        .D(n29572), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_6__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_6__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_6_ ( 
        .D(n29573), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_5__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_5__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_5_ ( 
        .D(n29570), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_4__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_4__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_4_ ( 
        .D(n29571), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_3__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_3__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_3_ ( 
        .D(n29584), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_2__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_2__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_2_ ( 
        .D(n29561), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_1__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_1__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_1_ ( 
        .D(n29544), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_0__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_0__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_0_ ( 
        .D(n29543), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[64]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[65]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[66]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[67]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[68]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[69]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[70]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[71]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[72]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[74]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[75]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[77]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[78]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[79]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[82]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[84]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[85]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[86]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[87]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[88]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[90]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[91]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[92]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[94]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[95]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[96]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[97]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[98]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[99]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[100]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[101]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[102]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[103]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[104]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[106]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[107]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[109]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[110]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[111]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[114]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[116]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[117]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[118]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[119]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[120]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[122]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[123]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[124]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[126]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[127]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[33]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[34]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[35]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[36]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[37]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[38]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[39]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[40]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[42]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[43]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[46]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[47]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[50]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[52]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[54]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[55]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[56]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[58]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[59]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[60]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[62]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[63]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[32]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[64]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[96]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[33]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[65]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[97]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[66]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[98]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[35]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[67]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[99]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[68]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[37]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[69]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[101]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[70]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[102]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[71]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[103]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[56]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[88]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[120]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[57]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[89]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[121]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[90]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[122]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[59]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[91]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[123]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[92]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[61]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[93]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[125]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[94]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[126]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[95]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[127]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[40]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[72]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[104]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[41]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[73]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[105]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[74]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[106]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[43]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[75]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[107]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[76]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[45]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[77]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[109]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[78]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[110]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[79]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[111]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[48]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[80]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[112]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[49]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[81]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[113]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[82]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[114]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[51]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[83]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[115]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[84]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[53]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[85]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[117]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[86]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[118]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[87]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[119]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_2_ ( .D(
        j202_soc_core_ahb2apb_01_N130), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[66]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_3_ ( .D(
        j202_soc_core_ahb2apb_01_N131), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[67]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_4_ ( .D(
        j202_soc_core_ahb2apb_01_N132), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[68]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_5_ ( .D(
        j202_soc_core_ahb2apb_01_N133), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[69]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_6_ ( .D(
        j202_soc_core_ahb2apb_01_N134), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[70]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_7_ ( .D(
        j202_soc_core_ahb2apb_01_N135), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[71]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_11_ ( .D(
        j202_soc_core_ahb2apb_01_N139), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[75]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_15_ ( .D(
        j202_soc_core_ahb2apb_01_N143), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[79]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_20_ ( .D(
        j202_soc_core_ahb2apb_01_N148), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[84]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_21_ ( .D(
        j202_soc_core_ahb2apb_01_N149), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[85]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_22_ ( .D(
        j202_soc_core_ahb2apb_01_N150), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[86]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_23_ ( .D(
        j202_soc_core_ahb2apb_01_N151), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[87]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_01_N128), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[64]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_10_ ( .D(
        j202_soc_core_ahb2apb_01_N138), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[74]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_24_ ( .D(
        j202_soc_core_ahb2apb_01_N152), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[88]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_26_ ( .D(
        j202_soc_core_ahb2apb_01_N154), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[90]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_27_ ( .D(
        j202_soc_core_ahb2apb_01_N155), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[91]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_28_ ( .D(
        j202_soc_core_ahb2apb_01_N156), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[92]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_30_ ( .D(
        j202_soc_core_ahb2apb_01_N158), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[94]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_31_ ( .D(
        j202_soc_core_ahb2apb_01_N159), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[95]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_8_ ( .D(
        n29552), .DE(n30068), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_6_ ( 
        .D(j202_soc_core_qspi_wb_addr[8]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_8_ ( .D(
        n10567), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_8_ ( .D(
        n29552), .DE(n10998), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_CE__0_ ( .D(
        j202_soc_core_ahb2aqu_00_N97), .DE(j202_soc_core_ahb2aqu_00_N95), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_CE__0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_state_reg_1_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_wb_slave_00_nxt_state_1_), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_22_ ( 
        .D(n65), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_21_ ( 
        .D(n64), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_20_ ( 
        .D(n63), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_18_ ( 
        .D(n62), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_15_ ( 
        .D(n61), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_14_ ( 
        .D(n60), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_13_ ( 
        .D(n59), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_12_ ( 
        .D(n58), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_11_ ( 
        .D(n57), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_bldc_core_00_pwm_period[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_10_ ( 
        .D(n56), .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_bldc_core_00_pwm_period[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_8_ ( 
        .D(n55), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_pwm_period[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_7_ ( 
        .D(n54), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_pwm_period[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_6_ ( 
        .D(n53), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_bldc_core_00_pwm_period[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_5_ ( 
        .D(n52), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_pwm_period[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_4_ ( 
        .D(n51), .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_bldc_core_00_pwm_period[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_3_ ( 
        .D(n50), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_pwm_period[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_2_ ( 
        .D(n49), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_pwm_period[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_1_ ( 
        .D(n48), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_pwm_period[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_0_ ( 
        .D(n47), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_pwm_period[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_23_ ( 
        .D(n46), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bcr_00_reg_o_reg_0_ ( 
        .D(n45), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_pwm_en) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bcr_00_reg_o_reg_1_ ( 
        .D(n44), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_adc_en) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ccr_00_reg_o_reg_1_ ( 
        .D(n43), .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_bldc_core_00_comm[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ccr_00_reg_o_reg_0_ ( 
        .D(n42), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_comm[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ccr_00_reg_o_reg_2_ ( 
        .D(n41), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_comm[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_00_reg_o_reg_0_ ( 
        .D(n40), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_wen_1_reg ( 
        .D(n29585), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_wen) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_00_reg_o_reg_0_ ( 
        .D(n39), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_reg_0_ ( 
        .D(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_nxt_latch_status_0_), .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bldc_int_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_nxt_bldc_int), 
        .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_bldc_int) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_19_ ( 
        .D(n29586), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[19])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_16_ ( .D(
        j202_soc_core_j22_cpu_ml_N319), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_16_ ( .D(n29833), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_mach[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_16_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[16]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_16_ ( .D(
        j202_soc_core_j22_cpu_ml_N354), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ml_N412), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_16_ ( .D(
        j202_soc_core_j22_cpu_rf_N314), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__16_ ( 
        .D(n29503), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[16]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_16_ ( 
        .D(j202_soc_core_qspi_wb_wdat[16]), .CLK(wb_clk_i), .RESET_B(n29830), 
        .Q(j202_soc_core_bldc_core_00_wdata[16]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_16_ ( 
        .D(n38), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_0_ ( .D(n37), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_uart_div1[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_16_ ( 
        .D(j202_soc_core_qspi_wb_wdat[16]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_N713), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_16_ ( 
        .D(j202_soc_core_wbqspiflash_00_N683), .DE(n29754), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[112]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[80]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[48]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_16_ ( .D(
        j202_soc_core_ahb2apb_01_N144), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[80]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_17_ ( .D(
        j202_soc_core_j22_cpu_ml_N320), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_17_ ( .D(n29832), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_mach[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_17_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[17]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_17_ ( .D(
        j202_soc_core_j22_cpu_ml_N355), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ml_N413), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_17_ ( .D(
        j202_soc_core_j22_cpu_rf_N315), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3365), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3329), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3290), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2698), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2735), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[50]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2772), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[82]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2809), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[114]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2846), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[146]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2883), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[178]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2920), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[210]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2957), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[242]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2994), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[274]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3031), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[306]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3068), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[337]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3105), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[369]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3142), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[401]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3179), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[433]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3216), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[465]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3253), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[497]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_18_ ( .D(n13104), 
        .DE(j202_soc_core_j22_cpu_rf_N2668), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3367), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3331), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3292), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2700), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2737), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[52]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2774), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[84]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2811), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[116]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2848), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[148]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2885), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[180]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2922), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[212]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2959), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[244]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2996), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[276]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3033), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[308]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3070), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[339]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3107), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[371]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3144), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[403]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3181), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[435]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3218), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[467]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3255), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[499]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_20_ ( .D(n13105), 
        .DE(j202_soc_core_j22_cpu_rf_N2668), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3366), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3330), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3291), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2699), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2736), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[51]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2773), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[83]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2810), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[115]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2847), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[147]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2884), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[179]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2921), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[211]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2958), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[243]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2995), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[275]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3032), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[307]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3069), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[338]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3106), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[370]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3143), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[402]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3180), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[434]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3217), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[466]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3254), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[498]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_19_ ( .D(n13100), 
        .DE(j202_soc_core_j22_cpu_rf_N2668), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_19_ ( .D(
        j202_soc_core_j22_cpu_ml_N357), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ml_N415), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_19_ ( .D(
        j202_soc_core_j22_cpu_rf_N317), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__19_ ( 
        .D(n29506), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[19]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_19_ ( 
        .D(j202_soc_core_qspi_wb_wdat[19]), .CLK(wb_clk_i), .RESET_B(n12069), 
        .Q(j202_soc_core_bldc_core_00_wdata[19]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_19_ ( 
        .D(n36), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_3_ ( .D(n35), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_uart_div1[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_19_ ( 
        .D(j202_soc_core_qspi_wb_wdat[19]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_N716), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_19_ ( 
        .D(j202_soc_core_wbqspiflash_00_N686), .DE(n29754), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[124]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[116]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[108]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[100]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[115]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[83]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[51]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_19_ ( .D(
        j202_soc_core_ahb2apb_01_N147), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[83]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_01_N129), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[65]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__17_ ( 
        .D(n29504), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[17]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_17_ ( 
        .D(j202_soc_core_qspi_wb_wdat[17]), .CLK(wb_clk_i), .RESET_B(n29827), 
        .Q(j202_soc_core_bldc_core_00_wdata[17]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_17_ ( 
        .D(n34), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_1_ ( .D(n33), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_uart_div1[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_17_ ( 
        .D(j202_soc_core_qspi_wb_wdat[17]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_N714), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_17_ ( 
        .D(j202_soc_core_wbqspiflash_00_N684), .DE(n29876), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[60]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[52]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[44]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[36]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[113]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[81]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[49]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_17_ ( .D(
        j202_soc_core_ahb2apb_01_N145), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[81]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_9_ ( .D(
        j202_soc_core_j22_cpu_rf_N307), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__25_ ( 
        .D(n29513), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_25_ ( 
        .D(j202_soc_core_qspi_wb_wdat[25]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[62]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[54]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[46]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[38]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[121]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[89]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[57]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_25_ ( .D(
        j202_soc_core_ahb2apb_01_N153), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[89]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__9_ ( .D(
        n29527), .DE(n30189), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_9_ ( 
        .D(j202_soc_core_qspi_wb_wdat[9]), .CLK(wb_clk_i), .RESET_B(n29827), 
        .Q(j202_soc_core_bldc_core_00_wdata[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_9_ ( 
        .D(n32), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_pwm_period[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld_reg ( 
        .D(n31), .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_9_ ( 
        .D(j202_soc_core_qspi_wb_wdat[9]), .CLK(wb_clk_i), .RESET_B(n29827), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_9_ ( 
        .D(n30), .CLK(wb_clk_i), .RESET_B(n29828), .Q(
        j202_soc_core_cmt_core_00_const1[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_9_ ( 
        .D(n29), .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_cmt_core_00_const0[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[9]), .CLK(wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_cmt_core_00_cnt0[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[9]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmf0_o_reg ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt0_to1), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmf0) );
  sky130_fd_sc_hd__dfstp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[0]), .CLK(wb_clk_i), .SET_B(n29827), .Q(j202_soc_core_cmt_core_00_cnt0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[0]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[0]), .CLK(wb_clk_i), 
        .RESET_B(n29745), .Q(j202_soc_core_prdata[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_00_N128), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[96]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[1]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cnt0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[1]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[1]), .CLK(wb_clk_i), 
        .RESET_B(n29830), .Q(j202_soc_core_prdata[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_00_N129), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[97]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[2]), .CLK(wb_clk_i), .RESET_B(n29828), .Q(j202_soc_core_cmt_core_00_cnt0[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[2]), .CLK(wb_clk_i), .RESET_B(n29828), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[2]), .CLK(wb_clk_i), 
        .RESET_B(n29828), .Q(j202_soc_core_prdata[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_2_ ( .D(
        j202_soc_core_ahb2apb_00_N130), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[98]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[3]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cnt0[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[3]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[3]), .CLK(wb_clk_i), 
        .RESET_B(n29827), .Q(j202_soc_core_prdata[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_3_ ( .D(
        j202_soc_core_ahb2apb_00_N131), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[99]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[4]), .CLK(wb_clk_i), .RESET_B(n12069), .Q(j202_soc_core_cmt_core_00_cnt0[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[4]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[4]), .CLK(wb_clk_i), 
        .RESET_B(n29830), .Q(j202_soc_core_prdata[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_4_ ( .D(
        j202_soc_core_ahb2apb_00_N132), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[100])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[5]), .CLK(wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_cmt_core_00_cnt0[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[5]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[6]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cnt0[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[6]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[7]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cnt0[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[7]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[8]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cnt0[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[8]), .CLK(wb_clk_i), .RESET_B(n29828), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[10]), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cnt0[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[10]), .CLK(wb_clk_i), .RESET_B(
        n29827), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[11]), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cnt0[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[11]), .CLK(wb_clk_i), .RESET_B(
        n29827), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[12]), .CLK(
        wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_cmt_core_00_cnt0[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[12]), .CLK(wb_clk_i), .RESET_B(
        n29827), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[12]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_prdata[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_12_ ( .D(
        j202_soc_core_ahb2apb_00_N140), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[108])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[13]), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cnt0[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[13]), .CLK(wb_clk_i), .RESET_B(
        n29827), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[14]), .CLK(
        wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_cmt_core_00_cnt0[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[14]), .CLK(wb_clk_i), .RESET_B(
        n29827), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[15]), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cnt0[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[15]), .CLK(wb_clk_i), .RESET_B(
        n29828), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_9_ ( 
        .D(j202_soc_core_qspi_wb_wdat[9]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_9_ ( .D(
        n10566), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[58]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[50]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[42]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[34]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[105]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[73]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[41]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_9_ ( .D(
        j202_soc_core_ahb2apb_01_N137), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[73]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_15_ ( .D(
        j202_soc_core_j22_cpu_ml_N427), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_32_ ( .D(
        j202_soc_core_j22_cpu_ml_N429), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[32]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_15_ ( .D(
        j202_soc_core_j22_cpu_rf_N313), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_15_ ( 
        .D(n29550), .DE(n30067), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_13_ ( 
        .D(j202_soc_core_qspi_wb_addr[15]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_15_ ( .D(
        n29550), .DE(n30030), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_13_ ( .D(
        j202_soc_core_j22_cpu_ml_N316), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_13_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[13]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_13_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[13]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_13_ ( .D(
        j202_soc_core_j22_cpu_rf_N311), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__29_ ( 
        .D(n29517), .DE(n30189), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[29]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_5_ ( .D(n28), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_uart_div0[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_clr_reg ( .D(
        j202_soc_core_uart_BRG_N21), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps_clr) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_0_ ( .D(
        j202_soc_core_uart_BRG_N12), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_1_ ( .D(
        j202_soc_core_uart_BRG_N13), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_2_ ( .D(
        j202_soc_core_uart_BRG_N14), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_3_ ( .D(
        j202_soc_core_uart_BRG_N15), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_4_ ( .D(
        j202_soc_core_uart_BRG_N16), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_5_ ( .D(
        j202_soc_core_uart_BRG_N17), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_6_ ( .D(
        j202_soc_core_uart_BRG_N18), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_7_ ( .D(
        j202_soc_core_uart_BRG_N19), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_1_ ( .D(
        j202_soc_core_uart_BRG_N36), .DE(n10716), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_br_clr_reg ( .D(
        j202_soc_core_uart_BRG_N47), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_clr) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_x4_r_reg ( .D(
        j202_soc_core_uart_BRG_br_clr), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_sio_ce_x4_r) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_0_ ( .D(
        j202_soc_core_uart_BRG_N35), .DE(n10716), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_2_ ( .D(
        j202_soc_core_uart_BRG_N37), .DE(n10716), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_3_ ( .D(
        j202_soc_core_uart_BRG_N38), .DE(n10716), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_4_ ( .D(
        j202_soc_core_uart_BRG_N39), .DE(n10716), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_5_ ( .D(
        j202_soc_core_uart_BRG_N40), .DE(n10716), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_6_ ( .D(
        j202_soc_core_uart_BRG_N41), .DE(n10716), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_7_ ( .D(
        j202_soc_core_uart_BRG_N42), .DE(n10716), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_x4_t_reg ( .D(n29601), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_BRG_sio_ce_x4_t) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_x4_reg ( .D(
        j202_soc_core_uart_BRG_sio_ce_x4_t), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_sio_ce_x4) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_change_reg ( .D(
        j202_soc_core_uart_TOP_N102), .DE(j202_soc_core_uart_TOP_N101), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_change) );
  sky130_fd_sc_hd__dfstp_1 j202_soc_core_uart_TOP_dpll_state_reg_0_ ( .D(n27), 
        .CLK(wb_clk_i), .SET_B(n29830), .Q(
        j202_soc_core_uart_TOP_dpll_state[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_sio_ce_r1_reg ( .D(n29607), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_sio_ce_r1) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_sio_ce_r2_reg ( .D(
        j202_soc_core_uart_TOP_rx_sio_ce_r1), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_sio_ce_r2) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_sio_ce_reg ( .D(
        j202_soc_core_uart_TOP_N118), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_sio_ce) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_9_ ( .D(
        j202_soc_core_uart_TOP_rxd_s), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_8_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_7_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_6_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_5_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_4_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_3_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_2_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_bit_cnt_reg_0_ ( .D(
        n29742), .DE(j202_soc_core_uart_TOP_N85), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_bit_cnt[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_bit_cnt_reg_1_ ( .D(
        j202_soc_core_uart_TOP_N87), .DE(j202_soc_core_uart_TOP_N85), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_bit_cnt[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_bit_cnt_reg_2_ ( .D(
        j202_soc_core_uart_TOP_N88), .DE(j202_soc_core_uart_TOP_N85), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_bit_cnt[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_bit_cnt_reg_3_ ( .D(
        j202_soc_core_uart_TOP_N89), .DE(j202_soc_core_uart_TOP_N85), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_bit_cnt[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_go_reg ( .D(
        j202_soc_core_uart_TOP_N128), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_go) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_valid_reg ( .D(n10949), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_valid) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_valid_r_reg ( .D(
        j202_soc_core_uart_TOP_rx_valid), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_valid_r) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_rx_fifo_wp_reg_0_ ( .D(n26), 
        .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_uart_TOP_rx_fifo_wp[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_rx_fifo_wp_reg_1_ ( .D(n25), 
        .CLK(wb_clk_i), .RESET_B(n29830), .Q(
        j202_soc_core_uart_TOP_rx_fifo_wp[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_gb_reg ( .D(
        j202_soc_core_uart_TOP_rx_fifo_N42), .DE(
        j202_soc_core_uart_TOP_rx_fifo_N41), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_gb) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__0_ ( .D(
        j202_soc_core_uart_TOP_rxr[2]), .DE(n29723), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__7_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(n29723), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__6_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(n29723), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__5_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(n29723), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__4_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(n29723), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__3_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(n29723), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__2_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(n29723), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__1_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(n29723), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__0_ ( .D(
        j202_soc_core_uart_TOP_rxr[2]), .DE(n29869), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__7_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(n29869), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__6_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(n29869), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__5_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(n29869), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__4_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(n29869), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__3_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(n29869), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__2_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(n29869), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__1_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(n29869), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__0_ ( .D(
        j202_soc_core_uart_TOP_rxr[2]), .DE(n29870), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__7_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(n29870), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__6_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(n29870), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__5_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(n29870), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__4_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(n29870), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__3_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(n29870), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__2_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(n29870), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__1_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(n29870), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__0_ ( .D(
        j202_soc_core_uart_TOP_rxr[2]), .DE(n29868), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__7_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(n29868), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__6_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(n29868), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__5_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(n29868), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__4_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(n29868), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__3_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(n29868), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__2_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(n29868), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__1_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(n29868), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[25]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_dpll_state_reg_1_ ( .D(n24), 
        .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_uart_TOP_dpll_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_cnt_reg_0_ ( .D(n29602), 
        .DE(j202_soc_core_uart_BRG_N55), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_cnt[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_cnt_reg_1_ ( .D(
        j202_soc_core_uart_BRG_N57), .DE(j202_soc_core_uart_BRG_N55), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_BRG_cnt[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_r_reg ( .D(n29609), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_BRG_sio_ce_r) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_reg ( .D(
        j202_soc_core_uart_BRG_N59), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_sio_ce) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_txf_empty_r_reg ( .D(
        j202_soc_core_uart_TOP_N16), .DE(n10717), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_txf_empty_r) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_load_reg ( .D(
        j202_soc_core_uart_TOP_N137), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_load) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_bit_cnt_reg_1_ ( .D(
        n29740), .DE(j202_soc_core_uart_TOP_N57), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_bit_cnt[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_bit_cnt_reg_3_ ( .D(
        j202_soc_core_uart_TOP_N61), .DE(j202_soc_core_uart_TOP_N57), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_bit_cnt[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_shift_en_reg ( .D(
        j202_soc_core_uart_TOP_N123), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_shift_en) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_shift_en_r_reg ( .D(n29494), 
        .DE(n10717), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_shift_en_r) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_bit_cnt_reg_0_ ( .D(
        j202_soc_core_uart_TOP_N58), .DE(j202_soc_core_uart_TOP_N57), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_bit_cnt[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_bit_cnt_reg_2_ ( .D(
        n29731), .DE(j202_soc_core_uart_TOP_N57), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_bit_cnt[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_tx_fifo_rp_reg_0_ ( .D(n23), 
        .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_uart_TOP_tx_fifo_rp[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_tx_fifo_rp_reg_1_ ( .D(n22), 
        .CLK(wb_clk_i), .RESET_B(n29827), .Q(
        j202_soc_core_uart_TOP_tx_fifo_rp[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_gb_reg ( .D(
        j202_soc_core_uart_TOP_tx_fifo_N42), .DE(
        j202_soc_core_uart_TOP_tx_fifo_N41), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_gb) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_8_ ( .D(
        j202_soc_core_uart_TOP_N33), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_7_ ( .D(
        j202_soc_core_uart_TOP_N32), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_6_ ( .D(
        j202_soc_core_uart_TOP_N31), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_5_ ( .D(
        j202_soc_core_uart_TOP_N30), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_4_ ( .D(
        j202_soc_core_uart_TOP_N29), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_3_ ( .D(
        j202_soc_core_uart_TOP_N28), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_2_ ( .D(
        j202_soc_core_uart_TOP_N27), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_1_ ( .D(
        j202_soc_core_uart_TOP_N26), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_0_ ( .D(
        j202_soc_core_uart_TOP_N25), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_txd_o_reg ( .D(
        j202_soc_core_uart_TOP_N43), .DE(n10717), .CLK(wb_clk_i), .Q(io_out[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_29_ ( 
        .D(j202_soc_core_qspi_wb_wdat[29]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[63]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[55]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[47]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[39]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[125]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[93]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[61]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_29_ ( .D(
        j202_soc_core_ahb2apb_01_N157), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[93]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_6_ ( .D(
        n29529), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_13_ ( .D(
        n29536), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[13])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_12_ ( .D(
        n29535), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[12])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_5_ ( .D(
        n29596), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_4_ ( .D(
        n29528), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_13_ ( 
        .D(n29474), .DE(n30067), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_11_ ( 
        .D(j202_soc_core_qspi_wb_addr[13]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_13_ ( .D(
        n29474), .DE(n10998), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_02_state_reg_0_ ( .D(
        j202_soc_core_ahb2apb_02_N89), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_02_state[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_02_state_reg_2_ ( .D(n29743), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2apb_02_state[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_02_state_reg_1_ ( .D(n29730), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2apb_02_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_2_ ( 
        .D(n29873), .DE(n10600), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_02_N23), .DE(n30052), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_hsize_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_02_N57), .DE(n30053), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_02_hsize_buf[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_hsize_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_02_N56), .DE(n30052), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_02_hsize_buf[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_hwrite_buf_reg ( .D(
        j202_soc_core_ahb2apb_02_N55), .DE(n30053), .CLK(wb_clk_i), .Q(
        j202_soc_core_pwrite[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_7_ ( .D(
        j202_soc_core_ahb2apb_02_N30), .DE(n30052), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_6_ ( .D(
        j202_soc_core_ahb2apb_02_N29), .DE(n30053), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_5_ ( .D(
        j202_soc_core_ahb2apb_02_N28), .DE(n30052), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_4_ ( .D(
        j202_soc_core_ahb2apb_02_N27), .DE(j202_soc_core_ahb2apb_02_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_reg_addr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_3_ ( .D(
        j202_soc_core_ahb2apb_02_N26), .DE(j202_soc_core_ahb2apb_02_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_reg_addr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_2_ ( .D(
        j202_soc_core_ahb2apb_02_N25), .DE(j202_soc_core_ahb2apb_02_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_reg_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_02_N24), .DE(j202_soc_core_ahb2apb_02_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_reg_addr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_31_ ( 
        .D(n29569), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_30_ ( 
        .D(n29449), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_29_ ( 
        .D(n29450), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_28_ ( 
        .D(n29568), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_27_ ( 
        .D(n29451), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_26_ ( 
        .D(n29452), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_25_ ( 
        .D(n29453), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_24_ ( 
        .D(n29454), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_23_ ( 
        .D(n29455), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_22_ ( 
        .D(n29456), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_21_ ( 
        .D(n29457), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_20_ ( 
        .D(n29458), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_19_ ( 
        .D(n29459), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_18_ ( 
        .D(n29460), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_17_ ( 
        .D(n29461), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_16_ ( 
        .D(n29462), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_15_ ( 
        .D(n29446), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_11_ ( 
        .D(n29447), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_10_ ( 
        .D(n29448), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_9_ ( 
        .D(n29463), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_8_ ( 
        .D(n29464), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_7_ ( 
        .D(n29465), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_6_ ( 
        .D(n29466), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_5_ ( 
        .D(n29467), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_4_ ( 
        .D(n29468), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_3_ ( 
        .D(n29469), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_2_ ( 
        .D(n29470), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_1_ ( 
        .D(n29471), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_0_ ( 
        .D(n29472), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_31_ ( 
        .D(n29569), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_30_ ( 
        .D(n29449), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_29_ ( 
        .D(n29450), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_28_ ( 
        .D(n29568), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_27_ ( 
        .D(n29451), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_26_ ( 
        .D(n29452), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_25_ ( 
        .D(n29453), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_24_ ( 
        .D(n29454), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_23_ ( 
        .D(n29455), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_22_ ( 
        .D(n29456), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_21_ ( 
        .D(n29457), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_20_ ( 
        .D(n29458), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_19_ ( 
        .D(n29459), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_18_ ( 
        .D(n29460), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_17_ ( 
        .D(n29461), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_16_ ( 
        .D(n29462), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_15_ ( 
        .D(n29446), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_11_ ( 
        .D(n29447), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_10_ ( 
        .D(n29448), .DE(n29824), .CLK(wb_clk_i), .Q(la_data_out[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_9_ ( 
        .D(n29463), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_8_ ( 
        .D(n29464), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_7_ ( 
        .D(n29465), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_6_ ( 
        .D(n29466), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_5_ ( 
        .D(n29467), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_4_ ( 
        .D(n29468), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_3_ ( 
        .D(n29469), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_2_ ( 
        .D(n29470), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_1_ ( 
        .D(n29471), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_0_ ( 
        .D(n29472), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_31_ ( 
        .D(n29569), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_30_ ( 
        .D(n29449), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_29_ ( 
        .D(n29450), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_28_ ( 
        .D(n29568), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_27_ ( 
        .D(n29451), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_26_ ( 
        .D(n29452), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_25_ ( 
        .D(n29453), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_24_ ( 
        .D(n29454), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_23_ ( 
        .D(n29455), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_22_ ( 
        .D(n29456), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_21_ ( 
        .D(n29457), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_20_ ( 
        .D(n29458), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_19_ ( 
        .D(n29459), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_18_ ( 
        .D(n29460), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_17_ ( 
        .D(n29461), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_16_ ( 
        .D(n29462), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_15_ ( 
        .D(n29446), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_11_ ( 
        .D(n29447), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_10_ ( 
        .D(n29448), .DE(n29825), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_9_ ( 
        .D(n29463), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_8_ ( 
        .D(n29464), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_7_ ( 
        .D(n29465), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_6_ ( 
        .D(n29466), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_5_ ( 
        .D(n29467), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_4_ ( 
        .D(n29468), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_3_ ( 
        .D(n29469), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_2_ ( 
        .D(n29470), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_1_ ( 
        .D(n29471), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_0_ ( 
        .D(n29472), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_10_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N50), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_15_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N55), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_31_ ( 
        .D(n29569), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_31_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N71), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_31_ ( .D(
        j202_soc_core_ahb2apb_02_N159), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[63]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_30_ ( 
        .D(n29449), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_30_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N70), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_30_ ( .D(
        j202_soc_core_ahb2apb_02_N158), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[62]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_29_ ( 
        .D(n29450), .DE(n10711), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_29_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N69), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_29_ ( .D(
        j202_soc_core_ahb2apb_02_N157), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[61]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_28_ ( 
        .D(n29568), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_28_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N68), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_28_ ( .D(
        j202_soc_core_ahb2apb_02_N156), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[60]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_27_ ( 
        .D(n29451), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_27_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N67), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_27_ ( .D(
        j202_soc_core_ahb2apb_02_N155), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[59]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_26_ ( 
        .D(n29452), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_26_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N66), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_26_ ( .D(
        j202_soc_core_ahb2apb_02_N154), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[58]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_25_ ( 
        .D(n29453), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_25_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N65), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_25_ ( .D(
        j202_soc_core_ahb2apb_02_N153), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[57]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_24_ ( 
        .D(n29454), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_24_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N64), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_24_ ( .D(
        j202_soc_core_ahb2apb_02_N152), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[56]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_23_ ( 
        .D(n29455), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_23_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N63), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_23_ ( .D(
        j202_soc_core_ahb2apb_02_N151), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[55]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_22_ ( 
        .D(n29456), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_22_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N62), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_22_ ( .D(
        j202_soc_core_ahb2apb_02_N150), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[54]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_21_ ( 
        .D(n29457), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_21_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N61), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_21_ ( .D(
        j202_soc_core_ahb2apb_02_N149), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[53]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_20_ ( 
        .D(n29458), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_20_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N60), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_20_ ( .D(
        j202_soc_core_ahb2apb_02_N148), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[52]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_19_ ( 
        .D(n29459), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_19_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N59), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_19_ ( .D(
        j202_soc_core_ahb2apb_02_N147), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[51]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_18_ ( 
        .D(n29460), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_18_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N58), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_18_ ( .D(
        j202_soc_core_ahb2apb_02_N146), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[50]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_17_ ( 
        .D(n29461), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_17_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N57), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_17_ ( .D(
        j202_soc_core_ahb2apb_02_N145), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[49]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_16_ ( 
        .D(n29462), .DE(n29826), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_16_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N56), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_16_ ( .D(
        j202_soc_core_ahb2apb_02_N144), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[48]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_9_ ( 
        .D(n29463), .DE(n10711), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_9_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N49), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_9_ ( .D(
        j202_soc_core_ahb2apb_02_N137), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[41]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_8_ ( 
        .D(n29464), .DE(n10711), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_8_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N48), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_8_ ( .D(
        j202_soc_core_ahb2apb_02_N136), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[40]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_7_ ( 
        .D(n29465), .DE(n10711), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_7_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N47), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_7_ ( .D(
        j202_soc_core_ahb2apb_02_N135), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[39]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_6_ ( 
        .D(n29466), .DE(n10711), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_6_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N46), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_6_ ( .D(
        j202_soc_core_ahb2apb_02_N134), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[38]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_5_ ( 
        .D(n29467), .DE(n10711), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_5_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N45), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_5_ ( .D(
        j202_soc_core_ahb2apb_02_N133), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[37]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_4_ ( 
        .D(n29468), .DE(n10711), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_4_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N44), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_4_ ( .D(
        j202_soc_core_ahb2apb_02_N132), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[36]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_3_ ( 
        .D(n29469), .DE(n10711), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_3_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N43), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_3_ ( .D(
        j202_soc_core_ahb2apb_02_N131), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[35]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_2_ ( 
        .D(n29470), .DE(n10711), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_2_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N42), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_2_ ( .D(
        j202_soc_core_ahb2apb_02_N130), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[34]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_1_ ( 
        .D(n29471), .DE(n10711), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_1_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N41), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_02_N129), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[33]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_0_ ( 
        .D(n29472), .DE(n10711), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N40), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_02_N128), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[32]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_11_ ( .D(
        n29538), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[11])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_10_ ( .D(
        n29591), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[10])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_3_ ( .D(
        n29531), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_2_ ( .D(
        n29592), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_9_ ( .D(
        n29600), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_8_ ( .D(
        n29539), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_1_ ( .D(
        n29533), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_29_ ( .D(
        j202_soc_core_j22_cpu_ml_N368), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_13_ ( .D(
        j202_soc_core_j22_cpu_ml_N425), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_6_ ( .D(
        j202_soc_core_j22_cpu_ml_N418), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3351), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2721), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[38]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2758), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[70]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2795), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[102]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2832), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[134]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2869), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[166]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2906), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[198]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2943), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[230]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2980), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[262]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3017), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[294]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3054), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[325]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3091), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[357]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3128), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[389]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3165), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[421]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3202), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[453]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_21_ ( .D(
        j202_soc_core_j22_cpu_ml_N360), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_21_ ( .D(
        j202_soc_core_j22_cpu_ml_N325), .DE(n29750), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_21_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[21]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3368), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3333), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3294), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2702), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2739), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[53]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2776), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[85]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2813), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[117]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2850), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[149]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2887), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[181]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2924), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[213]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2961), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[245]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2998), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[277]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3035), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[309]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3072), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[340]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3109), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[372]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3146), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[404]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3183), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[436]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3220), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[468]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3257), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[500]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_21_ ( .D(n12130), 
        .DE(j202_soc_core_j22_cpu_rf_N2668), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_21_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[21]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3350), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2720), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[37]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2757), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[69]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2794), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[101]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2831), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[133]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2868), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[165]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2905), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[197]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2942), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[229]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2979), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[261]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3016), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[293]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3053), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[324]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3090), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[356]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3127), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[388]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3164), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[420]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3201), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[452]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_5_ ( .D(
        j202_soc_core_j22_cpu_rf_N303), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3315), .DE(n13071), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3275), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2683), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3238), .DE(n29749), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[484]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_5_ ( .D(
        j202_soc_core_j22_cpu_ml_N417), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[6]), .CLK(wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_cmt_core_00_cnt1[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[6]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[6]), .CLK(wb_clk_i), 
        .RESET_B(n29830), .Q(j202_soc_core_prdata[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_6_ ( .D(
        j202_soc_core_ahb2apb_00_N134), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[102])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[7]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cnt1[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[7]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[8]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cnt1[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[8]), .CLK(wb_clk_i), .RESET_B(n29828), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[8]), .CLK(wb_clk_i), 
        .RESET_B(n29830), .Q(j202_soc_core_prdata[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_8_ ( .D(
        j202_soc_core_ahb2apb_00_N136), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[104])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[9]), .CLK(wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cnt1[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[9]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[9]), .CLK(wb_clk_i), 
        .RESET_B(n29830), .Q(j202_soc_core_prdata[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_9_ ( .D(
        j202_soc_core_ahb2apb_00_N137), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[105])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[10]), .CLK(
        wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_cmt_core_00_cnt1[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[10]), .CLK(wb_clk_i), .RESET_B(
        n29827), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[10]), .CLK(wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_prdata[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_10_ ( .D(
        j202_soc_core_ahb2apb_00_N138), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[106])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[11]), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cnt1[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[11]), .CLK(wb_clk_i), .RESET_B(
        n29827), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[11]), .CLK(wb_clk_i), .RESET_B(n29827), .Q(j202_soc_core_prdata[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_11_ ( .D(
        j202_soc_core_ahb2apb_00_N139), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[107])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[13]), .CLK(
        wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_cmt_core_00_cnt1[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[13]), .CLK(wb_clk_i), .RESET_B(
        n29827), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[13]), .CLK(wb_clk_i), .RESET_B(n29828), .Q(j202_soc_core_prdata[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_13_ ( .D(
        j202_soc_core_ahb2apb_00_N141), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[109])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[14]), .CLK(
        wb_clk_i), .RESET_B(n29830), .Q(j202_soc_core_cmt_core_00_cnt1[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[14]), .CLK(wb_clk_i), .RESET_B(
        n29745), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[14]), .CLK(wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_prdata[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_14_ ( .D(
        j202_soc_core_ahb2apb_00_N142), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[110])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[15]), .CLK(
        wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_cmt_core_00_cnt1[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[15]), .CLK(wb_clk_i), .RESET_B(
        n29827), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[15]), .CLK(wb_clk_i), .RESET_B(n29745), .Q(j202_soc_core_prdata[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_15_ ( .D(
        j202_soc_core_ahb2apb_00_N143), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[111])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_12_ ( 
        .D(j202_soc_core_qspi_wb_wdat[12]), .DE(n29752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_12_ ( 
        .D(n29475), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_12_ ( 
        .D(n29475), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_12_ ( 
        .D(n29475), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_12_ ( 
        .D(n29475), .DE(n10711), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_12_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N52), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_12_ ( .D(
        j202_soc_core_ahb2apb_02_N140), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[44]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[108]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[76]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[44]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_12_ ( .D(
        j202_soc_core_ahb2apb_01_N140), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[76]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_N670), .DE(n29876), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_N669), .DE(n29754), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_N668), .DE(n29876), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_24_ ( .D(
        n10551), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_25_ ( .D(
        n10550), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_26_ ( .D(
        n10549), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_22_ ( 
        .D(n12291), .DE(n13109), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_20_ ( 
        .D(j202_soc_core_qspi_wb_addr[22]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_8_ ( .D(
        j202_soc_core_ahb2apb_01_N136), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[72]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_23_ ( .D(
        j202_soc_core_j22_cpu_ml_N362), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_7_ ( .D(
        j202_soc_core_j22_cpu_ml_N419), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_23_ ( 
        .D(n12299), .DE(n13109), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_21_ ( 
        .D(j202_soc_core_qspi_wb_addr[23]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_27_ ( .D(
        j202_soc_core_j22_cpu_ml_N366), .DE(n29650), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_11_ ( .D(
        j202_soc_core_j22_cpu_ml_N423), .DE(j202_soc_core_j22_cpu_ml_N428), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_13_ ( .D(
        j202_soc_core_ahb2apb_01_N141), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[77]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_13_ ( 
        .D(n29477), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_13_ ( 
        .D(n29477), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_13_ ( 
        .D(n29477), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_13_ ( 
        .D(n29477), .DE(n10711), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_13_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N53), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_13_ ( .D(
        j202_soc_core_ahb2apb_02_N141), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[45]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_14_ ( .D(
        j202_soc_core_ahb2apb_01_N142), .DE(n29751), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[78]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_14_ ( 
        .D(n29478), .DE(n10714), .CLK(wb_clk_i), .Q(la_data_out[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_14_ ( 
        .D(n29478), .DE(n12082), .CLK(wb_clk_i), .Q(gpio_en_o[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_14_ ( 
        .D(n29478), .DE(n10712), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_14_ ( 
        .D(n29478), .DE(n10711), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_14_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N54), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_14_ ( .D(
        j202_soc_core_ahb2apb_02_N142), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[46]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__i__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3392), .DE(j202_soc_core_j22_cpu_rf_N3391), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__i__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_7_ ( .D(
        j202_soc_core_j22_cpu_rf_N305), .DE(n29748), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_11_ ( .D(
        j202_soc_core_ahb2apb_02_N139), .DE(j202_soc_core_ahb2apb_02_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[43]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_19_ ( 
        .D(n29479), .DE(n13109), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_17_ ( 
        .D(j202_soc_core_qspi_wb_addr[19]), .DE(n29630), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_29_ ( .D(
        n10546), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[29]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_nxt_latch_status_0_), 
        .CLK(wb_clk_i), .RESET_B(n29745), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[7]), .CLK(wb_clk_i), 
        .RESET_B(n29830), .Q(j202_soc_core_prdata[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_7_ ( .D(
        j202_soc_core_ahb2apb_00_N135), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[103])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N425), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N426), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N427), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N430), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N428), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N391), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N392), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N393), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N394), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N395), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_10_ ( .D(
        n10565), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_11_ ( .D(
        n10564), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_22_ ( .D(
        n10553), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_23_ ( .D(
        n10552), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_28_ ( .D(
        n10547), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_5_ ( .D(
        n10570), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N396), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N397), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_7_ ( .D(
        n10568), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N398), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_8_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N399), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_9_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N400), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_10_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N401), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_11_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N402), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_12_ ( .D(
        n10563), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_12_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N403), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_13_ ( .D(
        n10562), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_13_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N404), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_14_ ( .D(
        n10561), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_14_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N405), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_15_ ( .D(
        n10560), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_15_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N406), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_16_ ( .D(
        n10559), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_16_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N407), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_17_ ( .D(
        n10558), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_17_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N408), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_18_ ( .D(
        n10557), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_18_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N409), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_19_ ( .D(
        n10556), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_19_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N410), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_20_ ( .D(
        n10555), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_20_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N411), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_21_ ( .D(
        n10554), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_21_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N412), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_22_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N413), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_23_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N414), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_24_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N415), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_25_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N416), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_26_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N417), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_27_ ( .D(
        n10548), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_27_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N418), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_28_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N419), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_29_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N420), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_dat_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N317), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N315), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_30_ ( .D(
        n10545), .DE(n29877), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_30_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N421), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_31_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N422), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N390), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_dat_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N316), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N315), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_dat_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N319), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N315), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_dat_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N318), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N315), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[2]) );
  sky130_fd_sc_hd__fa_1 DP_OP_1508J1_126_2326_U6 ( .A(n29648), .B(
        DP_OP_1508J1_126_2326_n6), .CIN(DP_OP_1508J1_126_2326_n4), .COUT(
        DP_OP_1508J1_126_2326_n3), .SUM(U7_RSOP_1495_C3_DATA3_2) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_15_ ( .D(
        n29534), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[15])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_14_ ( .D(
        n29537), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[14])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[17]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_01_pstrb_o_reg_1_ ( .GATE(
        j202_soc_core_ahb2apb_01_N123), .D(n10784), .RESET_B(
        j202_soc_core_pwrite[1]), .Q(j202_soc_core_pstrb[5]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_02_pstrb_o_reg_1_ ( .GATE(
        j202_soc_core_ahb2apb_02_N123), .D(n10943), .RESET_B(
        j202_soc_core_pwrite[2]), .Q(j202_soc_core_pstrb[1]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_01_pstrb_o_reg_3_ ( .GATE(
        j202_soc_core_ahb2apb_01_N123), .D(n10786), .RESET_B(
        j202_soc_core_pwrite[1]), .Q(j202_soc_core_pstrb[7]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_02_pstrb_o_reg_2_ ( .GATE(
        j202_soc_core_ahb2apb_02_N123), .D(n10944), .RESET_B(
        j202_soc_core_pwrite[2]), .Q(j202_soc_core_pstrb[2]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_01_pstrb_o_reg_2_ ( .GATE(
        j202_soc_core_ahb2apb_01_N123), .D(n10785), .RESET_B(
        j202_soc_core_pwrite[1]), .Q(j202_soc_core_pstrb[6]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_02_pstrb_o_reg_3_ ( .GATE(
        j202_soc_core_ahb2apb_02_N123), .D(n10945), .RESET_B(
        j202_soc_core_pwrite[2]), .Q(j202_soc_core_pstrb[3]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_01_pstrb_o_reg_0_ ( .GATE(
        j202_soc_core_ahb2apb_01_N123), .D(n10783), .RESET_B(
        j202_soc_core_pwrite[1]), .Q(j202_soc_core_pstrb[4]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_02_pstrb_o_reg_0_ ( .GATE(
        j202_soc_core_ahb2apb_02_N123), .D(n10942), .RESET_B(
        j202_soc_core_pwrite[2]), .Q(j202_soc_core_pstrb[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_nega_o_reg ( 
        .D(n29849), .CLK(wb_clk_i), .RESET_B(n29830), .Q(io_out[17]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_posc_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posc), .CLK(wb_clk_i), .RESET_B(n29827), .Q(io_out[20]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_negb_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_negb), .CLK(wb_clk_i), .RESET_B(n29828), .Q(io_out[19]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_negc_o_reg ( 
        .D(n29608), .CLK(wb_clk_i), .RESET_B(n29827), .Q(io_out[21]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_posb_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posb), .CLK(wb_clk_i), .RESET_B(n29745), .Q(io_out[18]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_posa_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posa), .CLK(wb_clk_i), .RESET_B(n29830), .Q(io_out[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_wbqspiflash_00_spif_override_reg ( 
        .D(j202_soc_core_wbqspiflash_00_N742), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_override) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_4_ ( 
        .D(n29497), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__4_) );
  sky130_fd_sc_hd__dfxtp_2 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__0_ ( .D(
        j202_soc_core_j22_cpu_ml_N152), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[0]) );
  sky130_fd_sc_hd__dfxtp_2 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[8]) );
  sky130_fd_sc_hd__dfxtp_2 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[21]) );
  sky130_fd_sc_hd__dfxtp_2 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__1_ ( .D(
        j202_soc_core_j22_cpu_ml_N153), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_We__1_ ( 
        .D(n10641), .DE(n10645), .CLK(wb_clk_i), .Q(n12347), .Q_N(n12348) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3043), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(n12245), .Q_N() );
  sky130_fd_sc_hd__dfxtp_2 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__4_ ( .D(
        j202_soc_core_j22_cpu_ml_N156), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[4]) );
  sky130_fd_sc_hd__dfxtp_4 j202_soc_core_rst_reg ( .D(j202_soc_core_rst1), 
        .CLK(wb_clk_i), .Q(j202_soc_core_rst) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[32]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[53]) );
  sky130_fd_sc_hd__dfxtp_2 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__3_ ( .D(
        j202_soc_core_j22_cpu_ml_N155), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_00_state_reg_1_ ( .D(n29744), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2apb_00_state[1]) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rb__0_ ( 
        .D(n10619), .DE(n10609), .CLK(wb_clk_i), .Q(n12054), .Q_N() );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_rf_vbr_reg_12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3323), .DE(n13071), .CLK(wb_clk_i), .Q(
        n12042), .Q_N(n11095) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_MEM__2_ ( 
        .D(n10630), .DE(n10601), .CLK(wb_clk_i), .Q(n12040), .Q_N(n12041) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rn__0_ ( 
        .D(n10612), .DE(n13090), .CLK(wb_clk_i), .Q(n12036) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rn__3_ ( 
        .D(n10615), .DE(n13090), .CLK(wb_clk_i), .Q(n12034) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rn__2_ ( 
        .D(n10614), .DE(n30087), .CLK(wb_clk_i), .Q(n12032) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rn__1_ ( 
        .D(n10613), .DE(n30087), .CLK(wb_clk_i), .Q(n12030) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[45]) );
  sky130_fd_sc_hd__dfxtp_2 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__2_ ( .D(
        j202_soc_core_j22_cpu_ml_N154), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]) );
  sky130_fd_sc_hd__and2_1 U13325 ( .A(n27087), .B(n27856), .X(n13098) );
  sky130_fd_sc_hd__and2_1 U13326 ( .A(n10966), .B(n24178), .X(n29645) );
  sky130_fd_sc_hd__a21oi_2 U13328 ( .A1(n28442), .A2(n24291), .B1(n24290), .Y(
        n24292) );
  sky130_fd_sc_hd__inv_2 U13329 ( .A(n12260), .Y(n27586) );
  sky130_fd_sc_hd__inv_6 U13330 ( .A(n11083), .Y(n11084) );
  sky130_fd_sc_hd__inv_6 U13331 ( .A(n12375), .Y(n11134) );
  sky130_fd_sc_hd__o21a_1 U13332 ( .A1(n10957), .A2(n27990), .B1(n25147), .X(
        n25150) );
  sky130_fd_sc_hd__inv_2 U13334 ( .A(n23982), .Y(n11081) );
  sky130_fd_sc_hd__and2b_2 U13335 ( .B(n29548), .A_N(n25024), .X(n23980) );
  sky130_fd_sc_hd__and2_1 U13336 ( .A(n24790), .B(n24789), .X(n13054) );
  sky130_fd_sc_hd__inv_4 U13337 ( .A(n29823), .Y(n12375) );
  sky130_fd_sc_hd__nand2_1 U13338 ( .A(n25857), .B(n25861), .Y(n25856) );
  sky130_fd_sc_hd__inv_2 U13339 ( .A(n23977), .Y(n29821) );
  sky130_fd_sc_hd__inv_2 U13340 ( .A(n29823), .Y(n12374) );
  sky130_fd_sc_hd__nand2_1 U13341 ( .A(n23769), .B(n23768), .Y(n25989) );
  sky130_fd_sc_hd__nand2_1 U13342 ( .A(n23780), .B(n23779), .Y(n25985) );
  sky130_fd_sc_hd__nand2_1 U13343 ( .A(n23791), .B(n23790), .Y(n25979) );
  sky130_fd_sc_hd__nand2_1 U13344 ( .A(n23796), .B(n23795), .Y(n26894) );
  sky130_fd_sc_hd__nand2_1 U13345 ( .A(n23822), .B(n23821), .Y(n25987) );
  sky130_fd_sc_hd__nand2_1 U13346 ( .A(n23774), .B(n23773), .Y(n25984) );
  sky130_fd_sc_hd__nand2_1 U13347 ( .A(n23812), .B(n23811), .Y(n25988) );
  sky130_fd_sc_hd__nand2_1 U13348 ( .A(n11672), .B(n24424), .Y(n24699) );
  sky130_fd_sc_hd__nand2_1 U13349 ( .A(n28109), .B(n23501), .Y(n27847) );
  sky130_fd_sc_hd__nand2_1 U13351 ( .A(n25769), .B(n23563), .Y(n27119) );
  sky130_fd_sc_hd__inv_2 U13352 ( .A(n11181), .Y(n26896) );
  sky130_fd_sc_hd__clkbuf_1 U13353 ( .A(n29745), .X(n12069) );
  sky130_fd_sc_hd__nand2_1 U13355 ( .A(n22187), .B(n22186), .Y(n25626) );
  sky130_fd_sc_hd__nand2b_1 U13356 ( .A_N(n24592), .B(n10981), .Y(n24596) );
  sky130_fd_sc_hd__a22oi_1 U13359 ( .A1(j202_soc_core_j22_cpu_ml_mach[22]), 
        .A2(n23041), .B1(n22185), .B2(n24452), .Y(n22186) );
  sky130_fd_sc_hd__clkbuf_1 U13360 ( .A(n11006), .X(n28267) );
  sky130_fd_sc_hd__clkbuf_1 U13362 ( .A(n27991), .X(n11444) );
  sky130_fd_sc_hd__and4_1 U13364 ( .A(n23477), .B(n23476), .C(n23479), .D(
        n23478), .X(n23468) );
  sky130_fd_sc_hd__and2_0 U13366 ( .A(n28384), .B(n29746), .X(n13074) );
  sky130_fd_sc_hd__clkbuf_1 U13367 ( .A(n23508), .X(n26169) );
  sky130_fd_sc_hd__nand2_1 U13368 ( .A(n23346), .B(n23345), .Y(n24376) );
  sky130_fd_sc_hd__nor2_1 U13369 ( .A(n24563), .B(n12778), .Y(n23394) );
  sky130_fd_sc_hd__nand2_1 U13370 ( .A(n12229), .B(n12622), .Y(n23597) );
  sky130_fd_sc_hd__nand3_1 U13371 ( .A(n17087), .B(n14590), .C(n17085), .Y(
        n29436) );
  sky130_fd_sc_hd__inv_2 U13373 ( .A(n26916), .Y(n11123) );
  sky130_fd_sc_hd__o22a_1 U13374 ( .A1(n21934), .A2(n12862), .B1(n11149), .B2(
        n24068), .X(n11851) );
  sky130_fd_sc_hd__nand2_1 U13376 ( .A(n11852), .B(n11205), .Y(n11850) );
  sky130_fd_sc_hd__o22a_1 U13378 ( .A1(n24931), .A2(n26936), .B1(n28532), .B2(
        n26932), .X(n21721) );
  sky130_fd_sc_hd__clkbuf_1 U13379 ( .A(n22002), .X(n29490) );
  sky130_fd_sc_hd__nand2_1 U13380 ( .A(n17093), .B(io_in[14]), .Y(n17094) );
  sky130_fd_sc_hd__buf_2 U13381 ( .A(n28914), .X(n29745) );
  sky130_fd_sc_hd__o21a_1 U13382 ( .A1(n26166), .A2(n17053), .B1(n17052), .X(
        n17095) );
  sky130_fd_sc_hd__nand3_1 U13388 ( .A(n16739), .B(n20454), .C(n21917), .Y(
        n12875) );
  sky130_fd_sc_hd__o21ai_1 U13391 ( .A1(n22071), .A2(n22335), .B1(n22070), .Y(
        n22543) );
  sky130_fd_sc_hd__nand3_1 U13393 ( .A(n12742), .B(n17218), .C(n21919), .Y(
        n12630) );
  sky130_fd_sc_hd__o21ai_1 U13394 ( .A1(n16558), .A2(n16557), .B1(n16556), .Y(
        n25806) );
  sky130_fd_sc_hd__nor2_1 U13395 ( .A(n13007), .B(n13002), .Y(n13001) );
  sky130_fd_sc_hd__nor2_1 U13396 ( .A(n19066), .B(n19065), .Y(n22915) );
  sky130_fd_sc_hd__inv_2 U13397 ( .A(n21925), .Y(n11186) );
  sky130_fd_sc_hd__nor2_1 U13398 ( .A(n18833), .B(n18832), .Y(n28056) );
  sky130_fd_sc_hd__fa_2 U13400 ( .A(n19008), .B(n19007), .CIN(n19006), .COUT(
        n19028), .SUM(n19016) );
  sky130_fd_sc_hd__fa_1 U13401 ( .A(n18949), .B(n18948), .CIN(n18947), .COUT(
        n19054), .SUM(n19046) );
  sky130_fd_sc_hd__fa_1 U13402 ( .A(n17363), .B(n17362), .CIN(n17361), .COUT(
        n17385), .SUM(n17422) );
  sky130_fd_sc_hd__fa_2 U13403 ( .A(n18067), .B(n18066), .CIN(n18065), .COUT(
        n18303), .SUM(n18093) );
  sky130_fd_sc_hd__fa_1 U13405 ( .A(n17568), .B(n17567), .CIN(n17566), .COUT(
        n17589), .SUM(n17571) );
  sky130_fd_sc_hd__nand3_1 U13406 ( .A(n12119), .B(n15920), .C(n15919), .Y(
        n27809) );
  sky130_fd_sc_hd__fa_1 U13407 ( .A(n17963), .B(n17962), .CIN(n17961), .COUT(
        n17952), .SUM(n18057) );
  sky130_fd_sc_hd__o22ai_1 U13409 ( .A1(n18989), .A2(n18987), .B1(n18967), 
        .B2(n18986), .Y(n19027) );
  sky130_fd_sc_hd__fa_2 U13410 ( .A(n18049), .B(n18048), .CIN(n18047), .COUT(
        n18073), .SUM(n18269) );
  sky130_fd_sc_hd__fa_1 U13411 ( .A(n17645), .B(n17644), .CIN(n17643), .COUT(
        n18568), .SUM(n17670) );
  sky130_fd_sc_hd__fa_2 U13412 ( .A(n17792), .B(n17791), .CIN(n17790), .COUT(
        n17775), .SUM(n17911) );
  sky130_fd_sc_hd__a21oi_1 U13413 ( .A1(n18889), .A2(n16523), .B1(n14570), .Y(
        n26311) );
  sky130_fd_sc_hd__nand3_1 U13414 ( .A(n15066), .B(n15065), .C(n13096), .Y(
        n28499) );
  sky130_fd_sc_hd__nand3_1 U13416 ( .A(n14455), .B(n14454), .C(n12105), .Y(
        n27111) );
  sky130_fd_sc_hd__and2_2 U13417 ( .A(n23493), .B(
        j202_soc_core_j22_cpu_ml_macl[31]), .X(n13087) );
  sky130_fd_sc_hd__nand2_1 U13418 ( .A(n17340), .B(n18989), .Y(n18986) );
  sky130_fd_sc_hd__buf_2 U13419 ( .A(n11967), .X(n11455) );
  sky130_fd_sc_hd__and2_4 U13420 ( .A(n13478), .B(n13513), .X(n13053) );
  sky130_fd_sc_hd__inv_4 U13421 ( .A(n12224), .Y(n11967) );
  sky130_fd_sc_hd__inv_2 U13422 ( .A(n13957), .Y(n11124) );
  sky130_fd_sc_hd__or2_1 U13423 ( .A(n13294), .B(n23788), .X(n12086) );
  sky130_fd_sc_hd__buf_4 U13424 ( .A(j202_soc_core_j22_cpu_ml_bufa[27]), .X(
        n23571) );
  sky130_fd_sc_hd__buf_4 U13425 ( .A(j202_soc_core_j22_cpu_ml_bufa[23]), .X(
        n22087) );
  sky130_fd_sc_hd__nand2_2 U13427 ( .A(n17450), .B(n30022), .Y(n18189) );
  sky130_fd_sc_hd__nand2_1 U13428 ( .A(n13436), .B(n13429), .Y(n16491) );
  sky130_fd_sc_hd__nand2_1 U13429 ( .A(n13179), .B(n20464), .Y(n15685) );
  sky130_fd_sc_hd__buf_2 U13430 ( .A(j202_soc_core_j22_cpu_ml_bufb[14]), .X(
        n18966) );
  sky130_fd_sc_hd__buf_2 U13431 ( .A(j202_soc_core_j22_cpu_ml_bufb[11]), .X(
        n18941) );
  sky130_fd_sc_hd__buf_2 U13432 ( .A(j202_soc_core_j22_cpu_ml_bufb[9]), .X(
        n18999) );
  sky130_fd_sc_hd__buf_2 U13433 ( .A(j202_soc_core_j22_cpu_ml_bufb[32]), .X(
        n22024) );
  sky130_fd_sc_hd__buf_2 U13434 ( .A(j202_soc_core_j22_cpu_ml_bufb[12]), .X(
        n18971) );
  sky130_fd_sc_hd__buf_4 U13435 ( .A(j202_soc_core_j22_cpu_ml_bufa[31]), .X(
        n25777) );
  sky130_fd_sc_hd__buf_2 U13436 ( .A(j202_soc_core_j22_cpu_ml_bufb[8]), .X(
        n18964) );
  sky130_fd_sc_hd__buf_2 U13437 ( .A(j202_soc_core_j22_cpu_ml_bufb[4]), .X(
        n18377) );
  sky130_fd_sc_hd__buf_2 U13438 ( .A(j202_soc_core_j22_cpu_ml_bufb[5]), .X(
        n18387) );
  sky130_fd_sc_hd__buf_2 U13439 ( .A(j202_soc_core_j22_cpu_ml_bufb[7]), .X(
        n18366) );
  sky130_fd_sc_hd__buf_2 U13440 ( .A(j202_soc_core_j22_cpu_ml_bufb[3]), .X(
        n18371) );
  sky130_fd_sc_hd__buf_2 U13441 ( .A(j202_soc_core_j22_cpu_ml_bufb[6]), .X(
        n18367) );
  sky130_fd_sc_hd__clkbuf_1 U13443 ( .A(j202_soc_core_bootrom_00_address_w[10]), .X(n18764) );
  sky130_fd_sc_hd__buf_4 U13444 ( .A(j202_soc_core_j22_cpu_ml_bufb[1]), .X(
        n18363) );
  sky130_fd_sc_hd__inv_6 U13445 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .Y(n13179) );
  sky130_fd_sc_hd__inv_1 U13447 ( .A(n12395), .Y(n12216) );
  sky130_fd_sc_hd__and2_1 U13448 ( .A(n24574), .B(n29587), .X(n12152) );
  sky130_fd_sc_hd__inv_2 U13449 ( .A(n24471), .Y(n29773) );
  sky130_fd_sc_hd__nand2_1 U13451 ( .A(n22264), .B(n27355), .Y(n22265) );
  sky130_fd_sc_hd__nand2_2 U13453 ( .A(n11982), .B(n11987), .Y(n29746) );
  sky130_fd_sc_hd__nand2_1 U13455 ( .A(n12466), .B(n12090), .Y(n28062) );
  sky130_fd_sc_hd__nand2_4 U13456 ( .A(n24358), .B(n27047), .Y(n28477) );
  sky130_fd_sc_hd__inv_4 U13457 ( .A(n12372), .Y(n11131) );
  sky130_fd_sc_hd__o21a_1 U13460 ( .A1(n27648), .A2(n25425), .B1(n25424), .X(
        n25426) );
  sky130_fd_sc_hd__fah_1 U13463 ( .A(n18985), .B(n18984), .CI(n18983), .COUT(
        n19038), .SUM(n19006) );
  sky130_fd_sc_hd__a21o_1 U13464 ( .A1(n12048), .A2(n18205), .B1(n17718), .X(
        n17714) );
  sky130_fd_sc_hd__and2_1 U13465 ( .A(n25313), .B(n27856), .X(n13092) );
  sky130_fd_sc_hd__inv_2 U13467 ( .A(n12045), .Y(n12046) );
  sky130_fd_sc_hd__nor2_2 U13469 ( .A(n23602), .B(n24124), .Y(n24423) );
  sky130_fd_sc_hd__o21ai_1 U13472 ( .A1(n22563), .A2(n19087), .B1(n19088), .Y(
        n21964) );
  sky130_fd_sc_hd__nor2_1 U13473 ( .A(n22562), .B(n19087), .Y(n21960) );
  sky130_fd_sc_hd__nor2_1 U13475 ( .A(n11533), .B(n23451), .Y(n28118) );
  sky130_fd_sc_hd__and2_1 U13477 ( .A(n25383), .B(n27856), .X(n12130) );
  sky130_fd_sc_hd__nand3_1 U13478 ( .A(n12029), .B(n15482), .C(n21917), .Y(
        n20426) );
  sky130_fd_sc_hd__a21o_1 U13482 ( .A1(n18530), .A2(n18533), .B1(n17365), .X(
        n17400) );
  sky130_fd_sc_hd__a21o_1 U13484 ( .A1(n18486), .A2(n18483), .B1(n18345), .X(
        n18392) );
  sky130_fd_sc_hd__and2b_1 U13485 ( .B(n18470), .A_N(n18486), .X(n17939) );
  sky130_fd_sc_hd__nand4_2 U13487 ( .A(n12955), .B(n21695), .C(n21694), .D(
        n12799), .Y(n12798) );
  sky130_fd_sc_hd__a21o_1 U13489 ( .A1(n18471), .A2(n18474), .B1(n17383), .X(
        n18956) );
  sky130_fd_sc_hd__o22ai_1 U13490 ( .A1(n23227), .A2(n23230), .B1(n23221), 
        .B2(n23222), .Y(n23175) );
  sky130_fd_sc_hd__or2_2 U13492 ( .A(n21704), .B(n21703), .X(n21706) );
  sky130_fd_sc_hd__buf_2 U13494 ( .A(n25148), .X(n10957) );
  sky130_fd_sc_hd__inv_1 U13496 ( .A(n18293), .Y(n18884) );
  sky130_fd_sc_hd__and4_1 U13497 ( .A(n27730), .B(n24552), .C(n11449), .D(
        n24551), .X(n24554) );
  sky130_fd_sc_hd__clkbuf_1 U13498 ( .A(n24543), .X(n12255) );
  sky130_fd_sc_hd__inv_1 U13499 ( .A(n23388), .Y(n22009) );
  sky130_fd_sc_hd__buf_2 U13500 ( .A(n23388), .X(n29595) );
  sky130_fd_sc_hd__inv_1 U13501 ( .A(n22786), .Y(n18920) );
  sky130_fd_sc_hd__nor2_1 U13502 ( .A(n22047), .B(n22786), .Y(n22050) );
  sky130_fd_sc_hd__inv_1 U13503 ( .A(n23228), .Y(n24386) );
  sky130_fd_sc_hd__nor2_2 U13504 ( .A(n17865), .B(n17866), .Y(n22953) );
  sky130_fd_sc_hd__o211ai_1 U13505 ( .A1(n12874), .A2(n12395), .B1(n12598), 
        .C1(n12572), .Y(n11650) );
  sky130_fd_sc_hd__nand2_1 U13506 ( .A(n11921), .B(n12572), .Y(n24619) );
  sky130_fd_sc_hd__nand4_1 U13507 ( .A(n11379), .B(n11649), .C(n24551), .D(
        n27734), .Y(n12658) );
  sky130_fd_sc_hd__inv_2 U13508 ( .A(n11660), .Y(n23408) );
  sky130_fd_sc_hd__nand2b_1 U13509 ( .A_N(n11660), .B(n11176), .Y(n12230) );
  sky130_fd_sc_hd__nor2_2 U13510 ( .A(n27743), .B(n12778), .Y(n24633) );
  sky130_fd_sc_hd__inv_1 U13512 ( .A(n10958), .Y(n12551) );
  sky130_fd_sc_hd__nand4_1 U13513 ( .A(n12552), .B(n12553), .C(n12554), .D(
        n12555), .Y(n10958) );
  sky130_fd_sc_hd__nand3_2 U13516 ( .A(n10959), .B(n17094), .C(n30029), .Y(
        n11980) );
  sky130_fd_sc_hd__buf_4 U13517 ( .A(n11001), .X(n29488) );
  sky130_fd_sc_hd__clkbuf_1 U13518 ( .A(n24563), .X(n10960) );
  sky130_fd_sc_hd__inv_1 U13519 ( .A(n11762), .Y(n11707) );
  sky130_fd_sc_hd__nand2_1 U13523 ( .A(n22008), .B(n12153), .Y(n10962) );
  sky130_fd_sc_hd__nand2_1 U13525 ( .A(n16567), .B(n17069), .Y(n16568) );
  sky130_fd_sc_hd__nand2_1 U13526 ( .A(n12727), .B(n12140), .Y(n17069) );
  sky130_fd_sc_hd__inv_1 U13527 ( .A(n24802), .Y(n22264) );
  sky130_fd_sc_hd__nand3_1 U13528 ( .A(n22263), .B(n22261), .C(n22262), .Y(
        n24802) );
  sky130_fd_sc_hd__clkbuf_1 U13532 ( .A(n30059), .X(n10965) );
  sky130_fd_sc_hd__nand2_1 U13534 ( .A(n10967), .B(n12902), .Y(n12940) );
  sky130_fd_sc_hd__nor2_1 U13535 ( .A(n12896), .B(n12897), .Y(n10967) );
  sky130_fd_sc_hd__nand3_2 U13536 ( .A(n24427), .B(n24426), .C(n24425), .Y(
        n12363) );
  sky130_fd_sc_hd__nand2_2 U13537 ( .A(n24415), .B(n24414), .Y(n24427) );
  sky130_fd_sc_hd__a21boi_2 U13538 ( .A1(n12769), .A2(n12768), .B1_N(n17333), 
        .Y(n23507) );
  sky130_fd_sc_hd__nand3_1 U13540 ( .A(n18797), .B(n23514), .C(n23505), .Y(
        n12360) );
  sky130_fd_sc_hd__nand3_1 U13542 ( .A(n12609), .B(n12600), .C(n20582), .Y(
        n21693) );
  sky130_fd_sc_hd__nand2_1 U13543 ( .A(n10968), .B(n12529), .Y(n12029) );
  sky130_fd_sc_hd__nor2_1 U13544 ( .A(n12528), .B(n12527), .Y(n10968) );
  sky130_fd_sc_hd__inv_2 U13545 ( .A(n12816), .Y(n12283) );
  sky130_fd_sc_hd__a21oi_2 U13547 ( .A1(n24772), .A2(n27152), .B1(n24774), .Y(
        n24770) );
  sky130_fd_sc_hd__clkbuf_1 U13548 ( .A(n12566), .X(n10969) );
  sky130_fd_sc_hd__o22ai_1 U13549 ( .A1(n22365), .A2(n22081), .B1(n18836), 
        .B2(n18224), .Y(n18174) );
  sky130_fd_sc_hd__clkbuf_1 U13551 ( .A(n30062), .X(n10971) );
  sky130_fd_sc_hd__clkbuf_1 U13553 ( .A(n21960), .X(n10972) );
  sky130_fd_sc_hd__nor2_1 U13554 ( .A(n24562), .B(n27742), .Y(n11446) );
  sky130_fd_sc_hd__a21oi_2 U13555 ( .A1(n26417), .A2(n17225), .B1(n16563), .Y(
        n17063) );
  sky130_fd_sc_hd__a21oi_2 U13557 ( .A1(n27152), .A2(n27773), .B1(n27778), .Y(
        n26964) );
  sky130_fd_sc_hd__nor2_1 U13562 ( .A(n11604), .B(n12924), .Y(n10975) );
  sky130_fd_sc_hd__nor2_2 U13563 ( .A(n20984), .B(n20982), .Y(n21030) );
  sky130_fd_sc_hd__inv_1 U13564 ( .A(n26917), .Y(n26961) );
  sky130_fd_sc_hd__nand2_2 U13565 ( .A(n24360), .B(n23587), .Y(n26968) );
  sky130_fd_sc_hd__nand2_1 U13566 ( .A(n18680), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .Y(n18832) );
  sky130_fd_sc_hd__nor2_2 U13567 ( .A(n21231), .B(n21230), .Y(n24769) );
  sky130_fd_sc_hd__inv_1 U13568 ( .A(n10976), .Y(n25133) );
  sky130_fd_sc_hd__nand4_1 U13569 ( .A(n25127), .B(n25126), .C(n25125), .D(
        n25124), .Y(n10976) );
  sky130_fd_sc_hd__nor2_1 U13570 ( .A(n11636), .B(n23613), .Y(n12205) );
  sky130_fd_sc_hd__nand2_1 U13571 ( .A(n10978), .B(n10977), .Y(n19015) );
  sky130_fd_sc_hd__nand2_1 U13572 ( .A(n18970), .B(n18969), .Y(n10977) );
  sky130_fd_sc_hd__o21ai_1 U13573 ( .A1(n18969), .A2(n18970), .B1(n18968), .Y(
        n10978) );
  sky130_fd_sc_hd__xnor2_1 U13574 ( .A(n18968), .B(n10979), .Y(n19009) );
  sky130_fd_sc_hd__xnor2_1 U13575 ( .A(n18969), .B(n18970), .Y(n10979) );
  sky130_fd_sc_hd__nand2_4 U13576 ( .A(n23553), .B(n11610), .Y(n11929) );
  sky130_fd_sc_hd__and3_1 U13577 ( .A(n28123), .B(n28122), .C(n28121), .X(
        n12150) );
  sky130_fd_sc_hd__mux2i_1 U13579 ( .A0(n23266), .A1(n23265), .S(n27322), .Y(
        n23368) );
  sky130_fd_sc_hd__inv_8 U13581 ( .A(n24515), .Y(n24516) );
  sky130_fd_sc_hd__o2bb2ai_1 U13582 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[20]), .B2(n26686), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[17]), .A2_N(n25578), .Y(n23185) );
  sky130_fd_sc_hd__nor2_2 U13585 ( .A(n30088), .B(n23382), .Y(n24593) );
  sky130_fd_sc_hd__a22oi_2 U13586 ( .A1(j202_soc_core_memory0_ram_dout0[20]), 
        .A2(n20457), .B1(n20456), .B2(j202_soc_core_memory0_ram_dout0[148]), 
        .Y(n15372) );
  sky130_fd_sc_hd__nand2_1 U13587 ( .A(n11608), .B(n11607), .Y(n10982) );
  sky130_fd_sc_hd__inv_4 U13589 ( .A(n12374), .Y(n11130) );
  sky130_fd_sc_hd__inv_6 U13590 ( .A(n11134), .Y(n11073) );
  sky130_fd_sc_hd__inv_2 U13595 ( .A(n23966), .Y(n29823) );
  sky130_fd_sc_hd__inv_6 U13598 ( .A(n11131), .Y(n11071) );
  sky130_fd_sc_hd__buf_8 U13599 ( .A(n12370), .X(n10983) );
  sky130_fd_sc_hd__buf_8 U13600 ( .A(n12370), .X(n10984) );
  sky130_fd_sc_hd__inv_4 U13603 ( .A(n11134), .Y(n11024) );
  sky130_fd_sc_hd__inv_4 U13604 ( .A(n11134), .Y(n11031) );
  sky130_fd_sc_hd__inv_4 U13605 ( .A(n11134), .Y(n11030) );
  sky130_fd_sc_hd__inv_4 U13606 ( .A(n11134), .Y(n11023) );
  sky130_fd_sc_hd__clkinv_2 U13612 ( .A(n11156), .Y(n11027) );
  sky130_fd_sc_hd__clkinv_2 U13614 ( .A(n11160), .Y(n11033) );
  sky130_fd_sc_hd__inv_4 U13617 ( .A(n11131), .Y(n11028) );
  sky130_fd_sc_hd__buf_8 U13619 ( .A(n11137), .X(n10989) );
  sky130_fd_sc_hd__buf_8 U13620 ( .A(n11137), .X(n12315) );
  sky130_fd_sc_hd__inv_4 U13623 ( .A(n11130), .Y(n11067) );
  sky130_fd_sc_hd__inv_4 U13625 ( .A(n11130), .Y(n11036) );
  sky130_fd_sc_hd__clkinv_2 U13627 ( .A(n11153), .Y(n11038) );
  sky130_fd_sc_hd__clkinv_2 U13628 ( .A(n11152), .Y(n11072) );
  sky130_fd_sc_hd__nand3_2 U13629 ( .A(n12016), .B(n12014), .C(n12019), .Y(
        n10994) );
  sky130_fd_sc_hd__and2_1 U13631 ( .A(n10966), .B(n29555), .X(n29639) );
  sky130_fd_sc_hd__and2_1 U13633 ( .A(n10966), .B(n29556), .X(n29643) );
  sky130_fd_sc_hd__and2_1 U13634 ( .A(n10966), .B(n29545), .X(n29637) );
  sky130_fd_sc_hd__and2_1 U13635 ( .A(n29492), .B(n29557), .X(n29641) );
  sky130_fd_sc_hd__and2_1 U13636 ( .A(n29492), .B(n29553), .X(n29642) );
  sky130_fd_sc_hd__and2_1 U13637 ( .A(n29492), .B(n29565), .X(n29636) );
  sky130_fd_sc_hd__and2_1 U13638 ( .A(n29492), .B(n29581), .X(n29640) );
  sky130_fd_sc_hd__nand3_1 U13640 ( .A(n12954), .B(n12953), .C(n12951), .Y(
        n29594) );
  sky130_fd_sc_hd__buf_2 U13641 ( .A(n22789), .X(n23021) );
  sky130_fd_sc_hd__nor2_1 U13643 ( .A(n11520), .B(n11517), .Y(n27979) );
  sky130_fd_sc_hd__a21oi_2 U13644 ( .A1(n23202), .A2(n23201), .B1(n23200), .Y(
        n27318) );
  sky130_fd_sc_hd__nand3_1 U13646 ( .A(n12518), .B(n12516), .C(n12514), .Y(
        n12513) );
  sky130_fd_sc_hd__and3_1 U13647 ( .A(n11578), .B(n29489), .C(n23550), .X(
        n23446) );
  sky130_fd_sc_hd__inv_4 U13649 ( .A(n12373), .Y(n11129) );
  sky130_fd_sc_hd__inv_6 U13650 ( .A(n11129), .Y(n11064) );
  sky130_fd_sc_hd__and2_4 U13652 ( .A(n28062), .B(n12107), .X(n10998) );
  sky130_fd_sc_hd__inv_4 U13658 ( .A(n11129), .Y(n11066) );
  sky130_fd_sc_hd__inv_4 U13659 ( .A(n11130), .Y(n11069) );
  sky130_fd_sc_hd__inv_4 U13660 ( .A(n11134), .Y(n11074) );
  sky130_fd_sc_hd__buf_8 U13665 ( .A(n12371), .X(n11127) );
  sky130_fd_sc_hd__buf_8 U13666 ( .A(n12371), .X(n11155) );
  sky130_fd_sc_hd__inv_6 U13667 ( .A(n11129), .Y(n11065) );
  sky130_fd_sc_hd__inv_6 U13668 ( .A(n11130), .Y(n11068) );
  sky130_fd_sc_hd__inv_6 U13669 ( .A(n11131), .Y(n11070) );
  sky130_fd_sc_hd__buf_8 U13674 ( .A(n12369), .X(n11136) );
  sky130_fd_sc_hd__nor2_1 U13676 ( .A(n23948), .B(n23950), .Y(n11000) );
  sky130_fd_sc_hd__nand3_1 U13677 ( .A(n11382), .B(n11015), .C(n21174), .Y(
        n11001) );
  sky130_fd_sc_hd__nor2_1 U13679 ( .A(n23947), .B(n12238), .Y(n11002) );
  sky130_fd_sc_hd__nor2_1 U13680 ( .A(n23947), .B(n12238), .Y(n12229) );
  sky130_fd_sc_hd__nand2_1 U13682 ( .A(n24605), .B(n30201), .Y(n10619) );
  sky130_fd_sc_hd__nand2_4 U13686 ( .A(n11183), .B(n25350), .Y(n28492) );
  sky130_fd_sc_hd__clkbuf_1 U13687 ( .A(n28116), .X(n11005) );
  sky130_fd_sc_hd__nor2_1 U13688 ( .A(n10957), .B(n23397), .Y(n11006) );
  sky130_fd_sc_hd__nor2_1 U13689 ( .A(n10957), .B(n23397), .Y(n24559) );
  sky130_fd_sc_hd__inv_1 U13690 ( .A(n24405), .Y(n11007) );
  sky130_fd_sc_hd__inv_1 U13691 ( .A(n12230), .Y(n11836) );
  sky130_fd_sc_hd__nand3_1 U13694 ( .A(n11782), .B(n11780), .C(n11778), .Y(
        n11008) );
  sky130_fd_sc_hd__clkbuf_1 U13695 ( .A(n23597), .X(n28344) );
  sky130_fd_sc_hd__nand4_1 U13698 ( .A(n11635), .B(n12629), .C(n12626), .D(
        n12627), .Y(n11634) );
  sky130_fd_sc_hd__nand2_1 U13700 ( .A(n12623), .B(n12630), .Y(n22003) );
  sky130_fd_sc_hd__nand2_1 U13701 ( .A(n12623), .B(n12630), .Y(n12325) );
  sky130_fd_sc_hd__a22oi_2 U13702 ( .A1(j202_soc_core_memory0_ram_dout0[39]), 
        .A2(n21633), .B1(n21640), .B2(j202_soc_core_memory0_ram_dout0[199]), 
        .Y(n17234) );
  sky130_fd_sc_hd__nand2_2 U13704 ( .A(n30132), .B(n23551), .Y(n28409) );
  sky130_fd_sc_hd__a22oi_2 U13706 ( .A1(j202_soc_core_memory0_ram_dout0[7]), 
        .A2(n21639), .B1(n21503), .B2(j202_soc_core_memory0_ram_dout0[295]), 
        .Y(n17235) );
  sky130_fd_sc_hd__nor2_1 U13707 ( .A(n30054), .B(n11883), .Y(n11012) );
  sky130_fd_sc_hd__nor3b_2 U13708 ( .C_N(n11906), .A(n28388), .B(n24619), .Y(
        n24622) );
  sky130_fd_sc_hd__nand2_1 U13709 ( .A(n23603), .B(n12417), .Y(n11013) );
  sky130_fd_sc_hd__nand2_1 U13710 ( .A(n12212), .B(n11014), .Y(n24691) );
  sky130_fd_sc_hd__nand2_1 U13713 ( .A(n11370), .B(n11369), .Y(n11015) );
  sky130_fd_sc_hd__nand2_1 U13714 ( .A(n11370), .B(n11369), .Y(n11661) );
  sky130_fd_sc_hd__inv_8 U13716 ( .A(n11087), .Y(n11089) );
  sky130_fd_sc_hd__inv_8 U13717 ( .A(n11087), .Y(n11016) );
  sky130_fd_sc_hd__inv_8 U13718 ( .A(n11087), .Y(n11017) );
  sky130_fd_sc_hd__inv_8 U13719 ( .A(n11087), .Y(n11088) );
  sky130_fd_sc_hd__inv_8 U13720 ( .A(n11087), .Y(n11018) );
  sky130_fd_sc_hd__inv_8 U13721 ( .A(n11087), .Y(n11019) );
  sky130_fd_sc_hd__inv_8 U13722 ( .A(n11087), .Y(n11090) );
  sky130_fd_sc_hd__buf_8 U13723 ( .A(n11084), .X(n11020) );
  sky130_fd_sc_hd__buf_8 U13724 ( .A(n11084), .X(n11021) );
  sky130_fd_sc_hd__buf_8 U13725 ( .A(n11084), .X(n11079) );
  sky130_fd_sc_hd__buf_8 U13728 ( .A(n11084), .X(n11163) );
  sky130_fd_sc_hd__inv_1 U13729 ( .A(n12374), .Y(n11152) );
  sky130_fd_sc_hd__inv_1 U13730 ( .A(n12373), .Y(n11154) );
  sky130_fd_sc_hd__inv_1 U13733 ( .A(n12386), .Y(n11160) );
  sky130_fd_sc_hd__inv_1 U13735 ( .A(n12374), .Y(n11153) );
  sky130_fd_sc_hd__inv_1 U13736 ( .A(n12373), .Y(n11157) );
  sky130_fd_sc_hd__inv_2 U13737 ( .A(n23984), .Y(n11167) );
  sky130_fd_sc_hd__inv_4 U13738 ( .A(n11167), .Y(n11040) );
  sky130_fd_sc_hd__inv_4 U13739 ( .A(n11167), .Y(n11041) );
  sky130_fd_sc_hd__inv_4 U13740 ( .A(n11167), .Y(n11042) );
  sky130_fd_sc_hd__inv_4 U13741 ( .A(n11167), .Y(n11043) );
  sky130_fd_sc_hd__inv_2 U13742 ( .A(n23983), .Y(n11165) );
  sky130_fd_sc_hd__inv_4 U13743 ( .A(n11165), .Y(n11044) );
  sky130_fd_sc_hd__inv_4 U13744 ( .A(n11165), .Y(n11045) );
  sky130_fd_sc_hd__inv_4 U13745 ( .A(n11165), .Y(n11046) );
  sky130_fd_sc_hd__inv_4 U13746 ( .A(n11165), .Y(n11047) );
  sky130_fd_sc_hd__inv_2 U13747 ( .A(n23988), .Y(n11166) );
  sky130_fd_sc_hd__inv_4 U13748 ( .A(n11166), .Y(n11048) );
  sky130_fd_sc_hd__inv_4 U13749 ( .A(n11166), .Y(n11049) );
  sky130_fd_sc_hd__inv_4 U13750 ( .A(n11166), .Y(n11050) );
  sky130_fd_sc_hd__inv_4 U13751 ( .A(n11166), .Y(n11051) );
  sky130_fd_sc_hd__inv_2 U13752 ( .A(n23985), .Y(n11168) );
  sky130_fd_sc_hd__inv_4 U13753 ( .A(n11168), .Y(n11052) );
  sky130_fd_sc_hd__inv_4 U13754 ( .A(n11168), .Y(n11053) );
  sky130_fd_sc_hd__inv_4 U13755 ( .A(n11168), .Y(n11054) );
  sky130_fd_sc_hd__inv_4 U13756 ( .A(n11168), .Y(n11055) );
  sky130_fd_sc_hd__inv_2 U13757 ( .A(n23987), .Y(n11169) );
  sky130_fd_sc_hd__inv_4 U13758 ( .A(n11169), .Y(n11056) );
  sky130_fd_sc_hd__inv_4 U13759 ( .A(n11169), .Y(n11057) );
  sky130_fd_sc_hd__inv_4 U13760 ( .A(n11169), .Y(n11058) );
  sky130_fd_sc_hd__inv_4 U13761 ( .A(n11169), .Y(n11059) );
  sky130_fd_sc_hd__buf_8 U13766 ( .A(n11084), .X(n11080) );
  sky130_fd_sc_hd__inv_6 U13767 ( .A(n11081), .Y(n11082) );
  sky130_fd_sc_hd__inv_2 U13768 ( .A(n23986), .Y(n11083) );
  sky130_fd_sc_hd__inv_2 U13769 ( .A(n11083), .Y(n11085) );
  sky130_fd_sc_hd__probe_p_8 U13770 ( .A(n11084), .X(n11086) );
  sky130_fd_sc_hd__clkinv_1 U13773 ( .A(n16757), .Y(n14628) );
  sky130_fd_sc_hd__clkinv_1 U13775 ( .A(n16679), .Y(n16648) );
  sky130_fd_sc_hd__clkinv_1 U13777 ( .A(n14646), .Y(n16850) );
  sky130_fd_sc_hd__clkinv_1 U13778 ( .A(n15597), .Y(n15149) );
  sky130_fd_sc_hd__clkinv_1 U13779 ( .A(n25389), .Y(n17673) );
  sky130_fd_sc_hd__clkinv_1 U13780 ( .A(n22811), .Y(n17727) );
  sky130_fd_sc_hd__clkinv_1 U13781 ( .A(n15595), .Y(n15562) );
  sky130_fd_sc_hd__clkinv_1 U13782 ( .A(n15294), .Y(n15310) );
  sky130_fd_sc_hd__clkinv_1 U13783 ( .A(n15221), .Y(n15499) );
  sky130_fd_sc_hd__clkinv_1 U13784 ( .A(n15696), .Y(n16346) );
  sky130_fd_sc_hd__clkinv_1 U13786 ( .A(n16161), .Y(n16819) );
  sky130_fd_sc_hd__clkinv_1 U13787 ( .A(n16981), .Y(n16623) );
  sky130_fd_sc_hd__clkinv_1 U13788 ( .A(n26943), .Y(n25685) );
  sky130_fd_sc_hd__clkinv_1 U13789 ( .A(n21280), .Y(n18022) );
  sky130_fd_sc_hd__o22ai_1 U13790 ( .A1(n18993), .A2(n18376), .B1(n18375), 
        .B2(n18990), .Y(n11876) );
  sky130_fd_sc_hd__inv_1 U13791 ( .A(n17661), .Y(n17658) );
  sky130_fd_sc_hd__buf_2 U13792 ( .A(j202_soc_core_j22_cpu_ml_bufb[10]), .X(
        n18962) );
  sky130_fd_sc_hd__inv_1 U13794 ( .A(n18615), .Y(n12677) );
  sky130_fd_sc_hd__buf_2 U13795 ( .A(j202_soc_core_j22_cpu_ml_bufb[15]), .X(
        n18925) );
  sky130_fd_sc_hd__clkinv_1 U13796 ( .A(n21595), .Y(n21358) );
  sky130_fd_sc_hd__clkinv_1 U13797 ( .A(n19125), .Y(n20304) );
  sky130_fd_sc_hd__clkinv_1 U13798 ( .A(n17251), .Y(n17243) );
  sky130_fd_sc_hd__clkinv_1 U13799 ( .A(n19615), .Y(n20347) );
  sky130_fd_sc_hd__clkinv_1 U13800 ( .A(n20561), .Y(n20739) );
  sky130_fd_sc_hd__clkinv_1 U13802 ( .A(n18946), .Y(n19034) );
  sky130_fd_sc_hd__fa_1 U13803 ( .A(n18548), .B(n18547), .CIN(n18546), .COUT(
        n18565), .SUM(n18580) );
  sky130_fd_sc_hd__clkinv_1 U13804 ( .A(n27618), .Y(n18110) );
  sky130_fd_sc_hd__clkinv_1 U13805 ( .A(n21530), .Y(n21125) );
  sky130_fd_sc_hd__inv_1 U13806 ( .A(n19507), .Y(n19738) );
  sky130_fd_sc_hd__clkinv_1 U13807 ( .A(n17265), .Y(n18742) );
  sky130_fd_sc_hd__clkinv_1 U13808 ( .A(n21075), .Y(n18711) );
  sky130_fd_sc_hd__clkinv_1 U13809 ( .A(n18730), .Y(n18752) );
  sky130_fd_sc_hd__clkinv_1 U13811 ( .A(n20484), .Y(n20610) );
  sky130_fd_sc_hd__clkinv_1 U13812 ( .A(n19581), .Y(n20380) );
  sky130_fd_sc_hd__clkinv_1 U13813 ( .A(n15413), .Y(n19719) );
  sky130_fd_sc_hd__clkinv_1 U13815 ( .A(n15435), .Y(n19770) );
  sky130_fd_sc_hd__clkinv_1 U13816 ( .A(n19795), .Y(n19825) );
  sky130_fd_sc_hd__clkinv_1 U13817 ( .A(n16960), .Y(n16631) );
  sky130_fd_sc_hd__clkinv_1 U13818 ( .A(n14636), .Y(n14657) );
  sky130_fd_sc_hd__clkinv_1 U13819 ( .A(j202_soc_core_bootrom_00_address_w[11]), .Y(n13182) );
  sky130_fd_sc_hd__clkinv_1 U13820 ( .A(n20296), .Y(n20338) );
  sky130_fd_sc_hd__buf_2 U13823 ( .A(j202_soc_core_j22_cpu_ml_bufb[2]), .X(
        n18372) );
  sky130_fd_sc_hd__inv_2 U13824 ( .A(n22030), .Y(n18912) );
  sky130_fd_sc_hd__clkinv_1 U13825 ( .A(n15106), .Y(n15577) );
  sky130_fd_sc_hd__clkinv_1 U13826 ( .A(n21074), .Y(n21132) );
  sky130_fd_sc_hd__clkinv_1 U13827 ( .A(n21380), .Y(n21389) );
  sky130_fd_sc_hd__clkinv_1 U13828 ( .A(n20046), .Y(n19895) );
  sky130_fd_sc_hd__clkinv_1 U13829 ( .A(n20023), .Y(n18728) );
  sky130_fd_sc_hd__clkinv_1 U13830 ( .A(n20393), .Y(n17102) );
  sky130_fd_sc_hd__clkinv_1 U13831 ( .A(n19654), .Y(n20317) );
  sky130_fd_sc_hd__clkinv_1 U13832 ( .A(n19319), .Y(n20363) );
  sky130_fd_sc_hd__clkinv_1 U13833 ( .A(n19322), .Y(n20392) );
  sky130_fd_sc_hd__inv_2 U13834 ( .A(n16986), .Y(n21103) );
  sky130_fd_sc_hd__inv_2 U13835 ( .A(n13182), .Y(n11150) );
  sky130_fd_sc_hd__clkinv_1 U13836 ( .A(n14378), .Y(n14255) );
  sky130_fd_sc_hd__clkinv_1 U13838 ( .A(n13482), .Y(n14095) );
  sky130_fd_sc_hd__clkinv_1 U13839 ( .A(n21395), .Y(n21603) );
  sky130_fd_sc_hd__clkinv_1 U13840 ( .A(n21150), .Y(n21598) );
  sky130_fd_sc_hd__clkinv_1 U13841 ( .A(j202_soc_core_j22_cpu_regop_other__2_), 
        .Y(n18860) );
  sky130_fd_sc_hd__inv_1 U13842 ( .A(n12844), .Y(n11179) );
  sky130_fd_sc_hd__clkinv_1 U13843 ( .A(n20227), .Y(n20038) );
  sky130_fd_sc_hd__clkinv_1 U13844 ( .A(n20100), .Y(n20152) );
  sky130_fd_sc_hd__or2_2 U13845 ( .A(n21088), .B(n19148), .X(n19726) );
  sky130_fd_sc_hd__clkinv_1 U13847 ( .A(n13457), .Y(n13958) );
  sky130_fd_sc_hd__clkinv_1 U13848 ( .A(n27806), .Y(n25872) );
  sky130_fd_sc_hd__clkinv_1 U13850 ( .A(n13337), .Y(n13431) );
  sky130_fd_sc_hd__clkinv_1 U13851 ( .A(n21412), .Y(n21617) );
  sky130_fd_sc_hd__clkinv_1 U13852 ( .A(n20235), .Y(n19839) );
  sky130_fd_sc_hd__inv_1 U13853 ( .A(n12515), .Y(n12514) );
  sky130_fd_sc_hd__clkinv_1 U13855 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[3]), 
        .Y(n26270) );
  sky130_fd_sc_hd__inv_2 U13856 ( .A(n12647), .Y(n12497) );
  sky130_fd_sc_hd__inv_2 U13857 ( .A(n23545), .Y(n23542) );
  sky130_fd_sc_hd__clkinv_1 U13858 ( .A(n26919), .Y(n27790) );
  sky130_fd_sc_hd__clkinv_1 U13860 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[2]), 
        .Y(n21709) );
  sky130_fd_sc_hd__clkinv_1 U13861 ( .A(n14775), .Y(n11202) );
  sky130_fd_sc_hd__clkinv_1 U13862 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[1]), 
        .Y(n26374) );
  sky130_fd_sc_hd__nand2_2 U13863 ( .A(n23095), .B(n23094), .Y(n23104) );
  sky130_fd_sc_hd__clkinv_1 U13865 ( .A(n25761), .Y(n17785) );
  sky130_fd_sc_hd__clkinv_1 U13866 ( .A(n18094), .Y(n22567) );
  sky130_fd_sc_hd__clkinv_1 U13867 ( .A(n13383), .Y(n13839) );
  sky130_fd_sc_hd__clkinv_1 U13868 ( .A(n13840), .Y(n13707) );
  sky130_fd_sc_hd__clkinv_1 U13870 ( .A(n24147), .Y(n24152) );
  sky130_fd_sc_hd__clkinv_1 U13873 ( .A(n23550), .Y(n11182) );
  sky130_fd_sc_hd__inv_2 U13875 ( .A(n25557), .Y(n25559) );
  sky130_fd_sc_hd__clkinv_1 U13880 ( .A(n12286), .Y(n12287) );
  sky130_fd_sc_hd__clkinv_1 U13881 ( .A(n24627), .Y(n11170) );
  sky130_fd_sc_hd__clkinv_1 U13882 ( .A(n23137), .Y(n23149) );
  sky130_fd_sc_hd__inv_2 U13885 ( .A(n16110), .Y(n12973) );
  sky130_fd_sc_hd__clkinv_1 U13886 ( .A(n26421), .Y(n28502) );
  sky130_fd_sc_hd__clkinv_1 U13887 ( .A(n23621), .Y(n23622) );
  sky130_fd_sc_hd__clkinv_1 U13888 ( .A(n25220), .Y(n22101) );
  sky130_fd_sc_hd__clkbuf_1 U13890 ( .A(n12039), .X(n12402) );
  sky130_fd_sc_hd__clkinv_1 U13891 ( .A(n12653), .Y(n11192) );
  sky130_fd_sc_hd__clkinv_1 U13892 ( .A(j202_soc_core_ahb2wbqspi_00_stb_o), 
        .Y(n28866) );
  sky130_fd_sc_hd__clkinv_1 U13894 ( .A(j202_soc_core_j22_cpu_macop_MAC_[1]), 
        .Y(n28053) );
  sky130_fd_sc_hd__clkinv_1 U13895 ( .A(j202_soc_core_intc_core_00_rg_ipr[23]), 
        .Y(n26688) );
  sky130_fd_sc_hd__clkinv_1 U13897 ( .A(j202_soc_core_intc_core_00_rg_ipr[63]), 
        .Y(n26759) );
  sky130_fd_sc_hd__clkinv_1 U13898 ( .A(j202_soc_core_intc_core_00_rg_ipr[37]), 
        .Y(n26726) );
  sky130_fd_sc_hd__clkinv_1 U13899 ( .A(j202_soc_core_intc_core_00_rg_ipr[69]), 
        .Y(n27151) );
  sky130_fd_sc_hd__clkinv_1 U13900 ( .A(j202_soc_core_intc_core_00_rg_ipr[1]), 
        .Y(n24809) );
  sky130_fd_sc_hd__clkinv_1 U13901 ( .A(n30050), .Y(n12262) );
  sky130_fd_sc_hd__clkinv_1 U13902 ( .A(n29169), .Y(n28564) );
  sky130_fd_sc_hd__nand2_1 U13903 ( .A(n28442), .B(n28432), .Y(n28535) );
  sky130_fd_sc_hd__clkinv_1 U13904 ( .A(n23749), .Y(n24832) );
  sky130_fd_sc_hd__inv_2 U13905 ( .A(n12431), .Y(n24788) );
  sky130_fd_sc_hd__clkinv_1 U13906 ( .A(n24901), .Y(n28480) );
  sky130_fd_sc_hd__nor2_1 U13907 ( .A(n24291), .B(n28425), .Y(n27615) );
  sky130_fd_sc_hd__buf_2 U13908 ( .A(n25240), .X(n25245) );
  sky130_fd_sc_hd__inv_2 U13909 ( .A(n12402), .Y(n27461) );
  sky130_fd_sc_hd__clkinv_1 U13910 ( .A(n24141), .Y(n11161) );
  sky130_fd_sc_hd__clkinv_1 U13911 ( .A(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n28896) );
  sky130_fd_sc_hd__nand2_2 U13912 ( .A(n28691), .B(n26466), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N390) );
  sky130_fd_sc_hd__clkbuf_1 U13913 ( .A(n10712), .X(n29825) );
  sky130_fd_sc_hd__nand2_1 U13915 ( .A(n28895), .B(n12069), .Y(n29753) );
  sky130_fd_sc_hd__nand3_1 U13916 ( .A(n26567), .B(n28721), .C(n23854), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N311) );
  sky130_fd_sc_hd__clkinv_1 U13918 ( .A(gpio_en_o[0]), .Y(io_oeb[0]) );
  sky130_fd_sc_hd__clkinv_1 U13919 ( .A(gpio_en_o[9]), .Y(io_oeb[29]) );
  sky130_fd_sc_hd__and2_1 U13921 ( .A(n13385), .B(n13390), .X(n11091) );
  sky130_fd_sc_hd__and2_1 U13922 ( .A(n12943), .B(n11560), .X(n11092) );
  sky130_fd_sc_hd__inv_4 U13923 ( .A(n13392), .Y(n14275) );
  sky130_fd_sc_hd__and2_1 U13925 ( .A(j202_soc_core_j22_cpu_regop_Rs__1_), .B(
        j202_soc_core_j22_cpu_regop_Rs__0_), .X(n11094) );
  sky130_fd_sc_hd__and2_1 U13926 ( .A(n21025), .B(n12771), .X(n11096) );
  sky130_fd_sc_hd__and2_1 U13929 ( .A(n23030), .B(n23035), .X(n11099) );
  sky130_fd_sc_hd__o21a_1 U13930 ( .A1(n22783), .A2(n22604), .B1(n22785), .X(
        n11100) );
  sky130_fd_sc_hd__and2_1 U13932 ( .A(n12751), .B(n19428), .X(n11102) );
  sky130_fd_sc_hd__and2_1 U13934 ( .A(n25561), .B(n25560), .X(n11104) );
  sky130_fd_sc_hd__and2_1 U13935 ( .A(n12355), .B(n12356), .X(n11105) );
  sky130_fd_sc_hd__and2_1 U13936 ( .A(n12346), .B(n12345), .X(n11106) );
  sky130_fd_sc_hd__and4_1 U13937 ( .A(n20413), .B(n20414), .C(n11670), .D(
        n20412), .X(n11107) );
  sky130_fd_sc_hd__nand2_2 U13938 ( .A(n20425), .B(n20426), .Y(n23378) );
  sky130_fd_sc_hd__nand2_2 U13939 ( .A(n20425), .B(n20426), .Y(n12220) );
  sky130_fd_sc_hd__and3_1 U13940 ( .A(n21838), .B(n21839), .C(n21840), .X(
        n11108) );
  sky130_fd_sc_hd__inv_4 U13941 ( .A(n12087), .Y(n27146) );
  sky130_fd_sc_hd__inv_1 U13942 ( .A(n26168), .Y(n12366) );
  sky130_fd_sc_hd__and4_1 U13943 ( .A(n24171), .B(n24170), .C(n24169), .D(
        n24168), .X(n11109) );
  sky130_fd_sc_hd__a21oi_2 U13944 ( .A1(n26025), .A2(n27152), .B1(n26027), .Y(
        n26023) );
  sky130_fd_sc_hd__inv_1 U13945 ( .A(n25962), .Y(n11181) );
  sky130_fd_sc_hd__nor2_1 U13946 ( .A(n26194), .B(n12361), .Y(n25962) );
  sky130_fd_sc_hd__and2_1 U13948 ( .A(n28378), .B(n24104), .X(n11110) );
  sky130_fd_sc_hd__o211ai_2 U13949 ( .A1(n12395), .A2(n12874), .B1(n12598), 
        .C1(n12572), .Y(n23552) );
  sky130_fd_sc_hd__inv_2 U13950 ( .A(n23552), .Y(n24958) );
  sky130_fd_sc_hd__and2_1 U13951 ( .A(n12326), .B(n12716), .X(n11111) );
  sky130_fd_sc_hd__and2_4 U13952 ( .A(n11436), .B(n28417), .X(n11112) );
  sky130_fd_sc_hd__and3_2 U13955 ( .A(n26066), .B(n26065), .C(n11530), .X(
        n11115) );
  sky130_fd_sc_hd__nand2_4 U13958 ( .A(n12534), .B(n29828), .Y(n12276) );
  sky130_fd_sc_hd__nand2_2 U13959 ( .A(n23400), .B(n23399), .Y(n11906) );
  sky130_fd_sc_hd__nor2_1 U13960 ( .A(n12220), .B(n30079), .Y(n11596) );
  sky130_fd_sc_hd__inv_1 U13961 ( .A(n24562), .Y(n22004) );
  sky130_fd_sc_hd__fah_1 U13966 ( .A(n22030), .B(n22029), .CI(n22028), .COUT(
        n22035), .SUM(n22032) );
  sky130_fd_sc_hd__inv_1 U13968 ( .A(n18276), .Y(n12179) );
  sky130_fd_sc_hd__nand3_1 U13969 ( .A(n20886), .B(n20888), .C(n20887), .Y(
        n29481) );
  sky130_fd_sc_hd__nand2_2 U13971 ( .A(n23398), .B(n12861), .Y(n24563) );
  sky130_fd_sc_hd__inv_1 U13972 ( .A(n27315), .Y(n27317) );
  sky130_fd_sc_hd__inv_1 U13973 ( .A(n22789), .Y(n22604) );
  sky130_fd_sc_hd__o21a_1 U13975 ( .A1(n28532), .A2(n26939), .B1(n26919), .X(
        n11775) );
  sky130_fd_sc_hd__o22a_1 U13976 ( .A1(n26322), .A2(n11186), .B1(n28532), .B2(
        n22743), .X(n20980) );
  sky130_fd_sc_hd__nor2_1 U13978 ( .A(n23550), .B(n12362), .Y(n11551) );
  sky130_fd_sc_hd__inv_2 U13980 ( .A(n17993), .Y(n11118) );
  sky130_fd_sc_hd__inv_4 U13981 ( .A(n11118), .Y(n11119) );
  sky130_fd_sc_hd__nand2_1 U13982 ( .A(n17454), .B(n17453), .Y(n17993) );
  sky130_fd_sc_hd__a21oi_2 U13984 ( .A1(n23075), .A2(n23074), .B1(n23073), .Y(
        n27325) );
  sky130_fd_sc_hd__nand2_1 U13985 ( .A(n23156), .B(n23155), .Y(n23160) );
  sky130_fd_sc_hd__inv_1 U13986 ( .A(n27910), .Y(n11633) );
  sky130_fd_sc_hd__a21oi_2 U13987 ( .A1(n23288), .A2(n23287), .B1(n23286), .Y(
        n27342) );
  sky130_fd_sc_hd__mux2i_1 U13988 ( .A0(j202_soc_core_intc_core_00_rg_ipr[37]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[33]), .S(n23104), .Y(n23127) );
  sky130_fd_sc_hd__o211ai_1 U13989 ( .A1(n28379), .A2(n12345), .B1(n24965), 
        .C1(n28349), .Y(n25902) );
  sky130_fd_sc_hd__inv_1 U13990 ( .A(n22007), .Y(n12278) );
  sky130_fd_sc_hd__nand3_2 U13992 ( .A(n21980), .B(n21981), .C(n21982), .Y(
        n24790) );
  sky130_fd_sc_hd__a21oi_1 U13993 ( .A1(n25375), .A2(n27052), .B1(n26926), .Y(
        n23545) );
  sky130_fd_sc_hd__a21oi_1 U13994 ( .A1(n22281), .A2(n24764), .B1(n22280), .Y(
        n25375) );
  sky130_fd_sc_hd__nand2_1 U13995 ( .A(n22521), .B(n12895), .Y(n29502) );
  sky130_fd_sc_hd__and2_1 U13996 ( .A(n25856), .B(n27856), .X(n12133) );
  sky130_fd_sc_hd__nand3_1 U13998 ( .A(n22521), .B(n22520), .C(n12894), .Y(
        n29520) );
  sky130_fd_sc_hd__inv_2 U13999 ( .A(n29761), .Y(n12369) );
  sky130_fd_sc_hd__clkinv_1 U14001 ( .A(n25221), .Y(n25223) );
  sky130_fd_sc_hd__clkinv_1 U14002 ( .A(n24853), .Y(n12234) );
  sky130_fd_sc_hd__a21bo_2 U14003 ( .A1(n27617), .A2(n27152), .B1_N(n24682), 
        .X(n11475) );
  sky130_fd_sc_hd__nand3_1 U14004 ( .A(n22382), .B(n22381), .C(n22380), .Y(
        n27617) );
  sky130_fd_sc_hd__clkinv_1 U14005 ( .A(n12255), .Y(n24544) );
  sky130_fd_sc_hd__nand3_1 U14006 ( .A(n11170), .B(n11172), .C(n11110), .Y(
        n11632) );
  sky130_fd_sc_hd__inv_2 U14007 ( .A(n24421), .Y(n24424) );
  sky130_fd_sc_hd__and2_0 U14008 ( .A(n24146), .B(n24145), .X(n12107) );
  sky130_fd_sc_hd__and2_0 U14010 ( .A(n28268), .B(n11906), .X(n11905) );
  sky130_fd_sc_hd__inv_1 U14011 ( .A(n23950), .Y(n23951) );
  sky130_fd_sc_hd__clkinv_1 U14012 ( .A(n24422), .Y(n24116) );
  sky130_fd_sc_hd__nand2_1 U14013 ( .A(n24098), .B(n11646), .Y(n28090) );
  sky130_fd_sc_hd__nand2_1 U14015 ( .A(n11658), .B(n11656), .Y(n24406) );
  sky130_fd_sc_hd__inv_1 U14016 ( .A(n11517), .Y(n23406) );
  sky130_fd_sc_hd__clkinv_1 U14017 ( .A(n25029), .Y(n23053) );
  sky130_fd_sc_hd__inv_2 U14018 ( .A(n25855), .Y(n27389) );
  sky130_fd_sc_hd__inv_2 U14019 ( .A(n28470), .Y(n27897) );
  sky130_fd_sc_hd__buf_2 U14020 ( .A(n27572), .X(n12264) );
  sky130_fd_sc_hd__nor2_1 U14022 ( .A(n30063), .B(n12299), .Y(n17078) );
  sky130_fd_sc_hd__inv_2 U14023 ( .A(n25634), .Y(n25660) );
  sky130_fd_sc_hd__buf_2 U14024 ( .A(n12284), .X(n11442) );
  sky130_fd_sc_hd__clkinv_1 U14026 ( .A(n12094), .Y(n12726) );
  sky130_fd_sc_hd__nand2b_1 U14027 ( .A_N(n12351), .B(n12423), .Y(n27044) );
  sky130_fd_sc_hd__nand3_1 U14028 ( .A(n12751), .B(n19428), .C(n21919), .Y(
        n19543) );
  sky130_fd_sc_hd__clkinv_1 U14029 ( .A(n13365), .Y(n17048) );
  sky130_fd_sc_hd__and2_0 U14030 ( .A(n21318), .B(n22232), .X(n11795) );
  sky130_fd_sc_hd__inv_4 U14031 ( .A(n28379), .Y(n28417) );
  sky130_fd_sc_hd__nand2_1 U14032 ( .A(n28109), .B(n23753), .Y(n23841) );
  sky130_fd_sc_hd__clkinv_1 U14033 ( .A(n16718), .Y(n16719) );
  sky130_fd_sc_hd__inv_2 U14034 ( .A(n24879), .Y(n27616) );
  sky130_fd_sc_hd__or2_1 U14035 ( .A(n22475), .B(n11145), .X(n13046) );
  sky130_fd_sc_hd__nand3_1 U14036 ( .A(n14927), .B(n14926), .C(n12100), .Y(
        n25692) );
  sky130_fd_sc_hd__clkinv_1 U14037 ( .A(n26408), .Y(n28431) );
  sky130_fd_sc_hd__nand3_1 U14038 ( .A(n13525), .B(n12102), .C(n13524), .Y(
        n26378) );
  sky130_fd_sc_hd__a21oi_2 U14039 ( .A1(n19264), .A2(n16523), .B1(n13920), .Y(
        n26937) );
  sky130_fd_sc_hd__clkinv_1 U14040 ( .A(n15438), .Y(n19823) );
  sky130_fd_sc_hd__clkinv_1 U14041 ( .A(n21020), .Y(n11642) );
  sky130_fd_sc_hd__clkinv_1 U14042 ( .A(n19801), .Y(n15428) );
  sky130_fd_sc_hd__nand3_1 U14044 ( .A(n12167), .B(n28047), .C(n11146), .Y(
        n11562) );
  sky130_fd_sc_hd__clkinv_1 U14046 ( .A(n19434), .Y(n19512) );
  sky130_fd_sc_hd__clkinv_1 U14047 ( .A(n16694), .Y(n16642) );
  sky130_fd_sc_hd__clkinv_1 U14048 ( .A(n20815), .Y(n20766) );
  sky130_fd_sc_hd__clkinv_1 U14049 ( .A(n15593), .Y(n15230) );
  sky130_fd_sc_hd__inv_2 U14050 ( .A(n11148), .Y(n14798) );
  sky130_fd_sc_hd__clkinv_1 U14051 ( .A(n16654), .Y(n15666) );
  sky130_fd_sc_hd__nor2_1 U14052 ( .A(n18830), .B(n17358), .Y(n18678) );
  sky130_fd_sc_hd__inv_4 U14053 ( .A(n13726), .Y(n23787) );
  sky130_fd_sc_hd__inv_2 U14054 ( .A(n30190), .Y(n15951) );
  sky130_fd_sc_hd__inv_4 U14055 ( .A(n13725), .Y(n23792) );
  sky130_fd_sc_hd__or2_1 U14056 ( .A(n18535), .B(n18534), .X(n18541) );
  sky130_fd_sc_hd__inv_2 U14057 ( .A(n13958), .Y(n11125) );
  sky130_fd_sc_hd__clkinv_1 U14058 ( .A(n20850), .Y(n20630) );
  sky130_fd_sc_hd__clkinv_1 U14060 ( .A(n20210), .Y(n19910) );
  sky130_fd_sc_hd__clkinv_1 U14061 ( .A(n17564), .Y(n12481) );
  sky130_fd_sc_hd__clkinv_1 U14062 ( .A(n13425), .Y(n18870) );
  sky130_fd_sc_hd__clkinv_1 U14064 ( .A(n18731), .Y(n18763) );
  sky130_fd_sc_hd__and2_0 U14065 ( .A(n13287), .B(n13286), .X(n13347) );
  sky130_fd_sc_hd__clkinv_1 U14066 ( .A(j202_soc_core_ahb2apb_00_state[0]), 
        .Y(n21049) );
  sky130_fd_sc_hd__clkinv_1 U14067 ( .A(j202_soc_core_ahb2apb_00_state[1]), 
        .Y(n24724) );
  sky130_fd_sc_hd__clkinv_1 U14068 ( .A(j202_soc_core_memory0_ram_dout0_sel[7]), .Y(n15192) );
  sky130_fd_sc_hd__nand2_1 U14069 ( .A(n29527), .B(n11853), .Y(n24517) );
  sky130_fd_sc_hd__clkinv_1 U14071 ( .A(n25769), .Y(n23561) );
  sky130_fd_sc_hd__nand3_1 U14072 ( .A(n22737), .B(n21766), .C(n21767), .Y(
        n29526) );
  sky130_fd_sc_hd__nand2_1 U14073 ( .A(n23043), .B(n23042), .Y(n25464) );
  sky130_fd_sc_hd__and2_1 U14074 ( .A(n25131), .B(n25130), .X(n25132) );
  sky130_fd_sc_hd__inv_2 U14076 ( .A(n29492), .Y(n12843) );
  sky130_fd_sc_hd__inv_1 U14077 ( .A(n29597), .Y(n28200) );
  sky130_fd_sc_hd__o22ai_1 U14079 ( .A1(n23455), .A2(n28417), .B1(n11664), 
        .B2(n28114), .Y(n11502) );
  sky130_fd_sc_hd__inv_1 U14081 ( .A(n24924), .Y(n21765) );
  sky130_fd_sc_hd__nand3_1 U14082 ( .A(n11663), .B(n23454), .C(n11662), .Y(
        n11664) );
  sky130_fd_sc_hd__nand3_1 U14083 ( .A(n11665), .B(n11170), .C(n27910), .Y(
        n23548) );
  sky130_fd_sc_hd__inv_1 U14084 ( .A(n27016), .Y(n25937) );
  sky130_fd_sc_hd__o21a_1 U14085 ( .A1(n22780), .A2(n21729), .B1(n22799), .X(
        n22737) );
  sky130_fd_sc_hd__a21oi_1 U14086 ( .A1(n24904), .A2(n27152), .B1(n24907), .Y(
        n24913) );
  sky130_fd_sc_hd__nand3_1 U14087 ( .A(n25259), .B(n25260), .C(n25258), .Y(
        n25281) );
  sky130_fd_sc_hd__nand3_1 U14088 ( .A(n24682), .B(n22382), .C(n12913), .Y(
        n18857) );
  sky130_fd_sc_hd__nor2_1 U14089 ( .A(n23449), .B(n23450), .Y(n28115) );
  sky130_fd_sc_hd__inv_2 U14090 ( .A(n25770), .Y(n24853) );
  sky130_fd_sc_hd__nor2_1 U14091 ( .A(n11631), .B(n11632), .Y(n12346) );
  sky130_fd_sc_hd__and2_0 U14092 ( .A(n28269), .B(n11905), .X(n11904) );
  sky130_fd_sc_hd__nand2_1 U14093 ( .A(n23478), .B(n24452), .Y(n22382) );
  sky130_fd_sc_hd__inv_2 U14094 ( .A(n25024), .Y(n11138) );
  sky130_fd_sc_hd__inv_2 U14095 ( .A(n23463), .Y(n25770) );
  sky130_fd_sc_hd__clkinv_1 U14096 ( .A(n12251), .Y(n12211) );
  sky130_fd_sc_hd__inv_1 U14097 ( .A(n24553), .Y(n11604) );
  sky130_fd_sc_hd__clkinv_1 U14098 ( .A(n12821), .Y(n27731) );
  sky130_fd_sc_hd__o21ai_1 U14099 ( .A1(n19300), .A2(n12349), .B1(n19299), .Y(
        n19301) );
  sky130_fd_sc_hd__a21o_1 U14100 ( .A1(n27713), .A2(n23368), .B1(n23367), .X(
        n12093) );
  sky130_fd_sc_hd__o21a_1 U14101 ( .A1(n25658), .A2(n25664), .B1(n25657), .X(
        n25667) );
  sky130_fd_sc_hd__o21ai_1 U14102 ( .A1(n11866), .A2(n22273), .B1(n22272), .Y(
        n22274) );
  sky130_fd_sc_hd__inv_1 U14103 ( .A(n28262), .Y(n12966) );
  sky130_fd_sc_hd__nor2_1 U14104 ( .A(n24106), .B(n28090), .Y(n28151) );
  sky130_fd_sc_hd__clkinv_1 U14105 ( .A(n27905), .Y(n27906) );
  sky130_fd_sc_hd__a21oi_1 U14108 ( .A1(n27727), .A2(n28091), .B1(n27981), .Y(
        n12250) );
  sky130_fd_sc_hd__clkbuf_1 U14110 ( .A(n12583), .X(n11705) );
  sky130_fd_sc_hd__nand2_1 U14111 ( .A(n12922), .B(n28261), .Y(n23608) );
  sky130_fd_sc_hd__clkinv_1 U14112 ( .A(n11533), .Y(n23555) );
  sky130_fd_sc_hd__nand3_1 U14113 ( .A(n11910), .B(n10981), .C(n23444), .Y(
        n28416) );
  sky130_fd_sc_hd__nand3_1 U14114 ( .A(n11646), .B(n27979), .C(n12239), .Y(
        n24636) );
  sky130_fd_sc_hd__inv_1 U14115 ( .A(n24409), .Y(n28076) );
  sky130_fd_sc_hd__nand2_1 U14116 ( .A(n12326), .B(n11646), .Y(n11994) );
  sky130_fd_sc_hd__clkbuf_1 U14118 ( .A(n24399), .X(n24628) );
  sky130_fd_sc_hd__inv_1 U14119 ( .A(n11912), .Y(n11910) );
  sky130_fd_sc_hd__clkbuf_1 U14120 ( .A(n24550), .X(n11669) );
  sky130_fd_sc_hd__and2_0 U14121 ( .A(n12127), .B(n20899), .X(n12358) );
  sky130_fd_sc_hd__nand3_1 U14125 ( .A(n12201), .B(n12199), .C(n12197), .Y(
        n21865) );
  sky130_fd_sc_hd__nand2_1 U14126 ( .A(n25632), .B(n26916), .Y(n25352) );
  sky130_fd_sc_hd__nor2_2 U14127 ( .A(n24294), .B(n12351), .Y(n25433) );
  sky130_fd_sc_hd__nor2_1 U14128 ( .A(n24144), .B(n16100), .Y(n16571) );
  sky130_fd_sc_hd__inv_1 U14129 ( .A(n17058), .Y(n12334) );
  sky130_fd_sc_hd__and2_1 U14130 ( .A(n23955), .B(n12217), .X(n12218) );
  sky130_fd_sc_hd__clkinv_1 U14131 ( .A(n28027), .Y(n28036) );
  sky130_fd_sc_hd__and2_1 U14132 ( .A(n16307), .B(n12295), .X(n12140) );
  sky130_fd_sc_hd__a21oi_1 U14133 ( .A1(n23036), .A2(n19298), .B1(n19297), .Y(
        n19299) );
  sky130_fd_sc_hd__nand2_1 U14134 ( .A(n11536), .B(n22221), .Y(n11537) );
  sky130_fd_sc_hd__and2_0 U14137 ( .A(n12417), .B(n23421), .X(n12154) );
  sky130_fd_sc_hd__clkinv_1 U14138 ( .A(n24281), .Y(n26180) );
  sky130_fd_sc_hd__clkinv_1 U14139 ( .A(n11444), .Y(n12208) );
  sky130_fd_sc_hd__clkinv_1 U14140 ( .A(n27726), .Y(n27727) );
  sky130_fd_sc_hd__nand2_2 U14141 ( .A(n12066), .B(n23426), .Y(n12778) );
  sky130_fd_sc_hd__nand3_1 U14142 ( .A(n17066), .B(n16198), .C(n17064), .Y(
        n16199) );
  sky130_fd_sc_hd__and2_1 U14143 ( .A(n12495), .B(n21318), .X(n11796) );
  sky130_fd_sc_hd__a21oi_1 U14144 ( .A1(n27067), .A2(n17225), .B1(n16197), .Y(
        n17064) );
  sky130_fd_sc_hd__and2_0 U14145 ( .A(n11820), .B(n11811), .X(n11810) );
  sky130_fd_sc_hd__nand2_1 U14146 ( .A(n12417), .B(n28417), .Y(n11903) );
  sky130_fd_sc_hd__clkinv_1 U14147 ( .A(n11349), .Y(n21682) );
  sky130_fd_sc_hd__inv_2 U14150 ( .A(n11911), .Y(n11140) );
  sky130_fd_sc_hd__and2_0 U14152 ( .A(n16305), .B(n16306), .X(n12295) );
  sky130_fd_sc_hd__nand2_1 U14153 ( .A(n24357), .B(n22739), .Y(n12727) );
  sky130_fd_sc_hd__o211a_2 U14154 ( .A1(n26320), .A2(n11186), .B1(n21028), 
        .C1(n21027), .X(n21038) );
  sky130_fd_sc_hd__clkinv_1 U14155 ( .A(n11426), .Y(n22961) );
  sky130_fd_sc_hd__inv_2 U14156 ( .A(n29489), .Y(n11141) );
  sky130_fd_sc_hd__nand2_1 U14157 ( .A(n29848), .B(n22232), .Y(n11849) );
  sky130_fd_sc_hd__o2bb2ai_1 U14158 ( .B1(n25940), .B2(n24074), .A1_N(n25938), 
        .A2_N(n10965), .Y(n26192) );
  sky130_fd_sc_hd__a21oi_1 U14159 ( .A1(n11185), .A2(n11822), .B1(n11821), .Y(
        n11820) );
  sky130_fd_sc_hd__clkinv_1 U14160 ( .A(n10965), .Y(n26171) );
  sky130_fd_sc_hd__clkinv_1 U14161 ( .A(n17857), .Y(n12540) );
  sky130_fd_sc_hd__inv_1 U14162 ( .A(n12631), .Y(n20255) );
  sky130_fd_sc_hd__inv_1 U14164 ( .A(n25939), .Y(n29847) );
  sky130_fd_sc_hd__inv_2 U14165 ( .A(n29481), .Y(n11142) );
  sky130_fd_sc_hd__and2_0 U14166 ( .A(n21963), .B(n21961), .X(n21683) );
  sky130_fd_sc_hd__or2_0 U14167 ( .A(n24696), .B(n24411), .X(n13072) );
  sky130_fd_sc_hd__inv_2 U14168 ( .A(n22705), .Y(n21322) );
  sky130_fd_sc_hd__inv_1 U14169 ( .A(n19087), .Y(n19089) );
  sky130_fd_sc_hd__buf_4 U14170 ( .A(n14589), .X(n17225) );
  sky130_fd_sc_hd__clkinv_1 U14172 ( .A(n22193), .Y(n22194) );
  sky130_fd_sc_hd__inv_2 U14174 ( .A(n25985), .Y(n27842) );
  sky130_fd_sc_hd__inv_2 U14175 ( .A(n25977), .Y(n28061) );
  sky130_fd_sc_hd__inv_2 U14176 ( .A(n25988), .Y(n27845) );
  sky130_fd_sc_hd__inv_2 U14177 ( .A(n25987), .Y(n27844) );
  sky130_fd_sc_hd__inv_2 U14178 ( .A(n25980), .Y(n27835) );
  sky130_fd_sc_hd__inv_2 U14179 ( .A(n25984), .Y(n27840) );
  sky130_fd_sc_hd__nor2_2 U14180 ( .A(n18663), .B(n18664), .Y(n22199) );
  sky130_fd_sc_hd__inv_2 U14181 ( .A(n25989), .Y(n27846) );
  sky130_fd_sc_hd__clkinv_1 U14182 ( .A(n11403), .Y(n21755) );
  sky130_fd_sc_hd__nor2_1 U14183 ( .A(n11204), .B(n22222), .Y(n11369) );
  sky130_fd_sc_hd__nand2_1 U14184 ( .A(n26168), .B(n11205), .Y(n22115) );
  sky130_fd_sc_hd__inv_2 U14185 ( .A(n17053), .Y(n22739) );
  sky130_fd_sc_hd__nor2_1 U14186 ( .A(n17861), .B(n17862), .Y(n21268) );
  sky130_fd_sc_hd__inv_2 U14187 ( .A(n25978), .Y(n27834) );
  sky130_fd_sc_hd__inv_2 U14189 ( .A(n25983), .Y(n27838) );
  sky130_fd_sc_hd__inv_2 U14190 ( .A(n26894), .Y(n27839) );
  sky130_fd_sc_hd__clkinv_1 U14191 ( .A(n11471), .Y(n21875) );
  sky130_fd_sc_hd__inv_2 U14192 ( .A(n25979), .Y(n28112) );
  sky130_fd_sc_hd__inv_2 U14193 ( .A(n25986), .Y(n27843) );
  sky130_fd_sc_hd__and2_1 U14194 ( .A(n16887), .B(n12570), .X(n12143) );
  sky130_fd_sc_hd__o21ai_2 U14197 ( .A1(n22109), .A2(n18683), .B1(n18684), .Y(
        n21753) );
  sky130_fd_sc_hd__clkinv_1 U14198 ( .A(n19059), .Y(n19060) );
  sky130_fd_sc_hd__nor2_1 U14199 ( .A(n11630), .B(n11629), .Y(n12882) );
  sky130_fd_sc_hd__inv_1 U14200 ( .A(n22920), .Y(n21760) );
  sky130_fd_sc_hd__clkinv_1 U14201 ( .A(n20088), .Y(n20957) );
  sky130_fd_sc_hd__clkinv_1 U14202 ( .A(n21826), .Y(n11919) );
  sky130_fd_sc_hd__inv_1 U14203 ( .A(n20431), .Y(n20433) );
  sky130_fd_sc_hd__clkinv_1 U14204 ( .A(n20700), .Y(n20714) );
  sky130_fd_sc_hd__nand4_1 U14205 ( .A(n12736), .B(n12737), .C(n12733), .D(
        n12126), .Y(n11629) );
  sky130_fd_sc_hd__clkinv_1 U14206 ( .A(n16544), .Y(n17029) );
  sky130_fd_sc_hd__or2_0 U14207 ( .A(n22069), .B(n22175), .X(n22071) );
  sky130_fd_sc_hd__clkinv_1 U14208 ( .A(n22593), .Y(n23020) );
  sky130_fd_sc_hd__inv_1 U14209 ( .A(n22748), .Y(n22750) );
  sky130_fd_sc_hd__or2_0 U14210 ( .A(n25803), .B(n25804), .X(n25805) );
  sky130_fd_sc_hd__or2_0 U14211 ( .A(n18164), .B(n18165), .X(n12141) );
  sky130_fd_sc_hd__clkinv_1 U14212 ( .A(n17840), .Y(n17837) );
  sky130_fd_sc_hd__or2_0 U14214 ( .A(n22058), .B(n22059), .X(n22333) );
  sky130_fd_sc_hd__or2_0 U14215 ( .A(n22486), .B(n22487), .X(n22710) );
  sky130_fd_sc_hd__or2_0 U14216 ( .A(n22064), .B(n22065), .X(n22173) );
  sky130_fd_sc_hd__or2_0 U14218 ( .A(n22492), .B(n22493), .X(n22671) );
  sky130_fd_sc_hd__or2_0 U14219 ( .A(n22053), .B(n22054), .X(n22351) );
  sky130_fd_sc_hd__and2_0 U14220 ( .A(n22827), .B(n22825), .X(n11861) );
  sky130_fd_sc_hd__or2_0 U14221 ( .A(n22500), .B(n22501), .X(n22619) );
  sky130_fd_sc_hd__clkinv_1 U14223 ( .A(n18152), .Y(n18150) );
  sky130_fd_sc_hd__or2_0 U14224 ( .A(n22042), .B(n22043), .X(n22829) );
  sky130_fd_sc_hd__clkinv_1 U14225 ( .A(n28495), .Y(n25944) );
  sky130_fd_sc_hd__or2_0 U14226 ( .A(n22476), .B(n13046), .X(n22478) );
  sky130_fd_sc_hd__inv_1 U14227 ( .A(n12952), .Y(n12951) );
  sky130_fd_sc_hd__inv_2 U14228 ( .A(n26377), .Y(n11188) );
  sky130_fd_sc_hd__and2_0 U14229 ( .A(n22260), .B(n11205), .X(n22221) );
  sky130_fd_sc_hd__inv_2 U14230 ( .A(n26378), .Y(n11191) );
  sky130_fd_sc_hd__nand3_1 U14232 ( .A(n14233), .B(n13085), .C(n14232), .Y(
        n24879) );
  sky130_fd_sc_hd__nand4_2 U14233 ( .A(n13817), .B(n12092), .C(n13050), .D(
        n13816), .Y(n26377) );
  sky130_fd_sc_hd__inv_1 U14234 ( .A(n12654), .Y(n12498) );
  sky130_fd_sc_hd__nand3_1 U14235 ( .A(n13554), .B(n13541), .C(n13553), .Y(
        n22260) );
  sky130_fd_sc_hd__clkinv_1 U14236 ( .A(n16661), .Y(n16662) );
  sky130_fd_sc_hd__nand3_1 U14237 ( .A(n14812), .B(n14811), .C(n14810), .Y(
        n25271) );
  sky130_fd_sc_hd__nand3_1 U14238 ( .A(n11782), .B(n11780), .C(n11778), .Y(
        n21019) );
  sky130_fd_sc_hd__nand3_1 U14239 ( .A(n20975), .B(n20974), .C(n21022), .Y(
        n21690) );
  sky130_fd_sc_hd__clkinv_1 U14240 ( .A(n16608), .Y(n16615) );
  sky130_fd_sc_hd__inv_2 U14241 ( .A(n28529), .Y(n11144) );
  sky130_fd_sc_hd__clkinv_1 U14243 ( .A(n26276), .Y(n28475) );
  sky130_fd_sc_hd__clkinv_1 U14245 ( .A(n20808), .Y(n20812) );
  sky130_fd_sc_hd__a21o_1 U14246 ( .A1(n13347), .A2(n26189), .B1(n29746), .X(
        n13362) );
  sky130_fd_sc_hd__clkinv_1 U14247 ( .A(n20593), .Y(n20594) );
  sky130_fd_sc_hd__clkinv_1 U14248 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_N423), .Y(n26466) );
  sky130_fd_sc_hd__inv_1 U14249 ( .A(n11598), .Y(n20415) );
  sky130_fd_sc_hd__clkinv_1 U14250 ( .A(n21454), .Y(n21450) );
  sky130_fd_sc_hd__clkinv_1 U14252 ( .A(n15422), .Y(n19480) );
  sky130_fd_sc_hd__clkinv_1 U14253 ( .A(n13239), .Y(n19773) );
  sky130_fd_sc_hd__buf_6 U14254 ( .A(n18340), .X(n11145) );
  sky130_fd_sc_hd__clkinv_1 U14255 ( .A(n20367), .Y(n20369) );
  sky130_fd_sc_hd__clkinv_1 U14256 ( .A(n15211), .Y(n15502) );
  sky130_fd_sc_hd__or2_0 U14257 ( .A(n29266), .B(n26662), .X(
        j202_soc_core_wbqspiflash_00_lldriver_N315) );
  sky130_fd_sc_hd__clkinv_1 U14258 ( .A(n17005), .Y(n17008) );
  sky130_fd_sc_hd__clkinv_1 U14259 ( .A(n16653), .Y(n16656) );
  sky130_fd_sc_hd__and4_1 U14260 ( .A(n14832), .B(n14831), .C(n14830), .D(
        n14829), .X(n14833) );
  sky130_fd_sc_hd__clkinv_1 U14261 ( .A(n17943), .Y(n17903) );
  sky130_fd_sc_hd__clkinv_1 U14262 ( .A(n19754), .Y(n19798) );
  sky130_fd_sc_hd__clkinv_1 U14263 ( .A(n27316), .Y(n23172) );
  sky130_fd_sc_hd__clkinv_1 U14264 ( .A(n19465), .Y(n19739) );
  sky130_fd_sc_hd__clkinv_1 U14265 ( .A(n20206), .Y(n20163) );
  sky130_fd_sc_hd__clkinv_1 U14266 ( .A(n19879), .Y(n19959) );
  sky130_fd_sc_hd__clkinv_1 U14267 ( .A(n20056), .Y(n20119) );
  sky130_fd_sc_hd__clkinv_1 U14268 ( .A(n20297), .Y(n20353) );
  sky130_fd_sc_hd__clkinv_1 U14269 ( .A(n19764), .Y(n13240) );
  sky130_fd_sc_hd__or2_0 U14270 ( .A(n25180), .B(n28203), .X(n28177) );
  sky130_fd_sc_hd__clkinv_1 U14271 ( .A(n20350), .Y(n20334) );
  sky130_fd_sc_hd__clkinv_1 U14272 ( .A(n20291), .Y(n19544) );
  sky130_fd_sc_hd__clkinv_1 U14273 ( .A(n15546), .Y(n15596) );
  sky130_fd_sc_hd__clkinv_1 U14274 ( .A(n20390), .Y(n19554) );
  sky130_fd_sc_hd__or2_0 U14275 ( .A(n18243), .B(n18244), .X(n11416) );
  sky130_fd_sc_hd__nor2_2 U14276 ( .A(n15195), .B(n15198), .Y(n21489) );
  sky130_fd_sc_hd__clkinv_1 U14277 ( .A(n15280), .Y(n15152) );
  sky130_fd_sc_hd__clkinv_1 U14278 ( .A(n23107), .Y(n23128) );
  sky130_fd_sc_hd__nor2_2 U14279 ( .A(n15193), .B(n15198), .Y(n21639) );
  sky130_fd_sc_hd__and4_1 U14280 ( .A(n15021), .B(n15020), .C(n15019), .D(
        n15018), .X(n15022) );
  sky130_fd_sc_hd__clkinv_1 U14281 ( .A(n17002), .Y(n16700) );
  sky130_fd_sc_hd__clkinv_1 U14282 ( .A(n23104), .Y(n27332) );
  sky130_fd_sc_hd__and4_1 U14283 ( .A(n15051), .B(n15050), .C(n15049), .D(
        n15048), .X(n15052) );
  sky130_fd_sc_hd__clkinv_1 U14284 ( .A(n20013), .Y(n20052) );
  sky130_fd_sc_hd__inv_2 U14285 ( .A(n13958), .Y(n11194) );
  sky130_fd_sc_hd__inv_2 U14286 ( .A(n14107), .Y(n11195) );
  sky130_fd_sc_hd__inv_2 U14287 ( .A(n13957), .Y(n11196) );
  sky130_fd_sc_hd__inv_2 U14288 ( .A(n14106), .Y(n11197) );
  sky130_fd_sc_hd__inv_2 U14289 ( .A(n13946), .Y(n11193) );
  sky130_fd_sc_hd__nand2_1 U14290 ( .A(n18678), .B(n18679), .Y(n12167) );
  sky130_fd_sc_hd__clkinv_1 U14292 ( .A(n20362), .Y(n20292) );
  sky130_fd_sc_hd__clkinv_1 U14293 ( .A(n15277), .Y(n15138) );
  sky130_fd_sc_hd__clkinv_1 U14294 ( .A(n19813), .Y(n19708) );
  sky130_fd_sc_hd__clkinv_1 U14295 ( .A(n19432), .Y(n13220) );
  sky130_fd_sc_hd__nor2_2 U14296 ( .A(n26264), .B(n26048), .Y(n26916) );
  sky130_fd_sc_hd__clkinv_1 U14297 ( .A(n21567), .Y(n21129) );
  sky130_fd_sc_hd__clkinv_1 U14298 ( .A(n15096), .Y(n15153) );
  sky130_fd_sc_hd__clkinv_1 U14299 ( .A(n19809), .Y(n13241) );
  sky130_fd_sc_hd__clkinv_1 U14300 ( .A(n20199), .Y(n20030) );
  sky130_fd_sc_hd__clkinv_1 U14301 ( .A(n18755), .Y(n19999) );
  sky130_fd_sc_hd__and2_1 U14302 ( .A(n18223), .B(n12891), .X(n12117) );
  sky130_fd_sc_hd__clkinv_1 U14303 ( .A(n20268), .Y(n19559) );
  sky130_fd_sc_hd__clkinv_1 U14304 ( .A(n20371), .Y(n19608) );
  sky130_fd_sc_hd__clkinv_1 U14305 ( .A(n18249), .Y(n11464) );
  sky130_fd_sc_hd__or2_0 U14306 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[6]), .B(n28650), .X(n28653)
         );
  sky130_fd_sc_hd__or2_0 U14307 ( .A(n17577), .B(n17576), .X(n17637) );
  sky130_fd_sc_hd__o22ai_1 U14308 ( .A1(n19002), .A2(n17636), .B1(n17593), 
        .B2(n11967), .Y(n17614) );
  sky130_fd_sc_hd__nor2_1 U14309 ( .A(n21022), .B(n11203), .Y(n11639) );
  sky130_fd_sc_hd__or2_0 U14310 ( .A(n17487), .B(n17486), .X(n17490) );
  sky130_fd_sc_hd__inv_2 U14311 ( .A(n23493), .Y(n11146) );
  sky130_fd_sc_hd__nor2_1 U14312 ( .A(n13171), .B(n13172), .Y(n20458) );
  sky130_fd_sc_hd__or2_0 U14313 ( .A(n17789), .B(n17788), .X(n17791) );
  sky130_fd_sc_hd__or2_0 U14314 ( .A(n28648), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[5]), .X(n28650) );
  sky130_fd_sc_hd__o22ai_1 U14315 ( .A1(n19002), .A2(n17564), .B1(n17518), 
        .B2(n11967), .Y(n17542) );
  sky130_fd_sc_hd__or2_0 U14316 ( .A(n17523), .B(n17522), .X(n17567) );
  sky130_fd_sc_hd__clkinv_1 U14317 ( .A(n18699), .Y(n19505) );
  sky130_fd_sc_hd__clkinv_1 U14318 ( .A(n14677), .Y(n14643) );
  sky130_fd_sc_hd__inv_1 U14319 ( .A(n18958), .Y(n17389) );
  sky130_fd_sc_hd__a21oi_1 U14320 ( .A1(n23103), .A2(n23102), .B1(n23101), .Y(
        n27329) );
  sky130_fd_sc_hd__clkinv_1 U14321 ( .A(n14612), .Y(n16764) );
  sky130_fd_sc_hd__inv_2 U14322 ( .A(n13707), .Y(n11199) );
  sky130_fd_sc_hd__inv_2 U14323 ( .A(n14001), .Y(n11200) );
  sky130_fd_sc_hd__clkinv_1 U14324 ( .A(n24799), .Y(n18193) );
  sky130_fd_sc_hd__inv_2 U14325 ( .A(n13537), .Y(n11148) );
  sky130_fd_sc_hd__clkinv_1 U14327 ( .A(n18250), .Y(n11463) );
  sky130_fd_sc_hd__clkinv_1 U14328 ( .A(n18695), .Y(n17104) );
  sky130_fd_sc_hd__or2_0 U14329 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[4]), .B(n28645), .X(n28648)
         );
  sky130_fd_sc_hd__or2_0 U14330 ( .A(n26907), .B(n26906), .X(n28254) );
  sky130_fd_sc_hd__clkinv_1 U14331 ( .A(n21919), .Y(n11204) );
  sky130_fd_sc_hd__clkinv_1 U14333 ( .A(n18713), .Y(n18727) );
  sky130_fd_sc_hd__clkinv_1 U14334 ( .A(n13429), .Y(n13430) );
  sky130_fd_sc_hd__clkinv_1 U14335 ( .A(n13203), .Y(n21360) );
  sky130_fd_sc_hd__clkinv_1 U14336 ( .A(n21022), .Y(n11207) );
  sky130_fd_sc_hd__clkinv_1 U14337 ( .A(n22229), .Y(n11205) );
  sky130_fd_sc_hd__or2_0 U14338 ( .A(n13259), .B(n13258), .X(n20580) );
  sky130_fd_sc_hd__nand2b_1 U14340 ( .A_N(n17964), .B(n24675), .Y(n18834) );
  sky130_fd_sc_hd__clkinv_1 U14341 ( .A(n20455), .Y(n15197) );
  sky130_fd_sc_hd__clkinv_1 U14342 ( .A(n17250), .Y(n15675) );
  sky130_fd_sc_hd__o22ai_1 U14343 ( .A1(n18209), .A2(n18082), .B1(n18208), 
        .B2(n18206), .Y(n11860) );
  sky130_fd_sc_hd__clkinv_1 U14344 ( .A(n13479), .Y(n13478) );
  sky130_fd_sc_hd__buf_4 U14345 ( .A(n17453), .X(n18027) );
  sky130_fd_sc_hd__clkinv_1 U14346 ( .A(n22114), .Y(n11149) );
  sky130_fd_sc_hd__or2_0 U14347 ( .A(j202_soc_core_qspi_wb_addr[12]), .B(
        n23702), .X(n23704) );
  sky130_fd_sc_hd__clkinv_1 U14348 ( .A(n22087), .Y(n17455) );
  sky130_fd_sc_hd__or2_0 U14349 ( .A(j202_soc_core_qspi_wb_addr[9]), .B(n23698), .X(n23699) );
  sky130_fd_sc_hd__or2_0 U14350 ( .A(j202_soc_core_qspi_wb_addr[10]), .B(
        n23695), .X(n23697) );
  sky130_fd_sc_hd__clkinv_1 U14351 ( .A(n13390), .Y(n13391) );
  sky130_fd_sc_hd__or2_0 U14352 ( .A(j202_soc_core_qspi_wb_addr[14]), .B(
        n23691), .X(n23692) );
  sky130_fd_sc_hd__or2_0 U14353 ( .A(j202_soc_core_qspi_wb_addr[13]), .B(
        n23688), .X(n23690) );
  sky130_fd_sc_hd__or2_0 U14354 ( .A(j202_soc_core_qspi_wb_addr[3]), .B(n23860), .X(n23680) );
  sky130_fd_sc_hd__or2_0 U14356 ( .A(j202_soc_core_qspi_wb_addr[4]), .B(n23679), .X(n23678) );
  sky130_fd_sc_hd__or2_0 U14357 ( .A(j202_soc_core_qspi_wb_addr[5]), .B(n23676), .X(n23668) );
  sky130_fd_sc_hd__or2_0 U14358 ( .A(j202_soc_core_qspi_wb_addr[6]), .B(n23666), .X(n23665) );
  sky130_fd_sc_hd__or2_0 U14359 ( .A(j202_soc_core_qspi_wb_addr[7]), .B(n23663), .X(n23660) );
  sky130_fd_sc_hd__or2_0 U14360 ( .A(j202_soc_core_qspi_wb_addr[8]), .B(n23657), .X(n23658) );
  sky130_fd_sc_hd__or2_0 U14361 ( .A(j202_soc_core_qspi_wb_addr[15]), .B(
        n23655), .X(n23656) );
  sky130_fd_sc_hd__or2_0 U14362 ( .A(j202_soc_core_qspi_wb_addr[17]), .B(
        n23652), .X(n23654) );
  sky130_fd_sc_hd__or2_0 U14363 ( .A(j202_soc_core_qspi_wb_addr[19]), .B(
        n23649), .X(n23651) );
  sky130_fd_sc_hd__or2_0 U14364 ( .A(j202_soc_core_qspi_wb_addr[21]), .B(
        n23647), .X(n23648) );
  sky130_fd_sc_hd__or2_0 U14365 ( .A(j202_soc_core_qspi_wb_addr[11]), .B(
        n23705), .X(n23706) );
  sky130_fd_sc_hd__or2_0 U14366 ( .A(j202_soc_core_qspi_wb_addr[16]), .B(
        n23717), .X(n23719) );
  sky130_fd_sc_hd__or2_0 U14367 ( .A(j202_soc_core_qspi_wb_addr[18]), .B(
        n23724), .X(n23726) );
  sky130_fd_sc_hd__or2_0 U14368 ( .A(j202_soc_core_qspi_wb_addr[22]), .B(
        n23738), .X(n23740) );
  sky130_fd_sc_hd__or2_0 U14369 ( .A(j202_soc_core_qspi_wb_addr[20]), .B(
        n23731), .X(n23733) );
  sky130_fd_sc_hd__inv_2 U14370 ( .A(n17094), .Y(n11208) );
  sky130_fd_sc_hd__clkinv_1 U14371 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[3]), .Y(n28044) );
  sky130_fd_sc_hd__or2_0 U14373 ( .A(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[0]), .B(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[1]), .X(n13270) );
  sky130_fd_sc_hd__clkinv_1 U14374 ( .A(j202_soc_core_j22_cpu_macop_MAC_[4]), 
        .Y(n27763) );
  sky130_fd_sc_hd__clkinv_1 U14375 ( .A(j202_soc_core_intc_core_00_rg_ipr[47]), 
        .Y(n26122) );
  sky130_fd_sc_hd__clkinv_1 U14376 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .Y(n23860) );
  sky130_fd_sc_hd__or2_0 U14377 ( .A(start_n_reg[1]), .B(wb_rst_i), .X(n470)
         );
  sky130_fd_sc_hd__buf_2 U14378 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .X(n13199) );
  sky130_fd_sc_hd__inv_2 U14379 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .Y(n14597) );
  sky130_fd_sc_hd__and2_1 U14380 ( .A(n12030), .B(n12036), .X(n13449) );
  sky130_fd_sc_hd__xnor2_1 U14383 ( .A(j202_soc_core_j22_cpu_ml_bufa[11]), .B(
        j202_soc_core_j22_cpu_ml_bufa[12]), .Y(n17453) );
  sky130_fd_sc_hd__inv_2 U14385 ( .A(n24517), .Y(n11151) );
  sky130_fd_sc_hd__buf_4 U14386 ( .A(n24360), .X(n28055) );
  sky130_fd_sc_hd__nand3_1 U14387 ( .A(n26872), .B(n22617), .C(n22616), .Y(
        n29519) );
  sky130_fd_sc_hd__inv_4 U14388 ( .A(n25475), .Y(n27643) );
  sky130_fd_sc_hd__and2_1 U14389 ( .A(n25475), .B(n27856), .X(n12135) );
  sky130_fd_sc_hd__and2_0 U14390 ( .A(n25246), .B(n27856), .X(n12134) );
  sky130_fd_sc_hd__and2_1 U14392 ( .A(n26454), .B(n27856), .X(n29635) );
  sky130_fd_sc_hd__nand2_2 U14394 ( .A(n29526), .B(n11853), .Y(n24515) );
  sky130_fd_sc_hd__inv_2 U14395 ( .A(n24307), .Y(n29873) );
  sky130_fd_sc_hd__and2_1 U14396 ( .A(n24861), .B(n27856), .X(n12131) );
  sky130_fd_sc_hd__and2_1 U14397 ( .A(n25135), .B(n27856), .X(n13102) );
  sky130_fd_sc_hd__buf_4 U14398 ( .A(n26023), .X(n12343) );
  sky130_fd_sc_hd__clkinv_1 U14399 ( .A(n24828), .Y(n24831) );
  sky130_fd_sc_hd__buf_2 U14400 ( .A(n26023), .X(n26669) );
  sky130_fd_sc_hd__and2_0 U14401 ( .A(n27916), .B(n27917), .X(n12155) );
  sky130_fd_sc_hd__buf_4 U14402 ( .A(n27460), .X(n12471) );
  sky130_fd_sc_hd__and2_1 U14403 ( .A(n25709), .B(n27856), .X(n13100) );
  sky130_fd_sc_hd__nand2_2 U14406 ( .A(n25659), .B(n25667), .Y(n25662) );
  sky130_fd_sc_hd__and2_0 U14407 ( .A(n30203), .B(n12127), .X(n29438) );
  sky130_fd_sc_hd__o211ai_1 U14410 ( .A1(n26396), .A2(n27669), .B1(n11467), 
        .C1(n11466), .Y(j202_soc_core_j22_cpu_rf_N2626) );
  sky130_fd_sc_hd__nor2_2 U14411 ( .A(n25903), .B(n25902), .Y(n28081) );
  sky130_fd_sc_hd__nand2_1 U14415 ( .A(n23548), .B(n28417), .Y(n25149) );
  sky130_fd_sc_hd__nand3_1 U14416 ( .A(n22826), .B(n22556), .C(n11484), .Y(
        n29515) );
  sky130_fd_sc_hd__a21oi_1 U14417 ( .A1(n27462), .A2(n27152), .B1(n12329), .Y(
        n27460) );
  sky130_fd_sc_hd__nand2_2 U14418 ( .A(n12358), .B(n30203), .Y(n12275) );
  sky130_fd_sc_hd__buf_4 U14419 ( .A(n24913), .X(n27162) );
  sky130_fd_sc_hd__clkinv_1 U14420 ( .A(n25379), .Y(n22313) );
  sky130_fd_sc_hd__nand3_1 U14422 ( .A(n18857), .B(n18856), .C(n22266), .Y(
        n11472) );
  sky130_fd_sc_hd__inv_1 U14423 ( .A(n25128), .Y(n25106) );
  sky130_fd_sc_hd__clkinv_1 U14424 ( .A(n25768), .Y(n25774) );
  sky130_fd_sc_hd__clkinv_1 U14425 ( .A(n25775), .Y(n25780) );
  sky130_fd_sc_hd__inv_2 U14426 ( .A(n13054), .Y(n11164) );
  sky130_fd_sc_hd__clkinv_1 U14427 ( .A(n24904), .Y(n24909) );
  sky130_fd_sc_hd__nand2_1 U14429 ( .A(n22347), .B(n22346), .Y(n25665) );
  sky130_fd_sc_hd__and2_0 U14430 ( .A(n22425), .B(n22424), .X(n11566) );
  sky130_fd_sc_hd__nor2_1 U14433 ( .A(n11605), .B(n11606), .Y(n11572) );
  sky130_fd_sc_hd__clkinv_1 U14434 ( .A(n25676), .Y(n25678) );
  sky130_fd_sc_hd__nand2_2 U14435 ( .A(n24699), .B(n28417), .Y(n24425) );
  sky130_fd_sc_hd__nor2_1 U14436 ( .A(n11632), .B(n11633), .Y(n11359) );
  sky130_fd_sc_hd__inv_1 U14437 ( .A(n23449), .Y(n11663) );
  sky130_fd_sc_hd__clkinv_1 U14438 ( .A(n25222), .Y(n22102) );
  sky130_fd_sc_hd__inv_1 U14439 ( .A(n23577), .Y(n23580) );
  sky130_fd_sc_hd__clkinv_1 U14440 ( .A(n27020), .Y(n27022) );
  sky130_fd_sc_hd__nor2_1 U14441 ( .A(n28140), .B(n12215), .Y(n27749) );
  sky130_fd_sc_hd__clkinv_1 U14442 ( .A(n11440), .Y(n11439) );
  sky130_fd_sc_hd__and2_1 U14444 ( .A(n27731), .B(n11395), .X(n12215) );
  sky130_fd_sc_hd__inv_2 U14445 ( .A(n23471), .Y(n23472) );
  sky130_fd_sc_hd__clkbuf_1 U14446 ( .A(n23470), .X(n23577) );
  sky130_fd_sc_hd__and2_0 U14447 ( .A(n28385), .B(n30189), .X(n12090) );
  sky130_fd_sc_hd__a21o_1 U14448 ( .A1(n21900), .A2(n23044), .B1(n21899), .X(
        n21901) );
  sky130_fd_sc_hd__inv_1 U14449 ( .A(n28088), .Y(n28099) );
  sky130_fd_sc_hd__nand3_1 U14450 ( .A(n12492), .B(n12491), .C(n12490), .Y(
        n23477) );
  sky130_fd_sc_hd__inv_1 U14451 ( .A(n28342), .Y(n24659) );
  sky130_fd_sc_hd__clkinv_1 U14452 ( .A(n25211), .Y(n25213) );
  sky130_fd_sc_hd__a22oi_1 U14453 ( .A1(j202_soc_core_j22_cpu_ml_mach[20]), 
        .A2(n23041), .B1(n22345), .B2(n24452), .Y(n22346) );
  sky130_fd_sc_hd__and2_0 U14455 ( .A(n23959), .B(n12821), .X(n12128) );
  sky130_fd_sc_hd__inv_1 U14456 ( .A(n24624), .Y(n28078) );
  sky130_fd_sc_hd__inv_1 U14457 ( .A(n12925), .Y(n11515) );
  sky130_fd_sc_hd__clkinv_1 U14458 ( .A(n29540), .Y(n24597) );
  sky130_fd_sc_hd__clkinv_1 U14459 ( .A(n12093), .Y(n24370) );
  sky130_fd_sc_hd__clkinv_1 U14460 ( .A(n25991), .Y(n21900) );
  sky130_fd_sc_hd__nor2_1 U14461 ( .A(n23993), .B(n12944), .Y(n28029) );
  sky130_fd_sc_hd__inv_2 U14462 ( .A(n23450), .Y(n11662) );
  sky130_fd_sc_hd__clkinv_1 U14464 ( .A(n12249), .Y(n27890) );
  sky130_fd_sc_hd__nand3_1 U14465 ( .A(n12250), .B(n11543), .C(n27729), .Y(
        n28140) );
  sky130_fd_sc_hd__o21a_1 U14466 ( .A1(n11444), .A2(n27990), .B1(n27989), .X(
        n11528) );
  sky130_fd_sc_hd__nor2_1 U14468 ( .A(n24692), .B(n24100), .Y(n24631) );
  sky130_fd_sc_hd__clkinv_1 U14469 ( .A(n22448), .Y(n22449) );
  sky130_fd_sc_hd__o211a_1 U14470 ( .A1(n30139), .A2(n12244), .B1(n28344), 
        .C1(n24561), .X(n24567) );
  sky130_fd_sc_hd__nor2_1 U14472 ( .A(n11544), .B(n11111), .Y(n11543) );
  sky130_fd_sc_hd__clkbuf_1 U14473 ( .A(n12453), .X(n12251) );
  sky130_fd_sc_hd__inv_1 U14474 ( .A(n24545), .Y(n23404) );
  sky130_fd_sc_hd__clkinv_1 U14475 ( .A(n24596), .Y(n11945) );
  sky130_fd_sc_hd__nand3_1 U14477 ( .A(n28259), .B(n28416), .C(n11994), .Y(
        n11732) );
  sky130_fd_sc_hd__inv_2 U14478 ( .A(n11866), .Y(n11171) );
  sky130_fd_sc_hd__inv_4 U14480 ( .A(n11553), .Y(n12349) );
  sky130_fd_sc_hd__inv_1 U14481 ( .A(n11647), .Y(n28117) );
  sky130_fd_sc_hd__clkinv_1 U14482 ( .A(n26415), .Y(n26404) );
  sky130_fd_sc_hd__clkinv_1 U14483 ( .A(n27981), .Y(n27982) );
  sky130_fd_sc_hd__nand2_1 U14484 ( .A(n21872), .B(n27355), .Y(n21873) );
  sky130_fd_sc_hd__clkbuf_1 U14486 ( .A(n11648), .X(n11647) );
  sky130_fd_sc_hd__inv_2 U14487 ( .A(n12063), .Y(n12064) );
  sky130_fd_sc_hd__clkinv_1 U14488 ( .A(n11669), .Y(n24552) );
  sky130_fd_sc_hd__nor2_1 U14489 ( .A(n24423), .B(n24422), .Y(n11672) );
  sky130_fd_sc_hd__and2_0 U14491 ( .A(n11927), .B(n24591), .X(n11926) );
  sky130_fd_sc_hd__nand2_1 U14492 ( .A(n12820), .B(n11719), .Y(n23615) );
  sky130_fd_sc_hd__clkinv_1 U14494 ( .A(n24115), .Y(n23458) );
  sky130_fd_sc_hd__inv_2 U14495 ( .A(n24406), .Y(n11546) );
  sky130_fd_sc_hd__a2bb2oi_1 U14497 ( .B1(n25138), .B2(n27862), .A1_N(n27774), 
        .A2_N(n28448), .Y(n25136) );
  sky130_fd_sc_hd__inv_1 U14498 ( .A(n27885), .Y(n11173) );
  sky130_fd_sc_hd__nand3_1 U14499 ( .A(n11658), .B(n11656), .C(n11141), .Y(
        n11655) );
  sky130_fd_sc_hd__clkinv_1 U14500 ( .A(n12221), .Y(n21973) );
  sky130_fd_sc_hd__nor2_1 U14501 ( .A(n16569), .B(n16568), .Y(n16570) );
  sky130_fd_sc_hd__nand2_1 U14502 ( .A(n21865), .B(n21864), .Y(n12352) );
  sky130_fd_sc_hd__inv_2 U14504 ( .A(n24607), .Y(n11841) );
  sky130_fd_sc_hd__and3_1 U14505 ( .A(n25368), .B(n25367), .C(n25366), .X(
        n25369) );
  sky130_fd_sc_hd__inv_2 U14506 ( .A(n12238), .Y(n11174) );
  sky130_fd_sc_hd__inv_1 U14508 ( .A(n17069), .Y(n20892) );
  sky130_fd_sc_hd__inv_2 U14510 ( .A(n11114), .Y(n28448) );
  sky130_fd_sc_hd__inv_2 U14513 ( .A(n27739), .Y(n11175) );
  sky130_fd_sc_hd__clkinv_1 U14514 ( .A(n23560), .Y(n23052) );
  sky130_fd_sc_hd__inv_2 U14515 ( .A(n12337), .Y(n12227) );
  sky130_fd_sc_hd__inv_2 U14516 ( .A(n29436), .Y(n20895) );
  sky130_fd_sc_hd__nand2_1 U14517 ( .A(n12730), .B(n19257), .Y(n19258) );
  sky130_fd_sc_hd__nand3_1 U14518 ( .A(n11815), .B(n11819), .C(n11810), .Y(
        n21936) );
  sky130_fd_sc_hd__o211ai_1 U14520 ( .A1(n26162), .A2(n27785), .B1(n11843), 
        .C1(n11842), .Y(n11844) );
  sky130_fd_sc_hd__inv_2 U14521 ( .A(n26185), .Y(n24294) );
  sky130_fd_sc_hd__inv_2 U14522 ( .A(n23401), .Y(n11176) );
  sky130_fd_sc_hd__inv_2 U14523 ( .A(n12524), .Y(n23444) );
  sky130_fd_sc_hd__inv_4 U14524 ( .A(n28525), .Y(n25765) );
  sky130_fd_sc_hd__clkbuf_1 U14525 ( .A(n19304), .X(n21272) );
  sky130_fd_sc_hd__nor2_1 U14526 ( .A(n18335), .B(n21271), .Y(n18336) );
  sky130_fd_sc_hd__clkinv_1 U14527 ( .A(n24959), .Y(n25901) );
  sky130_fd_sc_hd__clkinv_1 U14528 ( .A(n24382), .Y(n24385) );
  sky130_fd_sc_hd__inv_2 U14529 ( .A(n24633), .Y(n11177) );
  sky130_fd_sc_hd__inv_2 U14530 ( .A(n27728), .Y(n11178) );
  sky130_fd_sc_hd__clkinv_1 U14531 ( .A(n27740), .Y(n27741) );
  sky130_fd_sc_hd__inv_2 U14532 ( .A(n30139), .Y(n27900) );
  sky130_fd_sc_hd__inv_1 U14533 ( .A(n21271), .Y(n22958) );
  sky130_fd_sc_hd__clkinv_1 U14534 ( .A(n29482), .Y(n21040) );
  sky130_fd_sc_hd__o211ai_1 U14535 ( .A1(n27786), .A2(n28470), .B1(n27788), 
        .C1(n11500), .Y(n12182) );
  sky130_fd_sc_hd__nand3_1 U14536 ( .A(n11829), .B(n11828), .C(n11827), .Y(
        n28528) );
  sky130_fd_sc_hd__inv_2 U14537 ( .A(n29440), .Y(n17058) );
  sky130_fd_sc_hd__clkinv_1 U14539 ( .A(n28408), .Y(n28380) );
  sky130_fd_sc_hd__clkinv_1 U14540 ( .A(n25476), .Y(n25477) );
  sky130_fd_sc_hd__clkinv_1 U14541 ( .A(n29546), .Y(n24719) );
  sky130_fd_sc_hd__inv_2 U14542 ( .A(n26195), .Y(n18807) );
  sky130_fd_sc_hd__clkinv_1 U14543 ( .A(n29473), .Y(n23050) );
  sky130_fd_sc_hd__nand2_1 U14544 ( .A(n11139), .B(n26162), .Y(n28459) );
  sky130_fd_sc_hd__o22a_1 U14545 ( .A1(n21683), .A2(n21682), .B1(n10972), .B2(
        n11565), .X(n11564) );
  sky130_fd_sc_hd__nand2_1 U14546 ( .A(n12542), .B(n26171), .Y(n24358) );
  sky130_fd_sc_hd__nand2_1 U14547 ( .A(n11549), .B(n26187), .Y(n28466) );
  sky130_fd_sc_hd__buf_4 U14548 ( .A(n24680), .X(n11180) );
  sky130_fd_sc_hd__nand2b_1 U14549 ( .A_N(n25941), .B(n26175), .Y(n28483) );
  sky130_fd_sc_hd__clkinv_1 U14551 ( .A(n24376), .Y(n27344) );
  sky130_fd_sc_hd__inv_2 U14552 ( .A(n24165), .Y(n25209) );
  sky130_fd_sc_hd__clkinv_1 U14553 ( .A(n29549), .Y(n25052) );
  sky130_fd_sc_hd__and2_0 U14554 ( .A(n12393), .B(n29593), .X(n12136) );
  sky130_fd_sc_hd__clkinv_1 U14555 ( .A(n29581), .Y(n27919) );
  sky130_fd_sc_hd__clkinv_1 U14556 ( .A(n11816), .Y(n11828) );
  sky130_fd_sc_hd__nand3_1 U14557 ( .A(n15645), .B(n13065), .C(n15644), .Y(
        n29440) );
  sky130_fd_sc_hd__clkinv_1 U14558 ( .A(n26364), .Y(n26367) );
  sky130_fd_sc_hd__clkinv_1 U14559 ( .A(n23029), .Y(n22550) );
  sky130_fd_sc_hd__nand2_1 U14560 ( .A(n18801), .B(n18800), .Y(n26195) );
  sky130_fd_sc_hd__nor2_1 U14561 ( .A(n21752), .B(n22869), .Y(n18334) );
  sky130_fd_sc_hd__clkinv_1 U14562 ( .A(n28384), .Y(n17054) );
  sky130_fd_sc_hd__clkinv_1 U14565 ( .A(n22869), .Y(n22871) );
  sky130_fd_sc_hd__clkinv_1 U14567 ( .A(n17060), .Y(n16738) );
  sky130_fd_sc_hd__inv_1 U14568 ( .A(n21730), .Y(n22884) );
  sky130_fd_sc_hd__clkbuf_1 U14569 ( .A(n19106), .X(n21193) );
  sky130_fd_sc_hd__clkinv_1 U14571 ( .A(n26261), .Y(n26263) );
  sky130_fd_sc_hd__inv_1 U14572 ( .A(n23368), .Y(n23274) );
  sky130_fd_sc_hd__nand2_1 U14573 ( .A(n29439), .B(n25392), .Y(n18801) );
  sky130_fd_sc_hd__clkinv_1 U14574 ( .A(n21192), .Y(n22195) );
  sky130_fd_sc_hd__and3_1 U14575 ( .A(n11825), .B(n11823), .C(n11818), .X(
        n11817) );
  sky130_fd_sc_hd__clkinv_1 U14576 ( .A(n12409), .Y(n29846) );
  sky130_fd_sc_hd__clkinv_1 U14577 ( .A(n23349), .Y(n23351) );
  sky130_fd_sc_hd__nand3_1 U14578 ( .A(n11825), .B(n11823), .C(n11824), .Y(
        n11816) );
  sky130_fd_sc_hd__clkinv_1 U14579 ( .A(n24589), .Y(
        j202_soc_core_j22_cpu_ifetch) );
  sky130_fd_sc_hd__clkinv_1 U14582 ( .A(n22398), .Y(n22143) );
  sky130_fd_sc_hd__clkinv_1 U14583 ( .A(n17059), .Y(n16566) );
  sky130_fd_sc_hd__nand2_1 U14584 ( .A(n18658), .B(n21960), .Y(n21192) );
  sky130_fd_sc_hd__clkinv_1 U14585 ( .A(n22269), .Y(n22271) );
  sky130_fd_sc_hd__clkinv_1 U14586 ( .A(n27333), .Y(n24377) );
  sky130_fd_sc_hd__clkinv_1 U14587 ( .A(n21683), .Y(n11563) );
  sky130_fd_sc_hd__clkinv_1 U14588 ( .A(n12331), .Y(n22957) );
  sky130_fd_sc_hd__inv_4 U14589 ( .A(n29587), .Y(n11610) );
  sky130_fd_sc_hd__clkinv_1 U14590 ( .A(n22802), .Y(n22805) );
  sky130_fd_sc_hd__clkinv_1 U14591 ( .A(n26169), .Y(n29495) );
  sky130_fd_sc_hd__clkinv_1 U14592 ( .A(n12435), .Y(n21868) );
  sky130_fd_sc_hd__clkinv_1 U14593 ( .A(n22711), .Y(n22073) );
  sky130_fd_sc_hd__clkinv_1 U14594 ( .A(n22566), .Y(n18882) );
  sky130_fd_sc_hd__clkinv_1 U14595 ( .A(n27751), .Y(n27912) );
  sky130_fd_sc_hd__clkinv_1 U14597 ( .A(n28031), .Y(n24663) );
  sky130_fd_sc_hd__clkbuf_1 U14598 ( .A(n22956), .X(n12331) );
  sky130_fd_sc_hd__nor2_1 U14599 ( .A(n22783), .B(n22602), .Y(n19086) );
  sky130_fd_sc_hd__clkinv_1 U14600 ( .A(n22210), .Y(n21867) );
  sky130_fd_sc_hd__inv_1 U14601 ( .A(n22830), .Y(n22790) );
  sky130_fd_sc_hd__inv_2 U14602 ( .A(n24027), .Y(n29848) );
  sky130_fd_sc_hd__clkinv_1 U14603 ( .A(n22231), .Y(n22235) );
  sky130_fd_sc_hd__inv_2 U14604 ( .A(n26174), .Y(n24091) );
  sky130_fd_sc_hd__clkinv_1 U14606 ( .A(n24653), .Y(n28357) );
  sky130_fd_sc_hd__clkinv_1 U14607 ( .A(n22215), .Y(n22217) );
  sky130_fd_sc_hd__inv_2 U14608 ( .A(n20965), .Y(n21183) );
  sky130_fd_sc_hd__nand2b_1 U14609 ( .A_N(n25939), .B(n22114), .Y(n22116) );
  sky130_fd_sc_hd__inv_1 U14610 ( .A(n22562), .Y(n22564) );
  sky130_fd_sc_hd__clkinv_1 U14611 ( .A(n21904), .Y(n21263) );
  sky130_fd_sc_hd__nor2_1 U14612 ( .A(n22953), .B(n22962), .Y(n17868) );
  sky130_fd_sc_hd__o21ai_2 U14613 ( .A1(n23835), .A2(n23813), .B1(n27845), .Y(
        j202_soc_core_j22_cpu_rf_N2857) );
  sky130_fd_sc_hd__o21ai_2 U14614 ( .A1(n23835), .A2(n23818), .B1(n27843), .Y(
        j202_soc_core_j22_cpu_rf_N3005) );
  sky130_fd_sc_hd__clkinv_1 U14615 ( .A(n24960), .Y(n25147) );
  sky130_fd_sc_hd__o21ai_2 U14616 ( .A1(n23829), .A2(n23834), .B1(n27840), .Y(
        j202_soc_core_j22_cpu_rf_N2746) );
  sky130_fd_sc_hd__clkinv_1 U14617 ( .A(n28406), .Y(n28396) );
  sky130_fd_sc_hd__clkinv_1 U14618 ( .A(n22873), .Y(n22874) );
  sky130_fd_sc_hd__inv_2 U14619 ( .A(n22017), .Y(n22602) );
  sky130_fd_sc_hd__clkinv_1 U14620 ( .A(n24411), .Y(n24413) );
  sky130_fd_sc_hd__o21ai_2 U14621 ( .A1(n23813), .A2(n23829), .B1(n28061), .Y(
        j202_soc_core_j22_cpu_rf_N2894) );
  sky130_fd_sc_hd__clkbuf_1 U14622 ( .A(n25349), .X(n26190) );
  sky130_fd_sc_hd__o21ai_2 U14623 ( .A1(n23850), .A2(n23818), .B1(n27842), .Y(
        j202_soc_core_j22_cpu_rf_N3116) );
  sky130_fd_sc_hd__clkinv_1 U14624 ( .A(n27577), .Y(n27156) );
  sky130_fd_sc_hd__o21ai_2 U14625 ( .A1(n23801), .A2(n23834), .B1(n27846), .Y(
        j202_soc_core_j22_cpu_rf_N2783) );
  sky130_fd_sc_hd__inv_1 U14626 ( .A(n22207), .Y(n22208) );
  sky130_fd_sc_hd__o21ai_2 U14627 ( .A1(n23829), .A2(n23818), .B1(n27837), .Y(
        j202_soc_core_j22_cpu_rf_N3042) );
  sky130_fd_sc_hd__inv_2 U14628 ( .A(n22745), .Y(n22702) );
  sky130_fd_sc_hd__nor2_1 U14629 ( .A(n18325), .B(n18324), .Y(n22211) );
  sky130_fd_sc_hd__o21a_1 U14630 ( .A1(n22175), .A2(n22335), .B1(n22174), .X(
        n22176) );
  sky130_fd_sc_hd__clkinv_1 U14631 ( .A(n24090), .Y(n29845) );
  sky130_fd_sc_hd__o21ai_2 U14632 ( .A1(n23801), .A2(n23818), .B1(n27838), .Y(
        j202_soc_core_j22_cpu_rf_N3079) );
  sky130_fd_sc_hd__o21a_1 U14633 ( .A1(n21462), .A2(n21833), .B1(n21461), .X(
        n21486) );
  sky130_fd_sc_hd__clkinv_1 U14634 ( .A(n19303), .Y(n21275) );
  sky130_fd_sc_hd__inv_1 U14636 ( .A(n21268), .Y(n21270) );
  sky130_fd_sc_hd__o21ai_2 U14637 ( .A1(n23813), .A2(n23850), .B1(n27834), .Y(
        j202_soc_core_j22_cpu_rf_N2968) );
  sky130_fd_sc_hd__clkinv_1 U14638 ( .A(n21273), .Y(n21274) );
  sky130_fd_sc_hd__o21ai_2 U14639 ( .A1(n23849), .A2(n23801), .B1(n28112), .Y(
        j202_soc_core_j22_cpu_rf_N3227) );
  sky130_fd_sc_hd__clkinv_1 U14640 ( .A(n16924), .Y(n16928) );
  sky130_fd_sc_hd__o21ai_2 U14641 ( .A1(n23829), .A2(n23849), .B1(n27836), .Y(
        j202_soc_core_j22_cpu_rf_N3190) );
  sky130_fd_sc_hd__o21ai_2 U14642 ( .A1(n23813), .A2(n23801), .B1(n27839), .Y(
        j202_soc_core_j22_cpu_rf_N2931) );
  sky130_fd_sc_hd__clkinv_1 U14643 ( .A(n21752), .Y(n22875) );
  sky130_fd_sc_hd__inv_2 U14646 ( .A(n16557), .Y(n17040) );
  sky130_fd_sc_hd__o21ai_2 U14647 ( .A1(n23850), .A2(n23834), .B1(n27835), .Y(
        j202_soc_core_j22_cpu_rf_N2820) );
  sky130_fd_sc_hd__nand2_1 U14648 ( .A(n26164), .B(n22739), .Y(n17087) );
  sky130_fd_sc_hd__clkinv_1 U14650 ( .A(n29747), .Y(n24542) );
  sky130_fd_sc_hd__o21ai_2 U14651 ( .A1(n23835), .A2(n23849), .B1(n27844), .Y(
        j202_soc_core_j22_cpu_rf_N3153) );
  sky130_fd_sc_hd__a21oi_2 U14652 ( .A1(n19062), .A2(n19061), .B1(n19060), .Y(
        n22921) );
  sky130_fd_sc_hd__nand2_1 U14653 ( .A(n11588), .B(n20424), .Y(n11587) );
  sky130_fd_sc_hd__clkinv_1 U14654 ( .A(n28394), .Y(n28397) );
  sky130_fd_sc_hd__inv_1 U14657 ( .A(n22353), .Y(n22354) );
  sky130_fd_sc_hd__clkinv_1 U14659 ( .A(n21235), .Y(n21237) );
  sky130_fd_sc_hd__clkinv_1 U14660 ( .A(n27191), .Y(n26595) );
  sky130_fd_sc_hd__clkinv_1 U14662 ( .A(n27986), .Y(n28198) );
  sky130_fd_sc_hd__clkinv_1 U14663 ( .A(n12692), .Y(n22241) );
  sky130_fd_sc_hd__clkinv_1 U14664 ( .A(n27772), .Y(n26981) );
  sky130_fd_sc_hd__clkinv_1 U14665 ( .A(n21961), .Y(n21962) );
  sky130_fd_sc_hd__inv_1 U14666 ( .A(n21957), .Y(n21959) );
  sky130_fd_sc_hd__clkinv_1 U14667 ( .A(n21681), .Y(n21963) );
  sky130_fd_sc_hd__clkinv_1 U14668 ( .A(n28127), .Y(n23455) );
  sky130_fd_sc_hd__clkinv_1 U14669 ( .A(n28155), .Y(n24602) );
  sky130_fd_sc_hd__clkinv_1 U14670 ( .A(n26510), .Y(n26528) );
  sky130_fd_sc_hd__clkinv_1 U14671 ( .A(n28352), .Y(n28353) );
  sky130_fd_sc_hd__clkinv_1 U14672 ( .A(n28125), .Y(n24412) );
  sky130_fd_sc_hd__inv_1 U14673 ( .A(n21753), .Y(n21754) );
  sky130_fd_sc_hd__nor2_1 U14674 ( .A(n21460), .B(
        j202_soc_core_memory0_ram_dout0[484]), .Y(n21833) );
  sky130_fd_sc_hd__inv_2 U14675 ( .A(n22743), .Y(n22701) );
  sky130_fd_sc_hd__inv_1 U14676 ( .A(n20443), .Y(n21788) );
  sky130_fd_sc_hd__nor2_1 U14677 ( .A(n11686), .B(n11685), .Y(n11684) );
  sky130_fd_sc_hd__nand3_1 U14679 ( .A(n21649), .B(n21648), .C(n21647), .Y(
        n21920) );
  sky130_fd_sc_hd__clkinv_1 U14680 ( .A(j202_soc_core_j22_cpu_rf_N2627), .Y(
        n26865) );
  sky130_fd_sc_hd__nand3_2 U14681 ( .A(n13365), .B(n13379), .C(n13443), .Y(
        n14588) );
  sky130_fd_sc_hd__and2_1 U14682 ( .A(n29484), .B(n29746), .X(n29647) );
  sky130_fd_sc_hd__and2_0 U14683 ( .A(n21318), .B(n21919), .X(n12022) );
  sky130_fd_sc_hd__clkinv_1 U14684 ( .A(n27576), .Y(n27582) );
  sky130_fd_sc_hd__nand3_1 U14685 ( .A(n12882), .B(n11624), .C(n12883), .Y(
        n11622) );
  sky130_fd_sc_hd__clkinv_1 U14686 ( .A(n27580), .Y(n27154) );
  sky130_fd_sc_hd__clkinv_1 U14687 ( .A(n15635), .Y(n15638) );
  sky130_fd_sc_hd__xnor2_1 U14688 ( .A(n18450), .B(n13028), .Y(n18664) );
  sky130_fd_sc_hd__clkinv_1 U14689 ( .A(n15636), .Y(n15637) );
  sky130_fd_sc_hd__and2_0 U14690 ( .A(n13086), .B(n22105), .X(n12099) );
  sky130_fd_sc_hd__inv_1 U14691 ( .A(n11856), .Y(n21194) );
  sky130_fd_sc_hd__clkinv_1 U14692 ( .A(n29073), .Y(n26864) );
  sky130_fd_sc_hd__nor2_1 U14693 ( .A(n18286), .B(n18287), .Y(n22971) );
  sky130_fd_sc_hd__clkinv_1 U14694 ( .A(n21232), .Y(n21233) );
  sky130_fd_sc_hd__nor2_1 U14695 ( .A(n11704), .B(n11702), .Y(n11701) );
  sky130_fd_sc_hd__inv_1 U14696 ( .A(n19105), .Y(n21195) );
  sky130_fd_sc_hd__clkinv_1 U14697 ( .A(n27225), .Y(n26596) );
  sky130_fd_sc_hd__clkinv_1 U14699 ( .A(n21055), .Y(n16919) );
  sky130_fd_sc_hd__clkinv_1 U14700 ( .A(n29879), .Y(n24652) );
  sky130_fd_sc_hd__clkinv_1 U14701 ( .A(n19109), .Y(n21234) );
  sky130_fd_sc_hd__clkinv_1 U14702 ( .A(n16186), .Y(n16187) );
  sky130_fd_sc_hd__clkinv_1 U14703 ( .A(n24704), .Y(n24705) );
  sky130_fd_sc_hd__o21ai_2 U14704 ( .A1(j202_soc_core_j22_cpu_regop_M_Wm__1_), 
        .A2(n23839), .B1(n23749), .Y(j202_soc_core_j22_cpu_rf_N3301) );
  sky130_fd_sc_hd__and2_0 U14705 ( .A(n21001), .B(n21919), .X(n12110) );
  sky130_fd_sc_hd__clkinv_1 U14706 ( .A(n21969), .Y(n21971) );
  sky130_fd_sc_hd__clkinv_1 U14707 ( .A(n26164), .Y(n26172) );
  sky130_fd_sc_hd__clkinv_1 U14708 ( .A(n26860), .Y(n27578) );
  sky130_fd_sc_hd__clkinv_1 U14709 ( .A(n26177), .Y(n26182) );
  sky130_fd_sc_hd__clkinv_1 U14711 ( .A(n26554), .Y(n26556) );
  sky130_fd_sc_hd__clkinv_1 U14712 ( .A(n22108), .Y(n22110) );
  sky130_fd_sc_hd__clkinv_1 U14713 ( .A(n21974), .Y(n21685) );
  sky130_fd_sc_hd__nor2_1 U14714 ( .A(n17864), .B(n17863), .Y(n22962) );
  sky130_fd_sc_hd__clkinv_1 U14715 ( .A(n17848), .Y(n11434) );
  sky130_fd_sc_hd__xnor2_1 U14716 ( .A(n18448), .B(n18449), .Y(n13028) );
  sky130_fd_sc_hd__clkinv_1 U14717 ( .A(n28084), .Y(n28087) );
  sky130_fd_sc_hd__nand2_1 U14718 ( .A(n21440), .B(n21629), .Y(n21777) );
  sky130_fd_sc_hd__and3_1 U14719 ( .A(n15479), .B(n15470), .C(n15476), .X(
        n15471) );
  sky130_fd_sc_hd__inv_1 U14720 ( .A(n21285), .Y(n18263) );
  sky130_fd_sc_hd__and2_0 U14721 ( .A(n19852), .B(n21919), .X(n13083) );
  sky130_fd_sc_hd__inv_2 U14722 ( .A(n17440), .Y(n19061) );
  sky130_fd_sc_hd__clkinv_1 U14723 ( .A(n27753), .Y(n25812) );
  sky130_fd_sc_hd__clkinv_1 U14724 ( .A(n26934), .Y(n26046) );
  sky130_fd_sc_hd__clkinv_1 U14725 ( .A(n22541), .Y(n22546) );
  sky130_fd_sc_hd__inv_1 U14726 ( .A(n17222), .Y(n20435) );
  sky130_fd_sc_hd__clkinv_1 U14727 ( .A(n15380), .Y(n15488) );
  sky130_fd_sc_hd__clkinv_1 U14728 ( .A(n10603), .Y(n24028) );
  sky130_fd_sc_hd__nand2_1 U14729 ( .A(n28109), .B(n23755), .Y(n23826) );
  sky130_fd_sc_hd__clkinv_1 U14730 ( .A(n15620), .Y(n13008) );
  sky130_fd_sc_hd__nand2_1 U14731 ( .A(n28109), .B(n24305), .Y(n13364) );
  sky130_fd_sc_hd__nor2_1 U14732 ( .A(n15083), .B(n15380), .Y(n16545) );
  sky130_fd_sc_hd__nand2b_1 U14733 ( .A_N(n19851), .B(n23511), .Y(n11749) );
  sky130_fd_sc_hd__clkinv_1 U14734 ( .A(n23136), .Y(n23258) );
  sky130_fd_sc_hd__clkinv_1 U14735 ( .A(n24919), .Y(n24920) );
  sky130_fd_sc_hd__clkinv_1 U14736 ( .A(n21260), .Y(n19294) );
  sky130_fd_sc_hd__clkinv_1 U14738 ( .A(n26392), .Y(n26156) );
  sky130_fd_sc_hd__clkinv_1 U14739 ( .A(n24372), .Y(n24373) );
  sky130_fd_sc_hd__nor2_1 U14740 ( .A(n17828), .B(n11777), .Y(n18683) );
  sky130_fd_sc_hd__inv_1 U14741 ( .A(n23251), .Y(n23237) );
  sky130_fd_sc_hd__clkinv_1 U14742 ( .A(n23150), .Y(n23138) );
  sky130_fd_sc_hd__clkinv_1 U14743 ( .A(n22544), .Y(n22545) );
  sky130_fd_sc_hd__clkinv_1 U14744 ( .A(n23334), .Y(n23347) );
  sky130_fd_sc_hd__or2_1 U14745 ( .A(n21933), .B(n21934), .X(n11824) );
  sky130_fd_sc_hd__nand2_1 U14746 ( .A(n18332), .B(n18333), .Y(n22109) );
  sky130_fd_sc_hd__clkinv_1 U14747 ( .A(n18282), .Y(n11482) );
  sky130_fd_sc_hd__clkinv_1 U14748 ( .A(n23267), .Y(n23269) );
  sky130_fd_sc_hd__clkinv_1 U14749 ( .A(n23019), .Y(n19085) );
  sky130_fd_sc_hd__inv_1 U14750 ( .A(n21029), .Y(n14579) );
  sky130_fd_sc_hd__clkinv_1 U14751 ( .A(n20964), .Y(n20968) );
  sky130_fd_sc_hd__inv_1 U14752 ( .A(n21030), .Y(n14572) );
  sky130_fd_sc_hd__inv_1 U14753 ( .A(n21698), .Y(n21700) );
  sky130_fd_sc_hd__clkinv_1 U14754 ( .A(n26933), .Y(n24884) );
  sky130_fd_sc_hd__clkinv_1 U14755 ( .A(n16896), .Y(n16295) );
  sky130_fd_sc_hd__clkinv_1 U14756 ( .A(n25840), .Y(n25829) );
  sky130_fd_sc_hd__clkinv_1 U14757 ( .A(n25844), .Y(n25838) );
  sky130_fd_sc_hd__inv_1 U14758 ( .A(n23254), .Y(n23255) );
  sky130_fd_sc_hd__clkinv_1 U14759 ( .A(n19229), .Y(n19230) );
  sky130_fd_sc_hd__clkinv_1 U14760 ( .A(n27817), .Y(n27039) );
  sky130_fd_sc_hd__nor2_1 U14761 ( .A(n19067), .B(n19068), .Y(n21260) );
  sky130_fd_sc_hd__nand3_1 U14762 ( .A(n12023), .B(n22230), .C(n27785), .Y(
        n11819) );
  sky130_fd_sc_hd__inv_2 U14763 ( .A(n19278), .Y(n21283) );
  sky130_fd_sc_hd__nand2_1 U14764 ( .A(n18920), .B(n22784), .Y(n12108) );
  sky130_fd_sc_hd__clkinv_1 U14765 ( .A(n19425), .Y(n19413) );
  sky130_fd_sc_hd__clkinv_1 U14766 ( .A(n16892), .Y(n16296) );
  sky130_fd_sc_hd__clkinv_1 U14767 ( .A(n21902), .Y(n19073) );
  sky130_fd_sc_hd__clkinv_1 U14768 ( .A(n20966), .Y(n20967) );
  sky130_fd_sc_hd__clkinv_1 U14769 ( .A(n16720), .Y(n16722) );
  sky130_fd_sc_hd__inv_1 U14770 ( .A(n17213), .Y(n17215) );
  sky130_fd_sc_hd__clkinv_1 U14771 ( .A(n21341), .Y(n21344) );
  sky130_fd_sc_hd__nand2_1 U14772 ( .A(n12886), .B(n12885), .Y(n21286) );
  sky130_fd_sc_hd__inv_1 U14773 ( .A(n21342), .Y(n21343) );
  sky130_fd_sc_hd__clkinv_1 U14774 ( .A(n16893), .Y(n16894) );
  sky130_fd_sc_hd__clkinv_1 U14775 ( .A(n26936), .Y(n21949) );
  sky130_fd_sc_hd__inv_1 U14776 ( .A(n24392), .Y(n27341) );
  sky130_fd_sc_hd__inv_1 U14777 ( .A(n20984), .Y(n20986) );
  sky130_fd_sc_hd__clkinv_1 U14778 ( .A(n26089), .Y(n26087) );
  sky130_fd_sc_hd__clkinv_1 U14779 ( .A(n20938), .Y(n21181) );
  sky130_fd_sc_hd__clkinv_1 U14780 ( .A(n21785), .Y(n21786) );
  sky130_fd_sc_hd__clkinv_1 U14781 ( .A(n21032), .Y(n21034) );
  sky130_fd_sc_hd__and2_0 U14782 ( .A(n24392), .B(n29480), .X(n12157) );
  sky130_fd_sc_hd__o211a_2 U14783 ( .A1(n27616), .A2(n18843), .B1(n18842), 
        .C1(n18841), .X(n12116) );
  sky130_fd_sc_hd__clkinv_1 U14784 ( .A(n16723), .Y(n16091) );
  sky130_fd_sc_hd__inv_1 U14785 ( .A(n20995), .Y(n20983) );
  sky130_fd_sc_hd__clkinv_1 U14786 ( .A(n16299), .Y(n16895) );
  sky130_fd_sc_hd__clkinv_1 U14787 ( .A(n20982), .Y(n20996) );
  sky130_fd_sc_hd__inv_1 U14788 ( .A(n21663), .Y(n21665) );
  sky130_fd_sc_hd__inv_1 U14789 ( .A(n22880), .Y(n22882) );
  sky130_fd_sc_hd__nor2_1 U14790 ( .A(n15489), .B(n15384), .Y(n15181) );
  sky130_fd_sc_hd__clkinv_1 U14791 ( .A(n16730), .Y(n16732) );
  sky130_fd_sc_hd__clkinv_1 U14792 ( .A(n16901), .Y(n16903) );
  sky130_fd_sc_hd__inv_1 U14793 ( .A(n21789), .Y(n21791) );
  sky130_fd_sc_hd__clkinv_1 U14794 ( .A(n15896), .Y(n15263) );
  sky130_fd_sc_hd__clkinv_1 U14796 ( .A(n22689), .Y(n22690) );
  sky130_fd_sc_hd__clkinv_1 U14797 ( .A(n22753), .Y(n18816) );
  sky130_fd_sc_hd__clkinv_1 U14798 ( .A(n16013), .Y(n14816) );
  sky130_fd_sc_hd__clkinv_1 U14799 ( .A(n20710), .Y(n20711) );
  sky130_fd_sc_hd__clkinv_1 U14800 ( .A(n20963), .Y(n21009) );
  sky130_fd_sc_hd__clkinv_1 U14801 ( .A(n20442), .Y(n21787) );
  sky130_fd_sc_hd__clkinv_1 U14802 ( .A(n15384), .Y(n15386) );
  sky130_fd_sc_hd__clkinv_1 U14803 ( .A(n15639), .Y(n15641) );
  sky130_fd_sc_hd__clkinv_1 U14804 ( .A(n22831), .Y(n22045) );
  sky130_fd_sc_hd__clkinv_1 U14805 ( .A(n22885), .Y(n21731) );
  sky130_fd_sc_hd__clkinv_1 U14806 ( .A(n21007), .Y(n21008) );
  sky130_fd_sc_hd__clkinv_1 U14807 ( .A(n15184), .Y(n15186) );
  sky130_fd_sc_hd__clkinv_1 U14808 ( .A(n21180), .Y(n20939) );
  sky130_fd_sc_hd__clkinv_1 U14809 ( .A(n22592), .Y(n22049) );
  sky130_fd_sc_hd__inv_1 U14810 ( .A(n17219), .Y(n17221) );
  sky130_fd_sc_hd__xnor2_1 U14811 ( .A(n11957), .B(n17839), .Y(n17829) );
  sky130_fd_sc_hd__inv_1 U14812 ( .A(n21325), .Y(n21327) );
  sky130_fd_sc_hd__clkinv_1 U14813 ( .A(n21340), .Y(n22691) );
  sky130_fd_sc_hd__clkinv_1 U14814 ( .A(n17041), .Y(n17043) );
  sky130_fd_sc_hd__clkinv_1 U14816 ( .A(n21011), .Y(n21013) );
  sky130_fd_sc_hd__clkinv_1 U14817 ( .A(n17031), .Y(n17032) );
  sky130_fd_sc_hd__clkinv_1 U14818 ( .A(n20940), .Y(n20942) );
  sky130_fd_sc_hd__clkinv_1 U14819 ( .A(n16194), .Y(n17033) );
  sky130_fd_sc_hd__nand2b_1 U14820 ( .A_N(n27330), .B(n23127), .Y(n23130) );
  sky130_fd_sc_hd__clkinv_1 U14821 ( .A(n15069), .Y(n14585) );
  sky130_fd_sc_hd__clkinv_1 U14822 ( .A(n22928), .Y(n22495) );
  sky130_fd_sc_hd__clkinv_1 U14823 ( .A(n22618), .Y(n22502) );
  sky130_fd_sc_hd__clkinv_1 U14824 ( .A(n22620), .Y(n22503) );
  sky130_fd_sc_hd__nor2_1 U14825 ( .A(n18219), .B(n18220), .Y(n22880) );
  sky130_fd_sc_hd__clkinv_1 U14826 ( .A(n21702), .Y(n13867) );
  sky130_fd_sc_hd__clkinv_1 U14827 ( .A(n17849), .Y(n11433) );
  sky130_fd_sc_hd__clkinv_1 U14828 ( .A(n22621), .Y(n22540) );
  sky130_fd_sc_hd__or2_1 U14829 ( .A(n19083), .B(n19084), .X(n12098) );
  sky130_fd_sc_hd__xnor2_1 U14830 ( .A(n17840), .B(n17841), .Y(n11957) );
  sky130_fd_sc_hd__clkinv_1 U14831 ( .A(n17809), .Y(n17747) );
  sky130_fd_sc_hd__clkinv_1 U14832 ( .A(n23026), .Y(n23028) );
  sky130_fd_sc_hd__clkinv_1 U14833 ( .A(n22670), .Y(n22494) );
  sky130_fd_sc_hd__clkinv_1 U14834 ( .A(n22709), .Y(n22488) );
  sky130_fd_sc_hd__clkinv_1 U14835 ( .A(n22712), .Y(n22489) );
  sky130_fd_sc_hd__clkinv_1 U14836 ( .A(n23264), .Y(n23266) );
  sky130_fd_sc_hd__clkinv_1 U14837 ( .A(n22332), .Y(n22060) );
  sky130_fd_sc_hd__clkinv_1 U14838 ( .A(n23220), .Y(n23252) );
  sky130_fd_sc_hd__clkinv_1 U14839 ( .A(n22800), .Y(n22061) );
  sky130_fd_sc_hd__clkinv_1 U14840 ( .A(n22350), .Y(n22055) );
  sky130_fd_sc_hd__clkinv_1 U14841 ( .A(n22828), .Y(n22044) );
  sky130_fd_sc_hd__clkinv_1 U14842 ( .A(n22714), .Y(n22483) );
  sky130_fd_sc_hd__clkinv_1 U14843 ( .A(n22238), .Y(n22240) );
  sky130_fd_sc_hd__clkinv_1 U14844 ( .A(n21214), .Y(n21216) );
  sky130_fd_sc_hd__nor2_1 U14845 ( .A(n13931), .B(n13932), .Y(n21663) );
  sky130_fd_sc_hd__clkinv_1 U14846 ( .A(n22338), .Y(n22801) );
  sky130_fd_sc_hd__clkinv_1 U14847 ( .A(n15771), .Y(n15779) );
  sky130_fd_sc_hd__clkinv_1 U14848 ( .A(n17010), .Y(n17011) );
  sky130_fd_sc_hd__inv_1 U14849 ( .A(n18624), .Y(n11345) );
  sky130_fd_sc_hd__clkinv_1 U14850 ( .A(n22172), .Y(n22066) );
  sky130_fd_sc_hd__clkinv_1 U14851 ( .A(n22268), .Y(n22067) );
  sky130_fd_sc_hd__inv_1 U14852 ( .A(n18625), .Y(n11344) );
  sky130_fd_sc_hd__clkinv_1 U14853 ( .A(n17553), .Y(n17550) );
  sky130_fd_sc_hd__clkinv_1 U14854 ( .A(n25832), .Y(n25823) );
  sky130_fd_sc_hd__clkinv_1 U14855 ( .A(n25097), .Y(n25069) );
  sky130_fd_sc_hd__clkinv_1 U14856 ( .A(n27425), .Y(n27418) );
  sky130_fd_sc_hd__clkinv_1 U14857 ( .A(n25096), .Y(n24808) );
  sky130_fd_sc_hd__clkinv_1 U14858 ( .A(n28231), .Y(n25075) );
  sky130_fd_sc_hd__clkinv_1 U14859 ( .A(n26425), .Y(n24887) );
  sky130_fd_sc_hd__clkinv_1 U14860 ( .A(n26434), .Y(n26437) );
  sky130_fd_sc_hd__clkinv_1 U14861 ( .A(n26293), .Y(n26420) );
  sky130_fd_sc_hd__clkinv_1 U14862 ( .A(n23519), .Y(n23522) );
  sky130_fd_sc_hd__inv_1 U14863 ( .A(n19236), .Y(n12567) );
  sky130_fd_sc_hd__clkinv_1 U14864 ( .A(n22178), .Y(n11187) );
  sky130_fd_sc_hd__clkinv_1 U14865 ( .A(n26308), .Y(n24935) );
  sky130_fd_sc_hd__clkinv_1 U14866 ( .A(n26992), .Y(n24974) );
  sky130_fd_sc_hd__clkinv_1 U14867 ( .A(n18268), .Y(n11459) );
  sky130_fd_sc_hd__clkinv_1 U14868 ( .A(n26102), .Y(n26101) );
  sky130_fd_sc_hd__nor2_1 U14869 ( .A(n18141), .B(n18142), .Y(n21214) );
  sky130_fd_sc_hd__clkinv_1 U14870 ( .A(n17824), .Y(n11493) );
  sky130_fd_sc_hd__clkinv_1 U14871 ( .A(n18844), .Y(n18820) );
  sky130_fd_sc_hd__clkinv_1 U14872 ( .A(n23523), .Y(n18821) );
  sky130_fd_sc_hd__clkinv_1 U14873 ( .A(n27587), .Y(n24181) );
  sky130_fd_sc_hd__or2_1 U14874 ( .A(n18844), .B(n18845), .X(n25688) );
  sky130_fd_sc_hd__clkinv_1 U14875 ( .A(n22599), .Y(n22601) );
  sky130_fd_sc_hd__and2_0 U14876 ( .A(n12525), .B(n22260), .X(n12159) );
  sky130_fd_sc_hd__clkinv_1 U14877 ( .A(n28515), .Y(n26135) );
  sky130_fd_sc_hd__clkinv_1 U14878 ( .A(n20807), .Y(n20853) );
  sky130_fd_sc_hd__clkinv_1 U14879 ( .A(n22486), .Y(n22016) );
  sky130_fd_sc_hd__clkinv_1 U14880 ( .A(n28499), .Y(n26281) );
  sky130_fd_sc_hd__clkinv_1 U14881 ( .A(n13350), .Y(n13356) );
  sky130_fd_sc_hd__clkinv_1 U14882 ( .A(n22062), .Y(n22059) );
  sky130_fd_sc_hd__clkinv_1 U14883 ( .A(n28463), .Y(n27065) );
  sky130_fd_sc_hd__clkinv_1 U14884 ( .A(n25692), .Y(n28513) );
  sky130_fd_sc_hd__clkinv_1 U14885 ( .A(n28471), .Y(n27851) );
  sky130_fd_sc_hd__inv_1 U14886 ( .A(n27033), .Y(n26296) );
  sky130_fd_sc_hd__clkinv_1 U14887 ( .A(n24929), .Y(n28481) );
  sky130_fd_sc_hd__clkinv_1 U14888 ( .A(n27548), .Y(n26982) );
  sky130_fd_sc_hd__clkinv_1 U14889 ( .A(n26479), .Y(n26480) );
  sky130_fd_sc_hd__o211a_2 U14890 ( .A1(n19727), .A2(n19726), .B1(n19725), 
        .C1(n19724), .X(n19840) );
  sky130_fd_sc_hd__clkinv_1 U14891 ( .A(n22492), .Y(n22491) );
  sky130_fd_sc_hd__clkinv_1 U14892 ( .A(n28541), .Y(n26265) );
  sky130_fd_sc_hd__clkinv_1 U14893 ( .A(n25138), .Y(n25139) );
  sky130_fd_sc_hd__clkinv_1 U14894 ( .A(n28446), .Y(n26275) );
  sky130_fd_sc_hd__clkinv_1 U14895 ( .A(n22500), .Y(n22499) );
  sky130_fd_sc_hd__and2_0 U14896 ( .A(n26945), .B(n27785), .X(n24952) );
  sky130_fd_sc_hd__clkinv_1 U14897 ( .A(n22020), .Y(n22065) );
  sky130_fd_sc_hd__clkinv_1 U14898 ( .A(n28519), .Y(n26272) );
  sky130_fd_sc_hd__clkinv_1 U14899 ( .A(n28478), .Y(n26215) );
  sky130_fd_sc_hd__clkinv_1 U14900 ( .A(n22058), .Y(n22057) );
  sky130_fd_sc_hd__clkinv_1 U14901 ( .A(n22490), .Y(n22487) );
  sky130_fd_sc_hd__clkinv_1 U14902 ( .A(n22504), .Y(n22501) );
  sky130_fd_sc_hd__clkinv_1 U14903 ( .A(n22064), .Y(n22063) );
  sky130_fd_sc_hd__and2_0 U14904 ( .A(n22260), .B(n22230), .X(n22227) );
  sky130_fd_sc_hd__clkinv_1 U14905 ( .A(n25825), .Y(n28457) );
  sky130_fd_sc_hd__clkinv_1 U14906 ( .A(n25230), .Y(n28487) );
  sky130_fd_sc_hd__clkinv_1 U14907 ( .A(n28050), .Y(n28043) );
  sky130_fd_sc_hd__fa_1 U14908 ( .A(n18940), .B(n18939), .CIN(n18938), .COUT(
        n18954), .SUM(n19053) );
  sky130_fd_sc_hd__clkinv_1 U14909 ( .A(n24716), .Y(n23746) );
  sky130_fd_sc_hd__nand2_1 U14910 ( .A(n21019), .B(n11096), .Y(n11645) );
  sky130_fd_sc_hd__clkinv_1 U14911 ( .A(n28493), .Y(n26277) );
  sky130_fd_sc_hd__inv_1 U14912 ( .A(n26330), .Y(n26435) );
  sky130_fd_sc_hd__clkinv_1 U14913 ( .A(n22056), .Y(n22053) );
  sky130_fd_sc_hd__clkinv_1 U14914 ( .A(n22510), .Y(n22505) );
  sky130_fd_sc_hd__clkinv_1 U14915 ( .A(n28489), .Y(n26309) );
  sky130_fd_sc_hd__clkinv_1 U14916 ( .A(n25081), .Y(n25082) );
  sky130_fd_sc_hd__clkinv_1 U14917 ( .A(n29413), .Y(n29416) );
  sky130_fd_sc_hd__clkinv_1 U14918 ( .A(n25945), .Y(n26867) );
  sky130_fd_sc_hd__clkinv_1 U14919 ( .A(n16967), .Y(n16318) );
  sky130_fd_sc_hd__clkinv_1 U14920 ( .A(n15716), .Y(n15708) );
  sky130_fd_sc_hd__clkinv_1 U14921 ( .A(n25465), .Y(n25471) );
  sky130_fd_sc_hd__clkinv_1 U14922 ( .A(n22451), .Y(n22455) );
  sky130_fd_sc_hd__nand4_1 U14923 ( .A(n13963), .B(n13041), .C(n13040), .D(
        n13042), .Y(n26941) );
  sky130_fd_sc_hd__clkinv_1 U14924 ( .A(n27760), .Y(n27761) );
  sky130_fd_sc_hd__clkinv_1 U14925 ( .A(n22383), .Y(n22386) );
  sky130_fd_sc_hd__clkinv_1 U14926 ( .A(n22395), .Y(n22396) );
  sky130_fd_sc_hd__clkinv_1 U14927 ( .A(n26937), .Y(n28521) );
  sky130_fd_sc_hd__nand3_1 U14928 ( .A(n14785), .B(n14784), .C(n13094), .Y(
        n24929) );
  sky130_fd_sc_hd__clkinv_1 U14929 ( .A(n28728), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N392) );
  sky130_fd_sc_hd__clkinv_1 U14930 ( .A(n28740), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N393) );
  sky130_fd_sc_hd__clkinv_1 U14931 ( .A(n29142), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N394) );
  sky130_fd_sc_hd__nand3_1 U14932 ( .A(n14094), .B(n12095), .C(n14093), .Y(
        n26009) );
  sky130_fd_sc_hd__clkinv_1 U14933 ( .A(n22427), .Y(n22430) );
  sky130_fd_sc_hd__clkinv_1 U14934 ( .A(n21983), .Y(n21995) );
  sky130_fd_sc_hd__o2bb2ai_1 U14935 ( .B1(n22655), .B2(n18536), .A1_N(n25679), 
        .A2_N(j202_soc_core_j22_cpu_ml_mach[10]), .Y(n17598) );
  sky130_fd_sc_hd__clkinv_1 U14936 ( .A(n16701), .Y(n15748) );
  sky130_fd_sc_hd__clkinv_1 U14937 ( .A(n25171), .Y(n26097) );
  sky130_fd_sc_hd__clkinv_1 U14938 ( .A(n20308), .Y(n20299) );
  sky130_fd_sc_hd__nand3_1 U14939 ( .A(n13786), .B(n13785), .C(n13784), .Y(
        n28529) );
  sky130_fd_sc_hd__clkinv_1 U14940 ( .A(n28667), .Y(n28668) );
  sky130_fd_sc_hd__clkinv_1 U14941 ( .A(n16223), .Y(n14626) );
  sky130_fd_sc_hd__o21ai_0 U14942 ( .A1(n26939), .A2(n26937), .B1(n26919), .Y(
        n12158) );
  sky130_fd_sc_hd__clkinv_1 U14943 ( .A(n24588), .Y(n29882) );
  sky130_fd_sc_hd__clkinv_1 U14944 ( .A(n24931), .Y(n28484) );
  sky130_fd_sc_hd__inv_2 U14945 ( .A(n22260), .Y(n11189) );
  sky130_fd_sc_hd__clkinv_1 U14946 ( .A(n21366), .Y(n21408) );
  sky130_fd_sc_hd__clkinv_1 U14947 ( .A(n21611), .Y(n21352) );
  sky130_fd_sc_hd__clkinv_1 U14948 ( .A(n19979), .Y(n19953) );
  sky130_fd_sc_hd__o22ai_1 U14949 ( .A1(n24854), .A2(n18937), .B1(n22522), 
        .B2(n18536), .Y(n12683) );
  sky130_fd_sc_hd__nand3_2 U14950 ( .A(n13493), .B(n12097), .C(n13492), .Y(
        n27115) );
  sky130_fd_sc_hd__clkinv_1 U14951 ( .A(n10600), .Y(n28383) );
  sky130_fd_sc_hd__clkinv_1 U14952 ( .A(n16586), .Y(n16591) );
  sky130_fd_sc_hd__clkinv_1 U14953 ( .A(n19175), .Y(n19176) );
  sky130_fd_sc_hd__clkinv_1 U14954 ( .A(n25406), .Y(n27715) );
  sky130_fd_sc_hd__inv_2 U14955 ( .A(n26334), .Y(n11190) );
  sky130_fd_sc_hd__clkinv_1 U14956 ( .A(n27816), .Y(n28473) );
  sky130_fd_sc_hd__clkinv_1 U14957 ( .A(n21565), .Y(n21409) );
  sky130_fd_sc_hd__clkinv_1 U14958 ( .A(n25451), .Y(n28454) );
  sky130_fd_sc_hd__inv_1 U14959 ( .A(n25973), .Y(n28449) );
  sky130_fd_sc_hd__clkinv_1 U14960 ( .A(n26285), .Y(n28526) );
  sky130_fd_sc_hd__and4_1 U14961 ( .A(n23883), .B(n29746), .C(n15646), .D(
        n28367), .X(n13361) );
  sky130_fd_sc_hd__clkinv_1 U14962 ( .A(n20855), .Y(n20642) );
  sky130_fd_sc_hd__clkinv_1 U14963 ( .A(n20628), .Y(n20679) );
  sky130_fd_sc_hd__o31a_1 U14964 ( .A1(n20624), .A2(n20651), .A3(n20808), .B1(
        n20804), .X(n20855) );
  sky130_fd_sc_hd__nor2_1 U14965 ( .A(n11696), .B(n11691), .Y(n11690) );
  sky130_fd_sc_hd__clkinv_1 U14966 ( .A(n15737), .Y(n16644) );
  sky130_fd_sc_hd__clkinv_1 U14967 ( .A(n14888), .Y(n14897) );
  sky130_fd_sc_hd__clkinv_1 U14968 ( .A(n20294), .Y(n19557) );
  sky130_fd_sc_hd__clkinv_1 U14969 ( .A(n28698), .Y(n24280) );
  sky130_fd_sc_hd__clkinv_1 U14970 ( .A(n26104), .Y(n26095) );
  sky130_fd_sc_hd__clkinv_1 U14971 ( .A(n20246), .Y(n20247) );
  sky130_fd_sc_hd__clkinv_1 U14972 ( .A(n25013), .Y(n27480) );
  sky130_fd_sc_hd__clkinv_1 U14973 ( .A(n24532), .Y(n24529) );
  sky130_fd_sc_hd__clkinv_1 U14974 ( .A(n28548), .Y(n24538) );
  sky130_fd_sc_hd__clkinv_1 U14975 ( .A(n27471), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[1]) );
  sky130_fd_sc_hd__clkinv_1 U14976 ( .A(n16225), .Y(n16231) );
  sky130_fd_sc_hd__clkinv_1 U14977 ( .A(n13612), .Y(n13613) );
  sky130_fd_sc_hd__nor2_1 U14978 ( .A(n11626), .B(n11625), .Y(n11624) );
  sky130_fd_sc_hd__clkinv_1 U14979 ( .A(n24862), .Y(n24863) );
  sky130_fd_sc_hd__clkinv_1 U14981 ( .A(n16227), .Y(n16228) );
  sky130_fd_sc_hd__clkinv_1 U14982 ( .A(n21549), .Y(n21560) );
  sky130_fd_sc_hd__clkinv_1 U14983 ( .A(n26651), .Y(n23639) );
  sky130_fd_sc_hd__clkinv_1 U14984 ( .A(n20022), .Y(n20027) );
  sky130_fd_sc_hd__clkinv_1 U14985 ( .A(n16657), .Y(n16658) );
  sky130_fd_sc_hd__clkinv_1 U14986 ( .A(n20789), .Y(n20661) );
  sky130_fd_sc_hd__clkinv_1 U14987 ( .A(n29746), .Y(n28275) );
  sky130_fd_sc_hd__clkinv_1 U14988 ( .A(n20136), .Y(n19997) );
  sky130_fd_sc_hd__clkinv_1 U14989 ( .A(n20763), .Y(n20535) );
  sky130_fd_sc_hd__clkinv_1 U14990 ( .A(n19759), .Y(n15391) );
  sky130_fd_sc_hd__clkinv_1 U14991 ( .A(n15476), .Y(n15477) );
  sky130_fd_sc_hd__clkinv_1 U14992 ( .A(n17326), .Y(n17327) );
  sky130_fd_sc_hd__clkinv_1 U14993 ( .A(n17047), .Y(n25862) );
  sky130_fd_sc_hd__clkinv_1 U14994 ( .A(n25247), .Y(n25250) );
  sky130_fd_sc_hd__clkinv_1 U14995 ( .A(n17210), .Y(n17211) );
  sky130_fd_sc_hd__clkinv_1 U14996 ( .A(n16772), .Y(n16773) );
  sky130_fd_sc_hd__clkinv_1 U14997 ( .A(n11626), .Y(n19220) );
  sky130_fd_sc_hd__clkinv_1 U14998 ( .A(n19519), .Y(n19474) );
  sky130_fd_sc_hd__clkinv_1 U14999 ( .A(n24673), .Y(n23892) );
  sky130_fd_sc_hd__clkinv_1 U15000 ( .A(n20053), .Y(n20209) );
  sky130_fd_sc_hd__clkinv_1 U15001 ( .A(n24764), .Y(n25439) );
  sky130_fd_sc_hd__clkinv_1 U15002 ( .A(n16976), .Y(n16979) );
  sky130_fd_sc_hd__clkinv_1 U15003 ( .A(n19576), .Y(n19552) );
  sky130_fd_sc_hd__clkinv_1 U15004 ( .A(n21827), .Y(n21830) );
  sky130_fd_sc_hd__nand2_1 U15005 ( .A(n24673), .B(n23753), .Y(n13308) );
  sky130_fd_sc_hd__a21oi_2 U15006 ( .A1(n22777), .A2(n16523), .B1(n14541), .Y(
        n28532) );
  sky130_fd_sc_hd__clkinv_1 U15007 ( .A(n18788), .Y(n18789) );
  sky130_fd_sc_hd__clkinv_1 U15008 ( .A(n16786), .Y(n16817) );
  sky130_fd_sc_hd__clkinv_1 U15009 ( .A(n20332), .Y(n20337) );
  sky130_fd_sc_hd__or2_0 U15010 ( .A(n26783), .B(n23632), .X(n12085) );
  sky130_fd_sc_hd__clkinv_1 U15011 ( .A(n16944), .Y(n16947) );
  sky130_fd_sc_hd__clkinv_1 U15012 ( .A(n15730), .Y(n16314) );
  sky130_fd_sc_hd__clkinv_1 U15013 ( .A(n17134), .Y(n17135) );
  sky130_fd_sc_hd__nand3_1 U15014 ( .A(n11986), .B(n11984), .C(n11983), .Y(
        n24673) );
  sky130_fd_sc_hd__clkinv_1 U15015 ( .A(n15275), .Y(n15100) );
  sky130_fd_sc_hd__nand4_1 U15016 ( .A(n20264), .B(n20265), .C(n20263), .D(
        n20260), .Y(n11589) );
  sky130_fd_sc_hd__inv_1 U15017 ( .A(n17446), .Y(n18340) );
  sky130_fd_sc_hd__clkinv_1 U15018 ( .A(n28884), .Y(n28885) );
  sky130_fd_sc_hd__clkinv_1 U15019 ( .A(n20146), .Y(n19892) );
  sky130_fd_sc_hd__clkinv_1 U15020 ( .A(n21599), .Y(n21423) );
  sky130_fd_sc_hd__clkinv_1 U15021 ( .A(n21821), .Y(n19924) );
  sky130_fd_sc_hd__clkinv_1 U15022 ( .A(n21414), .Y(n21418) );
  sky130_fd_sc_hd__clkinv_1 U15023 ( .A(n27764), .Y(n27382) );
  sky130_fd_sc_hd__clkinv_1 U15024 ( .A(n20219), .Y(n20202) );
  sky130_fd_sc_hd__clkinv_1 U15025 ( .A(n17155), .Y(n19371) );
  sky130_fd_sc_hd__clkinv_1 U15026 ( .A(n13856), .Y(n13857) );
  sky130_fd_sc_hd__clkinv_1 U15027 ( .A(n21605), .Y(n21608) );
  sky130_fd_sc_hd__clkinv_1 U15028 ( .A(n19373), .Y(n19564) );
  sky130_fd_sc_hd__clkinv_1 U15029 ( .A(n13205), .Y(n19517) );
  sky130_fd_sc_hd__clkinv_1 U15030 ( .A(n19516), .Y(n13188) );
  sky130_fd_sc_hd__clkinv_1 U15031 ( .A(n20777), .Y(n20529) );
  sky130_fd_sc_hd__clkinv_1 U15032 ( .A(n20844), .Y(n20525) );
  sky130_fd_sc_hd__clkinv_1 U15033 ( .A(n19666), .Y(n19669) );
  sky130_fd_sc_hd__clkinv_1 U15034 ( .A(n19683), .Y(n19684) );
  sky130_fd_sc_hd__clkinv_1 U15035 ( .A(n14383), .Y(n14384) );
  sky130_fd_sc_hd__clkinv_1 U15036 ( .A(n20595), .Y(n20471) );
  sky130_fd_sc_hd__clkinv_1 U15037 ( .A(n20019), .Y(n20028) );
  sky130_fd_sc_hd__nand3_1 U15038 ( .A(n12634), .B(n29883), .C(n29884), .Y(
        n21021) );
  sky130_fd_sc_hd__clkinv_1 U15039 ( .A(n21552), .Y(n21538) );
  sky130_fd_sc_hd__nand3_1 U15040 ( .A(n24852), .B(n18834), .C(n11146), .Y(
        n24764) );
  sky130_fd_sc_hd__clkinv_1 U15041 ( .A(n13243), .Y(n13244) );
  sky130_fd_sc_hd__clkinv_1 U15042 ( .A(n21562), .Y(n21564) );
  sky130_fd_sc_hd__clkinv_1 U15044 ( .A(n15430), .Y(n13236) );
  sky130_fd_sc_hd__o211a_2 U15045 ( .A1(n13641), .A2(n16444), .B1(n13540), 
        .C1(n13539), .X(n13541) );
  sky130_fd_sc_hd__inv_1 U15046 ( .A(n19698), .Y(n19720) );
  sky130_fd_sc_hd__clkinv_1 U15047 ( .A(n20744), .Y(n19147) );
  sky130_fd_sc_hd__clkinv_1 U15048 ( .A(n28742), .Y(n10572) );
  sky130_fd_sc_hd__clkinv_1 U15049 ( .A(n20601), .Y(n19204) );
  sky130_fd_sc_hd__clkinv_1 U15050 ( .A(n16788), .Y(n16794) );
  sky130_fd_sc_hd__clkinv_1 U15051 ( .A(n21522), .Y(n21410) );
  sky130_fd_sc_hd__clkinv_1 U15052 ( .A(n25666), .Y(n25672) );
  sky130_fd_sc_hd__clkinv_1 U15053 ( .A(n18004), .Y(n11506) );
  sky130_fd_sc_hd__clkinv_1 U15054 ( .A(n17206), .Y(n17209) );
  sky130_fd_sc_hd__clkinv_1 U15055 ( .A(n28733), .Y(n10571) );
  sky130_fd_sc_hd__clkinv_1 U15056 ( .A(n28741), .Y(n10569) );
  sky130_fd_sc_hd__clkinv_1 U15057 ( .A(n20327), .Y(n17103) );
  sky130_fd_sc_hd__nand4_1 U15058 ( .A(n19216), .B(n19217), .C(n19218), .D(
        n19219), .Y(n11625) );
  sky130_fd_sc_hd__clkinv_1 U15059 ( .A(n19664), .Y(n20335) );
  sky130_fd_sc_hd__clkinv_1 U15060 ( .A(n19732), .Y(n19736) );
  sky130_fd_sc_hd__clkinv_1 U15061 ( .A(n20737), .Y(n20608) );
  sky130_fd_sc_hd__clkinv_1 U15062 ( .A(n19511), .Y(n19746) );
  sky130_fd_sc_hd__clkinv_1 U15063 ( .A(n19761), .Y(n19762) );
  sky130_fd_sc_hd__clkinv_1 U15064 ( .A(n20663), .Y(n20819) );
  sky130_fd_sc_hd__clkinv_1 U15066 ( .A(n24535), .Y(n24534) );
  sky130_fd_sc_hd__clkinv_1 U15067 ( .A(n16609), .Y(n16614) );
  sky130_fd_sc_hd__clkinv_1 U15068 ( .A(n23238), .Y(n23239) );
  sky130_fd_sc_hd__clkinv_1 U15069 ( .A(n16696), .Y(n16308) );
  sky130_fd_sc_hd__clkinv_1 U15070 ( .A(n15533), .Y(n15588) );
  sky130_fd_sc_hd__clkinv_1 U15071 ( .A(n16689), .Y(n15758) );
  sky130_fd_sc_hd__clkinv_1 U15072 ( .A(n15424), .Y(n19774) );
  sky130_fd_sc_hd__clkinv_1 U15073 ( .A(n16814), .Y(n14649) );
  sky130_fd_sc_hd__and2_0 U15074 ( .A(n16689), .B(n16959), .X(n16690) );
  sky130_fd_sc_hd__clkinv_1 U15075 ( .A(n15526), .Y(n15319) );
  sky130_fd_sc_hd__clkinv_1 U15076 ( .A(n18785), .Y(n18787) );
  sky130_fd_sc_hd__clkinv_1 U15077 ( .A(n16191), .Y(n27064) );
  sky130_fd_sc_hd__clkinv_1 U15078 ( .A(n15329), .Y(n15498) );
  sky130_fd_sc_hd__clkinv_1 U15079 ( .A(n26662), .Y(n26663) );
  sky130_fd_sc_hd__clkinv_1 U15080 ( .A(n24651), .Y(n28346) );
  sky130_fd_sc_hd__clkinv_1 U15081 ( .A(n20221), .Y(n20185) );
  sky130_fd_sc_hd__clkinv_1 U15082 ( .A(n23242), .Y(n23244) );
  sky130_fd_sc_hd__clkinv_1 U15083 ( .A(n26497), .Y(n26499) );
  sky130_fd_sc_hd__clkinv_1 U15084 ( .A(n16162), .Y(n16163) );
  sky130_fd_sc_hd__clkinv_1 U15085 ( .A(n23133), .Y(n23135) );
  sky130_fd_sc_hd__clkinv_1 U15086 ( .A(n23227), .Y(n23229) );
  sky130_fd_sc_hd__inv_1 U15087 ( .A(n23224), .Y(n23226) );
  sky130_fd_sc_hd__clkinv_1 U15088 ( .A(n25595), .Y(n25599) );
  sky130_fd_sc_hd__clkinv_1 U15089 ( .A(n16969), .Y(n16645) );
  sky130_fd_sc_hd__clkinv_1 U15090 ( .A(n15472), .Y(n15475) );
  sky130_fd_sc_hd__clkinv_1 U15091 ( .A(n23319), .Y(n23320) );
  sky130_fd_sc_hd__clkinv_1 U15092 ( .A(n23328), .Y(n23329) );
  sky130_fd_sc_hd__clkinv_1 U15094 ( .A(n15393), .Y(n15395) );
  sky130_fd_sc_hd__clkinv_1 U15095 ( .A(n23142), .Y(n23144) );
  sky130_fd_sc_hd__clkinv_1 U15096 ( .A(n16697), .Y(n16651) );
  sky130_fd_sc_hd__clkinv_1 U15097 ( .A(n16575), .Y(n16311) );
  sky130_fd_sc_hd__clkinv_1 U15098 ( .A(n15495), .Y(n15117) );
  sky130_fd_sc_hd__clkinv_1 U15099 ( .A(n21139), .Y(n21085) );
  sky130_fd_sc_hd__clkinv_1 U15100 ( .A(n20242), .Y(n20245) );
  sky130_fd_sc_hd__clkinv_1 U15101 ( .A(n19482), .Y(n19472) );
  sky130_fd_sc_hd__clkinv_1 U15102 ( .A(n20474), .Y(n20843) );
  sky130_fd_sc_hd__clkinv_1 U15103 ( .A(n25710), .Y(n25713) );
  sky130_fd_sc_hd__clkinv_1 U15104 ( .A(n15293), .Y(n15228) );
  sky130_fd_sc_hd__clkinv_1 U15105 ( .A(n21593), .Y(n21600) );
  sky130_fd_sc_hd__clkinv_1 U15106 ( .A(n19797), .Y(n19802) );
  sky130_fd_sc_hd__clkinv_1 U15107 ( .A(n16804), .Y(n16215) );
  sky130_fd_sc_hd__clkinv_1 U15108 ( .A(n19699), .Y(n19744) );
  sky130_fd_sc_hd__clkinv_1 U15109 ( .A(n15774), .Y(n15775) );
  sky130_fd_sc_hd__clkinv_1 U15110 ( .A(n19881), .Y(n19882) );
  sky130_fd_sc_hd__clkinv_1 U15111 ( .A(n26455), .Y(n26459) );
  sky130_fd_sc_hd__clkinv_1 U15112 ( .A(n20653), .Y(n20654) );
  sky130_fd_sc_hd__or2_0 U15113 ( .A(n29184), .B(n29263), .X(
        j202_soc_core_wbqspiflash_00_lldriver_N356) );
  sky130_fd_sc_hd__clkinv_1 U15114 ( .A(n19344), .Y(n20271) );
  sky130_fd_sc_hd__clkinv_1 U15115 ( .A(n19340), .Y(n19558) );
  sky130_fd_sc_hd__clkinv_1 U15116 ( .A(n19807), .Y(n19808) );
  sky130_fd_sc_hd__clkinv_1 U15118 ( .A(n19970), .Y(n20120) );
  sky130_fd_sc_hd__clkinv_1 U15119 ( .A(n19821), .Y(n19822) );
  sky130_fd_sc_hd__clkinv_1 U15120 ( .A(n16686), .Y(n16375) );
  sky130_fd_sc_hd__clkinv_1 U15121 ( .A(n23231), .Y(n23233) );
  sky130_fd_sc_hd__clkinv_1 U15122 ( .A(n16672), .Y(n16603) );
  sky130_fd_sc_hd__clkinv_1 U15123 ( .A(n21384), .Y(n21076) );
  sky130_fd_sc_hd__clkinv_1 U15125 ( .A(n20015), .Y(n19889) );
  sky130_fd_sc_hd__clkinv_1 U15126 ( .A(n15699), .Y(n16335) );
  sky130_fd_sc_hd__clkinv_1 U15127 ( .A(n16183), .Y(n16184) );
  sky130_fd_sc_hd__o22ai_1 U15128 ( .A1(n11464), .A2(n11463), .B1(n11462), 
        .B2(n11461), .Y(n18277) );
  sky130_fd_sc_hd__clkinv_1 U15129 ( .A(n16983), .Y(n16984) );
  sky130_fd_sc_hd__clkinv_1 U15130 ( .A(n20923), .Y(n20924) );
  sky130_fd_sc_hd__clkinv_1 U15131 ( .A(n21124), .Y(n17290) );
  sky130_fd_sc_hd__clkinv_1 U15132 ( .A(n19955), .Y(n20021) );
  sky130_fd_sc_hd__clkinv_1 U15133 ( .A(n20633), .Y(n19162) );
  sky130_fd_sc_hd__clkinv_1 U15134 ( .A(n20645), .Y(n20802) );
  sky130_fd_sc_hd__clkinv_1 U15135 ( .A(n20612), .Y(n20665) );
  sky130_fd_sc_hd__clkinv_1 U15136 ( .A(n27469), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[0]) );
  sky130_fd_sc_hd__clkinv_1 U15137 ( .A(n28583), .Y(n29171) );
  sky130_fd_sc_hd__clkinv_1 U15138 ( .A(n16576), .Y(n15755) );
  sky130_fd_sc_hd__clkinv_1 U15139 ( .A(n19600), .Y(n19601) );
  sky130_fd_sc_hd__clkinv_1 U15140 ( .A(n17282), .Y(n21413) );
  sky130_fd_sc_hd__clkinv_1 U15141 ( .A(n20683), .Y(n20607) );
  sky130_fd_sc_hd__clkinv_1 U15142 ( .A(n19943), .Y(n18765) );
  sky130_fd_sc_hd__clkinv_1 U15143 ( .A(n16842), .Y(n16844) );
  sky130_fd_sc_hd__clkinv_1 U15144 ( .A(n16687), .Y(n16683) );
  sky130_fd_sc_hd__clkinv_1 U15145 ( .A(n16826), .Y(n16790) );
  sky130_fd_sc_hd__clkinv_1 U15146 ( .A(n28654), .Y(n28661) );
  sky130_fd_sc_hd__clkinv_1 U15147 ( .A(n16831), .Y(n14641) );
  sky130_fd_sc_hd__clkinv_1 U15148 ( .A(n20037), .Y(n20039) );
  sky130_fd_sc_hd__clkinv_1 U15149 ( .A(n16987), .Y(n16599) );
  sky130_fd_sc_hd__clkinv_1 U15150 ( .A(n23318), .Y(n23322) );
  sky130_fd_sc_hd__clkinv_1 U15151 ( .A(n14703), .Y(n14700) );
  sky130_fd_sc_hd__clkinv_1 U15152 ( .A(n25971), .Y(n25972) );
  sky130_fd_sc_hd__clkinv_1 U15153 ( .A(n20344), .Y(n19613) );
  sky130_fd_sc_hd__clkinv_1 U15154 ( .A(n19398), .Y(n17158) );
  sky130_fd_sc_hd__clkinv_1 U15155 ( .A(n20769), .Y(n20519) );
  sky130_fd_sc_hd__clkinv_1 U15156 ( .A(n27863), .Y(n27849) );
  sky130_fd_sc_hd__clkinv_1 U15158 ( .A(n25896), .Y(n25897) );
  sky130_fd_sc_hd__clkinv_1 U15159 ( .A(n20220), .Y(n20107) );
  sky130_fd_sc_hd__clkinv_1 U15160 ( .A(n20774), .Y(n20483) );
  sky130_fd_sc_hd__clkinv_1 U15161 ( .A(n28696), .Y(n28697) );
  sky130_fd_sc_hd__clkinv_1 U15162 ( .A(n14642), .Y(n14623) );
  sky130_fd_sc_hd__clkinv_1 U15163 ( .A(n20312), .Y(n19657) );
  sky130_fd_sc_hd__clkinv_1 U15164 ( .A(n16856), .Y(n16861) );
  sky130_fd_sc_hd__clkinv_1 U15165 ( .A(n23077), .Y(n23084) );
  sky130_fd_sc_hd__clkinv_1 U15167 ( .A(n25423), .Y(n25428) );
  sky130_fd_sc_hd__clkinv_1 U15168 ( .A(n28045), .Y(n23041) );
  sky130_fd_sc_hd__clkinv_1 U15169 ( .A(n19680), .Y(n19681) );
  sky130_fd_sc_hd__clkinv_1 U15170 ( .A(n19700), .Y(n19702) );
  sky130_fd_sc_hd__clkinv_1 U15171 ( .A(n15341), .Y(n15273) );
  sky130_fd_sc_hd__clkinv_1 U15172 ( .A(n16832), .Y(n14674) );
  sky130_fd_sc_hd__clkinv_1 U15173 ( .A(n20703), .Y(n20705) );
  sky130_fd_sc_hd__clkinv_1 U15174 ( .A(n23323), .Y(n23326) );
  sky130_fd_sc_hd__clkinv_1 U15175 ( .A(n29563), .Y(n25204) );
  sky130_fd_sc_hd__clkinv_1 U15176 ( .A(n13229), .Y(n13230) );
  sky130_fd_sc_hd__clkinv_1 U15177 ( .A(n17814), .Y(n11429) );
  sky130_fd_sc_hd__clkinv_1 U15178 ( .A(n20954), .Y(n20079) );
  sky130_fd_sc_hd__clkinv_1 U15179 ( .A(n19494), .Y(n19439) );
  sky130_fd_sc_hd__clkinv_1 U15180 ( .A(n28367), .Y(n24696) );
  sky130_fd_sc_hd__clkinv_1 U15181 ( .A(n23121), .Y(n23122) );
  sky130_fd_sc_hd__clkinv_1 U15182 ( .A(n15599), .Y(n15519) );
  sky130_fd_sc_hd__clkinv_1 U15183 ( .A(n21771), .Y(n21774) );
  sky130_fd_sc_hd__clkinv_1 U15184 ( .A(n20213), .Y(n20217) );
  sky130_fd_sc_hd__clkinv_1 U15185 ( .A(n20230), .Y(n19985) );
  sky130_fd_sc_hd__clkinv_1 U15186 ( .A(n20031), .Y(n19984) );
  sky130_fd_sc_hd__clkinv_1 U15187 ( .A(n16147), .Y(n16148) );
  sky130_fd_sc_hd__clkinv_1 U15188 ( .A(n20646), .Y(n20494) );
  sky130_fd_sc_hd__clkinv_1 U15189 ( .A(n16655), .Y(n15309) );
  sky130_fd_sc_hd__clkinv_1 U15190 ( .A(n16150), .Y(n14672) );
  sky130_fd_sc_hd__clkinv_1 U15191 ( .A(n23124), .Y(n23126) );
  sky130_fd_sc_hd__clkinv_1 U15193 ( .A(n15508), .Y(n15594) );
  sky130_fd_sc_hd__clkinv_1 U15194 ( .A(n20829), .Y(n20463) );
  sky130_fd_sc_hd__clkinv_1 U15195 ( .A(n16610), .Y(n16612) );
  sky130_fd_sc_hd__clkinv_1 U15196 ( .A(n28847), .Y(n28751) );
  sky130_fd_sc_hd__clkinv_1 U15197 ( .A(n23176), .Y(n23184) );
  sky130_fd_sc_hd__clkinv_1 U15198 ( .A(n18003), .Y(n11507) );
  sky130_fd_sc_hd__or2_0 U15199 ( .A(n18454), .B(n18453), .X(n17437) );
  sky130_fd_sc_hd__clkinv_1 U15200 ( .A(n19706), .Y(n19448) );
  sky130_fd_sc_hd__clkinv_1 U15201 ( .A(n15697), .Y(n16578) );
  sky130_fd_sc_hd__clkinv_1 U15203 ( .A(n21601), .Y(n21393) );
  sky130_fd_sc_hd__clkinv_1 U15204 ( .A(n29270), .Y(n28702) );
  sky130_fd_sc_hd__clkinv_1 U15205 ( .A(n20036), .Y(n20118) );
  sky130_fd_sc_hd__clkinv_1 U15206 ( .A(n19562), .Y(n20270) );
  sky130_fd_sc_hd__a2bb2oi_1 U15207 ( .B1(n14378), .B2(
        j202_soc_core_j22_cpu_regop_imm__2_), .A1_N(n19265), .A2_N(n16525), 
        .Y(n13916) );
  sky130_fd_sc_hd__clkinv_1 U15208 ( .A(n15751), .Y(n16374) );
  sky130_fd_sc_hd__clkinv_1 U15209 ( .A(j202_soc_core_wbqspiflash_00_N710), 
        .Y(n28022) );
  sky130_fd_sc_hd__clkinv_1 U15210 ( .A(n21457), .Y(n21449) );
  sky130_fd_sc_hd__a2bb2oi_1 U15211 ( .B1(n14378), .B2(
        j202_soc_core_j22_cpu_regop_imm__0_), .A1_N(n21671), .A2_N(n16525), 
        .Y(n13853) );
  sky130_fd_sc_hd__clkinv_1 U15212 ( .A(n20765), .Y(n20768) );
  sky130_fd_sc_hd__clkinv_1 U15213 ( .A(n15198), .Y(n15093) );
  sky130_fd_sc_hd__clkinv_1 U15214 ( .A(n27756), .Y(n24671) );
  sky130_fd_sc_hd__clkinv_1 U15215 ( .A(n21707), .Y(n26003) );
  sky130_fd_sc_hd__clkinv_1 U15216 ( .A(n21127), .Y(n21379) );
  sky130_fd_sc_hd__clkinv_1 U15218 ( .A(n21452), .Y(n21772) );
  sky130_fd_sc_hd__clkinv_1 U15219 ( .A(n21817), .Y(n19923) );
  sky130_fd_sc_hd__clkinv_1 U15220 ( .A(n19414), .Y(n19420) );
  sky130_fd_sc_hd__clkinv_1 U15221 ( .A(n21525), .Y(n21570) );
  sky130_fd_sc_hd__clkinv_1 U15222 ( .A(n19753), .Y(n19484) );
  sky130_fd_sc_hd__and2_0 U15223 ( .A(n16577), .B(n16677), .X(n12118) );
  sky130_fd_sc_hd__clkinv_1 U15224 ( .A(n19956), .Y(n20006) );
  sky130_fd_sc_hd__clkinv_1 U15225 ( .A(n20799), .Y(n20800) );
  sky130_fd_sc_hd__clkinv_1 U15226 ( .A(n20172), .Y(n18729) );
  sky130_fd_sc_hd__clkinv_1 U15227 ( .A(n16945), .Y(n16946) );
  sky130_fd_sc_hd__clkinv_1 U15228 ( .A(n21556), .Y(n17259) );
  sky130_fd_sc_hd__clkinv_1 U15229 ( .A(n16782), .Y(n16751) );
  sky130_fd_sc_hd__clkinv_1 U15230 ( .A(n16759), .Y(n16136) );
  sky130_fd_sc_hd__clkinv_1 U15231 ( .A(n15304), .Y(n15305) );
  sky130_fd_sc_hd__clkinv_1 U15232 ( .A(n14667), .Y(n14629) );
  sky130_fd_sc_hd__clkinv_1 U15233 ( .A(n14678), .Y(n16803) );
  sky130_fd_sc_hd__clkinv_1 U15234 ( .A(n15532), .Y(n15347) );
  sky130_fd_sc_hd__clkinv_1 U15235 ( .A(n20360), .Y(n20361) );
  sky130_fd_sc_hd__clkinv_1 U15236 ( .A(n16859), .Y(n16116) );
  sky130_fd_sc_hd__clkinv_1 U15237 ( .A(n16808), .Y(n16810) );
  sky130_fd_sc_hd__clkinv_1 U15238 ( .A(n16805), .Y(n16807) );
  sky130_fd_sc_hd__clkinv_1 U15239 ( .A(n19370), .Y(n19404) );
  sky130_fd_sc_hd__clkinv_1 U15240 ( .A(n15733), .Y(n16639) );
  sky130_fd_sc_hd__clkinv_1 U15241 ( .A(n20372), .Y(n19324) );
  sky130_fd_sc_hd__clkinv_1 U15242 ( .A(n19929), .Y(n19927) );
  sky130_fd_sc_hd__clkinv_1 U15243 ( .A(n19574), .Y(n20333) );
  sky130_fd_sc_hd__clkinv_1 U15244 ( .A(n20326), .Y(n20328) );
  sky130_fd_sc_hd__clkinv_1 U15245 ( .A(n20047), .Y(n19880) );
  sky130_fd_sc_hd__clkinv_1 U15246 ( .A(n15718), .Y(n15736) );
  sky130_fd_sc_hd__clkinv_1 U15247 ( .A(n20656), .Y(n16587) );
  sky130_fd_sc_hd__clkinv_1 U15248 ( .A(n16214), .Y(n16165) );
  sky130_fd_sc_hd__clkinv_1 U15249 ( .A(n16663), .Y(n16309) );
  sky130_fd_sc_hd__clkinv_1 U15250 ( .A(n20293), .Y(n20295) );
  sky130_fd_sc_hd__clkinv_1 U15251 ( .A(n26974), .Y(n26976) );
  sky130_fd_sc_hd__clkinv_1 U15252 ( .A(n24835), .Y(n24837) );
  sky130_fd_sc_hd__clkinv_1 U15253 ( .A(n17291), .Y(n21355) );
  sky130_fd_sc_hd__clkinv_1 U15254 ( .A(n22418), .Y(n22419) );
  sky130_fd_sc_hd__o2bb2ai_1 U15255 ( .B1(n21243), .B2(n16525), .A1_N(n14378), 
        .A2_N(j202_soc_core_j22_cpu_regop_imm__3_), .Y(n13717) );
  sky130_fd_sc_hd__clkinv_1 U15256 ( .A(n21426), .Y(n17287) );
  sky130_fd_sc_hd__clkinv_1 U15257 ( .A(n24092), .Y(n27776) );
  sky130_fd_sc_hd__clkinv_1 U15258 ( .A(n16273), .Y(n16276) );
  sky130_fd_sc_hd__clkinv_1 U15259 ( .A(n19597), .Y(n19599) );
  sky130_fd_sc_hd__clkinv_1 U15260 ( .A(n26653), .Y(n24278) );
  sky130_fd_sc_hd__clkinv_1 U15261 ( .A(n16204), .Y(n16209) );
  sky130_fd_sc_hd__clkinv_1 U15262 ( .A(n16818), .Y(n16217) );
  sky130_fd_sc_hd__clkinv_1 U15263 ( .A(n28161), .Y(n28165) );
  sky130_fd_sc_hd__clkinv_1 U15264 ( .A(n20077), .Y(n20072) );
  sky130_fd_sc_hd__buf_2 U15265 ( .A(n18678), .X(n28045) );
  sky130_fd_sc_hd__clkinv_1 U15266 ( .A(n25725), .Y(n25726) );
  sky130_fd_sc_hd__clkinv_1 U15267 ( .A(n20598), .Y(n19142) );
  sky130_fd_sc_hd__clkinv_1 U15268 ( .A(n13325), .Y(n28441) );
  sky130_fd_sc_hd__clkinv_1 U15269 ( .A(n21146), .Y(n21555) );
  sky130_fd_sc_hd__clkinv_1 U15270 ( .A(n27194), .Y(n26491) );
  sky130_fd_sc_hd__clkinv_1 U15271 ( .A(n16660), .Y(n16704) );
  sky130_fd_sc_hd__clkinv_1 U15272 ( .A(n19783), .Y(n19784) );
  sky130_fd_sc_hd__a2bb2oi_1 U15273 ( .B1(n14378), .B2(
        j202_soc_core_j22_cpu_regop_imm__11_), .A1_N(n21292), .A2_N(n16525), 
        .Y(n14012) );
  sky130_fd_sc_hd__clkinv_1 U15274 ( .A(n19733), .Y(n19740) );
  sky130_fd_sc_hd__clkinv_1 U15275 ( .A(n20736), .Y(n20549) );
  sky130_fd_sc_hd__clkinv_1 U15276 ( .A(n29176), .Y(n28619) );
  sky130_fd_sc_hd__a2bb2oi_1 U15277 ( .B1(n14378), .B2(
        j202_soc_core_j22_cpu_regop_imm__10_), .A1_N(n19282), .A2_N(n16525), 
        .Y(n14348) );
  sky130_fd_sc_hd__clkinv_1 U15278 ( .A(n16670), .Y(n16671) );
  sky130_fd_sc_hd__clkinv_1 U15279 ( .A(n19667), .Y(n19668) );
  sky130_fd_sc_hd__clkinv_1 U15280 ( .A(n18248), .Y(n11461) );
  sky130_fd_sc_hd__a2bb2oi_1 U15281 ( .B1(n14378), .B2(
        j202_soc_core_j22_cpu_regop_imm__9_), .A1_N(n22891), .A2_N(n16525), 
        .Y(n14380) );
  sky130_fd_sc_hd__clkinv_1 U15282 ( .A(n20841), .Y(n20677) );
  sky130_fd_sc_hd__clkinv_1 U15283 ( .A(n19693), .Y(n15412) );
  sky130_fd_sc_hd__clkinv_1 U15284 ( .A(n16303), .Y(n25286) );
  sky130_fd_sc_hd__clkinv_1 U15285 ( .A(n29115), .Y(n28547) );
  sky130_fd_sc_hd__clkinv_1 U15286 ( .A(n25109), .Y(n25266) );
  sky130_fd_sc_hd__clkinv_1 U15287 ( .A(n19656), .Y(n19621) );
  sky130_fd_sc_hd__clkinv_1 U15288 ( .A(n27787), .Y(n25682) );
  sky130_fd_sc_hd__clkinv_1 U15289 ( .A(n21162), .Y(n21168) );
  sky130_fd_sc_hd__clkinv_1 U15290 ( .A(n25015), .Y(n25012) );
  sky130_fd_sc_hd__clkinv_1 U15291 ( .A(n19765), .Y(n19435) );
  sky130_fd_sc_hd__clkinv_1 U15292 ( .A(n21399), .Y(n17260) );
  sky130_fd_sc_hd__clkinv_1 U15293 ( .A(n17322), .Y(n17329) );
  sky130_fd_sc_hd__clkinv_1 U15295 ( .A(n15257), .Y(n15631) );
  sky130_fd_sc_hd__clkinv_1 U15296 ( .A(n26574), .Y(n26579) );
  sky130_fd_sc_hd__clkinv_1 U15297 ( .A(n16275), .Y(n14608) );
  sky130_fd_sc_hd__clkinv_1 U15298 ( .A(n24070), .Y(n25933) );
  sky130_fd_sc_hd__and4_1 U15299 ( .A(n14912), .B(n14911), .C(n14910), .D(
        n14909), .X(n14913) );
  sky130_fd_sc_hd__nand2_1 U15300 ( .A(n12734), .B(n12735), .Y(n11630) );
  sky130_fd_sc_hd__clkinv_1 U15301 ( .A(n28106), .Y(n28107) );
  sky130_fd_sc_hd__clkinv_1 U15302 ( .A(n15580), .Y(n15581) );
  sky130_fd_sc_hd__clkinv_1 U15303 ( .A(n16243), .Y(n16247) );
  sky130_fd_sc_hd__clkinv_1 U15304 ( .A(n23004), .Y(n21747) );
  sky130_fd_sc_hd__clkinv_1 U15305 ( .A(n16246), .Y(n14620) );
  sky130_fd_sc_hd__clkinv_1 U15306 ( .A(n16943), .Y(n16605) );
  sky130_fd_sc_hd__clkinv_1 U15307 ( .A(n20389), .Y(n17111) );
  sky130_fd_sc_hd__clkinv_1 U15308 ( .A(n15560), .Y(n15528) );
  sky130_fd_sc_hd__clkinv_1 U15309 ( .A(n16258), .Y(n14696) );
  sky130_fd_sc_hd__clkinv_1 U15310 ( .A(n19612), .Y(n17138) );
  sky130_fd_sc_hd__clkinv_1 U15311 ( .A(n24540), .Y(n16930) );
  sky130_fd_sc_hd__clkinv_1 U15312 ( .A(n16216), .Y(n14655) );
  sky130_fd_sc_hd__clkinv_1 U15313 ( .A(n14596), .Y(n14706) );
  sky130_fd_sc_hd__clkinv_1 U15314 ( .A(n26616), .Y(n23875) );
  sky130_fd_sc_hd__clkinv_1 U15315 ( .A(n16746), .Y(n16849) );
  sky130_fd_sc_hd__clkinv_1 U15316 ( .A(n16747), .Y(n16271) );
  sky130_fd_sc_hd__clkinv_1 U15317 ( .A(n17101), .Y(n14673) );
  sky130_fd_sc_hd__clkinv_1 U15318 ( .A(n25166), .Y(n26991) );
  sky130_fd_sc_hd__clkinv_1 U15319 ( .A(n16274), .Y(n16126) );
  sky130_fd_sc_hd__clkinv_1 U15320 ( .A(n21003), .Y(n20978) );
  sky130_fd_sc_hd__clkinv_1 U15321 ( .A(n16698), .Y(n16699) );
  sky130_fd_sc_hd__clkinv_1 U15322 ( .A(n26035), .Y(n26037) );
  sky130_fd_sc_hd__clkinv_1 U15323 ( .A(n19584), .Y(n19642) );
  sky130_fd_sc_hd__clkinv_1 U15324 ( .A(n15130), .Y(n15344) );
  sky130_fd_sc_hd__clkinv_1 U15325 ( .A(n29170), .Y(n27515) );
  sky130_fd_sc_hd__and2_0 U15326 ( .A(n20199), .B(n14597), .X(n12115) );
  sky130_fd_sc_hd__clkinv_1 U15327 ( .A(n28162), .Y(n28163) );
  sky130_fd_sc_hd__clkinv_1 U15328 ( .A(n20076), .Y(n20078) );
  sky130_fd_sc_hd__clkinv_1 U15329 ( .A(n28202), .Y(n22761) );
  sky130_fd_sc_hd__clkinv_1 U15330 ( .A(n16334), .Y(n16680) );
  sky130_fd_sc_hd__clkinv_1 U15332 ( .A(n16376), .Y(n16367) );
  sky130_fd_sc_hd__clkinv_1 U15333 ( .A(n22285), .Y(n22990) );
  sky130_fd_sc_hd__clkinv_1 U15334 ( .A(n16349), .Y(n15727) );
  sky130_fd_sc_hd__clkinv_1 U15336 ( .A(n16573), .Y(n15671) );
  sky130_fd_sc_hd__clkinv_1 U15337 ( .A(n15535), .Y(n15605) );
  sky130_fd_sc_hd__clkinv_1 U15338 ( .A(n21571), .Y(n21109) );
  sky130_fd_sc_hd__clkinv_1 U15339 ( .A(n15676), .Y(n15672) );
  sky130_fd_sc_hd__clkinv_1 U15340 ( .A(n21453), .Y(n21448) );
  sky130_fd_sc_hd__clkinv_1 U15341 ( .A(n16921), .Y(n16922) );
  sky130_fd_sc_hd__clkinv_1 U15342 ( .A(n16809), .Y(n14631) );
  sky130_fd_sc_hd__clkinv_1 U15343 ( .A(n16226), .Y(n16775) );
  sky130_fd_sc_hd__clkinv_1 U15344 ( .A(n16789), .Y(n16791) );
  sky130_fd_sc_hd__clkinv_1 U15345 ( .A(n27610), .Y(n27611) );
  sky130_fd_sc_hd__clkinv_1 U15346 ( .A(n28432), .Y(n23627) );
  sky130_fd_sc_hd__clkinv_1 U15347 ( .A(n27486), .Y(n27482) );
  sky130_fd_sc_hd__clkinv_1 U15348 ( .A(n23563), .Y(n23495) );
  sky130_fd_sc_hd__clkinv_1 U15349 ( .A(n28340), .Y(n28341) );
  sky130_fd_sc_hd__clkinv_1 U15350 ( .A(n25009), .Y(n25005) );
  sky130_fd_sc_hd__clkinv_1 U15351 ( .A(n15583), .Y(n15300) );
  sky130_fd_sc_hd__clkinv_1 U15352 ( .A(n15274), .Y(n15525) );
  sky130_fd_sc_hd__clkinv_1 U15353 ( .A(n15394), .Y(n15269) );
  sky130_fd_sc_hd__clkinv_1 U15354 ( .A(n19504), .Y(n15159) );
  sky130_fd_sc_hd__clkinv_1 U15355 ( .A(n16745), .Y(n16762) );
  sky130_fd_sc_hd__inv_2 U15356 ( .A(n26048), .Y(n26426) );
  sky130_fd_sc_hd__clkinv_1 U15357 ( .A(n26640), .Y(n25344) );
  sky130_fd_sc_hd__clkinv_1 U15358 ( .A(n29267), .Y(n26569) );
  sky130_fd_sc_hd__clkinv_1 U15359 ( .A(n22998), .Y(n22722) );
  sky130_fd_sc_hd__clkinv_1 U15360 ( .A(n26593), .Y(n26603) );
  sky130_fd_sc_hd__clkinv_1 U15361 ( .A(n24034), .Y(n13378) );
  sky130_fd_sc_hd__clkinv_1 U15362 ( .A(n20687), .Y(n20827) );
  sky130_fd_sc_hd__clkinv_1 U15363 ( .A(n20741), .Y(n20487) );
  sky130_fd_sc_hd__clkinv_1 U15364 ( .A(n20490), .Y(n20491) );
  sky130_fd_sc_hd__clkinv_1 U15365 ( .A(n20528), .Y(n19202) );
  sky130_fd_sc_hd__clkinv_1 U15366 ( .A(n20652), .Y(n20482) );
  sky130_fd_sc_hd__clkinv_1 U15367 ( .A(n20559), .Y(n20509) );
  sky130_fd_sc_hd__clkinv_1 U15368 ( .A(n20731), .Y(n20521) );
  sky130_fd_sc_hd__clkinv_1 U15369 ( .A(n20675), .Y(n19157) );
  sky130_fd_sc_hd__clkinv_1 U15370 ( .A(n20486), .Y(n20466) );
  sky130_fd_sc_hd__clkinv_1 U15371 ( .A(n26464), .Y(n26463) );
  sky130_fd_sc_hd__clkinv_1 U15372 ( .A(n26520), .Y(n27186) );
  sky130_fd_sc_hd__clkinv_1 U15373 ( .A(n19397), .Y(n17127) );
  sky130_fd_sc_hd__clkinv_1 U15374 ( .A(n21521), .Y(n21524) );
  sky130_fd_sc_hd__and2_0 U15375 ( .A(n20371), .B(n20348), .X(n17133) );
  sky130_fd_sc_hd__clkinv_1 U15376 ( .A(n21536), .Y(n21532) );
  sky130_fd_sc_hd__clkinv_1 U15377 ( .A(n21421), .Y(n17294) );
  sky130_fd_sc_hd__clkinv_1 U15378 ( .A(n18716), .Y(n20166) );
  sky130_fd_sc_hd__clkinv_1 U15379 ( .A(n21415), .Y(n21138) );
  sky130_fd_sc_hd__clkinv_1 U15380 ( .A(n17146), .Y(n20617) );
  sky130_fd_sc_hd__clkinv_1 U15381 ( .A(n19981), .Y(n19982) );
  sky130_fd_sc_hd__clkinv_1 U15382 ( .A(n19561), .Y(n19622) );
  sky130_fd_sc_hd__clkinv_1 U15383 ( .A(n17267), .Y(n17271) );
  sky130_fd_sc_hd__clkinv_1 U15384 ( .A(n20364), .Y(n17152) );
  sky130_fd_sc_hd__clkinv_1 U15385 ( .A(n17150), .Y(n17151) );
  sky130_fd_sc_hd__clkinv_1 U15386 ( .A(n20182), .Y(n18723) );
  sky130_fd_sc_hd__inv_1 U15387 ( .A(n20060), .Y(n19897) );
  sky130_fd_sc_hd__clkinv_1 U15388 ( .A(n19369), .Y(n17148) );
  sky130_fd_sc_hd__clkinv_1 U15389 ( .A(n17272), .Y(n21615) );
  sky130_fd_sc_hd__clkinv_1 U15390 ( .A(n24697), .Y(n23418) );
  sky130_fd_sc_hd__clkinv_1 U15391 ( .A(n21354), .Y(n21082) );
  sky130_fd_sc_hd__clkinv_1 U15392 ( .A(n16780), .Y(n16132) );
  sky130_fd_sc_hd__clkinv_1 U15393 ( .A(n21527), .Y(n21090) );
  sky130_fd_sc_hd__clkinv_1 U15394 ( .A(n19812), .Y(n19487) );
  sky130_fd_sc_hd__clkinv_1 U15395 ( .A(n26511), .Y(n23634) );
  sky130_fd_sc_hd__clkinv_1 U15396 ( .A(n21576), .Y(n21114) );
  sky130_fd_sc_hd__clkinv_1 U15397 ( .A(n20376), .Y(n20378) );
  sky130_fd_sc_hd__clkinv_1 U15398 ( .A(n21550), .Y(n21122) );
  sky130_fd_sc_hd__clkinv_1 U15399 ( .A(n16154), .Y(n16155) );
  sky130_fd_sc_hd__clkinv_1 U15400 ( .A(n20137), .Y(n18768) );
  sky130_fd_sc_hd__clkinv_1 U15401 ( .A(n19951), .Y(n19946) );
  sky130_fd_sc_hd__clkinv_1 U15402 ( .A(n25152), .Y(n21320) );
  sky130_fd_sc_hd__clkinv_1 U15403 ( .A(n21573), .Y(n21427) );
  sky130_fd_sc_hd__clkinv_1 U15404 ( .A(n20173), .Y(n18714) );
  sky130_fd_sc_hd__and2_0 U15405 ( .A(n20268), .B(n20348), .X(n17106) );
  sky130_fd_sc_hd__clkinv_1 U15406 ( .A(n20306), .Y(n17107) );
  sky130_fd_sc_hd__clkinv_1 U15407 ( .A(n21142), .Y(n21147) );
  sky130_fd_sc_hd__clkinv_1 U15408 ( .A(n15598), .Y(n15137) );
  sky130_fd_sc_hd__clkinv_1 U15409 ( .A(n19827), .Y(n19828) );
  sky130_fd_sc_hd__clkinv_1 U15410 ( .A(n20029), .Y(n20112) );
  sky130_fd_sc_hd__clkinv_1 U15411 ( .A(n14610), .Y(n16262) );
  sky130_fd_sc_hd__clkinv_1 U15412 ( .A(n19206), .Y(n19207) );
  sky130_fd_sc_hd__clkinv_1 U15413 ( .A(n20828), .Y(n19126) );
  sky130_fd_sc_hd__clkinv_1 U15414 ( .A(n18504), .Y(n11409) );
  sky130_fd_sc_hd__nor2_1 U15415 ( .A(n18249), .B(n18250), .Y(n11462) );
  sky130_fd_sc_hd__clkinv_1 U15416 ( .A(n23000), .Y(n22639) );
  sky130_fd_sc_hd__clkinv_1 U15417 ( .A(n20814), .Y(n20816) );
  sky130_fd_sc_hd__nand2_2 U15418 ( .A(n13327), .B(n28047), .Y(n13325) );
  sky130_fd_sc_hd__clkinv_1 U15419 ( .A(n20033), .Y(n19957) );
  sky130_fd_sc_hd__clkinv_1 U15420 ( .A(n23272), .Y(n23276) );
  sky130_fd_sc_hd__clkinv_1 U15421 ( .A(n14684), .Y(n14685) );
  sky130_fd_sc_hd__clkinv_1 U15422 ( .A(n17288), .Y(n16611) );
  sky130_fd_sc_hd__clkinv_1 U15423 ( .A(n15431), .Y(n15403) );
  sky130_fd_sc_hd__clkinv_1 U15424 ( .A(n20603), .Y(n20604) );
  sky130_fd_sc_hd__clkinv_1 U15425 ( .A(n16619), .Y(n16620) );
  sky130_fd_sc_hd__clkinv_1 U15426 ( .A(n16988), .Y(n16601) );
  sky130_fd_sc_hd__clkinv_1 U15427 ( .A(n19781), .Y(n15420) );
  sky130_fd_sc_hd__clkinv_1 U15428 ( .A(n24075), .Y(n24905) );
  sky130_fd_sc_hd__clkinv_1 U15429 ( .A(n28617), .Y(n28620) );
  sky130_fd_sc_hd__clkinv_1 U15430 ( .A(n20790), .Y(n20624) );
  sky130_fd_sc_hd__clkinv_1 U15431 ( .A(n20055), .Y(n20145) );
  sky130_fd_sc_hd__clkinv_1 U15432 ( .A(n25658), .Y(n25868) );
  sky130_fd_sc_hd__nand2b_1 U15433 ( .A_N(n19463), .B(n15685), .Y(n19693) );
  sky130_fd_sc_hd__inv_2 U15434 ( .A(n27318), .Y(n23212) );
  sky130_fd_sc_hd__clkinv_1 U15435 ( .A(n24032), .Y(n23891) );
  sky130_fd_sc_hd__clkinv_1 U15436 ( .A(n20301), .Y(n20302) );
  sky130_fd_sc_hd__nor2_4 U15437 ( .A(n13163), .B(n13162), .Y(n21503) );
  sky130_fd_sc_hd__and2_0 U15438 ( .A(n29603), .B(n25534), .X(n29704) );
  sky130_fd_sc_hd__and2_0 U15439 ( .A(n29603), .B(n25548), .X(n29703) );
  sky130_fd_sc_hd__clkinv_1 U15440 ( .A(n24450), .Y(n21749) );
  sky130_fd_sc_hd__and2_0 U15441 ( .A(n29603), .B(n25550), .X(n29708) );
  sky130_fd_sc_hd__and2_0 U15442 ( .A(n29603), .B(n25532), .X(n29717) );
  sky130_fd_sc_hd__clkinv_1 U15443 ( .A(n16815), .Y(n16848) );
  sky130_fd_sc_hd__clkinv_1 U15444 ( .A(n19605), .Y(n13273) );
  sky130_fd_sc_hd__clkinv_1 U15445 ( .A(n27754), .Y(n27755) );
  sky130_fd_sc_hd__clkinv_1 U15446 ( .A(n28848), .Y(n26512) );
  sky130_fd_sc_hd__clkinv_1 U15447 ( .A(n27431), .Y(n26516) );
  sky130_fd_sc_hd__and2_0 U15448 ( .A(n29603), .B(n25536), .X(n29700) );
  sky130_fd_sc_hd__and2_0 U15449 ( .A(n29603), .B(n25538), .X(n29699) );
  sky130_fd_sc_hd__clkinv_1 U15450 ( .A(n20138), .Y(n18745) );
  sky130_fd_sc_hd__clkinv_1 U15451 ( .A(n25342), .Y(n28849) );
  sky130_fd_sc_hd__clkinv_1 U15452 ( .A(n26514), .Y(n26597) );
  sky130_fd_sc_hd__clkinv_1 U15453 ( .A(n28656), .Y(n27220) );
  sky130_fd_sc_hd__and2_0 U15454 ( .A(n29603), .B(n25546), .X(n29716) );
  sky130_fd_sc_hd__and2_0 U15455 ( .A(n29603), .B(n25540), .X(n29698) );
  sky130_fd_sc_hd__and2_0 U15456 ( .A(n29603), .B(n25542), .X(n29697) );
  sky130_fd_sc_hd__and2_0 U15457 ( .A(n29603), .B(n25544), .X(n29696) );
  sky130_fd_sc_hd__clkinv_1 U15458 ( .A(n23018), .Y(n22732) );
  sky130_fd_sc_hd__clkinv_1 U15459 ( .A(n28836), .Y(n26529) );
  sky130_fd_sc_hd__clkinv_1 U15460 ( .A(n28677), .Y(n25341) );
  sky130_fd_sc_hd__clkinv_1 U15461 ( .A(n28730), .Y(n28857) );
  sky130_fd_sc_hd__clkinv_1 U15462 ( .A(n27297), .Y(n26489) );
  sky130_fd_sc_hd__and2_0 U15463 ( .A(n29603), .B(n25514), .X(n29713) );
  sky130_fd_sc_hd__clkinv_1 U15464 ( .A(n28814), .Y(n23991) );
  sky130_fd_sc_hd__clkinv_1 U15465 ( .A(n16638), .Y(n15665) );
  sky130_fd_sc_hd__and2_0 U15466 ( .A(n29603), .B(n25516), .X(n29701) );
  sky130_fd_sc_hd__and2_0 U15467 ( .A(n29603), .B(n25518), .X(n29712) );
  sky130_fd_sc_hd__clkinv_1 U15468 ( .A(n20103), .Y(n18773) );
  sky130_fd_sc_hd__and2_0 U15469 ( .A(n29603), .B(n25520), .X(n29721) );
  sky130_fd_sc_hd__and2_0 U15471 ( .A(n29603), .B(n25522), .X(n29711) );
  sky130_fd_sc_hd__clkinv_1 U15472 ( .A(n27259), .Y(n28869) );
  sky130_fd_sc_hd__clkinv_1 U15473 ( .A(n19394), .Y(n16159) );
  sky130_fd_sc_hd__and2_0 U15474 ( .A(n29603), .B(n25524), .X(n29718) );
  sky130_fd_sc_hd__clkinv_1 U15475 ( .A(n27245), .Y(n27247) );
  sky130_fd_sc_hd__clkinv_1 U15476 ( .A(n16268), .Y(n16114) );
  sky130_fd_sc_hd__and2_0 U15477 ( .A(n29603), .B(n25526), .X(n29710) );
  sky130_fd_sc_hd__clkinv_1 U15478 ( .A(n27429), .Y(n26533) );
  sky130_fd_sc_hd__and2_0 U15479 ( .A(n29603), .B(n25528), .X(n29720) );
  sky130_fd_sc_hd__and2_0 U15480 ( .A(n29276), .B(n12069), .X(n29651) );
  sky130_fd_sc_hd__and2_0 U15481 ( .A(n29603), .B(n25530), .X(n29709) );
  sky130_fd_sc_hd__clkinv_1 U15482 ( .A(n16763), .Y(n14644) );
  sky130_fd_sc_hd__clkinv_1 U15483 ( .A(n16820), .Y(n14676) );
  sky130_fd_sc_hd__clkinv_1 U15484 ( .A(n19593), .Y(n28164) );
  sky130_fd_sc_hd__clkinv_1 U15485 ( .A(n24416), .Y(n23416) );
  sky130_fd_sc_hd__clkinv_1 U15486 ( .A(n13787), .Y(n13788) );
  sky130_fd_sc_hd__clkinv_1 U15487 ( .A(n14665), .Y(n14666) );
  sky130_fd_sc_hd__clkinv_1 U15488 ( .A(n11876), .Y(n11874) );
  sky130_fd_sc_hd__clkinv_1 U15489 ( .A(n29181), .Y(n12) );
  sky130_fd_sc_hd__inv_2 U15490 ( .A(n22365), .Y(n22979) );
  sky130_fd_sc_hd__clkinv_1 U15491 ( .A(n20515), .Y(n20674) );
  sky130_fd_sc_hd__clkinv_1 U15492 ( .A(n26781), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N34) );
  sky130_fd_sc_hd__clkinv_1 U15493 ( .A(n21097), .Y(n17284) );
  sky130_fd_sc_hd__clkinv_1 U15494 ( .A(n25830), .Y(n18806) );
  sky130_fd_sc_hd__clkinv_1 U15495 ( .A(n20516), .Y(n19122) );
  sky130_fd_sc_hd__clkinv_1 U15496 ( .A(n19145), .Y(n19123) );
  sky130_fd_sc_hd__clkinv_1 U15497 ( .A(n22230), .Y(n21934) );
  sky130_fd_sc_hd__clkinv_1 U15498 ( .A(n19180), .Y(n17122) );
  sky130_fd_sc_hd__clkinv_1 U15499 ( .A(n16755), .Y(n14705) );
  sky130_fd_sc_hd__clkinv_1 U15500 ( .A(n19183), .Y(n19186) );
  sky130_fd_sc_hd__and2_0 U15501 ( .A(n29603), .B(n25552), .X(n29695) );
  sky130_fd_sc_hd__clkinv_1 U15502 ( .A(n26901), .Y(n26902) );
  sky130_fd_sc_hd__and2_0 U15503 ( .A(n29603), .B(n28023), .X(n29707) );
  sky130_fd_sc_hd__and2_0 U15504 ( .A(n29603), .B(n28893), .X(n29706) );
  sky130_fd_sc_hd__inv_1 U15505 ( .A(n12668), .Y(n12667) );
  sky130_fd_sc_hd__clkinv_1 U15506 ( .A(n19949), .Y(n18741) );
  sky130_fd_sc_hd__clkinv_1 U15507 ( .A(n28102), .Y(n28105) );
  sky130_fd_sc_hd__clkinv_1 U15508 ( .A(n21613), .Y(n21614) );
  sky130_fd_sc_hd__clkinv_1 U15509 ( .A(n29405), .Y(n29399) );
  sky130_fd_sc_hd__clkinv_1 U15510 ( .A(n29147), .Y(n29475) );
  sky130_fd_sc_hd__clkinv_1 U15511 ( .A(n26594), .Y(n25337) );
  sky130_fd_sc_hd__clkinv_1 U15512 ( .A(n14602), .Y(n14595) );
  sky130_fd_sc_hd__clkinv_1 U15513 ( .A(n16135), .Y(n14682) );
  sky130_fd_sc_hd__clkinv_1 U15514 ( .A(n19874), .Y(n19863) );
  sky130_fd_sc_hd__clkinv_1 U15515 ( .A(n26150), .Y(n25808) );
  sky130_fd_sc_hd__clkinv_1 U15516 ( .A(n21394), .Y(n21526) );
  sky130_fd_sc_hd__clkinv_1 U15517 ( .A(n24750), .Y(n24752) );
  sky130_fd_sc_hd__clkinv_1 U15518 ( .A(n23372), .Y(n23373) );
  sky130_fd_sc_hd__clkinv_1 U15519 ( .A(n20058), .Y(n20101) );
  sky130_fd_sc_hd__clkinv_1 U15520 ( .A(n22760), .Y(n19594) );
  sky130_fd_sc_hd__clkinv_1 U15521 ( .A(n15120), .Y(n15097) );
  sky130_fd_sc_hd__clkinv_1 U15522 ( .A(n15683), .Y(n21102) );
  sky130_fd_sc_hd__clkinv_1 U15523 ( .A(n16095), .Y(n21026) );
  sky130_fd_sc_hd__o22ai_1 U15524 ( .A1(n18213), .A2(n18194), .B1(n18193), 
        .B2(n12538), .Y(n12891) );
  sky130_fd_sc_hd__o22ai_1 U15525 ( .A1(n18213), .A2(n18021), .B1(n18081), 
        .B2(n12538), .Y(n18077) );
  sky130_fd_sc_hd__clkinv_1 U15526 ( .A(n27922), .Y(n27920) );
  sky130_fd_sc_hd__clkinv_1 U15527 ( .A(n23278), .Y(n21054) );
  sky130_fd_sc_hd__clkinv_1 U15528 ( .A(n19712), .Y(n19713) );
  sky130_fd_sc_hd__clkinv_1 U15529 ( .A(n26157), .Y(n24911) );
  sky130_fd_sc_hd__clkinv_1 U15530 ( .A(n29276), .Y(n26652) );
  sky130_fd_sc_hd__clkinv_1 U15531 ( .A(n27434), .Y(n27437) );
  sky130_fd_sc_hd__clkinv_1 U15532 ( .A(n20034), .Y(n19820) );
  sky130_fd_sc_hd__inv_2 U15533 ( .A(n15747), .Y(n20531) );
  sky130_fd_sc_hd__clkinv_1 U15534 ( .A(n24539), .Y(n24183) );
  sky130_fd_sc_hd__clkinv_1 U15535 ( .A(n16851), .Y(n14601) );
  sky130_fd_sc_hd__clkinv_1 U15536 ( .A(n29157), .Y(n29465) );
  sky130_fd_sc_hd__clkinv_1 U15537 ( .A(n28615), .Y(n28612) );
  sky130_fd_sc_hd__clkinv_1 U15538 ( .A(n29159), .Y(n29467) );
  sky130_fd_sc_hd__clkinv_1 U15539 ( .A(n19694), .Y(n19444) );
  sky130_fd_sc_hd__clkinv_1 U15540 ( .A(n27257), .Y(n28744) );
  sky130_fd_sc_hd__clkinv_1 U15541 ( .A(n15568), .Y(n15301) );
  sky130_fd_sc_hd__clkinv_1 U15542 ( .A(n27395), .Y(n29568) );
  sky130_fd_sc_hd__and2_0 U15543 ( .A(n29603), .B(n25506), .X(n29715) );
  sky130_fd_sc_hd__clkinv_1 U15544 ( .A(n21206), .Y(n25822) );
  sky130_fd_sc_hd__clkinv_1 U15545 ( .A(n24979), .Y(n24024) );
  sky130_fd_sc_hd__clkinv_1 U15546 ( .A(n27208), .Y(n27248) );
  sky130_fd_sc_hd__and2_0 U15547 ( .A(n29603), .B(
        j202_soc_core_wbqspiflash_00_spi_spd), .X(n28695) );
  sky130_fd_sc_hd__clkinv_1 U15548 ( .A(n28692), .Y(n28714) );
  sky130_fd_sc_hd__clkinv_1 U15549 ( .A(n13190), .Y(n13191) );
  sky130_fd_sc_hd__and2_0 U15550 ( .A(n29603), .B(n25508), .X(n29719) );
  sky130_fd_sc_hd__clkinv_1 U15551 ( .A(n22452), .Y(n22417) );
  sky130_fd_sc_hd__clkinv_1 U15552 ( .A(n15710), .Y(n15711) );
  sky130_fd_sc_hd__clkinv_1 U15554 ( .A(n26495), .Y(n26630) );
  sky130_fd_sc_hd__and2_0 U15555 ( .A(n29603), .B(n25512), .X(n29705) );
  sky130_fd_sc_hd__clkinv_1 U15556 ( .A(n18923), .Y(n18928) );
  sky130_fd_sc_hd__clkinv_1 U15557 ( .A(n28210), .Y(n24739) );
  sky130_fd_sc_hd__clkinv_1 U15558 ( .A(n25494), .Y(n29450) );
  sky130_fd_sc_hd__and2_0 U15559 ( .A(n29603), .B(n25504), .X(n29702) );
  sky130_fd_sc_hd__clkinv_1 U15560 ( .A(n28863), .Y(n26487) );
  sky130_fd_sc_hd__ha_1 U15562 ( .A(n18025), .B(n18024), .COUT(n18017), .SUM(
        n18043) );
  sky130_fd_sc_hd__and2_0 U15564 ( .A(n29603), .B(n25510), .X(n29714) );
  sky130_fd_sc_hd__clkinv_1 U15565 ( .A(n27172), .Y(n29453) );
  sky130_fd_sc_hd__clkinv_1 U15566 ( .A(n25614), .Y(n29456) );
  sky130_fd_sc_hd__inv_2 U15567 ( .A(n14052), .Y(n15991) );
  sky130_fd_sc_hd__o22ai_1 U15568 ( .A1(n18496), .A2(n17412), .B1(n18341), 
        .B2(n17410), .Y(n18416) );
  sky130_fd_sc_hd__clkinv_1 U15569 ( .A(n25582), .Y(n29457) );
  sky130_fd_sc_hd__clkinv_1 U15570 ( .A(n23248), .Y(n23249) );
  sky130_fd_sc_hd__clkinv_1 U15571 ( .A(n29156), .Y(n29448) );
  sky130_fd_sc_hd__clkinv_1 U15572 ( .A(n23344), .Y(n23345) );
  sky130_fd_sc_hd__clkinv_1 U15573 ( .A(n24304), .Y(n22089) );
  sky130_fd_sc_hd__clkinv_1 U15574 ( .A(n18706), .Y(n20043) );
  sky130_fd_sc_hd__clkinv_1 U15575 ( .A(n23973), .Y(n24299) );
  sky130_fd_sc_hd__clkinv_1 U15576 ( .A(n25940), .Y(n25392) );
  sky130_fd_sc_hd__clkinv_1 U15577 ( .A(n22950), .Y(n21729) );
  sky130_fd_sc_hd__clkinv_1 U15578 ( .A(n28157), .Y(n28158) );
  sky130_fd_sc_hd__clkinv_1 U15579 ( .A(n23750), .Y(n23751) );
  sky130_fd_sc_hd__inv_1 U15580 ( .A(n23788), .Y(n23789) );
  sky130_fd_sc_hd__clkinv_1 U15581 ( .A(n26347), .Y(n26143) );
  sky130_fd_sc_hd__clkinv_1 U15582 ( .A(n18724), .Y(n18725) );
  sky130_fd_sc_hd__clkinv_1 U15583 ( .A(n20885), .Y(n19861) );
  sky130_fd_sc_hd__clkinv_1 U15584 ( .A(n21173), .Y(n19860) );
  sky130_fd_sc_hd__clkinv_1 U15585 ( .A(n29155), .Y(n29447) );
  sky130_fd_sc_hd__clkinv_1 U15586 ( .A(n24394), .Y(n28359) );
  sky130_fd_sc_hd__clkinv_1 U15587 ( .A(n19966), .Y(n19967) );
  sky130_fd_sc_hd__clkinv_1 U15588 ( .A(n22897), .Y(n22989) );
  sky130_fd_sc_hd__clkinv_1 U15589 ( .A(n29154), .Y(n29446) );
  sky130_fd_sc_hd__inv_2 U15590 ( .A(n16491), .Y(n16532) );
  sky130_fd_sc_hd__clkinv_1 U15591 ( .A(n24702), .Y(n23419) );
  sky130_fd_sc_hd__clkinv_1 U15592 ( .A(n29144), .Y(n29478) );
  sky130_fd_sc_hd__clkinv_1 U15593 ( .A(n17254), .Y(n17268) );
  sky130_fd_sc_hd__and2_0 U15594 ( .A(n24910), .B(n26295), .X(n26362) );
  sky130_fd_sc_hd__clkinv_1 U15595 ( .A(n20833), .Y(n20632) );
  sky130_fd_sc_hd__clkinv_1 U15596 ( .A(n28841), .Y(n25345) );
  sky130_fd_sc_hd__clkinv_1 U15597 ( .A(n20929), .Y(n22698) );
  sky130_fd_sc_hd__clkinv_1 U15598 ( .A(n27231), .Y(n26608) );
  sky130_fd_sc_hd__and2_0 U15599 ( .A(io_in[32]), .B(n12069), .X(n29671) );
  sky130_fd_sc_hd__and2_0 U15600 ( .A(io_in[29]), .B(n12069), .X(n29673) );
  sky130_fd_sc_hd__clkinv_1 U15601 ( .A(n29145), .Y(n29477) );
  sky130_fd_sc_hd__clkinv_1 U15602 ( .A(n27183), .Y(n28669) );
  sky130_fd_sc_hd__and2_0 U15603 ( .A(io_in[28]), .B(n12069), .X(n29674) );
  sky130_fd_sc_hd__clkinv_1 U15604 ( .A(n27201), .Y(n28871) );
  sky130_fd_sc_hd__and2_0 U15605 ( .A(io_in[7]), .B(n12069), .X(n29677) );
  sky130_fd_sc_hd__clkinv_1 U15606 ( .A(n28688), .Y(n27267) );
  sky130_fd_sc_hd__and2_0 U15607 ( .A(io_in[3]), .B(n12069), .X(n29679) );
  sky130_fd_sc_hd__and2_0 U15608 ( .A(io_in[1]), .B(n12069), .X(n29681) );
  sky130_fd_sc_hd__clkinv_1 U15609 ( .A(io_out[8]), .Y(n26633) );
  sky130_fd_sc_hd__clkinv_1 U15610 ( .A(n20858), .Y(n20505) );
  sky130_fd_sc_hd__clkinv_1 U15611 ( .A(n27601), .Y(n29569) );
  sky130_fd_sc_hd__clkinv_1 U15612 ( .A(n24773), .Y(n20447) );
  sky130_fd_sc_hd__clkinv_1 U15613 ( .A(n18679), .Y(n18681) );
  sky130_fd_sc_hd__clkinv_1 U15614 ( .A(n28895), .Y(n24031) );
  sky130_fd_sc_hd__clkinv_1 U15615 ( .A(n17160), .Y(n17161) );
  sky130_fd_sc_hd__inv_2 U15616 ( .A(n14482), .Y(n11201) );
  sky130_fd_sc_hd__clkinv_1 U15617 ( .A(n27310), .Y(n24257) );
  sky130_fd_sc_hd__clkinv_1 U15618 ( .A(n26790), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N33) );
  sky130_fd_sc_hd__clkinv_1 U15619 ( .A(n26764), .Y(n29874) );
  sky130_fd_sc_hd__clkinv_1 U15620 ( .A(n26798), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N32) );
  sky130_fd_sc_hd__clkinv_1 U15621 ( .A(n21405), .Y(n21545) );
  sky130_fd_sc_hd__clkinv_1 U15622 ( .A(n26819), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N28) );
  sky130_fd_sc_hd__clkinv_1 U15623 ( .A(n26842), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N24) );
  sky130_fd_sc_hd__clkinv_1 U15624 ( .A(n29023), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N20) );
  sky130_fd_sc_hd__and2_0 U15625 ( .A(n12069), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15]), .X(n29735) );
  sky130_fd_sc_hd__clkinv_1 U15626 ( .A(n28986), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N15) );
  sky130_fd_sc_hd__clkinv_1 U15627 ( .A(n18855), .Y(n23969) );
  sky130_fd_sc_hd__and2_0 U15628 ( .A(n12069), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]), .X(n29727) );
  sky130_fd_sc_hd__and2_0 U15629 ( .A(n12069), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[2]), .X(n29736) );
  sky130_fd_sc_hd__clkinv_1 U15630 ( .A(n20225), .Y(n18720) );
  sky130_fd_sc_hd__clkinv_1 U15631 ( .A(n19146), .Y(n19128) );
  sky130_fd_sc_hd__clkinv_1 U15632 ( .A(n19235), .Y(n18796) );
  sky130_fd_sc_hd__clkinv_1 U15634 ( .A(n19001), .Y(n11966) );
  sky130_fd_sc_hd__clkinv_1 U15635 ( .A(n27280), .Y(n27221) );
  sky130_fd_sc_hd__clkinv_1 U15636 ( .A(n22983), .Y(n18872) );
  sky130_fd_sc_hd__clkinv_1 U15637 ( .A(n24029), .Y(n26664) );
  sky130_fd_sc_hd__clkinv_1 U15638 ( .A(n25518), .Y(n25519) );
  sky130_fd_sc_hd__clkinv_1 U15639 ( .A(n25520), .Y(n25521) );
  sky130_fd_sc_hd__clkinv_1 U15640 ( .A(n26340), .Y(n26419) );
  sky130_fd_sc_hd__clkinv_1 U15641 ( .A(n25522), .Y(n25523) );
  sky130_fd_sc_hd__clkinv_1 U15642 ( .A(n25524), .Y(n25525) );
  sky130_fd_sc_hd__clkinv_1 U15643 ( .A(n25526), .Y(n25527) );
  sky130_fd_sc_hd__clkinv_1 U15645 ( .A(n25528), .Y(n25529) );
  sky130_fd_sc_hd__clkinv_1 U15646 ( .A(n28401), .Y(n15651) );
  sky130_fd_sc_hd__clkinv_1 U15647 ( .A(n25530), .Y(n25531) );
  sky130_fd_sc_hd__clkinv_1 U15648 ( .A(n25532), .Y(n25533) );
  sky130_fd_sc_hd__clkinv_1 U15649 ( .A(n25534), .Y(n25535) );
  sky130_fd_sc_hd__clkinv_1 U15650 ( .A(n28623), .Y(n29174) );
  sky130_fd_sc_hd__clkinv_1 U15651 ( .A(n25516), .Y(n25517) );
  sky130_fd_sc_hd__clkinv_1 U15652 ( .A(n25737), .Y(n29875) );
  sky130_fd_sc_hd__clkinv_1 U15653 ( .A(n25536), .Y(n25537) );
  sky130_fd_sc_hd__clkinv_1 U15654 ( .A(n15516), .Y(n13183) );
  sky130_fd_sc_hd__inv_1 U15655 ( .A(n23824), .Y(n23825) );
  sky130_fd_sc_hd__clkinv_1 U15656 ( .A(n23819), .Y(n23820) );
  sky130_fd_sc_hd__clkinv_1 U15657 ( .A(n25538), .Y(n25539) );
  sky130_fd_sc_hd__inv_1 U15658 ( .A(n23777), .Y(n23778) );
  sky130_fd_sc_hd__inv_1 U15659 ( .A(n23797), .Y(n23798) );
  sky130_fd_sc_hd__clkinv_1 U15660 ( .A(n29165), .Y(n29472) );
  sky130_fd_sc_hd__clkinv_1 U15661 ( .A(n29163), .Y(n29471) );
  sky130_fd_sc_hd__inv_1 U15662 ( .A(n23782), .Y(n23783) );
  sky130_fd_sc_hd__clkinv_1 U15663 ( .A(n23814), .Y(n23815) );
  sky130_fd_sc_hd__clkinv_1 U15664 ( .A(n28610), .Y(n28613) );
  sky130_fd_sc_hd__clkinv_1 U15665 ( .A(n23756), .Y(n23757) );
  sky130_fd_sc_hd__clkinv_1 U15666 ( .A(n23793), .Y(n23794) );
  sky130_fd_sc_hd__inv_1 U15667 ( .A(n23803), .Y(n23804) );
  sky130_fd_sc_hd__clkinv_1 U15668 ( .A(n25540), .Y(n25541) );
  sky130_fd_sc_hd__clkinv_1 U15669 ( .A(n23809), .Y(n23810) );
  sky130_fd_sc_hd__inv_1 U15670 ( .A(n23761), .Y(n23762) );
  sky130_fd_sc_hd__clkinv_1 U15671 ( .A(n29161), .Y(n29469) );
  sky130_fd_sc_hd__o22ai_1 U15672 ( .A1(n18486), .A2(n17692), .B1(n17745), 
        .B2(n18483), .Y(n17709) );
  sky130_fd_sc_hd__clkinv_1 U15673 ( .A(n25542), .Y(n25543) );
  sky130_fd_sc_hd__clkinv_1 U15674 ( .A(n29160), .Y(n29468) );
  sky130_fd_sc_hd__clkinv_1 U15675 ( .A(n27185), .Y(n27188) );
  sky130_fd_sc_hd__clkinv_1 U15676 ( .A(n25504), .Y(n25505) );
  sky130_fd_sc_hd__clkinv_1 U15677 ( .A(n16996), .Y(n16997) );
  sky130_fd_sc_hd__clkinv_1 U15678 ( .A(n25506), .Y(n25507) );
  sky130_fd_sc_hd__clkinv_1 U15680 ( .A(n25508), .Y(n25509) );
  sky130_fd_sc_hd__clkinv_1 U15681 ( .A(n25510), .Y(n25511) );
  sky130_fd_sc_hd__clkinv_1 U15682 ( .A(n25512), .Y(n25513) );
  sky130_fd_sc_hd__clkinv_1 U15683 ( .A(n25514), .Y(n25515) );
  sky130_fd_sc_hd__clkinv_1 U15684 ( .A(n29177), .Y(n29178) );
  sky130_fd_sc_hd__clkinv_1 U15685 ( .A(n23771), .Y(n23772) );
  sky130_fd_sc_hd__clkinv_1 U15686 ( .A(n25550), .Y(n25551) );
  sky130_fd_sc_hd__clkinv_1 U15687 ( .A(n29150), .Y(n29459) );
  sky130_fd_sc_hd__clkinv_1 U15688 ( .A(n29152), .Y(n29458) );
  sky130_fd_sc_hd__clkinv_1 U15689 ( .A(n29485), .Y(n24026) );
  sky130_fd_sc_hd__clkinv_1 U15690 ( .A(n27633), .Y(n29455) );
  sky130_fd_sc_hd__clkinv_1 U15691 ( .A(n14635), .Y(n14621) );
  sky130_fd_sc_hd__clkinv_1 U15692 ( .A(n27655), .Y(n29454) );
  sky130_fd_sc_hd__clkinv_1 U15693 ( .A(n25552), .Y(n25553) );
  sky130_fd_sc_hd__clkinv_1 U15694 ( .A(n27078), .Y(n29451) );
  sky130_fd_sc_hd__clkinv_1 U15695 ( .A(n28023), .Y(n28024) );
  sky130_fd_sc_hd__clkinv_1 U15696 ( .A(n27536), .Y(n27539) );
  sky130_fd_sc_hd__clkinv_1 U15697 ( .A(n28002), .Y(n29449) );
  sky130_fd_sc_hd__clkinv_1 U15698 ( .A(n28893), .Y(n28894) );
  sky130_fd_sc_hd__clkinv_1 U15699 ( .A(n14591), .Y(n14592) );
  sky130_fd_sc_hd__clkinv_1 U15700 ( .A(n28684), .Y(n28687) );
  sky130_fd_sc_hd__clkinv_1 U15701 ( .A(n25263), .Y(n23517) );
  sky130_fd_sc_hd__clkinv_1 U15702 ( .A(n29398), .Y(n29400) );
  sky130_fd_sc_hd__clkinv_1 U15703 ( .A(n16255), .Y(n16840) );
  sky130_fd_sc_hd__clkinv_1 U15704 ( .A(n26099), .Y(n26106) );
  sky130_fd_sc_hd__clkinv_1 U15705 ( .A(n27479), .Y(n27483) );
  sky130_fd_sc_hd__clkinv_1 U15706 ( .A(n23530), .Y(n24888) );
  sky130_fd_sc_hd__clkinv_1 U15707 ( .A(n13155), .Y(n13156) );
  sky130_fd_sc_hd__clkinv_1 U15708 ( .A(n16160), .Y(n14632) );
  sky130_fd_sc_hd__clkinv_1 U15709 ( .A(n15685), .Y(n16338) );
  sky130_fd_sc_hd__clkinv_1 U15710 ( .A(n29146), .Y(n29464) );
  sky130_fd_sc_hd__clkinv_1 U15711 ( .A(n28538), .Y(n28524) );
  sky130_fd_sc_hd__clkinv_1 U15712 ( .A(n25548), .Y(n25549) );
  sky130_fd_sc_hd__clkinv_1 U15713 ( .A(n29151), .Y(n29462) );
  sky130_fd_sc_hd__clkinv_1 U15714 ( .A(n29149), .Y(n29461) );
  sky130_fd_sc_hd__nor2_2 U15715 ( .A(n21359), .B(n16985), .Y(n19124) );
  sky130_fd_sc_hd__clkinv_1 U15716 ( .A(n29153), .Y(n29460) );
  sky130_fd_sc_hd__clkinv_1 U15717 ( .A(n23766), .Y(n23767) );
  sky130_fd_sc_hd__clkinv_1 U15719 ( .A(n29158), .Y(n29466) );
  sky130_fd_sc_hd__clkinv_1 U15720 ( .A(n29148), .Y(n29463) );
  sky130_fd_sc_hd__clkinv_1 U15721 ( .A(n25546), .Y(n25547) );
  sky130_fd_sc_hd__clkinv_1 U15722 ( .A(n25544), .Y(n25545) );
  sky130_fd_sc_hd__clkinv_1 U15723 ( .A(n27251), .Y(n27252) );
  sky130_fd_sc_hd__clkinv_1 U15724 ( .A(n27210), .Y(n27212) );
  sky130_fd_sc_hd__clkinv_1 U15725 ( .A(n27537), .Y(n27532) );
  sky130_fd_sc_hd__clkinv_1 U15726 ( .A(n28859), .Y(n28850) );
  sky130_fd_sc_hd__and2_0 U15727 ( .A(n29827), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[27]), .X(n29577) );
  sky130_fd_sc_hd__clkinv_1 U15728 ( .A(n28838), .Y(n28839) );
  sky130_fd_sc_hd__o21ai_2 U15729 ( .A1(n24296), .A2(n23894), .B1(n29745), .Y(
        j202_soc_core_ahb2apb_02_N127) );
  sky130_fd_sc_hd__clkinv_1 U15730 ( .A(n24665), .Y(n24666) );
  sky130_fd_sc_hd__clkinv_1 U15731 ( .A(n29576), .Y(n26749) );
  sky130_fd_sc_hd__and2_0 U15732 ( .A(n11150), .B(n19148), .X(n17240) );
  sky130_fd_sc_hd__clkinv_1 U15733 ( .A(n15175), .Y(n15176) );
  sky130_fd_sc_hd__clkinv_1 U15734 ( .A(n26661), .Y(n26465) );
  sky130_fd_sc_hd__inv_1 U15735 ( .A(n26555), .Y(n20899) );
  sky130_fd_sc_hd__clkinv_1 U15736 ( .A(n24720), .Y(n24723) );
  sky130_fd_sc_hd__and2_0 U15737 ( .A(io_in[0]), .B(n29827), .X(n29682) );
  sky130_fd_sc_hd__clkinv_1 U15738 ( .A(n29541), .Y(n24721) );
  sky130_fd_sc_hd__clkinv_1 U15739 ( .A(n26904), .Y(n23881) );
  sky130_fd_sc_hd__clkinv_1 U15740 ( .A(n26910), .Y(n23632) );
  sky130_fd_sc_hd__clkinv_1 U15741 ( .A(n27875), .Y(n29452) );
  sky130_fd_sc_hd__clkinv_1 U15742 ( .A(n13115), .Y(n13116) );
  sky130_fd_sc_hd__clkinv_1 U15743 ( .A(n22779), .Y(n22862) );
  sky130_fd_sc_hd__clkinv_1 U15744 ( .A(n29162), .Y(n29470) );
  sky130_fd_sc_hd__nand3_2 U15745 ( .A(n20900), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_sck), .C(n26568), .Y(n28895) );
  sky130_fd_sc_hd__and2_0 U15746 ( .A(n25202), .B(n29828), .X(n23854) );
  sky130_fd_sc_hd__clkinv_1 U15747 ( .A(n25202), .Y(n25203) );
  sky130_fd_sc_hd__clkinv_1 U15748 ( .A(n26600), .Y(n26570) );
  sky130_fd_sc_hd__clkinv_1 U15749 ( .A(n24285), .Y(n13319) );
  sky130_fd_sc_hd__clkinv_1 U15750 ( .A(n25030), .Y(n25031) );
  sky130_fd_sc_hd__clkinv_1 U15751 ( .A(n19098), .Y(n21660) );
  sky130_fd_sc_hd__clkinv_1 U15752 ( .A(n26634), .Y(n23878) );
  sky130_fd_sc_hd__clkinv_1 U15753 ( .A(n28402), .Y(n24395) );
  sky130_fd_sc_hd__clkinv_1 U15754 ( .A(n23836), .Y(n23842) );
  sky130_fd_sc_hd__clkinv_1 U15755 ( .A(n29125), .Y(n29849) );
  sky130_fd_sc_hd__clkinv_1 U15756 ( .A(n26483), .Y(n27228) );
  sky130_fd_sc_hd__clkinv_1 U15757 ( .A(n27181), .Y(n27184) );
  sky130_fd_sc_hd__clkinv_1 U15758 ( .A(n28870), .Y(n27232) );
  sky130_fd_sc_hd__clkinv_1 U15759 ( .A(n26295), .Y(n26298) );
  sky130_fd_sc_hd__clkinv_1 U15760 ( .A(n26266), .Y(n26140) );
  sky130_fd_sc_hd__clkinv_1 U15761 ( .A(n23532), .Y(n26424) );
  sky130_fd_sc_hd__clkinv_1 U15762 ( .A(n25089), .Y(n25085) );
  sky130_fd_sc_hd__clkinv_1 U15763 ( .A(n25086), .Y(n29402) );
  sky130_fd_sc_hd__clkinv_1 U15764 ( .A(n26612), .Y(n26647) );
  sky130_fd_sc_hd__clkinv_1 U15765 ( .A(n27279), .Y(n26484) );
  sky130_fd_sc_hd__clkinv_1 U15766 ( .A(n18825), .Y(n25818) );
  sky130_fd_sc_hd__nor2_1 U15767 ( .A(j202_soc_core_memory0_ram_dout0_sel[11]), 
        .B(n13153), .Y(n13155) );
  sky130_fd_sc_hd__clkinv_1 U15769 ( .A(n16457), .Y(n13587) );
  sky130_fd_sc_hd__clkinv_1 U15770 ( .A(n13275), .Y(n13276) );
  sky130_fd_sc_hd__clkinv_1 U15771 ( .A(n27293), .Y(n26544) );
  sky130_fd_sc_hd__clkinv_1 U15772 ( .A(n21200), .Y(n18838) );
  sky130_fd_sc_hd__clkinv_1 U15773 ( .A(n29575), .Y(n26720) );
  sky130_fd_sc_hd__clkinv_1 U15774 ( .A(n23275), .Y(n21053) );
  sky130_fd_sc_hd__and2_0 U15775 ( .A(n29830), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]), .X(n29739) );
  sky130_fd_sc_hd__clkinv_1 U15776 ( .A(n23117), .Y(n21051) );
  sky130_fd_sc_hd__clkinv_1 U15777 ( .A(n23307), .Y(n23308) );
  sky130_fd_sc_hd__and2_0 U15778 ( .A(n29827), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]), .X(n29737) );
  sky130_fd_sc_hd__clkinv_1 U15779 ( .A(n21201), .Y(n25827) );
  sky130_fd_sc_hd__clkinv_1 U15780 ( .A(n20823), .Y(n20508) );
  sky130_fd_sc_hd__clkinv_1 U15781 ( .A(n23119), .Y(n21052) );
  sky130_fd_sc_hd__clkinv_1 U15782 ( .A(n26189), .Y(n26179) );
  sky130_fd_sc_hd__clkinv_1 U15783 ( .A(n27430), .Y(n25554) );
  sky130_fd_sc_hd__and2_0 U15784 ( .A(io_in[26]), .B(n29827), .X(n29676) );
  sky130_fd_sc_hd__clkinv_1 U15785 ( .A(n26513), .Y(n26559) );
  sky130_fd_sc_hd__and2_0 U15786 ( .A(io_in[27]), .B(n29827), .X(n29675) );
  sky130_fd_sc_hd__clkinv_1 U15787 ( .A(n29562), .Y(n25183) );
  sky130_fd_sc_hd__and2_0 U15788 ( .A(io_in[30]), .B(n29830), .X(n29672) );
  sky130_fd_sc_hd__clkinv_1 U15789 ( .A(n24284), .Y(n23626) );
  sky130_fd_sc_hd__and2_0 U15790 ( .A(io_in[36]), .B(n29827), .X(n29667) );
  sky130_fd_sc_hd__clkinv_1 U15791 ( .A(n29037), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N22) );
  sky130_fd_sc_hd__and2_0 U15792 ( .A(n29745), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[18]), .X(n29604) );
  sky130_fd_sc_hd__clkinv_1 U15793 ( .A(n26144), .Y(n25831) );
  sky130_fd_sc_hd__clkinv_1 U15794 ( .A(n24020), .Y(n23903) );
  sky130_fd_sc_hd__clkinv_1 U15795 ( .A(n27286), .Y(n26486) );
  sky130_fd_sc_hd__clkinv_1 U15796 ( .A(n27268), .Y(n23633) );
  sky130_fd_sc_hd__clkinv_1 U15797 ( .A(n27219), .Y(n26575) );
  sky130_fd_sc_hd__clkinv_1 U15798 ( .A(n28072), .Y(n20429) );
  sky130_fd_sc_hd__clkinv_1 U15799 ( .A(n27285), .Y(n27278) );
  sky130_fd_sc_hd__nor2_1 U15800 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[1]), 
        .B(n26266), .Y(n26149) );
  sky130_fd_sc_hd__clkinv_1 U15801 ( .A(n24022), .Y(n24023) );
  sky130_fd_sc_hd__and2_0 U15802 ( .A(n29827), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14]), .X(n29729) );
  sky130_fd_sc_hd__clkinv_1 U15803 ( .A(n27125), .Y(n17226) );
  sky130_fd_sc_hd__clkinv_1 U15804 ( .A(n17675), .Y(n11959) );
  sky130_fd_sc_hd__clkinv_1 U15805 ( .A(n18743), .Y(n18698) );
  sky130_fd_sc_hd__clkinv_1 U15806 ( .A(n29543), .Y(n24812) );
  sky130_fd_sc_hd__clkinv_1 U15807 ( .A(n25068), .Y(n25064) );
  sky130_fd_sc_hd__clkinv_1 U15808 ( .A(n17636), .Y(n11961) );
  sky130_fd_sc_hd__inv_1 U15809 ( .A(n24674), .Y(n24676) );
  sky130_fd_sc_hd__clkinv_1 U15810 ( .A(n29096), .Y(n29607) );
  sky130_fd_sc_hd__clkinv_1 U15811 ( .A(n29601), .Y(n28597) );
  sky130_fd_sc_hd__clkinv_1 U15813 ( .A(n13474), .Y(n13352) );
  sky130_fd_sc_hd__clkinv_1 U15814 ( .A(n18700), .Y(n19865) );
  sky130_fd_sc_hd__clkinv_1 U15815 ( .A(j202_soc_core_uart_TOP_N24), .Y(n29306) );
  sky130_fd_sc_hd__clkinv_1 U15816 ( .A(n23972), .Y(n23962) );
  sky130_fd_sc_hd__clkinv_1 U15817 ( .A(n28608), .Y(n28605) );
  sky130_fd_sc_hd__clkinv_1 U15818 ( .A(n16933), .Y(n16934) );
  sky130_fd_sc_hd__clkinv_1 U15819 ( .A(n29586), .Y(n27705) );
  sky130_fd_sc_hd__clkinv_1 U15821 ( .A(n29558), .Y(n25055) );
  sky130_fd_sc_hd__clkinv_1 U15822 ( .A(n27476), .Y(n27478) );
  sky130_fd_sc_hd__nand2_1 U15823 ( .A(n26555), .B(n28914), .Y(n10577) );
  sky130_fd_sc_hd__clkinv_1 U15824 ( .A(n29571), .Y(n26680) );
  sky130_fd_sc_hd__clkinv_1 U15825 ( .A(n29608), .Y(n29120) );
  sky130_fd_sc_hd__clkinv_1 U15826 ( .A(n29573), .Y(n26697) );
  sky130_fd_sc_hd__clkinv_1 U15827 ( .A(n29561), .Y(n25156) );
  sky130_fd_sc_hd__inv_4 U15828 ( .A(n29088), .Y(n29830) );
  sky130_fd_sc_hd__clkinv_1 U15829 ( .A(n28867), .Y(n26490) );
  sky130_fd_sc_hd__clkinv_1 U15830 ( .A(n29274), .Y(n26474) );
  sky130_fd_sc_hd__clkinv_1 U15831 ( .A(n20976), .Y(n20977) );
  sky130_fd_sc_hd__clkinv_1 U15832 ( .A(n23582), .Y(n22634) );
  sky130_fd_sc_hd__buf_4 U15833 ( .A(n17729), .X(n18496) );
  sky130_fd_sc_hd__clkinv_1 U15834 ( .A(n23294), .Y(n23296) );
  sky130_fd_sc_hd__and2_0 U15835 ( .A(io_in[33]), .B(n28914), .X(n29670) );
  sky130_fd_sc_hd__clkinv_1 U15836 ( .A(n23285), .Y(n23287) );
  sky130_fd_sc_hd__clkinv_1 U15837 ( .A(n28593), .Y(j202_soc_core_uart_TOP_N95) );
  sky130_fd_sc_hd__clkinv_1 U15838 ( .A(n26984), .Y(n24972) );
  sky130_fd_sc_hd__clkinv_1 U15839 ( .A(n23961), .Y(n15655) );
  sky130_fd_sc_hd__and2_0 U15840 ( .A(io_in[34]), .B(n29828), .X(n29669) );
  sky130_fd_sc_hd__clkinv_1 U15841 ( .A(n28722), .Y(n28717) );
  sky130_fd_sc_hd__clkinv_1 U15842 ( .A(n23871), .Y(n26543) );
  sky130_fd_sc_hd__clkinv_1 U15843 ( .A(n25316), .Y(n25317) );
  sky130_fd_sc_hd__clkinv_1 U15844 ( .A(n26268), .Y(n18828) );
  sky130_fd_sc_hd__nor2_1 U15845 ( .A(j202_soc_core_qspi_wb_ack), .B(n28866), 
        .Y(n26555) );
  sky130_fd_sc_hd__clkinv_1 U15846 ( .A(n26264), .Y(n22117) );
  sky130_fd_sc_hd__clkinv_1 U15847 ( .A(n26532), .Y(n23861) );
  sky130_fd_sc_hd__buf_4 U15848 ( .A(n17339), .X(n18989) );
  sky130_fd_sc_hd__inv_2 U15849 ( .A(n14597), .Y(n19148) );
  sky130_fd_sc_hd__and2_0 U15850 ( .A(n29828), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13]), .X(n29738) );
  sky130_fd_sc_hd__clkinv_1 U15851 ( .A(n20930), .Y(n20931) );
  sky130_fd_sc_hd__clkinv_1 U15852 ( .A(n23807), .Y(n23835) );
  sky130_fd_sc_hd__inv_4 U15853 ( .A(n29088), .Y(n29827) );
  sky130_fd_sc_hd__and2_0 U15854 ( .A(io_in[4]), .B(n28914), .X(n29678) );
  sky130_fd_sc_hd__clkinv_1 U15855 ( .A(n29411), .Y(n29401) );
  sky130_fd_sc_hd__clkinv_1 U15856 ( .A(n18794), .Y(n18795) );
  sky130_fd_sc_hd__clkinv_1 U15857 ( .A(n20445), .Y(n21781) );
  sky130_fd_sc_hd__clkinv_1 U15858 ( .A(n25802), .Y(n26345) );
  sky130_fd_sc_hd__clkinv_1 U15859 ( .A(n28594), .Y(n24261) );
  sky130_fd_sc_hd__clkinv_1 U15860 ( .A(n28840), .Y(n27284) );
  sky130_fd_sc_hd__nand2b_1 U15861 ( .A_N(n12298), .B(n13147), .Y(n11987) );
  sky130_fd_sc_hd__clkinv_1 U15862 ( .A(n13151), .Y(n13149) );
  sky130_fd_sc_hd__clkinv_1 U15863 ( .A(n25073), .Y(n25066) );
  sky130_fd_sc_hd__clkinv_1 U15864 ( .A(n26899), .Y(n23894) );
  sky130_fd_sc_hd__clkinv_1 U15865 ( .A(n23169), .Y(n23170) );
  sky130_fd_sc_hd__clkinv_1 U15866 ( .A(n28603), .Y(n28606) );
  sky130_fd_sc_hd__clkinv_1 U15867 ( .A(n24454), .Y(n24465) );
  sky130_fd_sc_hd__buf_4 U15869 ( .A(n17443), .X(n18486) );
  sky130_fd_sc_hd__clkinv_1 U15870 ( .A(n26208), .Y(n26145) );
  sky130_fd_sc_hd__clkinv_1 U15871 ( .A(n18827), .Y(n26148) );
  sky130_fd_sc_hd__inv_2 U15872 ( .A(n21219), .Y(n18115) );
  sky130_fd_sc_hd__clkinv_1 U15873 ( .A(n23093), .Y(n23094) );
  sky130_fd_sc_hd__clkinv_1 U15874 ( .A(n26094), .Y(n26096) );
  sky130_fd_sc_hd__clkinv_1 U15875 ( .A(n23065), .Y(n23066) );
  sky130_fd_sc_hd__inv_2 U15876 ( .A(n24366), .Y(n18098) );
  sky130_fd_sc_hd__clkinv_1 U15877 ( .A(n24829), .Y(n22770) );
  sky130_fd_sc_hd__clkinv_1 U15878 ( .A(n15649), .Y(n15650) );
  sky130_fd_sc_hd__clkinv_1 U15879 ( .A(n27264), .Y(n26521) );
  sky130_fd_sc_hd__clkinv_1 U15880 ( .A(n23192), .Y(n23193) );
  sky130_fd_sc_hd__clkinv_1 U15881 ( .A(n13428), .Y(n13302) );
  sky130_fd_sc_hd__clkinv_1 U15882 ( .A(n23341), .Y(n23342) );
  sky130_fd_sc_hd__and2_0 U15883 ( .A(n29828), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]), .X(n29734) );
  sky130_fd_sc_hd__clkinv_1 U15884 ( .A(n25205), .Y(n27287) );
  sky130_fd_sc_hd__clkinv_1 U15885 ( .A(n22299), .Y(n17758) );
  sky130_fd_sc_hd__and2_0 U15886 ( .A(n29828), .B(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .X(n20900) );
  sky130_fd_sc_hd__clkinv_1 U15887 ( .A(n28914), .Y(n12084) );
  sky130_fd_sc_hd__clkinv_1 U15888 ( .A(n17350), .Y(n13324) );
  sky130_fd_sc_hd__clkinv_1 U15889 ( .A(n13174), .Y(n13175) );
  sky130_fd_sc_hd__clkinv_1 U15890 ( .A(j202_soc_core_j22_cpu_rf_gpr[27]), .Y(
        n15936) );
  sky130_fd_sc_hd__clkinv_1 U15891 ( .A(j202_soc_core_j22_cpu_rf_vbr[25]), .Y(
        n15885) );
  sky130_fd_sc_hd__clkinv_1 U15892 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__1_), 
        .Y(n23770) );
  sky130_fd_sc_hd__clkinv_1 U15893 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[121]), .Y(n27564) );
  sky130_fd_sc_hd__clkinv_1 U15894 ( .A(j202_soc_core_j22_cpu_rf_gpr[16]), .Y(
        n14536) );
  sky130_fd_sc_hd__clkinv_1 U15895 ( .A(j202_soc_core_cmt_core_00_cks0[1]), 
        .Y(n24007) );
  sky130_fd_sc_hd__clkinv_1 U15897 ( .A(j202_soc_core_uart_sio_ce), .Y(n29099)
         );
  sky130_fd_sc_hd__clkinv_1 U15898 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[26]), .Y(n26809) );
  sky130_fd_sc_hd__clkinv_1 U15899 ( .A(j202_soc_core_j22_cpu_rf_vbr[2]), .Y(
        n19270) );
  sky130_fd_sc_hd__clkinv_1 U15900 ( .A(j202_soc_core_j22_cpu_rf_vbr[16]), .Y(
        n14533) );
  sky130_fd_sc_hd__clkinv_1 U15901 ( .A(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[2]), .Y(n17202) );
  sky130_fd_sc_hd__clkinv_1 U15902 ( .A(j202_soc_core_intc_core_00_rg_ipr[103]), .Y(n27561) );
  sky130_fd_sc_hd__clkinv_1 U15903 ( .A(j202_soc_core_uart_TOP_rx_fifo_gb), 
        .Y(n23896) );
  sky130_fd_sc_hd__clkinv_1 U15904 ( .A(j202_soc_core_j22_cpu_memop_MEM__0_), 
        .Y(n24587) );
  sky130_fd_sc_hd__clkinv_1 U15905 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[29]), .Y(n29260) );
  sky130_fd_sc_hd__clkinv_1 U15906 ( .A(j202_soc_core_ahb2apb_00_state[2]), 
        .Y(n24725) );
  sky130_fd_sc_hd__clkinv_1 U15907 ( .A(j202_soc_core_j22_cpu_rf_tmp[16]), .Y(
        n14534) );
  sky130_fd_sc_hd__clkinv_1 U15908 ( .A(j202_soc_core_j22_cpu_pc[1]), .Y(
        n24792) );
  sky130_fd_sc_hd__clkinv_1 U15909 ( .A(j202_soc_core_intc_core_00_rg_ipr[98]), 
        .Y(n28181) );
  sky130_fd_sc_hd__clkinv_1 U15910 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[7]), .Y(n23663) );
  sky130_fd_sc_hd__clkinv_1 U15911 ( .A(j202_soc_core_j22_cpu_pc[25]), .Y(
        n22905) );
  sky130_fd_sc_hd__clkinv_1 U15912 ( .A(j202_soc_core_cmt_core_00_cnt1[11]), 
        .Y(n26989) );
  sky130_fd_sc_hd__clkinv_1 U15913 ( .A(gpio_en_o[16]), .Y(io_oeb[36]) );
  sky130_fd_sc_hd__clkinv_1 U15914 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__3_), 
        .Y(n23752) );
  sky130_fd_sc_hd__clkinv_1 U15915 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[103]), .Y(n17306) );
  sky130_fd_sc_hd__clkinv_1 U15916 ( .A(j202_soc_core_j22_cpu_rf_gbr[15]), .Y(
        n14565) );
  sky130_fd_sc_hd__clkinv_1 U15917 ( .A(j202_soc_core_j22_cpu_rf_pr[3]), .Y(
        n21244) );
  sky130_fd_sc_hd__clkinv_1 U15918 ( .A(j202_soc_core_j22_cpu_rf_pr[25]), .Y(
        n15889) );
  sky130_fd_sc_hd__buf_4 U15919 ( .A(j202_soc_core_j22_cpu_ml_bufa[3]), .X(
        n21219) );
  sky130_fd_sc_hd__clkinv_1 U15920 ( .A(j202_soc_core_j22_cpu_memop_Ma__1_), 
        .Y(n13443) );
  sky130_fd_sc_hd__clkinv_1 U15921 ( .A(j202_soc_core_intc_core_00_rg_itgt[57]), .Y(n27420) );
  sky130_fd_sc_hd__clkinv_1 U15922 ( .A(j202_soc_core_j22_cpu_rf_gpr[9]), .Y(
        n14310) );
  sky130_fd_sc_hd__clkinv_1 U15923 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[71]), .Y(n17307) );
  sky130_fd_sc_hd__clkinv_1 U15924 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .Y(n24199) );
  sky130_fd_sc_hd__clkinv_1 U15925 ( .A(j202_soc_core_j22_cpu_regop_imm__1_), 
        .Y(n13883) );
  sky130_fd_sc_hd__clkinv_1 U15926 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[31]), .Y(n26782) );
  sky130_fd_sc_hd__clkinv_1 U15927 ( .A(j202_soc_core_j22_cpu_rf_pr[15]), .Y(
        n18891) );
  sky130_fd_sc_hd__clkinv_1 U15928 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[6]), .Y(n23666) );
  sky130_fd_sc_hd__clkinv_1 U15929 ( .A(j202_soc_core_j22_cpu_rf_tmp[15]), .Y(
        n18896) );
  sky130_fd_sc_hd__clkinv_1 U15930 ( .A(j202_soc_core_j22_cpu_rf_gpr[21]), .Y(
        n14998) );
  sky130_fd_sc_hd__clkinv_1 U15931 ( .A(j202_soc_core_j22_cpu_ml_macl[26]), 
        .Y(n22655) );
  sky130_fd_sc_hd__clkinv_1 U15932 ( .A(j202_soc_core_uart_TOP_rx_fifo_wp[0]), 
        .Y(n27955) );
  sky130_fd_sc_hd__clkinv_1 U15933 ( .A(j202_soc_core_j22_cpu_regop_imm__10_), 
        .Y(n13978) );
  sky130_fd_sc_hd__clkinv_1 U15934 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[3]), .Y(n27680) );
  sky130_fd_sc_hd__clkinv_1 U15935 ( .A(j202_soc_core_intc_core_00_rg_ipr[101]), .Y(n27412) );
  sky130_fd_sc_hd__clkinv_1 U15936 ( .A(j202_soc_core_j22_cpu_rf_gbr[25]), .Y(
        n22904) );
  sky130_fd_sc_hd__clkinv_1 U15937 ( .A(j202_soc_core_j22_cpu_rf_vbr[15]), .Y(
        n18895) );
  sky130_fd_sc_hd__clkinv_1 U15938 ( .A(j202_soc_core_j22_cpu_ml_macl[10]), 
        .Y(n19281) );
  sky130_fd_sc_hd__clkinv_1 U15939 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[0]), 
        .Y(n29172) );
  sky130_fd_sc_hd__clkinv_1 U15940 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__2_), 
        .Y(n23775) );
  sky130_fd_sc_hd__clkinv_1 U15941 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[23]), .Y(n26824) );
  sky130_fd_sc_hd__clkinv_1 U15942 ( .A(j202_soc_core_j22_cpu_ma_M_area[1]), 
        .Y(n13260) );
  sky130_fd_sc_hd__clkinv_1 U15943 ( .A(j202_soc_core_j22_cpu_ml_macl[6]), .Y(
        n22131) );
  sky130_fd_sc_hd__clkinv_1 U15944 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[11]), .Y(n27000) );
  sky130_fd_sc_hd__clkinv_1 U15945 ( .A(j202_soc_core_intc_core_00_rg_itgt[25]), .Y(n27499) );
  sky130_fd_sc_hd__clkinv_1 U15946 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd), .Y(n28726) );
  sky130_fd_sc_hd__clkinv_1 U15947 ( .A(j202_soc_core_intc_core_00_rg_ipr[88]), 
        .Y(n27654) );
  sky130_fd_sc_hd__clkinv_1 U15948 ( .A(j202_soc_core_j22_cpu_ml_mach[29]), 
        .Y(n22479) );
  sky130_fd_sc_hd__clkinv_1 U15949 ( .A(j202_soc_core_j22_cpu_rf_gpr[491]), 
        .Y(n21884) );
  sky130_fd_sc_hd__clkinv_1 U15950 ( .A(j202_soc_core_qspi_wb_addr[5]), .Y(
        n28737) );
  sky130_fd_sc_hd__clkinv_1 U15951 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[7]), .Y(n27558) );
  sky130_fd_sc_hd__clkinv_1 U15952 ( .A(j202_soc_core_j22_cpu_rf_tmp[1]), .Y(
        n21987) );
  sky130_fd_sc_hd__inv_4 U15953 ( .A(j202_soc_core_rst), .Y(n29828) );
  sky130_fd_sc_hd__clkinv_1 U15954 ( .A(j202_soc_core_j22_cpu_rf_vbr[22]), .Y(
        n15027) );
  sky130_fd_sc_hd__clkinv_1 U15955 ( .A(j202_soc_core_j22_cpu_rf_tmp[22]), .Y(
        n15028) );
  sky130_fd_sc_hd__clkinv_1 U15956 ( .A(j202_soc_core_j22_cpu_rf_gpr[30]), .Y(
        n16445) );
  sky130_fd_sc_hd__clkinv_1 U15958 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[4]), .Y(n27495) );
  sky130_fd_sc_hd__clkinv_1 U15959 ( .A(j202_soc_core_j22_cpu_rf_gpr[501]), 
        .Y(n15026) );
  sky130_fd_sc_hd__clkinv_1 U15960 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[21]), .Y(n26843) );
  sky130_fd_sc_hd__clkinv_1 U15961 ( .A(j202_soc_core_intc_core_00_rg_ipr[87]), 
        .Y(n27630) );
  sky130_fd_sc_hd__clkinv_1 U15962 ( .A(j202_soc_core_j22_cpu_ma_M_address[0]), 
        .Y(n19115) );
  sky130_fd_sc_hd__clkinv_1 U15963 ( .A(j202_soc_core_j22_cpu_ml_macl[22]), 
        .Y(n22148) );
  sky130_fd_sc_hd__clkinv_1 U15964 ( .A(j202_soc_core_bldc_core_00_wdata[2]), 
        .Y(n28178) );
  sky130_fd_sc_hd__clkinv_1 U15965 ( .A(j202_soc_core_j22_cpu_rf_tmp[12]), .Y(
        n14062) );
  sky130_fd_sc_hd__clkinv_1 U15966 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[6]), .Y(n29067) );
  sky130_fd_sc_hd__clkinv_1 U15967 ( .A(j202_soc_core_j22_cpu_rf_gpr[497]), 
        .Y(n13427) );
  sky130_fd_sc_hd__clkinv_1 U15968 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[4]), .Y(n29069) );
  sky130_fd_sc_hd__clkinv_1 U15969 ( .A(j202_soc_core_j22_cpu_ml_mach[8]), .Y(
        n21745) );
  sky130_fd_sc_hd__clkinv_1 U15970 ( .A(j202_soc_core_intc_core_00_rg_itgt[71]), .Y(n27995) );
  sky130_fd_sc_hd__clkinv_1 U15971 ( .A(j202_soc_core_intc_core_00_rg_ipr[86]), 
        .Y(n25611) );
  sky130_fd_sc_hd__clkinv_1 U15972 ( .A(
        j202_soc_core_bldc_core_00_pwm_duty[11]), .Y(n27622) );
  sky130_fd_sc_hd__clkinv_1 U15973 ( .A(j202_soc_core_intc_core_00_rg_itgt[37]), .Y(n25573) );
  sky130_fd_sc_hd__clkinv_1 U15974 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[15]), .Y(n23655) );
  sky130_fd_sc_hd__clkinv_1 U15975 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]), .Y(n26674) );
  sky130_fd_sc_hd__clkinv_1 U15976 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .Y(n23724) );
  sky130_fd_sc_hd__clkinv_1 U15977 ( .A(j202_soc_core_bldc_core_00_wdata[0]), 
        .Y(n28209) );
  sky130_fd_sc_hd__clkinv_1 U15978 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]), .Y(n23717) );
  sky130_fd_sc_hd__clkinv_1 U15979 ( .A(j202_soc_core_bldc_core_00_wdata[1]), 
        .Y(n28282) );
  sky130_fd_sc_hd__inv_2 U15980 ( .A(n12030), .Y(n12031) );
  sky130_fd_sc_hd__clkinv_1 U15981 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[24]), .Y(n29051) );
  sky130_fd_sc_hd__clkinv_1 U15982 ( .A(j202_soc_core_j22_cpu_rf_tmp[18]), .Y(
        n13433) );
  sky130_fd_sc_hd__clkinv_1 U15983 ( .A(j202_soc_core_j22_cpu_ifetchl), .Y(
        n24711) );
  sky130_fd_sc_hd__clkinv_1 U15984 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .Y(n27349) );
  sky130_fd_sc_hd__clkinv_1 U15985 ( .A(j202_soc_core_intc_core_00_rg_itgt[70]), .Y(n27868) );
  sky130_fd_sc_hd__clkinv_1 U15987 ( .A(j202_soc_core_j22_cpu_intack), .Y(
        n22013) );
  sky130_fd_sc_hd__clkinv_1 U15988 ( .A(j202_soc_core_intc_core_00_rg_ipr[85]), 
        .Y(n25579) );
  sky130_fd_sc_hd__clkinv_1 U15989 ( .A(j202_soc_core_j22_cpu_rf_pr[6]), .Y(
        n22152) );
  sky130_fd_sc_hd__inv_2 U15990 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), 
        .Y(n17355) );
  sky130_fd_sc_hd__clkinv_1 U15991 ( .A(j202_soc_core_j22_cpu_rf_vbr[18]), .Y(
        n13432) );
  sky130_fd_sc_hd__clkinv_1 U15992 ( .A(j202_soc_core_intc_core_00_rg_ie[14]), 
        .Y(n26753) );
  sky130_fd_sc_hd__clkinv_1 U15993 ( .A(j202_soc_core_intc_core_00_rg_itgt[69]), .Y(n25606) );
  sky130_fd_sc_hd__clkinv_1 U15994 ( .A(j202_soc_core_qspi_wb_wdat[15]), .Y(
        n29006) );
  sky130_fd_sc_hd__clkinv_1 U15995 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[21]), .Y(n26841) );
  sky130_fd_sc_hd__clkinv_1 U15996 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[0]), 
        .Y(n29278) );
  sky130_fd_sc_hd__clkinv_1 U15997 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[9]), .Y(n28911) );
  sky130_fd_sc_hd__clkinv_1 U15998 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[3]), .Y(n13263) );
  sky130_fd_sc_hd__clkinv_1 U15999 ( .A(j202_soc_core_intc_core_00_rg_ipr[84]), 
        .Y(n27369) );
  sky130_fd_sc_hd__clkinv_1 U16000 ( .A(j202_soc_core_cmt_core_00_str1), .Y(
        n28285) );
  sky130_fd_sc_hd__clkinv_1 U16001 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[0]), .Y(n28683) );
  sky130_fd_sc_hd__clkinv_1 U16002 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[101]), .Y(n27626) );
  sky130_fd_sc_hd__clkinv_1 U16003 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[1]), 
        .Y(n24000) );
  sky130_fd_sc_hd__clkinv_1 U16004 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[3]), .Y(n26478) );
  sky130_fd_sc_hd__clkinv_1 U16005 ( .A(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_wen), .Y(
        n27701) );
  sky130_fd_sc_hd__clkinv_1 U16006 ( .A(j202_soc_core_qspi_wb_wdat[25]), .Y(
        n27164) );
  sky130_fd_sc_hd__clkinv_1 U16007 ( .A(j202_soc_core_intc_core_00_rg_ipr[82]), 
        .Y(n26859) );
  sky130_fd_sc_hd__clkinv_1 U16008 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[15]), .Y(n29012) );
  sky130_fd_sc_hd__clkinv_1 U16009 ( .A(j202_soc_core_j22_cpu_ml_mach[22]), 
        .Y(n22014) );
  sky130_fd_sc_hd__clkinv_1 U16010 ( .A(j202_soc_core_j22_cpu_ml_mach[21]), 
        .Y(n22019) );
  sky130_fd_sc_hd__clkinv_1 U16011 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[3]), .Y(n28703) );
  sky130_fd_sc_hd__inv_2 U16012 ( .A(n12036), .Y(n12037) );
  sky130_fd_sc_hd__clkinv_1 U16013 ( .A(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[1]), .Y(n21050) );
  sky130_fd_sc_hd__clkinv_1 U16014 ( .A(j202_soc_core_uart_TOP_load), .Y(
        n24271) );
  sky130_fd_sc_hd__clkinv_1 U16015 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[27]), .Y(n29130) );
  sky130_fd_sc_hd__clkinv_1 U16016 ( .A(j202_soc_core_j22_cpu_rf_tmp[25]), .Y(
        n15887) );
  sky130_fd_sc_hd__clkinv_1 U16017 ( .A(j202_soc_core_j22_cpu_ml_mach[6]), .Y(
        n22112) );
  sky130_fd_sc_hd__clkinv_1 U16018 ( .A(j202_soc_core_intc_core_00_rg_itgt[88]), .Y(n28185) );
  sky130_fd_sc_hd__clkinv_1 U16019 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[4]), .Y(n13261) );
  sky130_fd_sc_hd__clkinv_1 U16020 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]), .Y(n13321) );
  sky130_fd_sc_hd__clkinv_1 U16021 ( .A(j202_soc_core_qspi_wb_wdat[13]), .Y(
        n28992) );
  sky130_fd_sc_hd__clkinv_1 U16022 ( .A(j202_soc_core_j22_cpu_ml_mach[23]), 
        .Y(n22015) );
  sky130_fd_sc_hd__clkinv_1 U16023 ( .A(j202_soc_core_j22_cpu_ml_mach[14]), 
        .Y(n24455) );
  sky130_fd_sc_hd__clkinv_1 U16024 ( .A(j202_soc_core_intc_core_00_rg_ipr[95]), 
        .Y(n27598) );
  sky130_fd_sc_hd__clkinv_1 U16025 ( .A(j202_soc_core_cmt_core_00_cnt1[9]), 
        .Y(n26988) );
  sky130_fd_sc_hd__clkinv_1 U16026 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[23]), .Y(n26830) );
  sky130_fd_sc_hd__clkinv_1 U16027 ( .A(j202_soc_core_j22_cpu_rf_gpr[29]), .Y(
        n16080) );
  sky130_fd_sc_hd__clkinv_1 U16028 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .Y(n13320) );
  sky130_fd_sc_hd__clkinv_1 U16029 ( .A(j202_soc_core_j22_cpu_ml_mach[30]), 
        .Y(n22475) );
  sky130_fd_sc_hd__clkinv_1 U16030 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[41]), .Y(n20619) );
  sky130_fd_sc_hd__clkinv_1 U16031 ( .A(j202_soc_core_intc_core_00_rg_itgt[31]), .Y(n27397) );
  sky130_fd_sc_hd__clkinv_1 U16032 ( .A(j202_soc_core_j22_cpu_ml_macl[7]), .Y(
        n18836) );
  sky130_fd_sc_hd__clkinv_1 U16033 ( .A(j202_soc_core_intc_core_00_rg_ipr[94]), 
        .Y(n27999) );
  sky130_fd_sc_hd__clkinv_1 U16035 ( .A(j202_soc_core_j22_cpu_rf_gpr[23]), .Y(
        n14799) );
  sky130_fd_sc_hd__clkinv_1 U16036 ( .A(j202_soc_core_intc_core_00_rg_ipr[92]), 
        .Y(n27394) );
  sky130_fd_sc_hd__clkinv_1 U16037 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]), .Y(n23731) );
  sky130_fd_sc_hd__clkinv_1 U16038 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[10]), .Y(n28912) );
  sky130_fd_sc_hd__clkinv_1 U16039 ( .A(j202_soc_core_qspi_wb_addr[8]), .Y(
        n28782) );
  sky130_fd_sc_hd__clkinv_1 U16040 ( .A(j202_soc_core_j22_cpu_macop_MAC_[3]), 
        .Y(n28042) );
  sky130_fd_sc_hd__clkinv_1 U16041 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[22]), .Y(n26836) );
  sky130_fd_sc_hd__clkinv_1 U16042 ( .A(j202_soc_core_intc_core_00_rg_itgt[30]), .Y(n27659) );
  sky130_fd_sc_hd__clkinv_1 U16043 ( .A(j202_soc_core_j22_cpu_macop_MAC_[2]), 
        .Y(n28424) );
  sky130_fd_sc_hd__clkinv_1 U16044 ( .A(j202_soc_core_aquc_WE_), .Y(n25034) );
  sky130_fd_sc_hd__clkinv_1 U16046 ( .A(j202_soc_core_intc_core_00_rg_ipr[91]), 
        .Y(n27075) );
  sky130_fd_sc_hd__clkinv_1 U16047 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[13]), .Y(n28998) );
  sky130_fd_sc_hd__clkinv_1 U16048 ( .A(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[1]), .Y(n22759) );
  sky130_fd_sc_hd__clkinv_1 U16049 ( .A(j202_soc_core_j22_cpu_ml_macl[23]), 
        .Y(n22081) );
  sky130_fd_sc_hd__clkinv_1 U16050 ( .A(j202_soc_core_wbqspiflash_00_state[3]), 
        .Y(n27224) );
  sky130_fd_sc_hd__clkinv_1 U16051 ( .A(
        j202_soc_core_bldc_core_00_pwm_duty[10]), .Y(n25624) );
  sky130_fd_sc_hd__clkinv_1 U16052 ( .A(j202_soc_core_bldc_core_00_pwm_duty[0]), .Y(n25182) );
  sky130_fd_sc_hd__clkinv_1 U16053 ( .A(j202_soc_core_bldc_core_00_pwm_duty[9]), .Y(n25570) );
  sky130_fd_sc_hd__clkinv_1 U16054 ( .A(j202_soc_core_qspi_wb_wdat[31]), .Y(
        n27593) );
  sky130_fd_sc_hd__clkinv_1 U16055 ( .A(j202_soc_core_bldc_core_00_pwm_duty[8]), .Y(n27381) );
  sky130_fd_sc_hd__clkinv_1 U16056 ( .A(
        j202_soc_core_wbqspiflash_00_w_qspi_sck), .Y(n29183) );
  sky130_fd_sc_hd__clkinv_1 U16057 ( .A(j202_soc_core_j22_cpu_rf_gbr[2]), .Y(
        n13915) );
  sky130_fd_sc_hd__clkinv_1 U16058 ( .A(j202_soc_core_intc_core_00_rg_itgt[26]), .Y(n27971) );
  sky130_fd_sc_hd__clkinv_1 U16059 ( .A(j202_soc_core_j22_cpu_ml_mach[28]), 
        .Y(n22484) );
  sky130_fd_sc_hd__clkinv_1 U16061 ( .A(j202_soc_core_bldc_core_00_pwm_duty[6]), .Y(n27143) );
  sky130_fd_sc_hd__clkinv_1 U16062 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[8]), .Y(n23657) );
  sky130_fd_sc_hd__clkinv_1 U16063 ( .A(j202_soc_core_intc_core_00_rg_itgt[24]), .Y(n28234) );
  sky130_fd_sc_hd__clkinv_1 U16064 ( .A(j202_soc_core_bldc_core_00_pwm_duty[3]), .Y(n26113) );
  sky130_fd_sc_hd__clkinv_1 U16065 ( .A(j202_soc_core_j22_cpu_rf_gpr[28]), .Y(
        n15912) );
  sky130_fd_sc_hd__clkinv_1 U16066 ( .A(j202_soc_core_bldc_core_00_pwm_duty[2]), .Y(n26879) );
  sky130_fd_sc_hd__clkinv_1 U16067 ( .A(j202_soc_core_intc_core_00_rg_ipr[90]), 
        .Y(n27872) );
  sky130_fd_sc_hd__clkinv_1 U16068 ( .A(j202_soc_core_bldc_core_00_pwm_duty[1]), .Y(n25782) );
  sky130_fd_sc_hd__clkinv_1 U16069 ( .A(j202_soc_core_intc_core_00_rg_itgt[68]), .Y(n27129) );
  sky130_fd_sc_hd__clkinv_1 U16070 ( .A(j202_soc_core_intc_core_00_rg_itgt[29]), .Y(n27371) );
  sky130_fd_sc_hd__inv_2 U16071 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[4]), 
        .Y(n18831) );
  sky130_fd_sc_hd__clkinv_1 U16072 ( .A(j202_soc_core_j22_cpu_rfuo_sr__s_), 
        .Y(n24668) );
  sky130_fd_sc_hd__clkinv_1 U16073 ( .A(j202_soc_core_j22_cpu_rf_gpr[8]), .Y(
        n14259) );
  sky130_fd_sc_hd__clkinv_1 U16074 ( .A(j202_soc_core_cmt_core_00_reg_addr[3]), 
        .Y(n28221) );
  sky130_fd_sc_hd__clkinv_1 U16075 ( .A(j202_soc_core_j22_cpu_ml_mach[4]), .Y(
        n17720) );
  sky130_fd_sc_hd__clkinv_1 U16076 ( .A(j202_soc_core_j22_cpu_rf_tmp[31]), .Y(
        n16486) );
  sky130_fd_sc_hd__clkinv_1 U16077 ( .A(j202_soc_core_intc_core_00_rg_itgt[19]), .Y(n25193) );
  sky130_fd_sc_hd__clkinv_1 U16078 ( .A(j202_soc_core_j22_cpu_rf_pr[9]), .Y(
        n22892) );
  sky130_fd_sc_hd__clkinv_1 U16079 ( .A(j202_soc_core_intc_core_00_rg_itgt[6]), 
        .Y(n26703) );
  sky130_fd_sc_hd__clkinv_1 U16080 ( .A(j202_soc_core_uart_TOP_dpll_state[1]), 
        .Y(n23047) );
  sky130_fd_sc_hd__clkinv_1 U16081 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[0]), .Y(n28218) );
  sky130_fd_sc_hd__clkinv_1 U16082 ( .A(j202_soc_core_intc_core_00_rg_itgt[41]), .Y(n27411) );
  sky130_fd_sc_hd__clkinv_1 U16083 ( .A(j202_soc_core_aquc_ADR__1_), .Y(n13267) );
  sky130_fd_sc_hd__clkinv_1 U16084 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[1]), .Y(n25736) );
  sky130_fd_sc_hd__clkinv_1 U16085 ( .A(j202_soc_core_j22_cpu_ml_macl[3]), .Y(
        n21221) );
  sky130_fd_sc_hd__clkinv_1 U16086 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[24]), .Y(n29135) );
  sky130_fd_sc_hd__clkinv_1 U16087 ( .A(j202_soc_core_j22_cpu_ml_macl[4]), .Y(
        n21849) );
  sky130_fd_sc_hd__clkinv_1 U16088 ( .A(j202_soc_core_intc_core_00_rg_itgt[27]), .Y(n25194) );
  sky130_fd_sc_hd__clkinv_1 U16089 ( .A(j202_soc_core_intc_core_00_rg_itgt[16]), .Y(n26765) );
  sky130_fd_sc_hd__clkinv_1 U16090 ( .A(j202_soc_core_j22_cpu_rf_gpr[22]), .Y(
        n14834) );
  sky130_fd_sc_hd__clkinv_1 U16091 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]), .Y(n23691) );
  sky130_fd_sc_hd__clkinv_1 U16092 ( .A(j202_soc_core_j22_cpu_rf_pr[2]), .Y(
        n19266) );
  sky130_fd_sc_hd__clkinv_1 U16093 ( .A(j202_soc_core_intc_core_00_rg_itgt[18]), .Y(n26858) );
  sky130_fd_sc_hd__clkinv_1 U16094 ( .A(j202_soc_core_j22_cpu_rf_vbr[26]), .Y(
        n15853) );
  sky130_fd_sc_hd__clkinv_1 U16095 ( .A(j202_soc_core_qspi_wb_wdat[0]), .Y(
        n28900) );
  sky130_fd_sc_hd__clkinv_1 U16096 ( .A(j202_soc_core_j22_cpu_ml_macl[19]), 
        .Y(n22815) );
  sky130_fd_sc_hd__clkinv_1 U16097 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[2]), .Y(n28171) );
  sky130_fd_sc_hd__clkinv_1 U16098 ( .A(j202_soc_core_j22_cpu_rf_gpr[25]), .Y(
        n15888) );
  sky130_fd_sc_hd__clkinv_1 U16099 ( .A(j202_soc_core_intc_core_00_rg_itgt[7]), 
        .Y(n26695) );
  sky130_fd_sc_hd__clkinv_1 U16100 ( .A(j202_soc_core_j22_cpu_rf_tmp[26]), .Y(
        n15854) );
  sky130_fd_sc_hd__clkinv_1 U16101 ( .A(j202_soc_core_aquc_ADR__2_), .Y(n13266) );
  sky130_fd_sc_hd__clkinv_1 U16102 ( .A(j202_soc_core_intc_core_00_rg_ipr[38]), 
        .Y(n26710) );
  sky130_fd_sc_hd__clkinv_1 U16103 ( .A(j202_soc_core_j22_cpu_rf_vbr[31]), .Y(
        n16485) );
  sky130_fd_sc_hd__clkinv_1 U16104 ( .A(j202_soc_core_j22_cpu_opst[3]), .Y(
        n20428) );
  sky130_fd_sc_hd__clkinv_1 U16105 ( .A(j202_soc_core_j22_cpu_rf_gpr[505]), 
        .Y(n15852) );
  sky130_fd_sc_hd__clkinv_1 U16106 ( .A(j202_soc_core_j22_cpu_rf_gpr[490]), 
        .Y(n21292) );
  sky130_fd_sc_hd__clkinv_1 U16107 ( .A(j202_soc_core_intc_core_00_rg_itgt[72]), .Y(n28180) );
  sky130_fd_sc_hd__clkinv_1 U16108 ( .A(j202_soc_core_j22_cpu_ml_macl[24]), 
        .Y(n18179) );
  sky130_fd_sc_hd__clkinv_1 U16109 ( .A(j202_soc_core_uart_TOP_dpll_state[0]), 
        .Y(n29092) );
  sky130_fd_sc_hd__clkinv_1 U16110 ( .A(j202_soc_core_intc_core_00_rg_itgt[80]), .Y(n28183) );
  sky130_fd_sc_hd__clkinv_1 U16111 ( .A(j202_soc_core_j22_cpu_istall), .Y(
        n15646) );
  sky130_fd_sc_hd__clkinv_1 U16112 ( .A(j202_soc_core_qspi_wb_addr[7]), .Y(
        n28748) );
  sky130_fd_sc_hd__clkinv_1 U16113 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[13]), .Y(n23688) );
  sky130_fd_sc_hd__clkinv_1 U16114 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16]), .Y(n29013) );
  sky130_fd_sc_hd__clkinv_1 U16115 ( .A(j202_soc_core_cmt_core_00_cnt1[2]), 
        .Y(n27524) );
  sky130_fd_sc_hd__clkinv_1 U16116 ( .A(j202_soc_core_j22_cpu_rf_gpr[31]), .Y(
        n16489) );
  sky130_fd_sc_hd__clkinv_1 U16117 ( .A(j202_soc_core_intc_core_00_rg_itgt[15]), .Y(n26743) );
  sky130_fd_sc_hd__clkinv_1 U16118 ( .A(j202_soc_core_j22_cpu_rf_gpr[488]), 
        .Y(n22891) );
  sky130_fd_sc_hd__clkinv_1 U16119 ( .A(j202_soc_core_j22_cpu_ml_macl[15]), 
        .Y(n18888) );
  sky130_fd_sc_hd__clkinv_1 U16120 ( .A(j202_soc_core_intc_core_00_rg_itgt[14]), .Y(n26745) );
  sky130_fd_sc_hd__clkinv_1 U16121 ( .A(j202_soc_core_j22_cpu_rf_gpr[503]), 
        .Y(n14774) );
  sky130_fd_sc_hd__clkinv_1 U16122 ( .A(j202_soc_core_j22_cpu_ml_macl[21]), 
        .Y(n22279) );
  sky130_fd_sc_hd__clkinv_1 U16123 ( .A(j202_soc_core_uart_TOP_rx_fifo_wp[1]), 
        .Y(n24002) );
  sky130_fd_sc_hd__clkinv_1 U16124 ( .A(j202_soc_core_j22_cpu_pc[27]), .Y(
        n22531) );
  sky130_fd_sc_hd__clkinv_1 U16125 ( .A(j202_soc_core_intc_core_00_rg_itgt[10]), .Y(n26732) );
  sky130_fd_sc_hd__clkinv_1 U16126 ( .A(j202_soc_core_j22_cpu_rf_gpr[14]), .Y(
        n14144) );
  sky130_fd_sc_hd__clkinv_1 U16127 ( .A(j202_soc_core_j22_cpu_rf_gpr[480]), 
        .Y(n21984) );
  sky130_fd_sc_hd__clkinv_1 U16128 ( .A(j202_soc_core_j22_cpu_ml_mach[31]), 
        .Y(n22474) );
  sky130_fd_sc_hd__clkinv_1 U16129 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[30]), .Y(n26789) );
  sky130_fd_sc_hd__clkinv_1 U16130 ( .A(j202_soc_core_qspi_wb_wdat[18]), .Y(
        n27128) );
  sky130_fd_sc_hd__clkinv_1 U16131 ( .A(j202_soc_core_intc_core_00_rg_itgt[64]), .Y(n28179) );
  sky130_fd_sc_hd__clkinv_1 U16132 ( .A(j202_soc_core_intc_core_00_rg_itgt[8]), 
        .Y(n26718) );
  sky130_fd_sc_hd__clkinv_1 U16133 ( .A(j202_soc_core_qspi_wb_wdat[20]), .Y(
        n27367) );
  sky130_fd_sc_hd__clkinv_1 U16134 ( .A(j202_soc_core_j22_cpu_rf_tmp[24]), .Y(
        n14777) );
  sky130_fd_sc_hd__clkinv_1 U16135 ( .A(j202_soc_core_intc_core_00_rg_itgt[13]), .Y(n26737) );
  sky130_fd_sc_hd__clkinv_1 U16136 ( .A(j202_soc_core_qspi_wb_wdat[10]), .Y(
        n28970) );
  sky130_fd_sc_hd__clkinv_1 U16137 ( .A(j202_soc_core_j22_cpu_pc[31]), .Y(
        n22463) );
  sky130_fd_sc_hd__clkinv_1 U16138 ( .A(j202_soc_core_intc_core_00_rg_itgt[9]), 
        .Y(n26712) );
  sky130_fd_sc_hd__clkinv_1 U16139 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]), .Y(n24525) );
  sky130_fd_sc_hd__clkinv_1 U16140 ( .A(j202_soc_core_qspi_wb_wdat[21]), .Y(
        n25572) );
  sky130_fd_sc_hd__clkinv_1 U16141 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[12]), .Y(n28987) );
  sky130_fd_sc_hd__clkinv_1 U16142 ( .A(j202_soc_core_cmt_core_00_reg_addr[5]), 
        .Y(n24019) );
  sky130_fd_sc_hd__clkinv_1 U16143 ( .A(j202_soc_core_uart_BRG_br_cnt[6]), .Y(
        n28630) );
  sky130_fd_sc_hd__clkinv_1 U16144 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[6]), .Y(n27465) );
  sky130_fd_sc_hd__clkinv_1 U16145 ( .A(j202_soc_core_cmt_core_00_cks0[0]), 
        .Y(n24009) );
  sky130_fd_sc_hd__clkinv_1 U16146 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[108]), .Y(n19921) );
  sky130_fd_sc_hd__clkinv_1 U16147 ( .A(j202_soc_core_intc_core_00_rg_itgt[5]), 
        .Y(n26679) );
  sky130_fd_sc_hd__clkinv_1 U16148 ( .A(j202_soc_core_j22_cpu_rf_gpr[26]), .Y(
        n15795) );
  sky130_fd_sc_hd__clkinv_1 U16149 ( .A(j202_soc_core_j22_cpu_rf_gpr[2]), .Y(
        n13914) );
  sky130_fd_sc_hd__clkinv_1 U16150 ( .A(j202_soc_core_intc_core_00_rg_itgt[76]), .Y(n27130) );
  sky130_fd_sc_hd__clkinv_1 U16151 ( .A(j202_soc_core_aquc_ADR__0_), .Y(n13268) );
  sky130_fd_sc_hd__clkinv_1 U16152 ( .A(j202_soc_core_j22_cpu_ml_mach[1]), .Y(
        n18360) );
  sky130_fd_sc_hd__clkinv_1 U16153 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[7]), .Y(n28561) );
  sky130_fd_sc_hd__clkinv_1 U16154 ( .A(j202_soc_core_intc_core_00_rg_itgt[1]), 
        .Y(n24825) );
  sky130_fd_sc_hd__clkinv_1 U16155 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[0]), .Y(n24005) );
  sky130_fd_sc_hd__clkinv_1 U16156 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[5]), .Y(n28558) );
  sky130_fd_sc_hd__clkinv_1 U16157 ( .A(j202_soc_core_j22_cpu_ml_mach[12]), 
        .Y(n21893) );
  sky130_fd_sc_hd__clkinv_1 U16158 ( .A(j202_soc_core_j22_cpu_pc_hold), .Y(
        n20427) );
  sky130_fd_sc_hd__clkinv_1 U16159 ( .A(j202_soc_core_cmt_core_00_reg_addr[4]), 
        .Y(n24018) );
  sky130_fd_sc_hd__clkinv_1 U16160 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[3]), .Y(n24266) );
  sky130_fd_sc_hd__clkinv_1 U16161 ( .A(j202_soc_core_j22_cpu_rf_gbr[26]), .Y(
        n22658) );
  sky130_fd_sc_hd__clkinv_1 U16162 ( .A(j202_soc_core_j22_cpu_ml_macl[17]), 
        .Y(n22844) );
  sky130_fd_sc_hd__clkinv_1 U16163 ( .A(j202_soc_core_intc_core_00_rg_itgt[45]), .Y(n25574) );
  sky130_fd_sc_hd__clkinv_1 U16164 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[9]), .Y(n23698) );
  sky130_fd_sc_hd__clkinv_1 U16165 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[1]), .Y(n24269) );
  sky130_fd_sc_hd__clkinv_1 U16166 ( .A(j202_soc_core_uart_BRG_br_cnt[4]), .Y(
        n28626) );
  sky130_fd_sc_hd__clkinv_1 U16167 ( .A(j202_soc_core_intc_core_00_rg_itgt[77]), .Y(n25607) );
  sky130_fd_sc_hd__clkinv_1 U16168 ( .A(j202_soc_core_j22_cpu_rf_tmp[2]), .Y(
        n19271) );
  sky130_fd_sc_hd__clkinv_1 U16169 ( .A(j202_soc_core_intc_core_00_rg_ipr[60]), 
        .Y(n26756) );
  sky130_fd_sc_hd__clkinv_1 U16170 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[10]), .Y(n23695) );
  sky130_fd_sc_hd__clkinv_1 U16171 ( .A(j202_soc_core_cmt_core_00_reg_addr[0]), 
        .Y(n23901) );
  sky130_fd_sc_hd__buf_4 U16172 ( .A(j202_soc_core_j22_cpu_ml_bufa[7]), .X(
        n27618) );
  sky130_fd_sc_hd__clkinv_1 U16173 ( .A(j202_soc_core_j22_cpu_rf_gpr[0]), .Y(
        n13794) );
  sky130_fd_sc_hd__clkinv_1 U16174 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[109]), .Y(n27627) );
  sky130_fd_sc_hd__clkinv_1 U16175 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[28]), .Y(n29256) );
  sky130_fd_sc_hd__clkinv_1 U16176 ( .A(j202_soc_core_cmt_core_00_reg_addr[6]), 
        .Y(n23900) );
  sky130_fd_sc_hd__clkinv_1 U16177 ( .A(j202_soc_core_j22_cpu_pc[26]), .Y(
        n22659) );
  sky130_fd_sc_hd__clkinv_1 U16178 ( .A(j202_soc_core_cmt_core_00_str0), .Y(
        n28213) );
  sky130_fd_sc_hd__clkinv_1 U16179 ( .A(j202_soc_core_j22_cpu_regop_imm__8_), 
        .Y(n14256) );
  sky130_fd_sc_hd__clkinv_1 U16180 ( .A(j202_soc_core_intc_core_00_rg_itgt[0]), 
        .Y(n24819) );
  sky130_fd_sc_hd__clkinv_1 U16181 ( .A(j202_soc_core_j22_cpu_memop_MEM__1_), 
        .Y(n24590) );
  sky130_fd_sc_hd__clkinv_1 U16182 ( .A(j202_soc_core_intr_vec__6_), .Y(n29066) );
  sky130_fd_sc_hd__clkinv_1 U16183 ( .A(j202_soc_core_uart_sio_ce_x4), .Y(
        n29095) );
  sky130_fd_sc_hd__clkinv_1 U16184 ( .A(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[0]), .Y(n23899) );
  sky130_fd_sc_hd__clkinv_1 U16185 ( .A(j202_soc_core_intc_core_00_rg_itgt[78]), .Y(n27869) );
  sky130_fd_sc_hd__clkinv_1 U16186 ( .A(j202_soc_core_j22_cpu_ml_mach[7]), .Y(
        n17488) );
  sky130_fd_sc_hd__clkinv_1 U16187 ( .A(j202_soc_core_j22_cpu_ml_mach[26]), 
        .Y(n22482) );
  sky130_fd_sc_hd__clkinv_1 U16188 ( .A(j202_soc_core_cmt_core_00_cnt1[0]), 
        .Y(n27516) );
  sky130_fd_sc_hd__and2_1 U16189 ( .A(n12032), .B(n12034), .X(n13447) );
  sky130_fd_sc_hd__clkinv_1 U16190 ( .A(j202_soc_core_j22_cpu_rf_pr[11]), .Y(
        n21293) );
  sky130_fd_sc_hd__clkinv_1 U16191 ( .A(j202_soc_core_intc_core_00_rg_itgt[3]), 
        .Y(n25188) );
  sky130_fd_sc_hd__clkinv_1 U16192 ( .A(j202_soc_core_intc_core_00_rg_itgt[79]), .Y(n27996) );
  sky130_fd_sc_hd__clkinv_1 U16193 ( .A(j202_soc_core_j22_cpu_ml_macl[20]), 
        .Y(n22318) );
  sky130_fd_sc_hd__inv_2 U16194 ( .A(j202_soc_core_bootrom_00_address_w[7]), 
        .Y(n18744) );
  sky130_fd_sc_hd__clkinv_1 U16195 ( .A(j202_soc_core_j22_cpu_rf_pr[0]), .Y(
        n21672) );
  sky130_fd_sc_hd__clkinv_1 U16196 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[105]), .Y(n27560) );
  sky130_fd_sc_hd__clkinv_1 U16197 ( .A(j202_soc_core_intc_core_00_rg_itgt[2]), 
        .Y(n25161) );
  sky130_fd_sc_hd__clkinv_1 U16198 ( .A(j202_soc_core_j22_cpu_ml_macl[8]), .Y(
        n21733) );
  sky130_fd_sc_hd__clkinv_1 U16199 ( .A(j202_soc_core_j22_cpu_opst[2]), .Y(
        n23420) );
  sky130_fd_sc_hd__clkinv_1 U16200 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[29]), .Y(n26799) );
  sky130_fd_sc_hd__clkinv_1 U16201 ( .A(j202_soc_core_uart_BRG_br_cnt[2]), .Y(
        n28632) );
  sky130_fd_sc_hd__clkinv_1 U16202 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[3]), .Y(n29072) );
  sky130_fd_sc_hd__clkinv_1 U16203 ( .A(j202_soc_core_intc_core_00_rg_itgt[11]), .Y(n25189) );
  sky130_fd_sc_hd__clkinv_1 U16204 ( .A(j202_soc_core_j22_cpu_rf_gpr[15]), .Y(
        n14564) );
  sky130_fd_sc_hd__clkinv_1 U16205 ( .A(j202_soc_core_j22_cpu_rf_gbr[11]), .Y(
        n14011) );
  sky130_fd_sc_hd__clkinv_1 U16206 ( .A(j202_soc_core_j22_cpu_ml_mach[16]), 
        .Y(n22027) );
  sky130_fd_sc_hd__clkinv_1 U16207 ( .A(j202_soc_core_j22_cpu_opst[1]), .Y(
        n28373) );
  sky130_fd_sc_hd__clkinv_1 U16208 ( .A(j202_soc_core_intc_core_00_rg_itgt[17]), .Y(n26762) );
  sky130_fd_sc_hd__clkinv_1 U16209 ( .A(j202_soc_core_qspi_wb_wdat[2]), .Y(
        n28915) );
  sky130_fd_sc_hd__clkinv_1 U16210 ( .A(j202_soc_core_intc_core_00_rg_itgt[86]), .Y(n27873) );
  sky130_fd_sc_hd__clkinv_1 U16211 ( .A(j202_soc_core_j22_cpu_rf_vbr[23]), .Y(
        n14862) );
  sky130_fd_sc_hd__clkinv_1 U16212 ( .A(j202_soc_core_qspi_wb_wdat[1]), .Y(
        n28902) );
  sky130_fd_sc_hd__clkinv_1 U16213 ( .A(j202_soc_core_j22_cpu_ml_mach[27]), 
        .Y(n22485) );
  sky130_fd_sc_hd__clkinv_1 U16214 ( .A(j202_soc_core_intc_core_00_rg_ipr[44]), 
        .Y(n25191) );
  sky130_fd_sc_hd__clkinv_1 U16215 ( .A(j202_soc_core_intc_core_00_rg_itgt[92]), .Y(n27133) );
  sky130_fd_sc_hd__clkinv_1 U16216 ( .A(j202_soc_core_j22_cpu_ml_macl[2]), .Y(
        n19244) );
  sky130_fd_sc_hd__clkinv_1 U16217 ( .A(j202_soc_core_j22_cpu_rf_tmp[23]), .Y(
        n14864) );
  sky130_fd_sc_hd__clkinv_1 U16218 ( .A(j202_soc_core_j22_cpu_rf_gbr[10]), .Y(
        n14347) );
  sky130_fd_sc_hd__clkinv_1 U16219 ( .A(j202_soc_core_intc_core_00_rg_ipr[118]), .Y(n25608) );
  sky130_fd_sc_hd__clkinv_1 U16220 ( .A(j202_soc_core_uart_BRG_br_clr), .Y(
        n28624) );
  sky130_fd_sc_hd__clkinv_1 U16221 ( .A(j202_soc_core_j22_cpu_ml_mach[9]), .Y(
        n18982) );
  sky130_fd_sc_hd__clkinv_1 U16222 ( .A(j202_soc_core_j22_cpu_rf_gpr[502]), 
        .Y(n14861) );
  sky130_fd_sc_hd__clkinv_1 U16223 ( .A(j202_soc_core_j22_cpu_rf_gpr[24]), .Y(
        n14742) );
  sky130_fd_sc_hd__clkinv_1 U16224 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .Y(n23738) );
  sky130_fd_sc_hd__clkinv_1 U16225 ( .A(j202_soc_core_intc_core_00_rg_itgt[87]), .Y(n28000) );
  sky130_fd_sc_hd__clkinv_1 U16226 ( .A(j202_soc_core_j22_cpu_ml_mach[24]), 
        .Y(n22480) );
  sky130_fd_sc_hd__clkinv_1 U16227 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[5]), .Y(n23676) );
  sky130_fd_sc_hd__clkinv_1 U16228 ( .A(j202_soc_core_wbqspiflash_00_state[1]), 
        .Y(n23640) );
  sky130_fd_sc_hd__clkinv_1 U16229 ( .A(j202_soc_core_j22_cpu_rf_gpr[493]), 
        .Y(n22572) );
  sky130_fd_sc_hd__inv_2 U16230 ( .A(j202_soc_core_j22_cpu_regop_other__0_), 
        .Y(n18869) );
  sky130_fd_sc_hd__clkinv_1 U16231 ( .A(j202_soc_core_aquc_SEL__0_), .Y(n22414) );
  sky130_fd_sc_hd__clkinv_1 U16232 ( .A(j202_soc_core_intc_core_00_rg_ipr[117]), .Y(n25575) );
  sky130_fd_sc_hd__clkinv_1 U16233 ( .A(j202_soc_core_intc_core_00_rg_ipr[12]), 
        .Y(n26671) );
  sky130_fd_sc_hd__clkinv_1 U16234 ( .A(j202_soc_core_j22_cpu_rf_gpr[489]), 
        .Y(n19282) );
  sky130_fd_sc_hd__clkinv_1 U16235 ( .A(j202_soc_core_wbqspiflash_00_state[4]), 
        .Y(n26580) );
  sky130_fd_sc_hd__clkinv_1 U16236 ( .A(j202_soc_core_j22_cpu_ml_macl[18]), 
        .Y(n22366) );
  sky130_fd_sc_hd__clkinv_1 U16237 ( .A(j202_soc_core_cmt_core_00_cnt1[13]), 
        .Y(n26080) );
  sky130_fd_sc_hd__clkinv_1 U16238 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[5]), .Y(n24749) );
  sky130_fd_sc_hd__clkinv_1 U16239 ( .A(j202_soc_core_intc_core_00_rg_ie[13]), 
        .Y(n25784) );
  sky130_fd_sc_hd__clkinv_1 U16240 ( .A(j202_soc_core_qspi_wb_wdat[4]), .Y(
        n28906) );
  sky130_fd_sc_hd__clkinv_1 U16241 ( .A(j202_soc_core_wbqspiflash_00_state[2]), 
        .Y(n26588) );
  sky130_fd_sc_hd__clkinv_1 U16242 ( .A(j202_soc_core_j22_cpu_rf_gpr[506]), 
        .Y(n16000) );
  sky130_fd_sc_hd__clkinv_1 U16243 ( .A(j202_soc_core_j22_cpu_rf_gbr[30]), .Y(
        n22581) );
  sky130_fd_sc_hd__clkinv_1 U16244 ( .A(j202_soc_core_j22_cpu_rf_tmp[27]), .Y(
        n16002) );
  sky130_fd_sc_hd__clkinv_1 U16245 ( .A(j202_soc_core_j22_cpu_rf_gpr[1]), .Y(
        n13882) );
  sky130_fd_sc_hd__clkinv_1 U16246 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[31]), .Y(n26780) );
  sky130_fd_sc_hd__clkinv_1 U16248 ( .A(j202_soc_core_j22_cpu_rf_gbr[16]), .Y(
        n22771) );
  sky130_fd_sc_hd__clkinv_1 U16249 ( .A(j202_soc_core_j22_cpu_rf_gpr[481]), 
        .Y(n19265) );
  sky130_fd_sc_hd__clkinv_1 U16251 ( .A(j202_soc_core_j22_cpu_rf_vbr[1]), .Y(
        n13777) );
  sky130_fd_sc_hd__clkinv_1 U16252 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[20]), .Y(n29043) );
  sky130_fd_sc_hd__clkinv_1 U16253 ( .A(j202_soc_core_uart_BRG_ps[6]), .Y(
        n28618) );
  sky130_fd_sc_hd__clkinv_1 U16254 ( .A(j202_soc_core_intc_core_00_rg_ie[12]), 
        .Y(n25187) );
  sky130_fd_sc_hd__clkinv_1 U16255 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[31]), .Y(n29133) );
  sky130_fd_sc_hd__clkinv_1 U16256 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[11]), .Y(n28913) );
  sky130_fd_sc_hd__clkinv_1 U16257 ( .A(j202_soc_core_cmt_core_00_cmf1), .Y(
        n24730) );
  sky130_fd_sc_hd__clkinv_1 U16258 ( .A(j202_soc_core_j22_cpu_ml_mach[2]), .Y(
        n18406) );
  sky130_fd_sc_hd__clkinv_1 U16259 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[11]), .Y(n23705) );
  sky130_fd_sc_hd__clkinv_1 U16260 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[7]), .Y(n27550) );
  sky130_fd_sc_hd__clkinv_1 U16261 ( .A(j202_soc_core_memory0_ram_dout0[498]), 
        .Y(n13178) );
  sky130_fd_sc_hd__clkinv_1 U16262 ( .A(j202_soc_core_j22_cpu_pc[12]), .Y(
        n20933) );
  sky130_fd_sc_hd__clkinv_1 U16263 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .Y(n23862) );
  sky130_fd_sc_hd__or2_0 U16264 ( .A(start_n_reg[0]), .B(wb_rst_i), .X(n4) );
  sky130_fd_sc_hd__clkinv_1 U16265 ( .A(j202_soc_core_j22_cpu_rf_pr[16]), .Y(
        n14535) );
  sky130_fd_sc_hd__clkinv_1 U16266 ( .A(j202_soc_core_intr_vec__0_), .Y(n27348) );
  sky130_fd_sc_hd__clkinv_1 U16267 ( .A(j202_soc_core_pwrite[0]), .Y(n24729)
         );
  sky130_fd_sc_hd__clkinv_1 U16268 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[4]), .Y(n24741) );
  sky130_fd_sc_hd__clkinv_1 U16269 ( .A(j202_soc_core_j22_cpu_rf_gpr[10]), .Y(
        n14346) );
  sky130_fd_sc_hd__clkinv_1 U16270 ( .A(j202_soc_core_j22_cpu_ml_macl[1]), .Y(
        n21942) );
  sky130_fd_sc_hd__clkinv_1 U16271 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[2]), .Y(n24200) );
  sky130_fd_sc_hd__clkinv_1 U16272 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[46]), .Y(n20098) );
  sky130_fd_sc_hd__clkinv_1 U16273 ( .A(j202_soc_core_j22_cpu_ml_macl[5]), .Y(
        n22245) );
  sky130_fd_sc_hd__clkinv_1 U16274 ( .A(j202_soc_core_qspi_wb_wdat[22]), .Y(
        n26834) );
  sky130_fd_sc_hd__clkinv_1 U16275 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[107]), .Y(n20760) );
  sky130_fd_sc_hd__clkinv_1 U16276 ( .A(j202_soc_core_j22_cpu_rf_vbr[9]), .Y(
        n14374) );
  sky130_fd_sc_hd__clkinv_1 U16277 ( .A(j202_soc_core_qspi_wb_wdat[3]), .Y(
        n28922) );
  sky130_fd_sc_hd__clkinv_1 U16278 ( .A(j202_soc_core_j22_cpu_rf_vbr[24]), .Y(
        n14776) );
  sky130_fd_sc_hd__clkinv_1 U16279 ( .A(j202_soc_core_wbqspiflash_00_spi_wr), 
        .Y(n26558) );
  sky130_fd_sc_hd__clkinv_1 U16280 ( .A(j202_soc_core_intr_level__3_), .Y(
        n16909) );
  sky130_fd_sc_hd__clkinv_1 U16281 ( .A(j202_soc_core_qspi_wb_wdat[23]), .Y(
        n27625) );
  sky130_fd_sc_hd__clkinv_1 U16282 ( .A(j202_soc_core_intr_level__2_), .Y(
        n16908) );
  sky130_fd_sc_hd__clkinv_1 U16283 ( .A(j202_soc_core_j22_cpu_ml_macl[31]), 
        .Y(n18475) );
  sky130_fd_sc_hd__clkinv_1 U16284 ( .A(j202_soc_core_wbqspiflash_00_spi_busy), 
        .Y(n26623) );
  sky130_fd_sc_hd__clkinv_1 U16285 ( .A(j202_soc_core_j22_cpu_rf_vbr[11]), .Y(
        n21297) );
  sky130_fd_sc_hd__clkinv_1 U16286 ( .A(j202_soc_core_j22_cpu_rf_gpr[492]), 
        .Y(n22981) );
  sky130_fd_sc_hd__clkinv_1 U16287 ( .A(j202_soc_core_intr_level__1_), .Y(
        n16910) );
  sky130_fd_sc_hd__clkinv_1 U16288 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[10]), .Y(n28976) );
  sky130_fd_sc_hd__clkinv_1 U16289 ( .A(j202_soc_core_j22_cpu_rf_tmp[17]), .Y(
        n14479) );
  sky130_fd_sc_hd__clkinv_1 U16290 ( .A(j202_soc_core_j22_cpu_rf_gbr[1]), .Y(
        n13781) );
  sky130_fd_sc_hd__clkinv_1 U16291 ( .A(j202_soc_core_j22_cpu_rf_vbr[17]), .Y(
        n14478) );
  sky130_fd_sc_hd__clkinv_1 U16292 ( .A(j202_soc_core_j22_cpu_rfuo_sr__m_), 
        .Y(n22895) );
  sky130_fd_sc_hd__clkinv_1 U16293 ( .A(j202_soc_core_j22_cpu_regop_imm__0_), 
        .Y(n13795) );
  sky130_fd_sc_hd__clkinv_1 U16294 ( .A(j202_soc_core_j22_cpu_rf_tmp[9]), .Y(
        n22896) );
  sky130_fd_sc_hd__clkinv_1 U16295 ( .A(j202_soc_core_intc_core_00_rg_itgt[95]), .Y(n28001) );
  sky130_fd_sc_hd__clkinv_1 U16296 ( .A(j202_soc_core_intc_core_00_rg_ipr[124]), .Y(n27392) );
  sky130_fd_sc_hd__clkinv_1 U16297 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[12]), .Y(n23702) );
  sky130_fd_sc_hd__clkinv_1 U16298 ( .A(j202_soc_core_intc_core_00_rg_itgt[84]), .Y(n27132) );
  sky130_fd_sc_hd__clkinv_1 U16299 ( .A(j202_soc_core_j22_cpu_rf_pr[17]), .Y(
        n14481) );
  sky130_fd_sc_hd__clkinv_1 U16300 ( .A(j202_soc_core_j22_cpu_id_opn_v_), .Y(
        n19429) );
  sky130_fd_sc_hd__clkinv_1 U16301 ( .A(j202_soc_core_j22_cpu_rf_gbr[17]), .Y(
        n22856) );
  sky130_fd_sc_hd__clkinv_1 U16302 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[9]), .Y(n24008) );
  sky130_fd_sc_hd__clkinv_1 U16303 ( .A(j202_soc_core_j22_cpu_rf_pr[31]), .Y(
        n16492) );
  sky130_fd_sc_hd__clkinv_1 U16304 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[30]), .Y(n26791) );
  sky130_fd_sc_hd__clkinv_1 U16305 ( .A(j202_soc_core_j22_cpu_rf_tmp[10]), .Y(
        n14344) );
  sky130_fd_sc_hd__clkinv_1 U16306 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[3]), .Y(n27674) );
  sky130_fd_sc_hd__clkinv_1 U16307 ( .A(j202_soc_core_j22_cpu_rf_tmp[11]), .Y(
        n21298) );
  sky130_fd_sc_hd__clkinv_1 U16308 ( .A(j202_soc_core_aquc_ADR__5_), .Y(n13264) );
  sky130_fd_sc_hd__clkinv_1 U16309 ( .A(j202_soc_core_intc_core_00_rg_itgt[94]), .Y(n27874) );
  sky130_fd_sc_hd__clkinv_1 U16310 ( .A(j202_soc_core_intc_core_00_rg_itgt[53]), .Y(n25580) );
  sky130_fd_sc_hd__clkinv_1 U16311 ( .A(j202_soc_core_intc_core_00_rg_ipr[122]), .Y(n27870) );
  sky130_fd_sc_hd__clkinv_1 U16312 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[1]), 
        .Y(n18689) );
  sky130_fd_sc_hd__clkinv_1 U16313 ( .A(j202_soc_core_cmt_core_00_cnt1[14]), 
        .Y(n26086) );
  sky130_fd_sc_hd__clkinv_1 U16314 ( .A(j202_soc_core_j22_cpu_rf_vbr[10]), .Y(
        n14343) );
  sky130_fd_sc_hd__clkinv_1 U16315 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[1]), 
        .Y(n24004) );
  sky130_fd_sc_hd__clkinv_1 U16316 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[125]), .Y(n27632) );
  sky130_fd_sc_hd__clkinv_1 U16317 ( .A(j202_soc_core_intc_core_00_rg_ipr[108]), .Y(n25190) );
  sky130_fd_sc_hd__clkinv_1 U16318 ( .A(j202_soc_core_j22_cpu_ml_mach[11]), 
        .Y(n18937) );
  sky130_fd_sc_hd__clkinv_1 U16319 ( .A(j202_soc_core_j22_cpu_ml_macl[25]), 
        .Y(n22889) );
  sky130_fd_sc_hd__clkinv_1 U16320 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__2_), 
        .Y(n24718) );
  sky130_fd_sc_hd__clkinv_1 U16321 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[0]), 
        .Y(n27921) );
  sky130_fd_sc_hd__clkinv_1 U16322 ( .A(j202_soc_core_intc_core_00_rg_itgt[85]), .Y(n25612) );
  sky130_fd_sc_hd__clkinv_1 U16323 ( .A(j202_soc_core_intc_core_00_rg_itgt[93]), .Y(n25613) );
  sky130_fd_sc_hd__clkinv_1 U16324 ( .A(j202_soc_core_j22_cpu_ml_mach[5]), .Y(
        n17762) );
  sky130_fd_sc_hd__clkinv_1 U16325 ( .A(j202_soc_core_j22_cpu_ml_mach[15]), 
        .Y(n19092) );
  sky130_fd_sc_hd__clkinv_1 U16326 ( .A(j202_soc_core_j22_cpu_ml_macl[9]), .Y(
        n18195) );
  sky130_fd_sc_hd__clkinv_1 U16327 ( .A(j202_soc_core_qspi_wb_wdat[7]), .Y(
        n28949) );
  sky130_fd_sc_hd__clkinv_1 U16328 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[4]), .Y(n23679) );
  sky130_fd_sc_hd__clkinv_1 U16329 ( .A(j202_soc_core_j22_cpu_pc[30]), .Y(
        n22582) );
  sky130_fd_sc_hd__clkinv_1 U16330 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[28]), .Y(n29058) );
  sky130_fd_sc_hd__clkinv_1 U16331 ( .A(j202_soc_core_qspi_wb_wdat[6]), .Y(
        n28942) );
  sky130_fd_sc_hd__clkinv_1 U16332 ( .A(j202_soc_core_j22_cpu_ml_mach[25]), 
        .Y(n22481) );
  sky130_fd_sc_hd__clkinv_1 U16333 ( .A(j202_soc_core_j22_cpu_rf_gbr[31]), .Y(
        n22462) );
  sky130_fd_sc_hd__clkinv_1 U16334 ( .A(wbs_dat_o[0]), .Y(n10525) );
  sky130_fd_sc_hd__clkinv_1 U16335 ( .A(j202_soc_core_intc_core_00_rg_itgt[61]), .Y(n25581) );
  sky130_fd_sc_hd__clkinv_1 U16336 ( .A(j202_soc_core_qspi_wb_wdat[5]), .Y(
        n28935) );
  sky130_fd_sc_hd__clkinv_1 U16337 ( .A(j202_soc_core_j22_cpu_rf_pr[10]), .Y(
        n19283) );
  sky130_fd_sc_hd__clkinv_1 U16338 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[117]), .Y(n27631) );
  sky130_fd_sc_hd__clkinv_1 U16339 ( .A(j202_soc_core_intc_core_00_rg_ipr[39]), 
        .Y(n26730) );
  sky130_fd_sc_hd__clkinv_1 U16340 ( .A(j202_soc_core_wbqspiflash_00_spi_in[4]), .Y(n29195) );
  sky130_fd_sc_hd__clkinv_1 U16341 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[0]), .Y(n28723) );
  sky130_fd_sc_hd__clkinv_1 U16342 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[10]), .Y(n24976) );
  sky130_fd_sc_hd__clkinv_1 U16343 ( .A(j202_soc_core_intc_core_00_rg_itgt[36]), .Y(n25742) );
  sky130_fd_sc_hd__clkinv_1 U16344 ( .A(j202_soc_core_intc_core_00_rg_ie[20]), 
        .Y(n27312) );
  sky130_fd_sc_hd__clkinv_1 U16345 ( .A(j202_soc_core_j22_cpu_rf_gpr[12]), .Y(
        n14032) );
  sky130_fd_sc_hd__clkinv_1 U16346 ( .A(j202_soc_core_intc_core_00_rg_ipr[51]), 
        .Y(n25323) );
  sky130_fd_sc_hd__clkinv_1 U16347 ( .A(j202_soc_core_intc_core_00_rg_ie[2]), 
        .Y(n25160) );
  sky130_fd_sc_hd__clkinv_1 U16348 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[11]), .Y(n26996) );
  sky130_fd_sc_hd__clkinv_1 U16349 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[5]), .Y(n27432) );
  sky130_fd_sc_hd__clkinv_1 U16351 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[13]), .Y(n27723) );
  sky130_fd_sc_hd__clkinv_1 U16352 ( .A(j202_soc_core_wbqspiflash_00_spi_spd), 
        .Y(n28727) );
  sky130_fd_sc_hd__inv_1 U16353 ( .A(j202_soc_core_intc_core_00_rg_ipr[49]), 
        .Y(n25745) );
  sky130_fd_sc_hd__clkinv_1 U16354 ( .A(j202_soc_core_qspi_wb_addr[11]), .Y(
        n28800) );
  sky130_fd_sc_hd__clkinv_1 U16355 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[14]), .Y(n26875) );
  sky130_fd_sc_hd__clkinv_1 U16356 ( .A(j202_soc_core_memory0_ram_dout0_sel[1]), .Y(n13165) );
  sky130_fd_sc_hd__clkinv_1 U16357 ( .A(
        j202_soc_core_bldc_core_00_hall_value[2]), .Y(n28159) );
  sky130_fd_sc_hd__clkinv_1 U16358 ( .A(j202_soc_core_memory0_ram_dout0_sel[3]), .Y(n13173) );
  sky130_fd_sc_hd__nand2_1 U16359 ( .A(j202_soc_core_memory0_ram_dout0[479]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12581) );
  sky130_fd_sc_hd__clkinv_1 U16360 ( .A(j202_soc_core_intc_core_00_rg_ie[17]), 
        .Y(n25741) );
  sky130_fd_sc_hd__clkinv_1 U16361 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[6]), .Y(n27459) );
  sky130_fd_sc_hd__clkinv_1 U16362 ( .A(j202_soc_core_memory0_ram_dout0_sel[2]), .Y(n13166) );
  sky130_fd_sc_hd__clkinv_1 U16363 ( .A(
        j202_soc_core_intc_core_00_in_intreq[17]), .Y(n25733) );
  sky130_fd_sc_hd__clkinv_1 U16364 ( .A(j202_soc_core_ahb2apb_02_state[0]), 
        .Y(n24260) );
  sky130_fd_sc_hd__clkinv_1 U16365 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[9]), .Y(n28964) );
  sky130_fd_sc_hd__clkinv_1 U16366 ( .A(j202_soc_core_intc_core_00_rg_itgt[39]), .Y(n25485) );
  sky130_fd_sc_hd__clkinv_1 U16367 ( .A(j202_soc_core_qspi_wb_addr[2]), .Y(
        n28739) );
  sky130_fd_sc_hd__clkinv_1 U16368 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[1]), .Y(n29084) );
  sky130_fd_sc_hd__clkinv_1 U16369 ( .A(j202_soc_core_wbqspiflash_00_spif_cmd), 
        .Y(n26534) );
  sky130_fd_sc_hd__clkinv_1 U16370 ( .A(j202_soc_core_intc_core_00_rg_ie[15]), 
        .Y(n26116) );
  sky130_fd_sc_hd__clkinv_1 U16371 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[2]), .Y(n29086) );
  sky130_fd_sc_hd__clkinv_1 U16372 ( .A(j202_soc_core_intc_core_00_rg_itgt[47]), .Y(n25486) );
  sky130_fd_sc_hd__clkinv_1 U16373 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[8]), .Y(n27964) );
  sky130_fd_sc_hd__clkinv_1 U16374 ( .A(j202_soc_core_j22_cpu_ml_macl[13]), 
        .Y(n24445) );
  sky130_fd_sc_hd__clkinv_1 U16375 ( .A(j202_soc_core_memory0_ram_dout0_sel[6]), .Y(n13164) );
  sky130_fd_sc_hd__clkinv_1 U16376 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[3]), .Y(n28798) );
  sky130_fd_sc_hd__clkinv_1 U16377 ( .A(j202_soc_core_qspi_wb_addr[3]), .Y(
        n26530) );
  sky130_fd_sc_hd__clkinv_1 U16378 ( .A(j202_soc_core_j22_cpu_ml_mach[10]), 
        .Y(n19307) );
  sky130_fd_sc_hd__clkinv_1 U16379 ( .A(j202_soc_core_intc_core_00_rg_itgt[62]), .Y(n27171) );
  sky130_fd_sc_hd__clkinv_1 U16380 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[7]), .Y(n28829) );
  sky130_fd_sc_hd__clkinv_1 U16381 ( .A(j202_soc_core_j22_cpu_rf_tmp[0]), .Y(
        n21674) );
  sky130_fd_sc_hd__clkinv_1 U16382 ( .A(j202_soc_core_intc_core_00_rg_itgt[55]), .Y(n25492) );
  sky130_fd_sc_hd__clkinv_1 U16383 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[93]), .Y(n15664) );
  sky130_fd_sc_hd__clkinv_1 U16384 ( .A(j202_soc_core_intc_core_00_rg_itgt[54]), .Y(n27170) );
  sky130_fd_sc_hd__clkinv_1 U16385 ( .A(j202_soc_core_memory0_ram_dout0_sel[4]), .Y(n13170) );
  sky130_fd_sc_hd__clkinv_1 U16386 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[32]), .Y(n19638) );
  sky130_fd_sc_hd__clkinv_1 U16387 ( .A(j202_soc_core_intc_core_00_rg_itgt[46]), .Y(n27166) );
  sky130_fd_sc_hd__clkinv_1 U16388 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[8]), .Y(n27968) );
  sky130_fd_sc_hd__clkinv_1 U16389 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[68]), .Y(n21447) );
  sky130_fd_sc_hd__clkinv_1 U16390 ( .A(j202_soc_core_j22_cpu_rf_gpr[19]), .Y(
        n14889) );
  sky130_fd_sc_hd__clkinv_1 U16391 ( .A(j202_soc_core_intc_core_00_rg_itgt[58]), .Y(n27938) );
  sky130_fd_sc_hd__clkinv_1 U16392 ( .A(j202_soc_core_j22_cpu_ml_macl[28]), 
        .Y(n22630) );
  sky130_fd_sc_hd__clkinv_1 U16393 ( .A(j202_soc_core_j22_cpu_rf_gpr[483]), 
        .Y(n21798) );
  sky130_fd_sc_hd__clkinv_1 U16394 ( .A(
        j202_soc_core_wbqspiflash_00_write_in_progress), .Y(n27614) );
  sky130_fd_sc_hd__clkinv_1 U16395 ( .A(j202_soc_core_intc_core_00_rg_ipr[27]), 
        .Y(n26708) );
  sky130_fd_sc_hd__clkinv_1 U16396 ( .A(j202_soc_core_j22_cpu_rf_vbr[4]), .Y(
        n21800) );
  sky130_fd_sc_hd__clkinv_1 U16397 ( .A(j202_soc_core_intc_core_00_rg_ie[11]), 
        .Y(n28068) );
  sky130_fd_sc_hd__clkinv_1 U16398 ( .A(j202_soc_core_intc_core_00_bs_addr[6]), 
        .Y(n29408) );
  sky130_fd_sc_hd__clkinv_1 U16399 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[7]), .Y(n28955) );
  sky130_fd_sc_hd__clkinv_1 U16400 ( .A(j202_soc_core_j22_cpu_rf_pr[8]), .Y(
        n21735) );
  sky130_fd_sc_hd__clkinv_1 U16401 ( .A(j202_soc_core_qspi_wb_wdat[9]), .Y(
        n28963) );
  sky130_fd_sc_hd__clkinv_1 U16402 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[3]), 
        .Y(n13287) );
  sky130_fd_sc_hd__clkinv_1 U16403 ( .A(j202_soc_core_intc_core_00_rg_itgt[38]), .Y(n27165) );
  sky130_fd_sc_hd__clkinv_1 U16404 ( .A(j202_soc_core_j22_cpu_id_opn_inst__12_), .Y(n19856) );
  sky130_fd_sc_hd__clkinv_1 U16405 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__0_), 
        .Y(n21801) );
  sky130_fd_sc_hd__clkinv_1 U16406 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[97]), .Y(n19360) );
  sky130_fd_sc_hd__clkinv_1 U16407 ( .A(j202_soc_core_intc_core_00_rg_ie[3]), 
        .Y(n27352) );
  sky130_fd_sc_hd__clkinv_1 U16408 ( .A(j202_soc_core_j22_cpu_rf_tmp[4]), .Y(
        n21802) );
  sky130_fd_sc_hd__clkinv_1 U16409 ( .A(j202_soc_core_j22_cpu_ml_macl[12]), 
        .Y(n21883) );
  sky130_fd_sc_hd__clkinv_1 U16410 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[9]), .Y(n28969) );
  sky130_fd_sc_hd__clkinv_1 U16411 ( .A(j202_soc_core_intc_core_00_rg_itgt[44]), .Y(n25743) );
  sky130_fd_sc_hd__clkinv_1 U16412 ( .A(j202_soc_core_pwrite[2]), .Y(n26898)
         );
  sky130_fd_sc_hd__clkinv_1 U16413 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[11]), .Y(n28978) );
  sky130_fd_sc_hd__clkinv_1 U16414 ( .A(j202_soc_core_uart_BRG_ps_clr), .Y(
        n28601) );
  sky130_fd_sc_hd__clkinv_1 U16415 ( .A(j202_soc_core_j22_cpu_rf_tmp[21]), .Y(
        n15058) );
  sky130_fd_sc_hd__clkinv_1 U16416 ( .A(j202_soc_core_j22_cpu_rf_vbr[6]), .Y(
        n13575) );
  sky130_fd_sc_hd__clkinv_1 U16417 ( .A(j202_soc_core_intc_core_00_rg_ie[19]), 
        .Y(n27710) );
  sky130_fd_sc_hd__clkinv_1 U16418 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[15]), .Y(n26134) );
  sky130_fd_sc_hd__clkinv_1 U16419 ( .A(j202_soc_core_cmt_core_00_cks1[1]), 
        .Y(n23906) );
  sky130_fd_sc_hd__clkinv_1 U16420 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[5]), .Y(n28575) );
  sky130_fd_sc_hd__clkinv_1 U16421 ( .A(j202_soc_core_intc_core_00_rg_ipr[77]), 
        .Y(n25791) );
  sky130_fd_sc_hd__clkinv_1 U16422 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[3]), .Y(n28571) );
  sky130_fd_sc_hd__clkinv_1 U16423 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[9]), .Y(n23907) );
  sky130_fd_sc_hd__clkinv_1 U16424 ( .A(j202_soc_core_cmt_core_00_cmf0), .Y(
        n27551) );
  sky130_fd_sc_hd__clkinv_1 U16425 ( .A(j202_soc_core_j22_cpu_rf_gpr[500]), 
        .Y(n15056) );
  sky130_fd_sc_hd__clkinv_1 U16426 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[7]), .Y(n28580) );
  sky130_fd_sc_hd__clkinv_1 U16427 ( .A(j202_soc_core_intc_core_00_rg_ipr[64]), 
        .Y(n28230) );
  sky130_fd_sc_hd__clkinv_1 U16428 ( .A(j202_soc_core_intc_core_00_rg_ie[1]), 
        .Y(n24822) );
  sky130_fd_sc_hd__clkinv_1 U16429 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[14]), .Y(n26893) );
  sky130_fd_sc_hd__clkinv_1 U16430 ( .A(j202_soc_core_j22_cpu_rf_pr[7]), .Y(
        n14290) );
  sky130_fd_sc_hd__clkinv_1 U16431 ( .A(j202_soc_core_j22_cpu_ml_macl[29]), 
        .Y(n18026) );
  sky130_fd_sc_hd__clkinv_1 U16432 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__2_), 
        .Y(n22154) );
  sky130_fd_sc_hd__clkinv_1 U16433 ( .A(j202_soc_core_cmt_core_00_cks1[0]), 
        .Y(n23908) );
  sky130_fd_sc_hd__clkinv_1 U16434 ( .A(j202_soc_core_j22_cpu_rf_tmp[6]), .Y(
        n22155) );
  sky130_fd_sc_hd__clkinv_1 U16435 ( .A(j202_soc_core_qspi_wb_wdat[11]), .Y(
        n28977) );
  sky130_fd_sc_hd__clkinv_1 U16436 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[10]), .Y(n28546) );
  sky130_fd_sc_hd__clkinv_1 U16437 ( .A(j202_soc_core_j22_cpu_rf_gbr[14]), .Y(
        n14145) );
  sky130_fd_sc_hd__clkinv_1 U16438 ( .A(j202_soc_core_bootrom_00_sel_w), .Y(
        n13147) );
  sky130_fd_sc_hd__clkinv_1 U16439 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[11]), .Y(n28983) );
  sky130_fd_sc_hd__clkinv_1 U16440 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[0]), .Y(n28228) );
  sky130_fd_sc_hd__clkinv_1 U16442 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[91]), .Y(n16111) );
  sky130_fd_sc_hd__clkinv_1 U16443 ( .A(j202_soc_core_memory0_ram_dout0_sel[8]), .Y(n13159) );
  sky130_fd_sc_hd__clkinv_1 U16444 ( .A(j202_soc_core_qspi_wb_addr[12]), .Y(
        n28808) );
  sky130_fd_sc_hd__clkinv_1 U16445 ( .A(j202_soc_core_j22_cpu_rf_pr[14]), .Y(
        n22573) );
  sky130_fd_sc_hd__clkinv_1 U16446 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[12]), .Y(n25170) );
  sky130_fd_sc_hd__clkinv_1 U16447 ( .A(j202_soc_core_bldc_core_00_comm[2]), 
        .Y(n29119) );
  sky130_fd_sc_hd__clkinv_1 U16448 ( .A(j202_soc_core_wbqspiflash_00_spif_ctrl), .Y(n26481) );
  sky130_fd_sc_hd__clkinv_1 U16449 ( .A(j202_soc_core_j22_cpu_rf_gpr[17]), .Y(
        n14480) );
  sky130_fd_sc_hd__clkinv_1 U16450 ( .A(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[1]), .Y(n19337) );
  sky130_fd_sc_hd__clkinv_1 U16451 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[4]), .Y(n28806) );
  sky130_fd_sc_hd__clkinv_1 U16452 ( .A(j202_soc_core_j22_cpu_rf_gpr[498]), 
        .Y(n14917) );
  sky130_fd_sc_hd__clkinv_1 U16453 ( .A(j202_soc_core_qspi_wb_wdat[17]), .Y(
        n25732) );
  sky130_fd_sc_hd__clkinv_1 U16454 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[26]), .Y(n26813) );
  sky130_fd_sc_hd__clkinv_1 U16455 ( .A(j202_soc_core_j22_cpu_rf_vbr[14]), .Y(
        n14141) );
  sky130_fd_sc_hd__clkinv_1 U16456 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[27]), .Y(n21309) );
  sky130_fd_sc_hd__clkinv_1 U16457 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[17]), .Y(n25757) );
  sky130_fd_sc_hd__clkinv_1 U16458 ( .A(j202_soc_core_j22_cpu_rf_tmp[19]), .Y(
        n14919) );
  sky130_fd_sc_hd__clkinv_1 U16459 ( .A(n30145), .Y(n19308) );
  sky130_fd_sc_hd__clkinv_1 U16460 ( .A(gpio_en_o[12]), .Y(io_oeb[32]) );
  sky130_fd_sc_hd__clkinv_1 U16461 ( .A(j202_soc_core_j22_cpu_ml_mach[3]), .Y(
        n17710) );
  sky130_fd_sc_hd__clkinv_1 U16462 ( .A(j202_soc_core_j22_cpu_rf_tmp[14]), .Y(
        n14142) );
  sky130_fd_sc_hd__clkinv_1 U16463 ( .A(j202_soc_core_intc_core_00_rg_itgt[60]), .Y(n25749) );
  sky130_fd_sc_hd__clkinv_1 U16464 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[1]), .Y(n26852) );
  sky130_fd_sc_hd__clkinv_1 U16465 ( .A(j202_soc_core_j22_cpu_rf_vbr[19]), .Y(
        n14918) );
  sky130_fd_sc_hd__clkinv_1 U16466 ( .A(j202_soc_core_j22_cpu_rf_gpr[482]), 
        .Y(n21243) );
  sky130_fd_sc_hd__clkinv_1 U16468 ( .A(j202_soc_core_intc_core_00_rg_ipr[19]), 
        .Y(n25324) );
  sky130_fd_sc_hd__clkinv_1 U16469 ( .A(j202_soc_core_j22_cpu_id_opn_inst__13_), .Y(n19858) );
  sky130_fd_sc_hd__clkinv_1 U16470 ( .A(j202_soc_core_j22_cpu_rf_tmp[3]), .Y(
        n21249) );
  sky130_fd_sc_hd__clkinv_1 U16471 ( .A(j202_soc_core_intc_core_00_rg_ipr[93]), 
        .Y(n25491) );
  sky130_fd_sc_hd__clkinv_1 U16472 ( .A(j202_soc_core_j22_cpu_rf_vbr[3]), .Y(
        n21248) );
  sky130_fd_sc_hd__clkinv_1 U16473 ( .A(j202_soc_core_memory0_ram_dout0_sel[5]), .Y(n13176) );
  sky130_fd_sc_hd__clkinv_1 U16474 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[5]), .Y(n11989) );
  sky130_fd_sc_hd__clkinv_1 U16475 ( .A(j202_soc_core_intc_core_00_rg_ipr[55]), 
        .Y(n26740) );
  sky130_fd_sc_hd__clkinv_1 U16476 ( .A(j202_soc_core_cmt_core_00_reg_addr[2]), 
        .Y(n28222) );
  sky130_fd_sc_hd__clkinv_1 U16477 ( .A(j202_soc_core_intc_core_00_rg_itgt[52]), .Y(n25748) );
  sky130_fd_sc_hd__clkinv_1 U16478 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[1]), .Y(n28725) );
  sky130_fd_sc_hd__clkinv_1 U16479 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[15]), .Y(n26093) );
  sky130_fd_sc_hd__clkinv_1 U16480 ( .A(j202_soc_core_j22_cpu_ml_mach[0]), .Y(
        n21687) );
  sky130_fd_sc_hd__clkinv_1 U16481 ( .A(j202_soc_core_intc_core_00_rg_ipr[125]), .Y(n25487) );
  sky130_fd_sc_hd__clkinv_1 U16482 ( .A(j202_soc_core_intc_core_00_rg_ipr[6]), 
        .Y(n25154) );
  sky130_fd_sc_hd__clkinv_1 U16483 ( .A(j202_soc_core_pwrite[1]), .Y(n25061)
         );
  sky130_fd_sc_hd__clkinv_1 U16484 ( .A(j202_soc_core_bldc_core_00_comm[0]), 
        .Y(n29126) );
  sky130_fd_sc_hd__clkinv_1 U16485 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[95]), .Y(n16333) );
  sky130_fd_sc_hd__clkinv_1 U16487 ( .A(j202_soc_core_qspi_wb_wdat[30]), .Y(
        n27993) );
  sky130_fd_sc_hd__clkinv_1 U16488 ( .A(j202_soc_core_gpio_core_00_reg_addr[3]), .Y(n26908) );
  sky130_fd_sc_hd__clkinv_1 U16489 ( .A(j202_soc_core_cmt_core_00_cnt0[3]), 
        .Y(n24977) );
  sky130_fd_sc_hd__clkinv_1 U16490 ( .A(j202_soc_core_intc_core_00_rg_ipr[15]), 
        .Y(n26123) );
  sky130_fd_sc_hd__clkinv_1 U16491 ( .A(j202_soc_core_intc_core_00_rg_ipr[11]), 
        .Y(n26672) );
  sky130_fd_sc_hd__clkinv_1 U16492 ( .A(j202_soc_core_intc_core_00_rg_ie[7]), 
        .Y(n26692) );
  sky130_fd_sc_hd__clkinv_1 U16493 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[9]), .Y(n26477) );
  sky130_fd_sc_hd__clkinv_1 U16494 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[14]), .Y(n29005) );
  sky130_fd_sc_hd__clkinv_1 U16495 ( .A(j202_soc_core_j22_cpu_ml_bufb[31]), 
        .Y(n28434) );
  sky130_fd_sc_hd__clkinv_1 U16496 ( .A(j202_soc_core_intc_core_00_rg_ipr[3]), 
        .Y(n27574) );
  sky130_fd_sc_hd__clkinv_1 U16497 ( .A(j202_soc_core_intc_core_00_bs_addr[5]), 
        .Y(n29414) );
  sky130_fd_sc_hd__clkinv_1 U16498 ( .A(j202_soc_core_j22_cpu_rf_gpr[479]), 
        .Y(n21671) );
  sky130_fd_sc_hd__clkinv_1 U16499 ( .A(j202_soc_core_intc_core_00_rg_ipr[14]), 
        .Y(n25155) );
  sky130_fd_sc_hd__clkinv_1 U16500 ( .A(
        j202_soc_core_memory0_ram_dout0_sel[11]), .Y(n13152) );
  sky130_fd_sc_hd__clkinv_1 U16501 ( .A(j202_soc_core_qspi_wb_wdat[28]), .Y(
        n27391) );
  sky130_fd_sc_hd__clkinv_1 U16502 ( .A(j202_soc_core_intc_core_00_rg_ipr[7]), 
        .Y(n27150) );
  sky130_fd_sc_hd__clkinv_1 U16503 ( .A(j202_soc_core_j22_cpu_rf_pr[5]), .Y(
        n22284) );
  sky130_fd_sc_hd__clkinv_1 U16504 ( .A(j202_soc_core_intc_core_00_bs_addr[7]), 
        .Y(n25084) );
  sky130_fd_sc_hd__clkinv_1 U16505 ( .A(j202_soc_core_j22_cpu_rf_gbr[20]), .Y(
        n22321) );
  sky130_fd_sc_hd__clkinv_1 U16506 ( .A(j202_soc_core_intc_core_00_bs_addr[8]), 
        .Y(n24780) );
  sky130_fd_sc_hd__clkinv_1 U16507 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__0_), 
        .Y(n13341) );
  sky130_fd_sc_hd__clkinv_1 U16508 ( .A(j202_soc_core_wbqspiflash_00_spi_valid), .Y(n27307) );
  sky130_fd_sc_hd__clkinv_1 U16509 ( .A(j202_soc_core_ahb2apb_01_state[1]), 
        .Y(n25037) );
  sky130_fd_sc_hd__clkinv_1 U16510 ( .A(j202_soc_core_qspi_wb_wdat[14]), .Y(
        n28999) );
  sky130_fd_sc_hd__clkinv_1 U16511 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[3]), .Y(n28927) );
  sky130_fd_sc_hd__clkinv_1 U16512 ( .A(j202_soc_core_j22_cpu_rf_tmp[5]), .Y(
        n22288) );
  sky130_fd_sc_hd__clkinv_1 U16513 ( .A(j202_soc_core_intc_core_00_rg_ie[5]), 
        .Y(n26676) );
  sky130_fd_sc_hd__clkinv_1 U16515 ( .A(j202_soc_core_j22_cpu_rf_pr[20]), .Y(
        n14974) );
  sky130_fd_sc_hd__clkinv_1 U16516 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[3]), .Y(n24521) );
  sky130_fd_sc_hd__clkinv_1 U16517 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__1_), 
        .Y(n22287) );
  sky130_fd_sc_hd__clkinv_1 U16518 ( .A(j202_soc_core_j22_cpu_rf_vbr[20]), .Y(
        n14972) );
  sky130_fd_sc_hd__clkinv_1 U16519 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[9]), .Y(n27928) );
  sky130_fd_sc_hd__clkinv_1 U16520 ( .A(gpio_en_o[6]), .Y(io_oeb[26]) );
  sky130_fd_sc_hd__clkinv_1 U16521 ( .A(j202_soc_core_qspi_wb_wdat[26]), .Y(
        n27867) );
  sky130_fd_sc_hd__inv_2 U16522 ( .A(j202_soc_core_bootrom_00_address_w[3]), 
        .Y(n19130) );
  sky130_fd_sc_hd__clkinv_1 U16523 ( .A(j202_soc_core_j22_cpu_rfuo_sr__t_), 
        .Y(n21717) );
  sky130_fd_sc_hd__clkinv_1 U16524 ( .A(j202_soc_core_ahb2apb_01_state[2]), 
        .Y(n25038) );
  sky130_fd_sc_hd__clkinv_1 U16525 ( .A(j202_soc_core_j22_cpu_rf_tmp[20]), .Y(
        n14973) );
  sky130_fd_sc_hd__clkinv_1 U16526 ( .A(j202_soc_core_j22_cpu_rf_vbr[5]), .Y(
        n22286) );
  sky130_fd_sc_hd__clkinv_1 U16527 ( .A(j202_soc_core_ahb2apb_01_state[0]), 
        .Y(n24431) );
  sky130_fd_sc_hd__clkinv_1 U16528 ( .A(j202_soc_core_intc_core_00_rg_ie[9]), 
        .Y(n26715) );
  sky130_fd_sc_hd__clkinv_1 U16529 ( .A(j202_soc_core_intc_core_00_rg_ie[6]), 
        .Y(n26701) );
  sky130_fd_sc_hd__clkinv_1 U16530 ( .A(j202_soc_core_j22_cpu_rf_gpr[484]), 
        .Y(n22283) );
  sky130_fd_sc_hd__clkinv_1 U16531 ( .A(j202_soc_core_cmt_core_00_cnt0[9]), 
        .Y(n25014) );
  sky130_fd_sc_hd__clkinv_1 U16532 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[0]), .Y(n28258) );
  sky130_fd_sc_hd__clkinv_1 U16533 ( .A(j202_soc_core_qspi_wb_wdat[24]), .Y(
        n27651) );
  sky130_fd_sc_hd__inv_1 U16534 ( .A(j202_soc_core_j22_cpu_regop_Rm__2_), .Y(
        n13380) );
  sky130_fd_sc_hd__clkinv_1 U16535 ( .A(j202_soc_core_j22_cpu_rf_gpr[494]), 
        .Y(n18890) );
  sky130_fd_sc_hd__clkinv_1 U16536 ( .A(j202_soc_core_j22_cpu_pc[0]), .Y(
        n13849) );
  sky130_fd_sc_hd__clkinv_1 U16537 ( .A(j202_soc_core_intc_core_00_rg_ie[18]), 
        .Y(n26855) );
  sky130_fd_sc_hd__nor2_1 U16538 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[3]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[5]), .Y(n26208) );
  sky130_fd_sc_hd__clkinv_1 U16539 ( .A(j202_soc_core_intc_core_00_rg_ipr[26]), 
        .Y(n26690) );
  sky130_fd_sc_hd__clkinv_1 U16540 ( .A(j202_soc_core_j22_cpu_rf_gpr[4]), .Y(
        n13751) );
  sky130_fd_sc_hd__clkinv_1 U16541 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[2]), .Y(n28921) );
  sky130_fd_sc_hd__clkinv_1 U16542 ( .A(j202_soc_core_j22_cpu_rf_pr[4]), .Y(
        n21799) );
  sky130_fd_sc_hd__clkinv_1 U16543 ( .A(j202_soc_core_j22_cpu_rf_tmp[8]), .Y(
        n21738) );
  sky130_fd_sc_hd__clkinv_1 U16544 ( .A(j202_soc_core_j22_cpu_regop_imm__4_), 
        .Y(n13599) );
  sky130_fd_sc_hd__clkinv_1 U16545 ( .A(j202_soc_core_intc_core_00_rg_ipr[121]), .Y(n27167) );
  sky130_fd_sc_hd__clkinv_1 U16546 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[2]), 
        .Y(n13286) );
  sky130_fd_sc_hd__clkinv_1 U16547 ( .A(j202_soc_core_intr_vec__2_), .Y(n24787) );
  sky130_fd_sc_hd__clkinv_1 U16548 ( .A(j202_soc_core_j22_cpu_rf_vbr[0]), .Y(
        n13848) );
  sky130_fd_sc_hd__clkinv_1 U16549 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .Y(n23898) );
  sky130_fd_sc_hd__clkinv_1 U16550 ( .A(j202_soc_core_intc_core_00_rg_ipr[89]), 
        .Y(n27169) );
  sky130_fd_sc_hd__clkinv_1 U16551 ( .A(j202_soc_core_intc_core_00_rg_ie[8]), 
        .Y(n26724) );
  sky130_fd_sc_hd__clkinv_1 U16552 ( .A(j202_soc_core_intc_core_00_rg_ipr[57]), 
        .Y(n26754) );
  sky130_fd_sc_hd__clkinv_1 U16553 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[1]), 
        .Y(n29277) );
  sky130_fd_sc_hd__clkinv_1 U16554 ( .A(j202_soc_core_j22_cpu_rf_gpr[6]), .Y(
        n13512) );
  sky130_fd_sc_hd__clkinv_1 U16555 ( .A(j202_soc_core_j22_cpu_ma_M_area[0]), 
        .Y(n13274) );
  sky130_fd_sc_hd__clkinv_1 U16556 ( .A(j202_soc_core_j22_cpu_rfuo_sr__q_), 
        .Y(n21737) );
  sky130_fd_sc_hd__clkinv_1 U16557 ( .A(j202_soc_core_intc_core_00_rg_itgt[50]), .Y(n27937) );
  sky130_fd_sc_hd__clkinv_1 U16558 ( .A(j202_soc_core_intc_core_00_rg_ipr[25]), 
        .Y(n26705) );
  sky130_fd_sc_hd__clkinv_1 U16559 ( .A(j202_soc_core_intc_core_00_rg_ipr[24]), 
        .Y(n26706) );
  sky130_fd_sc_hd__clkinv_1 U16560 ( .A(j202_soc_core_bldc_core_00_comm[1]), 
        .Y(n29121) );
  sky130_fd_sc_hd__clkinv_1 U16561 ( .A(j202_soc_core_j22_cpu_rf_vbr[8]), .Y(
        n14258) );
  sky130_fd_sc_hd__clkinv_1 U16562 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__0_), 
        .Y(n23765) );
  sky130_fd_sc_hd__clkinv_1 U16563 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]), .Y(n24531) );
  sky130_fd_sc_hd__clkinv_1 U16564 ( .A(j202_soc_core_j22_cpu_rf_gpr[487]), 
        .Y(n21734) );
  sky130_fd_sc_hd__clkinv_1 U16565 ( .A(j202_soc_core_intc_core_00_bs_addr[3]), 
        .Y(n29403) );
  sky130_fd_sc_hd__clkinv_1 U16566 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[102]), .Y(n21065) );
  sky130_fd_sc_hd__clkinv_1 U16567 ( .A(j202_soc_core_intc_core_00_bs_addr[2]), 
        .Y(n25072) );
  sky130_fd_sc_hd__clkinv_1 U16569 ( .A(j202_soc_core_intc_core_00_rg_itgt[42]), .Y(n27934) );
  sky130_fd_sc_hd__clkinv_1 U16570 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[0]), .Y(n28780) );
  sky130_fd_sc_hd__clkinv_1 U16571 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__1_), 
        .Y(n24717) );
  sky130_fd_sc_hd__clkinv_1 U16572 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[4]), .Y(n28928) );
  sky130_fd_sc_hd__clkinv_1 U16573 ( .A(
        j202_soc_core_memory0_ram_dout0_sel[13]), .Y(n13148) );
  sky130_fd_sc_hd__clkinv_1 U16574 ( .A(j202_soc_core_intc_core_00_rg_ie[10]), 
        .Y(n25059) );
  sky130_fd_sc_hd__clkinv_1 U16575 ( .A(j202_soc_core_j22_cpu_ml_macl[14]), 
        .Y(n24464) );
  sky130_fd_sc_hd__clkinv_1 U16576 ( .A(j202_soc_core_intc_core_00_bs_addr[9]), 
        .Y(n27414) );
  sky130_fd_sc_hd__clkinv_1 U16577 ( .A(j202_soc_core_j22_cpu_rf_gpr[3]), .Y(
        n13660) );
  sky130_fd_sc_hd__clkinv_1 U16578 ( .A(j202_soc_core_intc_core_00_rg_itgt[34]), .Y(n27933) );
  sky130_fd_sc_hd__buf_4 U16579 ( .A(j202_soc_core_j22_cpu_ml_bufa[32]), .X(
        n22023) );
  sky130_fd_sc_hd__clkinv_1 U16580 ( .A(j202_soc_core_intc_core_00_rg_ipr[4]), 
        .Y(n24827) );
  sky130_fd_sc_hd__clkinv_1 U16581 ( .A(j202_soc_core_intc_core_00_rg_ie[4]), 
        .Y(n26684) );
  sky130_fd_sc_hd__clkinv_1 U16582 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[8]), .Y(n23638) );
  sky130_fd_sc_hd__clkinv_1 U16583 ( .A(j202_soc_core_qspi_wb_wdat[27]), .Y(
        n27070) );
  sky130_fd_sc_hd__clkinv_1 U16584 ( .A(j202_soc_core_intr_vec__4_), .Y(n29068) );
  sky130_fd_sc_hd__clkinv_1 U16585 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[9]), .Y(n27932) );
  sky130_fd_sc_hd__clkinv_1 U16586 ( .A(j202_soc_core_cmt_core_00_cnt0[6]), 
        .Y(n24978) );
  sky130_fd_sc_hd__clkinv_1 U16587 ( .A(j202_soc_core_qspi_wb_wdat[29]), .Y(
        n25484) );
  sky130_fd_sc_hd__clkinv_1 U16588 ( .A(j202_soc_core_j22_cpu_ml_mach[13]), 
        .Y(n24440) );
  sky130_fd_sc_hd__clkinv_1 U16589 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[65]), .Y(n19361) );
  sky130_fd_sc_hd__clkinv_1 U16590 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[0]), 
        .Y(n18799) );
  sky130_fd_sc_hd__clkinv_1 U16591 ( .A(j202_soc_core_j22_cpu_regop_imm__6_), 
        .Y(n13514) );
  sky130_fd_sc_hd__clkinv_1 U16592 ( .A(j202_soc_core_gpio_core_00_reg_addr[0]), .Y(n26777) );
  sky130_fd_sc_hd__clkinv_1 U16593 ( .A(j202_soc_core_intc_core_00_rg_itgt[63]), .Y(n25493) );
  sky130_fd_sc_hd__clkinv_1 U16594 ( .A(j202_soc_core_j22_cpu_ml_macl[30]), 
        .Y(n22561) );
  sky130_fd_sc_hd__clkinv_1 U16595 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[2]), .Y(n28916) );
  sky130_fd_sc_hd__buf_2 U16596 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .X(n21145) );
  sky130_fd_sc_hd__clkinv_1 U16597 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld), .Y(n29117) );
  sky130_fd_sc_hd__clkinv_1 U16598 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[70]), .Y(n21066) );
  sky130_fd_sc_hd__clkinv_1 U16599 ( .A(j202_soc_core_intr_vec__1_), .Y(n28366) );
  sky130_fd_sc_hd__clkinv_1 U16600 ( .A(j202_soc_core_j22_cpu_rf_vbr[21]), .Y(
        n15057) );
  sky130_fd_sc_hd__clkinv_1 U16601 ( .A(j202_soc_core_intc_core_00_rg_ipr[30]), 
        .Y(n26689) );
  sky130_fd_sc_hd__clkinv_1 U16602 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[16]), .Y(n27108) );
  sky130_fd_sc_hd__clkinv_1 U16603 ( .A(j202_soc_core_intc_core_00_rg_ipr[75]), 
        .Y(n26767) );
  sky130_fd_sc_hd__clkinv_1 U16604 ( .A(j202_soc_core_intc_core_00_rg_ipr[58]), 
        .Y(n26742) );
  sky130_fd_sc_hd__clkinv_1 U16605 ( .A(j202_soc_core_j22_cpu_regop_We__2_), 
        .Y(n13305) );
  sky130_fd_sc_hd__clkinv_1 U16606 ( .A(j202_soc_core_j22_cpu_rf_gpr[13]), .Y(
        n14176) );
  sky130_fd_sc_hd__clkinv_1 U16607 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[1]), 
        .Y(n24722) );
  sky130_fd_sc_hd__clkinv_1 U16608 ( .A(j202_soc_core_j22_cpu_rf_tmp[7]), .Y(
        n18867) );
  sky130_fd_sc_hd__clkinv_1 U16609 ( .A(j202_soc_core_qspi_wb_wdat[19]), .Y(
        n25319) );
  sky130_fd_sc_hd__clkinv_1 U16610 ( .A(j202_soc_core_intc_core_00_rg_ipr[28]), 
        .Y(n26707) );
  sky130_fd_sc_hd__clkinv_1 U16611 ( .A(j202_soc_core_intc_core_00_rg_ipr[43]), 
        .Y(n26735) );
  sky130_fd_sc_hd__clkinv_1 U16612 ( .A(j202_soc_core_j22_cpu_regop_imm__7_), 
        .Y(n14225) );
  sky130_fd_sc_hd__clkinv_1 U16613 ( .A(j202_soc_core_j22_cpu_rf_gbr[13]), .Y(
        n14177) );
  sky130_fd_sc_hd__clkinv_1 U16614 ( .A(j202_soc_core_j22_cpu_rf_gpr[507]), 
        .Y(n15966) );
  sky130_fd_sc_hd__clkinv_1 U16615 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[2]), .Y(n13322) );
  sky130_fd_sc_hd__clkinv_1 U16616 ( .A(j202_soc_core_intc_core_00_rg_itgt[28]), .Y(n27100) );
  sky130_fd_sc_hd__clkinv_1 U16618 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[101]), .Y(n21518) );
  sky130_fd_sc_hd__clkinv_1 U16619 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]), .Y(n23646) );
  sky130_fd_sc_hd__clkinv_1 U16620 ( .A(j202_soc_core_j22_cpu_ml_macl[0]), .Y(
        n21708) );
  sky130_fd_sc_hd__clkinv_1 U16621 ( .A(j202_soc_core_intc_core_00_rg_eimk[6]), 
        .Y(n27450) );
  sky130_fd_sc_hd__clkinv_1 U16622 ( .A(j202_soc_core_j22_cpu_rf_gpr[18]), .Y(
        n13476) );
  sky130_fd_sc_hd__clkinv_1 U16623 ( .A(j202_soc_core_bldc_core_00_pwm_duty[7]), .Y(n25315) );
  sky130_fd_sc_hd__clkinv_1 U16624 ( .A(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled), .Y(n27296) );
  sky130_fd_sc_hd__clkinv_1 U16625 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[6]), .Y(n27445) );
  sky130_fd_sc_hd__clkinv_1 U16626 ( .A(j202_soc_core_intc_core_00_rg_itgt[20]), .Y(n27099) );
  sky130_fd_sc_hd__clkinv_1 U16627 ( .A(j202_soc_core_j22_cpu_rf_tmp[28]), .Y(
        n15968) );
  sky130_fd_sc_hd__clkinv_1 U16628 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]), .Y(n28956) );
  sky130_fd_sc_hd__clkinv_1 U16629 ( .A(j202_soc_core_intc_core_00_rg_ipr[76]), 
        .Y(n25192) );
  sky130_fd_sc_hd__clkinv_1 U16630 ( .A(j202_soc_core_intc_core_00_rg_ipr[42]), 
        .Y(n25070) );
  sky130_fd_sc_hd__clkinv_1 U16631 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[2]), .Y(n13278) );
  sky130_fd_sc_hd__clkinv_1 U16632 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]), .Y(n23652) );
  sky130_fd_sc_hd__clkinv_1 U16633 ( .A(gpio_en_o[7]), .Y(io_oeb[27]) );
  sky130_fd_sc_hd__clkinv_1 U16634 ( .A(j202_soc_core_uart_BRG_ps[2]), .Y(
        n28604) );
  sky130_fd_sc_hd__clkinv_1 U16635 ( .A(j202_soc_core_j22_cpu_rf_gpr[5]), .Y(
        n13641) );
  sky130_fd_sc_hd__clkinv_1 U16636 ( .A(
        j202_soc_core_bldc_core_00_hall_value[0]), .Y(n28207) );
  sky130_fd_sc_hd__clkinv_1 U16637 ( .A(j202_soc_core_j22_cpu_rf_gbr[29]), .Y(
        n22999) );
  sky130_fd_sc_hd__clkinv_1 U16638 ( .A(j202_soc_core_intc_core_00_rg_ipr[0]), 
        .Y(n24826) );
  sky130_fd_sc_hd__clkinv_1 U16639 ( .A(j202_soc_core_j22_cpu_rf_tmp[13]), .Y(
        n14174) );
  sky130_fd_sc_hd__clkinv_1 U16640 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[19]), .Y(n29036) );
  sky130_fd_sc_hd__clkinv_1 U16641 ( .A(j202_soc_core_intc_core_00_rg_itgt[12]), .Y(n26738) );
  sky130_fd_sc_hd__clkinv_1 U16642 ( .A(j202_soc_core_j22_cpu_memop_MEM__3_), 
        .Y(n24647) );
  sky130_fd_sc_hd__clkinv_1 U16643 ( .A(la_data_out[0]), .Y(n28253) );
  sky130_fd_sc_hd__clkinv_1 U16644 ( .A(j202_soc_core_intc_core_00_rg_ipr[56]), 
        .Y(n26755) );
  sky130_fd_sc_hd__clkinv_1 U16645 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[5]), .Y(n28941) );
  sky130_fd_sc_hd__clkinv_1 U16646 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[0]), .Y(n24030) );
  sky130_fd_sc_hd__clkinv_1 U16647 ( .A(j202_soc_core_intc_core_00_rg_ipr[71]), 
        .Y(n26766) );
  sky130_fd_sc_hd__clkinv_1 U16648 ( .A(j202_soc_core_j22_cpu_rf_vbr[28]), .Y(
        n15967) );
  sky130_fd_sc_hd__clkinv_1 U16649 ( .A(j202_soc_core_intc_core_00_rg_ipr[80]), 
        .Y(n27098) );
  sky130_fd_sc_hd__clkinv_1 U16650 ( .A(j202_soc_core_intc_core_00_rg_ipr[40]), 
        .Y(n26734) );
  sky130_fd_sc_hd__clkinv_1 U16651 ( .A(j202_soc_core_intc_core_00_rg_ipr[81]), 
        .Y(n25747) );
  sky130_fd_sc_hd__clkinv_1 U16652 ( .A(j202_soc_core_j22_cpu_rf_vbr[13]), .Y(
        n14173) );
  sky130_fd_sc_hd__clkinv_1 U16653 ( .A(j202_soc_core_intc_core_00_rg_itgt[4]), 
        .Y(n26685) );
  sky130_fd_sc_hd__inv_2 U16654 ( .A(j202_soc_core_intc_core_00_rg_ipr[61]), 
        .Y(n25488) );
  sky130_fd_sc_hd__clkinv_1 U16655 ( .A(j202_soc_core_j22_cpu_pc[29]), .Y(
        n23001) );
  sky130_fd_sc_hd__clkinv_1 U16656 ( .A(j202_soc_core_intc_core_00_rg_ipr[83]), 
        .Y(n25325) );
  sky130_fd_sc_hd__clkinv_1 U16657 ( .A(j202_soc_core_intc_core_00_rg_ipr[2]), 
        .Y(n27149) );
  sky130_fd_sc_hd__clkinv_1 U16658 ( .A(j202_soc_core_intc_core_00_rg_ipr[67]), 
        .Y(n27684) );
  sky130_fd_sc_hd__clkinv_1 U16659 ( .A(j202_soc_core_j22_cpu_rf_pr[29]), .Y(
        n16079) );
  sky130_fd_sc_hd__inv_1 U16660 ( .A(j202_soc_core_intc_core_00_rg_ipr[22]), 
        .Y(n25610) );
  sky130_fd_sc_hd__clkinv_1 U16661 ( .A(j202_soc_core_j22_cpu_ml_mach[18]), 
        .Y(n22021) );
  sky130_fd_sc_hd__clkinv_1 U16662 ( .A(j202_soc_core_intc_core_00_bs_addr[4]), 
        .Y(n27417) );
  sky130_fd_sc_hd__clkinv_1 U16663 ( .A(j202_soc_core_intc_core_00_rg_eimk[7]), 
        .Y(n27563) );
  sky130_fd_sc_hd__clkinv_1 U16664 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[66]), .Y(n17196) );
  sky130_fd_sc_hd__inv_2 U16665 ( .A(j202_soc_core_j22_cpu_regop_Rm__3_), .Y(
        n13413) );
  sky130_fd_sc_hd__clkinv_1 U16666 ( .A(j202_soc_core_j22_cpu_ml_macl[16]), 
        .Y(n22764) );
  sky130_fd_sc_hd__clkinv_1 U16667 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]), .Y(n23647) );
  sky130_fd_sc_hd__clkinv_1 U16668 ( .A(j202_soc_core_intc_core_00_rg_ipr[20]), 
        .Y(n26687) );
  sky130_fd_sc_hd__clkinv_1 U16669 ( .A(j202_soc_core_intc_core_00_rg_ipr[36]), 
        .Y(n26728) );
  sky130_fd_sc_hd__clkinv_1 U16670 ( .A(j202_soc_core_j22_cpu_rf_gbr[19]), .Y(
        n22818) );
  sky130_fd_sc_hd__clkinv_1 U16671 ( .A(j202_soc_core_j22_cpu_rf_gpr[11]), .Y(
        n14010) );
  sky130_fd_sc_hd__clkinv_1 U16672 ( .A(j202_soc_core_j22_cpu_rf_vbr[29]), .Y(
        n16076) );
  sky130_fd_sc_hd__clkinv_1 U16673 ( .A(j202_soc_core_intc_core_00_rg_eimk[0]), 
        .Y(n28232) );
  sky130_fd_sc_hd__clkinv_1 U16674 ( .A(j202_soc_core_cmt_core_00_cnt1[6]), 
        .Y(n23942) );
  sky130_fd_sc_hd__clkinv_1 U16675 ( .A(j202_soc_core_intc_core_00_rg_ipr[5]), 
        .Y(n24810) );
  sky130_fd_sc_hd__clkinv_1 U16676 ( .A(j202_soc_core_intr_vec__3_), .Y(n29071) );
  sky130_fd_sc_hd__clkinv_1 U16677 ( .A(j202_soc_core_j22_cpu_rf_tmp[29]), .Y(
        n16078) );
  sky130_fd_sc_hd__clkinv_1 U16678 ( .A(j202_soc_core_intc_core_00_rg_ipr[70]), 
        .Y(n26761) );
  sky130_fd_sc_hd__clkinv_1 U16679 ( .A(j202_soc_core_j22_cpu_regop_imm__5_), 
        .Y(n13542) );
  sky130_fd_sc_hd__clkinv_1 U16680 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[45]), .Y(n20071) );
  sky130_fd_sc_hd__clkinv_1 U16681 ( .A(j202_soc_core_qspi_wb_addr[13]), .Y(
        n28816) );
  sky130_fd_sc_hd__clkinv_1 U16682 ( .A(j202_soc_core_j22_cpu_rf_gpr[20]), .Y(
        n14975) );
  sky130_fd_sc_hd__clkinv_1 U16683 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[1]), .Y(n28307) );
  sky130_fd_sc_hd__clkinv_1 U16684 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[0]), .Y(n17189) );
  sky130_fd_sc_hd__clkinv_1 U16685 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[2]), .Y(n26568) );
  sky130_fd_sc_hd__clkinv_1 U16686 ( .A(j202_soc_core_cmt_core_00_cnt1[5]), 
        .Y(n27543) );
  sky130_fd_sc_hd__clkinv_1 U16687 ( .A(j202_soc_core_j22_cpu_rf_pr[13]), .Y(
        n22984) );
  sky130_fd_sc_hd__clkinv_1 U16688 ( .A(j202_soc_core_intc_core_00_rg_eimk[1]), 
        .Y(n29078) );
  sky130_fd_sc_hd__clkinv_1 U16689 ( .A(gpio_en_o[4]), .Y(io_oeb[4]) );
  sky130_fd_sc_hd__clkinv_1 U16690 ( .A(j202_soc_core_j22_cpu_ml_mach[19]), 
        .Y(n22022) );
  sky130_fd_sc_hd__clkinv_1 U16691 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .Y(n23649) );
  sky130_fd_sc_hd__clkinv_1 U16692 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[19]), .Y(n29038) );
  sky130_fd_sc_hd__clkinv_1 U16693 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[1]), .Y(n17190) );
  sky130_fd_sc_hd__clkinv_1 U16694 ( .A(j202_soc_core_j22_cpu_ml_mach[20]), 
        .Y(n22018) );
  sky130_fd_sc_hd__clkinv_1 U16695 ( .A(j202_soc_core_cmt_core_00_cnt0[4]), 
        .Y(n27489) );
  sky130_fd_sc_hd__nor2_1 U16696 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[1]), .B(
        j202_soc_core_j22_cpu_ma_M_MEM[0]), .Y(n11985) );
  sky130_fd_sc_hd__clkinv_1 U16697 ( .A(j202_soc_core_intc_core_00_rg_ie[16]), 
        .Y(n26763) );
  sky130_fd_sc_hd__clkinv_1 U16698 ( .A(j202_soc_core_j22_cpu_memop_Ma__0_), 
        .Y(n13379) );
  sky130_fd_sc_hd__clkinv_1 U16699 ( .A(
        j202_soc_core_wbqspiflash_00_write_protect), .Y(n27407) );
  sky130_fd_sc_hd__clkinv_1 U16700 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[10]), .Y(n28971) );
  sky130_fd_sc_hd__clkinv_1 U16701 ( .A(j202_soc_core_j22_cpu_pc[3]), .Y(
        n20446) );
  sky130_fd_sc_hd__clkinv_1 U16702 ( .A(j202_soc_core_cmt_core_00_cnt0[12]), 
        .Y(n25176) );
  sky130_fd_sc_hd__clkinv_1 U16703 ( .A(gpio_en_o[13]), .Y(io_oeb[33]) );
  sky130_fd_sc_hd__clkinv_1 U16704 ( .A(j202_soc_core_j22_cpu_rf_vbr[30]), .Y(
        n16527) );
  sky130_fd_sc_hd__clkinv_1 U16705 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[1]), .Y(n28566) );
  sky130_fd_sc_hd__clkinv_1 U16706 ( .A(gpio_en_o[15]), .Y(io_oeb[35]) );
  sky130_fd_sc_hd__clkinv_1 U16707 ( .A(j202_soc_core_j22_cpu_rf_tmp[30]), .Y(
        n16528) );
  sky130_fd_sc_hd__clkinv_1 U16708 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[18]), .Y(n27141) );
  sky130_fd_sc_hd__clkinv_1 U16709 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[69]), .Y(n21511) );
  sky130_fd_sc_hd__clkinv_1 U16710 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[0]), .Y(n23904) );
  sky130_fd_sc_hd__clkinv_1 U16711 ( .A(j202_soc_core_gpio_core_00_reg_addr[2]), .Y(n23856) );
  sky130_fd_sc_hd__clkinv_1 U16712 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__3_), 
        .Y(n23831) );
  sky130_fd_sc_hd__clkinv_1 U16713 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[1]), .Y(n28294) );
  sky130_fd_sc_hd__clkinv_1 U16714 ( .A(j202_soc_core_cmt_core_00_cnt0[10]), 
        .Y(n25019) );
  sky130_fd_sc_hd__clkinv_1 U16716 ( .A(j202_soc_core_j22_cpu_rf_gpr[509]), 
        .Y(n16526) );
  sky130_fd_sc_hd__clkinv_1 U16717 ( .A(j202_soc_core_intc_core_00_rg_ipr[35]), 
        .Y(n26729) );
  sky130_fd_sc_hd__clkinv_1 U16718 ( .A(j202_soc_core_j22_cpu_rf_gpr[486]), 
        .Y(n18871) );
  sky130_fd_sc_hd__clkinv_1 U16719 ( .A(j202_soc_core_intc_core_00_rg_ie[26]), 
        .Y(n27871) );
  sky130_fd_sc_hd__clkinv_1 U16720 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[0]), .Y(n28250) );
  sky130_fd_sc_hd__clkinv_1 U16721 ( .A(j202_soc_core_qspi_wb_cyc), .Y(n27226)
         );
  sky130_fd_sc_hd__clkinv_1 U16722 ( .A(j202_soc_core_j22_cpu_rf_gpr[485]), 
        .Y(n22151) );
  sky130_fd_sc_hd__clkinv_1 U16723 ( .A(j202_soc_core_intc_core_00_rg_ipr[73]), 
        .Y(n27936) );
  sky130_fd_sc_hd__clkinv_1 U16724 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[6]), .Y(n28948) );
  sky130_fd_sc_hd__clkinv_1 U16725 ( .A(j202_soc_core_j22_cpu_rf_gpr[7]), .Y(
        n18864) );
  sky130_fd_sc_hd__clkinv_1 U16726 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[20]), .Y(n27379) );
  sky130_fd_sc_hd__clkinv_1 U16727 ( .A(j202_soc_core_intc_core_00_rg_ipr[72]), 
        .Y(n27970) );
  sky130_fd_sc_hd__clkinv_1 U16728 ( .A(j202_soc_core_cmt_core_00_cnt0[14]), 
        .Y(n26105) );
  sky130_fd_sc_hd__clkinv_1 U16729 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[17]), .Y(n29024) );
  sky130_fd_sc_hd__clkinv_1 U16730 ( .A(j202_soc_core_wbqspiflash_00_spi_in[0]), .Y(n29139) );
  sky130_fd_sc_hd__clkinv_1 U16731 ( .A(j202_soc_core_j22_cpu_rf_gbr[7]), .Y(
        n14289) );
  sky130_fd_sc_hd__clkinv_1 U16732 ( .A(j202_soc_core_aquc_CE__1_), .Y(n22413)
         );
  sky130_fd_sc_hd__clkbuf_1 U16733 ( .A(j202_soc_core_j22_cpu_ml_bufa[14]), 
        .X(n24454) );
  sky130_fd_sc_hd__clkinv_1 U16734 ( .A(j202_soc_core_uart_BRG_ps[4]), .Y(
        n28611) );
  sky130_fd_sc_hd__clkinv_1 U16735 ( .A(
        j202_soc_core_bldc_core_00_hall_value[1]), .Y(n28279) );
  sky130_fd_sc_hd__clkinv_1 U16736 ( .A(j202_soc_core_bldc_core_00_pwm_duty[5]), .Y(n25759) );
  sky130_fd_sc_hd__clkinv_1 U16737 ( .A(j202_soc_core_j22_cpu_ml_mach[17]), 
        .Y(n22034) );
  sky130_fd_sc_hd__buf_4 U16738 ( .A(j202_soc_core_j22_cpu_ml_bufa[5]), .X(
        n24366) );
  sky130_fd_sc_hd__clkinv_1 U16739 ( .A(j202_soc_core_j22_cpu_ml_macl[27]), 
        .Y(n22522) );
  sky130_fd_sc_hd__clkinv_1 U16740 ( .A(gpio_en_o[14]), .Y(io_oeb[34]) );
  sky130_fd_sc_hd__clkinv_1 U16741 ( .A(j202_soc_core_cmt_core_00_cnt0[7]), 
        .Y(n25008) );
  sky130_fd_sc_hd__clkinv_1 U16742 ( .A(j202_soc_core_qspi_wb_we), .Y(n27238)
         );
  sky130_fd_sc_hd__clkinv_1 U16743 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[21]), .Y(n25591) );
  sky130_fd_sc_hd__clkinv_1 U16744 ( .A(j202_soc_core_intc_core_00_rg_ipr[68]), 
        .Y(n27497) );
  sky130_fd_sc_hd__clkinv_1 U16745 ( .A(j202_soc_core_intc_core_00_rg_eimk[4]), 
        .Y(n27498) );
  sky130_fd_sc_hd__clkinv_1 U16746 ( .A(j202_soc_core_gpio_core_00_reg_addr[4]), .Y(n26909) );
  sky130_fd_sc_hd__clkinv_1 U16747 ( .A(j202_soc_core_intc_core_00_rg_ipr[74]), 
        .Y(n25076) );
  sky130_fd_sc_hd__clkinv_1 U16748 ( .A(j202_soc_core_j22_cpu_rf_pr[1]), .Y(
        n21985) );
  sky130_fd_sc_hd__clkinv_1 U16749 ( .A(j202_soc_core_bldc_core_00_pwm_duty[4]), .Y(n27110) );
  sky130_fd_sc_hd__clkinv_1 U16750 ( .A(j202_soc_core_intc_core_00_rg_ipr[66]), 
        .Y(n28182) );
  sky130_fd_sc_hd__clkinv_1 U16751 ( .A(gpio_en_o[2]), .Y(io_oeb[2]) );
  sky130_fd_sc_hd__clkinv_1 U16752 ( .A(j202_soc_core_j22_cpu_regop_We__3_), 
        .Y(n23888) );
  sky130_fd_sc_hd__clkinv_1 U16753 ( .A(gpio_en_o[8]), .Y(io_oeb[28]) );
  sky130_fd_sc_hd__clkinv_1 U16754 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[19]), .Y(n25717) );
  sky130_fd_sc_hd__clkinv_1 U16755 ( .A(j202_soc_core_j22_cpu_rf_vbr[7]), .Y(
        n18874) );
  sky130_fd_sc_hd__clkinv_1 U16756 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__3_), 
        .Y(n18866) );
  sky130_fd_sc_hd__clkinv_1 U16757 ( .A(j202_soc_core_intc_core_00_rg_ipr[79]), 
        .Y(n26124) );
  sky130_fd_sc_hd__clkinv_1 U16758 ( .A(j202_soc_core_intc_core_00_rg_ipr[59]), 
        .Y(n26757) );
  sky130_fd_sc_hd__clkinv_1 U16761 ( .A(j202_soc_core_qspi_wb_wdat[16]), .Y(
        n27096) );
  sky130_fd_sc_hd__clkinv_1 U16762 ( .A(j202_soc_core_j22_cpu_ml_macl[11]), 
        .Y(n18078) );
  sky130_fd_sc_hd__clkinv_1 U16763 ( .A(j202_soc_core_intc_core_00_rg_ipr[78]), 
        .Y(n26883) );
  sky130_fd_sc_hd__clkinv_1 U16764 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[5]), .Y(n27409) );
  sky130_fd_sc_hd__clkinv_1 U16765 ( .A(j202_soc_core_intc_core_00_rg_eimk[3]), 
        .Y(n27686) );
  sky130_fd_sc_hd__clkinv_1 U16766 ( .A(j202_soc_core_intc_core_00_rg_ie[0]), 
        .Y(n24816) );
  sky130_fd_sc_hd__clkinv_1 U16767 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[0]), 
        .Y(n27957) );
  sky130_fd_sc_hd__clkinv_1 U16768 ( .A(gpio_en_o[5]), .Y(io_oeb[7]) );
  sky130_fd_sc_hd__and2_0 U16769 ( .A(j202_soc_core_j22_cpu_ml_M_macop_MAC_[3]), .B(j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .X(n13075) );
  sky130_fd_sc_hd__clkinv_1 U16770 ( .A(j202_soc_core_qspi_wb_addr[24]), .Y(
        n23644) );
  sky130_fd_sc_hd__clkinv_1 U16771 ( .A(j202_soc_core_intc_core_00_rg_eimk[5]), 
        .Y(n27419) );
  sky130_fd_sc_hd__or2_0 U16772 ( .A(io_in[37]), .B(wb_rst_i), .X(n3) );
  sky130_fd_sc_hd__nand2_1 U16899 ( .A(n11335), .B(n11334), .Y(n18390) );
  sky130_fd_sc_hd__nand2_1 U16900 ( .A(n18355), .B(n11336), .Y(n11334) );
  sky130_fd_sc_hd__o21ai_1 U16901 ( .A1(n11336), .A2(n18355), .B1(n18354), .Y(
        n11335) );
  sky130_fd_sc_hd__inv_2 U16902 ( .A(n11338), .Y(n11336) );
  sky130_fd_sc_hd__xor2_1 U16903 ( .A(n18354), .B(n11337), .X(n18409) );
  sky130_fd_sc_hd__xnor2_1 U16904 ( .A(n11338), .B(n18355), .Y(n11337) );
  sky130_fd_sc_hd__a2bb2oi_2 U16905 ( .B1(n11340), .B2(n11339), .A1_N(n18474), 
        .A2_N(n17429), .Y(n11338) );
  sky130_fd_sc_hd__inv_2 U16906 ( .A(n18356), .Y(n11339) );
  sky130_fd_sc_hd__inv_1 U16907 ( .A(n18471), .Y(n11340) );
  sky130_fd_sc_hd__fah_1 U16908 ( .A(n18447), .B(n18446), .CI(n18445), .COUT(
        n18456), .SUM(n18449) );
  sky130_fd_sc_hd__nand2_1 U16910 ( .A(n11342), .B(n11341), .Y(n18639) );
  sky130_fd_sc_hd__nand2_1 U16911 ( .A(n18624), .B(n18625), .Y(n11341) );
  sky130_fd_sc_hd__nand2_1 U16912 ( .A(n11347), .B(n11343), .Y(n11342) );
  sky130_fd_sc_hd__nand2_1 U16913 ( .A(n11345), .B(n11344), .Y(n11343) );
  sky130_fd_sc_hd__xnor2_1 U16914 ( .A(n11347), .B(n11346), .Y(n18633) );
  sky130_fd_sc_hd__xnor2_1 U16915 ( .A(n18625), .B(n18624), .Y(n11346) );
  sky130_fd_sc_hd__nand2_1 U16916 ( .A(n18612), .B(n18611), .Y(n11347) );
  sky130_fd_sc_hd__clkbuf_1 U16919 ( .A(j202_soc_core_j22_cpu_ml_bufa[13]), 
        .X(n11350) );
  sky130_fd_sc_hd__nand2_2 U16921 ( .A(n18686), .B(n18336), .Y(n18337) );
  sky130_fd_sc_hd__nand2_1 U16922 ( .A(n11353), .B(n11352), .Y(n18300) );
  sky130_fd_sc_hd__nand2_1 U16923 ( .A(n18063), .B(n18064), .Y(n11352) );
  sky130_fd_sc_hd__o21ai_1 U16924 ( .A1(n18063), .A2(n18064), .B1(n18062), .Y(
        n11353) );
  sky130_fd_sc_hd__xnor2_1 U16925 ( .A(n18062), .B(n11354), .Y(n18304) );
  sky130_fd_sc_hd__xnor2_1 U16926 ( .A(n18064), .B(n18063), .Y(n11354) );
  sky130_fd_sc_hd__xnor2_1 U16927 ( .A(n11350), .B(n17452), .Y(n17454) );
  sky130_fd_sc_hd__nand3_2 U16928 ( .A(n20973), .B(n21020), .C(n11712), .Y(
        n11711) );
  sky130_fd_sc_hd__nand3_2 U16929 ( .A(n12643), .B(n12635), .C(n12639), .Y(
        n20973) );
  sky130_fd_sc_hd__xnor2_1 U16932 ( .A(n17639), .B(n11355), .Y(n17685) );
  sky130_fd_sc_hd__xnor2_1 U16933 ( .A(n17641), .B(n17640), .Y(n11355) );
  sky130_fd_sc_hd__nand2_1 U16934 ( .A(n17659), .B(n17660), .Y(n12679) );
  sky130_fd_sc_hd__nand2_1 U16935 ( .A(n11357), .B(n11356), .Y(n17660) );
  sky130_fd_sc_hd__nand2_1 U16936 ( .A(n17640), .B(n17641), .Y(n11356) );
  sky130_fd_sc_hd__o21ai_1 U16937 ( .A1(n17640), .A2(n17641), .B1(n17639), .Y(
        n11357) );
  sky130_fd_sc_hd__nand2_1 U16940 ( .A(n11596), .B(n10981), .Y(n12822) );
  sky130_fd_sc_hd__inv_2 U16941 ( .A(n11358), .Y(n13035) );
  sky130_fd_sc_hd__nand3_2 U16942 ( .A(n11711), .B(n11710), .C(n19847), .Y(
        n11358) );
  sky130_fd_sc_hd__o21ai_1 U16943 ( .A1(n18592), .A2(n18593), .B1(n18591), .Y(
        n18595) );
  sky130_fd_sc_hd__nand2_1 U16944 ( .A(n11113), .B(n11359), .Y(n12052) );
  sky130_fd_sc_hd__o22ai_1 U16945 ( .A1(n18533), .A2(n17630), .B1(n17595), 
        .B2(n18530), .Y(n17610) );
  sky130_fd_sc_hd__a21oi_1 U16946 ( .A1(n22959), .A2(n17868), .B1(n17867), .Y(
        n17869) );
  sky130_fd_sc_hd__nor2_1 U16948 ( .A(n24543), .B(n23381), .Y(n28116) );
  sky130_fd_sc_hd__nand2_2 U16949 ( .A(n12324), .B(n23378), .Y(n23947) );
  sky130_fd_sc_hd__nand2_1 U16951 ( .A(n11361), .B(n11360), .Y(n17683) );
  sky130_fd_sc_hd__nand2_1 U16952 ( .A(n17607), .B(n17606), .Y(n11360) );
  sky130_fd_sc_hd__o21ai_1 U16953 ( .A1(n17606), .A2(n17607), .B1(n17605), .Y(
        n11361) );
  sky130_fd_sc_hd__xnor2_1 U16954 ( .A(n17605), .B(n11362), .Y(n17572) );
  sky130_fd_sc_hd__xnor2_1 U16955 ( .A(n17606), .B(n17607), .Y(n11362) );
  sky130_fd_sc_hd__nand4_1 U16956 ( .A(n12762), .B(n12754), .C(n12763), .D(
        n12753), .Y(n11364) );
  sky130_fd_sc_hd__nor2_1 U16957 ( .A(n11364), .B(n11363), .Y(n11365) );
  sky130_fd_sc_hd__nand2_1 U16959 ( .A(n11366), .B(n11365), .Y(n11370) );
  sky130_fd_sc_hd__nor2_1 U16960 ( .A(n11368), .B(n11367), .Y(n11366) );
  sky130_fd_sc_hd__nand4_1 U16961 ( .A(n12760), .B(n12752), .C(n12755), .D(
        n11738), .Y(n11367) );
  sky130_fd_sc_hd__nand4_1 U16962 ( .A(n11736), .B(n11737), .C(n12761), .D(
        n12802), .Y(n11368) );
  sky130_fd_sc_hd__nand4_1 U16963 ( .A(n12760), .B(n12763), .C(n12762), .D(
        n12761), .Y(n12759) );
  sky130_fd_sc_hd__nand4_1 U16964 ( .A(n12752), .B(n12755), .C(n12753), .D(
        n12754), .Y(n12764) );
  sky130_fd_sc_hd__nand4_1 U16966 ( .A(n11371), .B(n12129), .C(n12919), .D(
        n12512), .Y(n12511) );
  sky130_fd_sc_hd__nand2_1 U16968 ( .A(n12513), .B(n20462), .Y(n11371) );
  sky130_fd_sc_hd__inv_1 U16969 ( .A(n11373), .Y(n11909) );
  sky130_fd_sc_hd__nand2_1 U16970 ( .A(n12335), .B(n11373), .Y(n12001) );
  sky130_fd_sc_hd__o21a_1 U16971 ( .A1(n11424), .A2(n11373), .B1(n11372), .X(
        n27905) );
  sky130_fd_sc_hd__nand2_1 U16972 ( .A(n11002), .B(n24102), .Y(n11372) );
  sky130_fd_sc_hd__nand2_2 U16973 ( .A(n11532), .B(n12227), .Y(n11373) );
  sky130_fd_sc_hd__nor2b_1 U16978 ( .B_N(n23618), .A(n23620), .Y(n11437) );
  sky130_fd_sc_hd__nand4_1 U16979 ( .A(n24612), .B(n24410), .C(n28123), .D(
        n11375), .Y(n24415) );
  sky130_fd_sc_hd__nor2_1 U16980 ( .A(n27884), .B(n24408), .Y(n11375) );
  sky130_fd_sc_hd__nor2_2 U16981 ( .A(n28348), .B(n12288), .Y(n24612) );
  sky130_fd_sc_hd__nand2_1 U16984 ( .A(n12583), .B(n11449), .Y(n11377) );
  sky130_fd_sc_hd__nand2_2 U16985 ( .A(n23456), .B(n12239), .Y(n11449) );
  sky130_fd_sc_hd__inv_1 U16987 ( .A(n24610), .Y(n11379) );
  sky130_fd_sc_hd__a2bb2oi_2 U16988 ( .B1(n23399), .B2(n23400), .A1_N(n28409), 
        .A2_N(n24573), .Y(n27734) );
  sky130_fd_sc_hd__inv_2 U16989 ( .A(n11636), .Y(n11532) );
  sky130_fd_sc_hd__nand3_2 U16990 ( .A(n11728), .B(n12316), .C(n11580), .Y(
        n11636) );
  sky130_fd_sc_hd__nand2_1 U16991 ( .A(n12770), .B(n19851), .Y(n23509) );
  sky130_fd_sc_hd__nand3_1 U16992 ( .A(n11891), .B(n11887), .C(n11886), .Y(
        n12770) );
  sky130_fd_sc_hd__and2_1 U16994 ( .A(n20089), .B(n21917), .X(n11928) );
  sky130_fd_sc_hd__nand4_1 U16996 ( .A(n20871), .B(n20866), .C(n20867), .D(
        n11476), .Y(n11381) );
  sky130_fd_sc_hd__nand2_2 U16998 ( .A(n12283), .B(n21917), .Y(n11382) );
  sky130_fd_sc_hd__nor2_2 U16999 ( .A(n21681), .B(n21957), .Y(n18658) );
  sky130_fd_sc_hd__nand4_1 U17000 ( .A(n24617), .B(n11098), .C(n24401), .D(
        n24400), .Y(n24403) );
  sky130_fd_sc_hd__o22ai_1 U17001 ( .A1(n18474), .A2(n18473), .B1(n18472), 
        .B2(n18471), .Y(n18534) );
  sky130_fd_sc_hd__nand2_4 U17002 ( .A(n18474), .B(n17335), .Y(n18471) );
  sky130_fd_sc_hd__nor2_1 U17003 ( .A(n23550), .B(n11636), .Y(n24550) );
  sky130_fd_sc_hd__inv_2 U17004 ( .A(n24505), .Y(n24506) );
  sky130_fd_sc_hd__nand2_2 U17006 ( .A(j202_soc_core_memory0_ram_dout0[300]), 
        .B(n21503), .Y(n20903) );
  sky130_fd_sc_hd__clkinv_1 U17007 ( .A(n12273), .Y(n11608) );
  sky130_fd_sc_hd__nand3_1 U17008 ( .A(n12767), .B(n12765), .C(n12850), .Y(
        n11383) );
  sky130_fd_sc_hd__nand2_1 U17010 ( .A(n11385), .B(n24579), .Y(n23616) );
  sky130_fd_sc_hd__nor2_1 U17011 ( .A(n23608), .B(n11386), .Y(n11385) );
  sky130_fd_sc_hd__nand2_1 U17012 ( .A(n30073), .B(n24110), .Y(n11386) );
  sky130_fd_sc_hd__nand2_1 U17013 ( .A(n28037), .B(n12815), .Y(n23402) );
  sky130_fd_sc_hd__nand2_4 U17014 ( .A(n11387), .B(n12220), .Y(n24564) );
  sky130_fd_sc_hd__inv_2 U17015 ( .A(n12324), .Y(n11387) );
  sky130_fd_sc_hd__inv_1 U17016 ( .A(n24639), .Y(n11631) );
  sky130_fd_sc_hd__nand3_2 U17017 ( .A(n27991), .B(n23557), .C(n24968), .Y(
        n23397) );
  sky130_fd_sc_hd__nor2_1 U17018 ( .A(n12815), .B(n12236), .Y(n23379) );
  sky130_fd_sc_hd__nand2_1 U17019 ( .A(n23408), .B(n11006), .Y(n12236) );
  sky130_fd_sc_hd__inv_1 U17020 ( .A(n23387), .Y(n11580) );
  sky130_fd_sc_hd__nand3_2 U17024 ( .A(n12498), .B(n12496), .C(n12497), .Y(
        n25349) );
  sky130_fd_sc_hd__clkbuf_1 U17025 ( .A(n12064), .X(n11389) );
  sky130_fd_sc_hd__nand2_1 U17026 ( .A(n24640), .B(n11106), .Y(n11519) );
  sky130_fd_sc_hd__inv_1 U17027 ( .A(n11724), .Y(n23456) );
  sky130_fd_sc_hd__nand2_1 U17029 ( .A(n11390), .B(n20454), .Y(n12656) );
  sky130_fd_sc_hd__nand4_1 U17030 ( .A(n11396), .B(n12833), .C(n12831), .D(
        n12832), .Y(n11390) );
  sky130_fd_sc_hd__xnor2_1 U17031 ( .A(n17829), .B(n11391), .Y(n11777) );
  sky130_fd_sc_hd__xnor2_1 U17032 ( .A(n17830), .B(n17831), .Y(n11391) );
  sky130_fd_sc_hd__xnor3_1 U17033 ( .A(n17815), .B(n17813), .C(n11429), .X(
        n17830) );
  sky130_fd_sc_hd__clkbuf_1 U17034 ( .A(j202_soc_core_j22_cpu_ml_bufa[18]), 
        .X(n11392) );
  sky130_fd_sc_hd__nand2_2 U17036 ( .A(j202_soc_core_memory0_ram_dout0[268]), 
        .B(n21634), .Y(n20914) );
  sky130_fd_sc_hd__nand2b_4 U17037 ( .A_N(n11487), .B(n29595), .Y(n27739) );
  sky130_fd_sc_hd__nand3_2 U17038 ( .A(n23386), .B(n23387), .C(n11142), .Y(
        n11487) );
  sky130_fd_sc_hd__nor2_1 U17041 ( .A(n11394), .B(n11940), .Y(n11450) );
  sky130_fd_sc_hd__nand4_1 U17042 ( .A(n12450), .B(n12451), .C(n15662), .D(
        n15658), .Y(n11394) );
  sky130_fd_sc_hd__nand4_1 U17044 ( .A(n12866), .B(n12867), .C(n12868), .D(
        n15471), .Y(n12531) );
  sky130_fd_sc_hd__inv_2 U17045 ( .A(n11178), .Y(n12326) );
  sky130_fd_sc_hd__nor2_1 U17046 ( .A(n24621), .B(n12944), .Y(n12943) );
  sky130_fd_sc_hd__inv_2 U17048 ( .A(n25433), .Y(n25466) );
  sky130_fd_sc_hd__inv_2 U17051 ( .A(n12325), .Y(n23426) );
  sky130_fd_sc_hd__nand2_1 U17052 ( .A(j202_soc_core_memory0_ram_dout0[406]), 
        .B(n21496), .Y(n11396) );
  sky130_fd_sc_hd__nor2b_1 U17053 ( .B_N(n24618), .A(n23608), .Y(n12945) );
  sky130_fd_sc_hd__inv_1 U17054 ( .A(n11452), .Y(n11451) );
  sky130_fd_sc_hd__nand2_1 U17057 ( .A(n11399), .B(n11486), .Y(n22121) );
  sky130_fd_sc_hd__and2_0 U17059 ( .A(n22118), .B(n25263), .X(n11400) );
  sky130_fd_sc_hd__inv_8 U17060 ( .A(n23988), .Y(n29755) );
  sky130_fd_sc_hd__inv_8 U17061 ( .A(n23984), .Y(n29758) );
  sky130_fd_sc_hd__inv_8 U17062 ( .A(n23987), .Y(n29756) );
  sky130_fd_sc_hd__inv_8 U17063 ( .A(n23985), .Y(n29757) );
  sky130_fd_sc_hd__inv_8 U17064 ( .A(n23983), .Y(n29759) );
  sky130_fd_sc_hd__a21boi_2 U17065 ( .A1(n19243), .A2(n19241), .B1_N(n19240), 
        .Y(n21217) );
  sky130_fd_sc_hd__nand2_1 U17066 ( .A(n21939), .B(n11143), .Y(n11401) );
  sky130_fd_sc_hd__clkbuf_1 U17067 ( .A(n18923), .X(n11402) );
  sky130_fd_sc_hd__inv_1 U17068 ( .A(n24469), .Y(n26872) );
  sky130_fd_sc_hd__inv_2 U17069 ( .A(n17356), .Y(n17965) );
  sky130_fd_sc_hd__nand2_1 U17070 ( .A(n22937), .B(n24452), .Y(n25259) );
  sky130_fd_sc_hd__nand3_1 U17071 ( .A(n12390), .B(n25279), .C(n11414), .Y(
        n11413) );
  sky130_fd_sc_hd__inv_6 U17072 ( .A(n30080), .Y(n11866) );
  sky130_fd_sc_hd__nor2_1 U17073 ( .A(n11404), .B(n11918), .Y(n11917) );
  sky130_fd_sc_hd__nand4_1 U17074 ( .A(n20901), .B(n20902), .C(n20903), .D(
        n11919), .Y(n11404) );
  sky130_fd_sc_hd__o21ai_1 U17075 ( .A1(n11856), .A2(n21189), .B1(n21190), .Y(
        n22196) );
  sky130_fd_sc_hd__nor2_1 U17076 ( .A(n11405), .B(n12433), .Y(n23489) );
  sky130_fd_sc_hd__nand2_1 U17077 ( .A(n11477), .B(n23488), .Y(n11405) );
  sky130_fd_sc_hd__or2_0 U17078 ( .A(n12065), .B(n25397), .X(n26920) );
  sky130_fd_sc_hd__xnor2_1 U17079 ( .A(n18527), .B(n11406), .Y(n18606) );
  sky130_fd_sc_hd__xnor2_1 U17080 ( .A(n18529), .B(n18528), .Y(n11406) );
  sky130_fd_sc_hd__nand2_1 U17081 ( .A(n11408), .B(n11407), .Y(n18522) );
  sky130_fd_sc_hd__nand2_1 U17082 ( .A(n18505), .B(n11410), .Y(n11407) );
  sky130_fd_sc_hd__o21ai_1 U17083 ( .A1(n11410), .A2(n18505), .B1(n18504), .Y(
        n11408) );
  sky130_fd_sc_hd__xnor3_1 U17084 ( .A(n11410), .B(n18505), .C(n11409), .X(
        n18620) );
  sky130_fd_sc_hd__nand2_1 U17085 ( .A(n11412), .B(n11411), .Y(n11410) );
  sky130_fd_sc_hd__nand2_1 U17086 ( .A(n18528), .B(n18529), .Y(n11411) );
  sky130_fd_sc_hd__o21ai_1 U17087 ( .A1(n18529), .A2(n18528), .B1(n18527), .Y(
        n11412) );
  sky130_fd_sc_hd__nand2_1 U17088 ( .A(n26022), .B(n26021), .Y(n26027) );
  sky130_fd_sc_hd__nand3_1 U17089 ( .A(n23505), .B(n12410), .C(n23514), .Y(
        n26160) );
  sky130_fd_sc_hd__nand3_2 U17090 ( .A(n23504), .B(n23502), .C(n23503), .Y(
        n18797) );
  sky130_fd_sc_hd__nand2_1 U17091 ( .A(n26963), .B(n26962), .Y(n27778) );
  sky130_fd_sc_hd__inv_1 U17092 ( .A(n11413), .Y(n25284) );
  sky130_fd_sc_hd__nand2_2 U17093 ( .A(j202_soc_core_memory0_ram_dout0[332]), 
        .B(n21490), .Y(n20913) );
  sky130_fd_sc_hd__nand3_2 U17095 ( .A(n23443), .B(n23442), .C(n23441), .Y(
        n12288) );
  sky130_fd_sc_hd__nor2_2 U17096 ( .A(n24792), .B(n19430), .Y(n21919) );
  sky130_fd_sc_hd__nand2_1 U17098 ( .A(n11161), .B(n11415), .Y(n10538) );
  sky130_fd_sc_hd__nand2_1 U17099 ( .A(n24132), .B(n28417), .Y(n11415) );
  sky130_fd_sc_hd__nand2_1 U17100 ( .A(n25149), .B(n25147), .Y(n24141) );
  sky130_fd_sc_hd__nand3_1 U17101 ( .A(n23489), .B(n23491), .C(n23490), .Y(
        n23494) );
  sky130_fd_sc_hd__nand2_1 U17103 ( .A(n18242), .B(n11416), .Y(n12889) );
  sky130_fd_sc_hd__o21ai_1 U17104 ( .A1(n19279), .A2(n18265), .B1(n18264), .Y(
        n21880) );
  sky130_fd_sc_hd__clkbuf_1 U17105 ( .A(j202_soc_core_j22_cpu_ml_bufa[15]), 
        .X(n11417) );
  sky130_fd_sc_hd__xor2_1 U17106 ( .A(n11418), .B(n12476), .X(n18325) );
  sky130_fd_sc_hd__xnor2_1 U17107 ( .A(n17948), .B(n17947), .Y(n11418) );
  sky130_fd_sc_hd__nand2_1 U17108 ( .A(n11420), .B(n11419), .Y(n17807) );
  sky130_fd_sc_hd__nand2_1 U17109 ( .A(n17777), .B(n17776), .Y(n11419) );
  sky130_fd_sc_hd__o21ai_1 U17110 ( .A1(n17776), .A2(n17777), .B1(n17775), .Y(
        n11420) );
  sky130_fd_sc_hd__xnor2_1 U17111 ( .A(n17775), .B(n11421), .Y(n17874) );
  sky130_fd_sc_hd__xnor2_1 U17112 ( .A(n17776), .B(n17777), .Y(n11421) );
  sky130_fd_sc_hd__inv_1 U17113 ( .A(n12886), .Y(n18262) );
  sky130_fd_sc_hd__xnor3_1 U17114 ( .A(n18268), .B(n18267), .C(n18266), .X(
        n12886) );
  sky130_fd_sc_hd__nand4_1 U17115 ( .A(n16885), .B(n16882), .C(n16883), .D(
        n16884), .Y(n16886) );
  sky130_fd_sc_hd__inv_1 U17116 ( .A(n11422), .Y(n16572) );
  sky130_fd_sc_hd__nand3_1 U17117 ( .A(n12299), .B(n29479), .C(n29442), .Y(
        n11422) );
  sky130_fd_sc_hd__clkbuf_1 U17119 ( .A(n28130), .X(n11423) );
  sky130_fd_sc_hd__clkbuf_1 U17120 ( .A(n11610), .X(n11424) );
  sky130_fd_sc_hd__o21ai_1 U17121 ( .A1(n12417), .A2(n23421), .B1(n23947), .Y(
        n11719) );
  sky130_fd_sc_hd__nand2_1 U17122 ( .A(n11161), .B(n11425), .Y(n10537) );
  sky130_fd_sc_hd__nand2_1 U17123 ( .A(n24142), .B(n28417), .Y(n11425) );
  sky130_fd_sc_hd__buf_2 U17124 ( .A(n22007), .X(n29489) );
  sky130_fd_sc_hd__clkbuf_1 U17126 ( .A(n22959), .X(n11426) );
  sky130_fd_sc_hd__nor2_4 U17127 ( .A(n23448), .B(n11542), .Y(n28091) );
  sky130_fd_sc_hd__nand2_1 U17128 ( .A(n11428), .B(n11427), .Y(n17844) );
  sky130_fd_sc_hd__nand2_1 U17129 ( .A(n17814), .B(n17815), .Y(n11427) );
  sky130_fd_sc_hd__o21ai_1 U17130 ( .A1(n17815), .A2(n17814), .B1(n17813), .Y(
        n11428) );
  sky130_fd_sc_hd__nand2_1 U17131 ( .A(n11431), .B(n11430), .Y(n17857) );
  sky130_fd_sc_hd__nand2_1 U17132 ( .A(n17848), .B(n17849), .Y(n11430) );
  sky130_fd_sc_hd__nand2_1 U17133 ( .A(n17847), .B(n11432), .Y(n11431) );
  sky130_fd_sc_hd__nand2_1 U17134 ( .A(n11434), .B(n11433), .Y(n11432) );
  sky130_fd_sc_hd__xnor2_1 U17135 ( .A(n11435), .B(n17847), .Y(n17856) );
  sky130_fd_sc_hd__xnor2_1 U17136 ( .A(n17849), .B(n17848), .Y(n11435) );
  sky130_fd_sc_hd__fah_1 U17137 ( .A(n17600), .B(n17599), .CI(n17598), .COUT(
        n17627), .SUM(n17603) );
  sky130_fd_sc_hd__nand4_1 U17138 ( .A(n23619), .B(n12350), .C(n11437), .D(
        n23617), .Y(n11436) );
  sky130_fd_sc_hd__nand2_1 U17142 ( .A(n21316), .B(n11441), .Y(n11440) );
  sky130_fd_sc_hd__nor2b_1 U17143 ( .B_N(n21047), .A(n29482), .Y(n11441) );
  sky130_fd_sc_hd__nand3_2 U17144 ( .A(n11559), .B(n11621), .C(n12942), .Y(
        n11582) );
  sky130_fd_sc_hd__nand2_1 U17145 ( .A(n29512), .B(n12214), .Y(n24491) );
  sky130_fd_sc_hd__nand2_1 U17146 ( .A(n22737), .B(n22738), .Y(n29512) );
  sky130_fd_sc_hd__clkbuf_1 U17147 ( .A(n22799), .X(n11443) );
  sky130_fd_sc_hd__nand4_1 U17150 ( .A(n17319), .B(n17317), .C(n17318), .D(
        n17320), .Y(n11518) );
  sky130_fd_sc_hd__nor2_2 U17151 ( .A(n11445), .B(n11446), .Y(n24546) );
  sky130_fd_sc_hd__inv_1 U17152 ( .A(n11784), .Y(n11445) );
  sky130_fd_sc_hd__nor2_2 U17153 ( .A(n15196), .B(n15198), .Y(n21642) );
  sky130_fd_sc_hd__nand4_1 U17154 ( .A(n11447), .B(n21059), .C(n21057), .D(
        n21058), .Y(n21064) );
  sky130_fd_sc_hd__nand4_1 U17155 ( .A(n12192), .B(n12193), .C(n12191), .D(
        n11448), .Y(n12190) );
  sky130_fd_sc_hd__nand2_1 U17157 ( .A(j202_soc_core_memory0_ram_dout0[166]), 
        .B(n21487), .Y(n11447) );
  sky130_fd_sc_hd__nand2_1 U17158 ( .A(j202_soc_core_memory0_ram_dout0[404]), 
        .B(n21496), .Y(n11448) );
  sky130_fd_sc_hd__nand2_1 U17161 ( .A(n11450), .B(n11453), .Y(n12575) );
  sky130_fd_sc_hd__o21ai_1 U17162 ( .A1(n12430), .A2(n11451), .B1(n28089), .Y(
        n24616) );
  sky130_fd_sc_hd__nand2_1 U17163 ( .A(n23611), .B(n23383), .Y(n11452) );
  sky130_fd_sc_hd__nand3_2 U17165 ( .A(n12921), .B(n12920), .C(n20252), .Y(
        n12316) );
  sky130_fd_sc_hd__nand2_1 U17166 ( .A(n12511), .B(n20093), .Y(n12921) );
  sky130_fd_sc_hd__nor2_1 U17167 ( .A(n11939), .B(n11938), .Y(n11453) );
  sky130_fd_sc_hd__inv_1 U17168 ( .A(n11454), .Y(n11972) );
  sky130_fd_sc_hd__nand4_1 U17169 ( .A(n21061), .B(n21060), .C(n21063), .D(
        n21062), .Y(n11454) );
  sky130_fd_sc_hd__nand3_2 U17171 ( .A(n19263), .B(n27123), .C(n22266), .Y(
        n22437) );
  sky130_fd_sc_hd__o21ai_2 U17172 ( .A1(n18331), .A2(n19110), .B1(n18330), .Y(
        n18686) );
  sky130_fd_sc_hd__nand2_1 U17173 ( .A(n11457), .B(n11456), .Y(n18284) );
  sky130_fd_sc_hd__nand2_1 U17174 ( .A(n18267), .B(n18268), .Y(n11456) );
  sky130_fd_sc_hd__nand2_1 U17175 ( .A(n18266), .B(n11458), .Y(n11457) );
  sky130_fd_sc_hd__nand2b_1 U17176 ( .A_N(n18267), .B(n11459), .Y(n11458) );
  sky130_fd_sc_hd__clkbuf_1 U17177 ( .A(n27122), .X(n11460) );
  sky130_fd_sc_hd__xnor2_1 U17178 ( .A(n11465), .B(n18248), .Y(n18273) );
  sky130_fd_sc_hd__xnor2_1 U17179 ( .A(n18249), .B(n18250), .Y(n11465) );
  sky130_fd_sc_hd__nor2_4 U17180 ( .A(n27743), .B(n12524), .Y(n27728) );
  sky130_fd_sc_hd__nand2_1 U17181 ( .A(n26394), .B(n26393), .Y(n11466) );
  sky130_fd_sc_hd__nand2_1 U17182 ( .A(n11442), .B(n26395), .Y(n11467) );
  sky130_fd_sc_hd__xnor2_1 U17183 ( .A(n17910), .B(n11468), .Y(n18010) );
  sky130_fd_sc_hd__xnor2_1 U17184 ( .A(n17911), .B(n17912), .Y(n11468) );
  sky130_fd_sc_hd__fa_1 U17185 ( .A(n17920), .B(n17919), .CIN(n17918), .COUT(
        n17888), .SUM(n17970) );
  sky130_fd_sc_hd__nor2_2 U17187 ( .A(n13152), .B(n13153), .Y(n21495) );
  sky130_fd_sc_hd__nand2_1 U17189 ( .A(n11914), .B(n11917), .Y(n11913) );
  sky130_fd_sc_hd__nand2_1 U17191 ( .A(n28035), .B(n11689), .Y(n10539) );
  sky130_fd_sc_hd__nand4_1 U17193 ( .A(n24108), .B(n24631), .C(n28029), .D(
        n11470), .Y(n11469) );
  sky130_fd_sc_hd__inv_1 U17194 ( .A(n12338), .Y(n11470) );
  sky130_fd_sc_hd__clkbuf_1 U17195 ( .A(n22962), .X(n11471) );
  sky130_fd_sc_hd__nand2_1 U17196 ( .A(n11509), .B(n11101), .Y(n23574) );
  sky130_fd_sc_hd__nand2_1 U17197 ( .A(n11472), .B(n18880), .Y(n11529) );
  sky130_fd_sc_hd__clkbuf_1 U17200 ( .A(j202_soc_core_j22_cpu_ml_bufa[20]), 
        .X(n11474) );
  sky130_fd_sc_hd__inv_1 U17201 ( .A(n28038), .Y(n12063) );
  sky130_fd_sc_hd__nand2_1 U17202 ( .A(j202_soc_core_memory0_ram_dout0[75]), 
        .B(n21642), .Y(n11476) );
  sky130_fd_sc_hd__nor2_1 U17203 ( .A(n12659), .B(n12422), .Y(n12974) );
  sky130_fd_sc_hd__nand4_1 U17204 ( .A(n12660), .B(n12661), .C(n12662), .D(
        n12663), .Y(n12659) );
  sky130_fd_sc_hd__nor2_1 U17205 ( .A(n24453), .B(n23483), .Y(n11477) );
  sky130_fd_sc_hd__clkbuf_1 U17206 ( .A(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .X(n11478) );
  sky130_fd_sc_hd__nand2_1 U17208 ( .A(n11480), .B(n11479), .Y(n18289) );
  sky130_fd_sc_hd__nand2_1 U17209 ( .A(n18283), .B(n18282), .Y(n11479) );
  sky130_fd_sc_hd__nand2_1 U17210 ( .A(n18281), .B(n11481), .Y(n11480) );
  sky130_fd_sc_hd__nand2b_1 U17211 ( .A_N(n18283), .B(n11482), .Y(n11481) );
  sky130_fd_sc_hd__xnor2_1 U17212 ( .A(n18281), .B(n11483), .Y(n18287) );
  sky130_fd_sc_hd__xnor2_1 U17213 ( .A(n18282), .B(n18283), .Y(n11483) );
  sky130_fd_sc_hd__and2_0 U17214 ( .A(n22557), .B(n21255), .X(n11484) );
  sky130_fd_sc_hd__nand3_4 U17218 ( .A(n23505), .B(n12410), .C(n23514), .Y(
        n12351) );
  sky130_fd_sc_hd__nand2_1 U17219 ( .A(n25370), .B(n25642), .Y(n11485) );
  sky130_fd_sc_hd__nand4_1 U17220 ( .A(n12210), .B(n22116), .C(n22115), .D(
        n11191), .Y(n11486) );
  sky130_fd_sc_hd__a21o_1 U17221 ( .A1(n22147), .A2(n26426), .B1(n22146), .X(
        n12329) );
  sky130_fd_sc_hd__nor2_1 U17222 ( .A(n23948), .B(n23950), .Y(n11560) );
  sky130_fd_sc_hd__nand2_1 U17223 ( .A(n11497), .B(n11499), .Y(
        j202_soc_core_j22_cpu_rf_N3299) );
  sky130_fd_sc_hd__inv_2 U17224 ( .A(n11487), .Y(n24606) );
  sky130_fd_sc_hd__nor2_2 U17225 ( .A(n15192), .B(n15198), .Y(n21641) );
  sky130_fd_sc_hd__nand2_2 U17226 ( .A(j202_soc_core_memory0_ram_dout0[365]), 
        .B(n21495), .Y(n12801) );
  sky130_fd_sc_hd__nand2_2 U17227 ( .A(j202_soc_core_memory0_ram_dout0[429]), 
        .B(n12156), .Y(n12800) );
  sky130_fd_sc_hd__inv_2 U17229 ( .A(n11488), .Y(n23442) );
  sky130_fd_sc_hd__inv_2 U17230 ( .A(n23439), .Y(n11489) );
  sky130_fd_sc_hd__o22ai_1 U17231 ( .A1(n27859), .A2(n27586), .B1(n27858), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N3343) );
  sky130_fd_sc_hd__nand2_1 U17232 ( .A(n18334), .B(n22872), .Y(n21271) );
  sky130_fd_sc_hd__nand2_1 U17233 ( .A(n11490), .B(n28417), .Y(n24632) );
  sky130_fd_sc_hd__nand2_1 U17234 ( .A(n12053), .B(n24640), .Y(n11490) );
  sky130_fd_sc_hd__nand2_1 U17236 ( .A(n29500), .B(n11853), .Y(n24436) );
  sky130_fd_sc_hd__nand3_1 U17237 ( .A(n12408), .B(n22826), .C(n21255), .Y(
        n29500) );
  sky130_fd_sc_hd__o22ai_1 U17238 ( .A1(n27859), .A2(n25594), .B1(n27858), 
        .B2(n12267), .Y(j202_soc_core_j22_cpu_rf_N3333) );
  sky130_fd_sc_hd__nand2_1 U17239 ( .A(n11492), .B(n11491), .Y(n17839) );
  sky130_fd_sc_hd__nand2_1 U17240 ( .A(n17823), .B(n17824), .Y(n11491) );
  sky130_fd_sc_hd__o21ai_1 U17241 ( .A1(n17824), .A2(n17823), .B1(n17822), .Y(
        n11492) );
  sky130_fd_sc_hd__xnor3_1 U17242 ( .A(n11493), .B(n17823), .C(n17822), .X(
        n17812) );
  sky130_fd_sc_hd__nand2_1 U17243 ( .A(n23544), .B(n23545), .Y(n25561) );
  sky130_fd_sc_hd__clkbuf_1 U17244 ( .A(n23382), .X(n11494) );
  sky130_fd_sc_hd__nand3_2 U17245 ( .A(n13035), .B(n13036), .C(n13034), .Y(
        n12318) );
  sky130_fd_sc_hd__nand2_1 U17246 ( .A(n23396), .B(n12233), .Y(n23994) );
  sky130_fd_sc_hd__nand3_1 U17247 ( .A(n24968), .B(n27991), .C(n23557), .Y(
        n12233) );
  sky130_fd_sc_hd__inv_1 U17248 ( .A(n12273), .Y(n12282) );
  sky130_fd_sc_hd__nand4_1 U17250 ( .A(n20912), .B(n20913), .C(n20914), .D(
        n20904), .Y(n11916) );
  sky130_fd_sc_hd__nand3_2 U17253 ( .A(n20585), .B(n20584), .C(n20583), .Y(
        n23434) );
  sky130_fd_sc_hd__buf_6 U17254 ( .A(n23434), .X(n29593) );
  sky130_fd_sc_hd__nand2_2 U17255 ( .A(n26414), .B(n27828), .Y(n27355) );
  sky130_fd_sc_hd__nand4_1 U17256 ( .A(n12999), .B(n12998), .C(n12997), .D(
        n12996), .Y(n12995) );
  sky130_fd_sc_hd__inv_1 U17257 ( .A(n11742), .Y(n23504) );
  sky130_fd_sc_hd__inv_2 U17258 ( .A(n24503), .Y(n24504) );
  sky130_fd_sc_hd__nand3_2 U17259 ( .A(n18797), .B(n23514), .C(n23505), .Y(
        n12361) );
  sky130_fd_sc_hd__nand2b_1 U17261 ( .A_N(n27897), .B(n23749), .Y(n11497) );
  sky130_fd_sc_hd__nand2_1 U17262 ( .A(n12181), .B(n24832), .Y(n11499) );
  sky130_fd_sc_hd__nand2_1 U17263 ( .A(n28470), .B(n25397), .Y(n11500) );
  sky130_fd_sc_hd__nand4_1 U17264 ( .A(n12807), .B(n12808), .C(n12809), .D(
        n11501), .Y(n12806) );
  sky130_fd_sc_hd__nand2_1 U17265 ( .A(j202_soc_core_memory0_ram_dout0[370]), 
        .B(n21495), .Y(n11501) );
  sky130_fd_sc_hd__nand2_2 U17266 ( .A(n11634), .B(n12624), .Y(n12623) );
  sky130_fd_sc_hd__nand2_2 U17267 ( .A(n11502), .B(n27894), .Y(n10622) );
  sky130_fd_sc_hd__nor2_2 U17268 ( .A(n23611), .B(n12430), .Y(n27981) );
  sky130_fd_sc_hd__nand3_2 U17269 ( .A(n29595), .B(n29488), .C(n12599), .Y(
        n12598) );
  sky130_fd_sc_hd__nor2_2 U17271 ( .A(n30072), .B(n11177), .Y(n23439) );
  sky130_fd_sc_hd__nand2_1 U17272 ( .A(n23554), .B(n11547), .Y(n27737) );
  sky130_fd_sc_hd__nand2_1 U17273 ( .A(n11546), .B(n11545), .Y(n23554) );
  sky130_fd_sc_hd__nand4_1 U17274 ( .A(n12775), .B(n12774), .C(n12772), .D(
        n12773), .Y(n11783) );
  sky130_fd_sc_hd__nor2_2 U17275 ( .A(n11177), .B(n12230), .Y(n12781) );
  sky130_fd_sc_hd__nand2_1 U17276 ( .A(n11504), .B(n11503), .Y(n18009) );
  sky130_fd_sc_hd__nand2_1 U17277 ( .A(n18004), .B(n18003), .Y(n11503) );
  sky130_fd_sc_hd__nand2_1 U17278 ( .A(n18002), .B(n11505), .Y(n11504) );
  sky130_fd_sc_hd__nand2_1 U17279 ( .A(n11507), .B(n11506), .Y(n11505) );
  sky130_fd_sc_hd__xnor2_1 U17280 ( .A(n11508), .B(n18002), .Y(n18005) );
  sky130_fd_sc_hd__xnor2_1 U17281 ( .A(n18004), .B(n18003), .Y(n11508) );
  sky130_fd_sc_hd__inv_1 U17282 ( .A(n12847), .Y(n11514) );
  sky130_fd_sc_hd__a21boi_1 U17283 ( .A1(n23036), .A2(n21263), .B1_N(n21906), 
        .Y(n21264) );
  sky130_fd_sc_hd__nand2_1 U17284 ( .A(n24153), .B(n25679), .Y(n11509) );
  sky130_fd_sc_hd__nand2_2 U17286 ( .A(n25722), .B(n25310), .Y(n25313) );
  sky130_fd_sc_hd__nand2_4 U17287 ( .A(n11183), .B(n25291), .Y(n28525) );
  sky130_fd_sc_hd__nand2_1 U17288 ( .A(n11510), .B(n18578), .Y(n18617) );
  sky130_fd_sc_hd__nand2_1 U17289 ( .A(n18574), .B(n18575), .Y(n11510) );
  sky130_fd_sc_hd__xnor2_1 U17290 ( .A(n22598), .B(n11511), .Y(n24453) );
  sky130_fd_sc_hd__o21ai_1 U17291 ( .A1(n22597), .A2(n12349), .B1(n22596), .Y(
        n11511) );
  sky130_fd_sc_hd__nand3_2 U17292 ( .A(n25908), .B(n25907), .C(n25906), .Y(
        n27016) );
  sky130_fd_sc_hd__a21oi_2 U17293 ( .A1(n21964), .A2(n18658), .B1(n18657), .Y(
        n19106) );
  sky130_fd_sc_hd__nand2_1 U17294 ( .A(n11513), .B(n11512), .Y(n25309) );
  sky130_fd_sc_hd__o21a_1 U17295 ( .A1(n26285), .A2(n26939), .B1(n26919), .X(
        n11512) );
  sky130_fd_sc_hd__nand2_1 U17296 ( .A(n25765), .B(n26916), .Y(n11513) );
  sky130_fd_sc_hd__nor2_1 U17297 ( .A(n11515), .B(n11514), .Y(n11571) );
  sky130_fd_sc_hd__nand3_2 U17298 ( .A(n23505), .B(n12410), .C(n23514), .Y(
        n12279) );
  sky130_fd_sc_hd__o21ai_1 U17299 ( .A1(n12995), .A2(n12990), .B1(n20454), .Y(
        n11516) );
  sky130_fd_sc_hd__clkbuf_1 U17300 ( .A(n23397), .X(n11517) );
  sky130_fd_sc_hd__inv_2 U17301 ( .A(n28133), .Y(n28037) );
  sky130_fd_sc_hd__nand3b_1 U17303 ( .A_N(n11114), .B(n27786), .C(n26330), .Y(
        n25127) );
  sky130_fd_sc_hd__nand2_1 U17305 ( .A(n11519), .B(n28417), .Y(n24641) );
  sky130_fd_sc_hd__nand4_1 U17309 ( .A(n12522), .B(n21486), .C(n15375), .D(
        n12523), .Y(n12521) );
  sky130_fd_sc_hd__nand2_1 U17310 ( .A(n11522), .B(n27807), .Y(n24171) );
  sky130_fd_sc_hd__nand2_1 U17311 ( .A(n24157), .B(n11523), .Y(n11522) );
  sky130_fd_sc_hd__o21a_1 U17312 ( .A1(n28481), .A2(n26939), .B1(n26919), .X(
        n11523) );
  sky130_fd_sc_hd__nand3_2 U17313 ( .A(n11109), .B(n11525), .C(n11524), .Y(
        n26454) );
  sky130_fd_sc_hd__nand2_1 U17314 ( .A(n24172), .B(n24173), .Y(n11524) );
  sky130_fd_sc_hd__and2_1 U17315 ( .A(n24175), .B(n24174), .X(n11525) );
  sky130_fd_sc_hd__nand2_1 U17317 ( .A(n30073), .B(n11373), .Y(n24121) );
  sky130_fd_sc_hd__nand2_1 U17319 ( .A(n28081), .B(n11528), .Y(n10532) );
  sky130_fd_sc_hd__nand2_2 U17320 ( .A(n23507), .B(n23506), .Y(n23505) );
  sky130_fd_sc_hd__inv_1 U17321 ( .A(n30073), .Y(n28264) );
  sky130_fd_sc_hd__inv_1 U17323 ( .A(n11529), .Y(n22521) );
  sky130_fd_sc_hd__o21a_2 U17324 ( .A1(n29495), .A2(n12351), .B1(n30077), .X(
        n28442) );
  sky130_fd_sc_hd__a21boi_0 U17325 ( .A1(n27361), .A2(n12673), .B1_N(n26067), 
        .Y(n11530) );
  sky130_fd_sc_hd__inv_2 U17326 ( .A(n24471), .Y(n24472) );
  sky130_fd_sc_hd__nand2_2 U17327 ( .A(j202_soc_core_memory0_ram_dout0[461]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11531) );
  sky130_fd_sc_hd__nand3_2 U17328 ( .A(n11532), .B(n11182), .C(n11610), .Y(
        n24573) );
  sky130_fd_sc_hd__nand3_2 U17329 ( .A(n11532), .B(n29587), .C(n23549), .Y(
        n28378) );
  sky130_fd_sc_hd__inv_2 U17330 ( .A(n28378), .Y(n28411) );
  sky130_fd_sc_hd__clkbuf_1 U17331 ( .A(n12205), .X(n11533) );
  sky130_fd_sc_hd__inv_2 U17333 ( .A(n12336), .Y(n24405) );
  sky130_fd_sc_hd__nand3_2 U17334 ( .A(n11578), .B(n29489), .C(n11535), .Y(
        n12336) );
  sky130_fd_sc_hd__inv_2 U17335 ( .A(n12621), .Y(n11536) );
  sky130_fd_sc_hd__nand2_1 U17336 ( .A(n22231), .B(n22260), .Y(n11538) );
  sky130_fd_sc_hd__nand4_1 U17337 ( .A(n11540), .B(n11538), .C(n26916), .D(
        n11537), .Y(n22259) );
  sky130_fd_sc_hd__a21oi_2 U17340 ( .A1(n12575), .A2(n13082), .B1(n19862), .Y(
        n11607) );
  sky130_fd_sc_hd__inv_2 U17341 ( .A(n11542), .Y(n23614) );
  sky130_fd_sc_hd__nor2_2 U17342 ( .A(n12337), .B(n11542), .Y(n27885) );
  sky130_fd_sc_hd__nand2_2 U17343 ( .A(n11581), .B(n23955), .Y(n11542) );
  sky130_fd_sc_hd__nand2_2 U17344 ( .A(n12781), .B(n23557), .Y(n24695) );
  sky130_fd_sc_hd__nand2_1 U17345 ( .A(n12216), .B(n12218), .Y(n27729) );
  sky130_fd_sc_hd__nand2_1 U17346 ( .A(n27730), .B(n28261), .Y(n11544) );
  sky130_fd_sc_hd__inv_2 U17347 ( .A(n11141), .Y(n11545) );
  sky130_fd_sc_hd__nand2_1 U17348 ( .A(n23446), .B(n12620), .Y(n11547) );
  sky130_fd_sc_hd__nand2_1 U17349 ( .A(n11548), .B(n26941), .Y(n25932) );
  sky130_fd_sc_hd__o21ai_1 U17350 ( .A1(n11123), .A2(n28466), .B1(n26919), .Y(
        n11548) );
  sky130_fd_sc_hd__inv_1 U17351 ( .A(n12361), .Y(n11549) );
  sky130_fd_sc_hd__nand3_2 U17352 ( .A(n29489), .B(n11610), .C(n11551), .Y(
        n12395) );
  sky130_fd_sc_hd__inv_2 U17353 ( .A(n23549), .Y(n23550) );
  sky130_fd_sc_hd__nand3_1 U17354 ( .A(n11553), .B(n19086), .C(n23030), .Y(
        n12893) );
  sky130_fd_sc_hd__o211ai_1 U17355 ( .A1(n11565), .A2(n30080), .B1(n11564), 
        .C1(n11552), .Y(n24855) );
  sky130_fd_sc_hd__nand3_1 U17356 ( .A(n11553), .B(n11563), .C(n10972), .Y(
        n11552) );
  sky130_fd_sc_hd__inv_2 U17357 ( .A(n11554), .Y(n13024) );
  sky130_fd_sc_hd__nand2_1 U17358 ( .A(n11555), .B(n23494), .Y(n11554) );
  sky130_fd_sc_hd__nand3_1 U17359 ( .A(n23467), .B(n23468), .C(n23466), .Y(
        n11555) );
  sky130_fd_sc_hd__nand3_1 U17360 ( .A(n11555), .B(n23494), .C(n23563), .Y(
        n24360) );
  sky130_fd_sc_hd__nor2_2 U17361 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[0]), .B(n17359), .Y(n23493) );
  sky130_fd_sc_hd__nor2_4 U17363 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .B(n17356), .Y(n18679) );
  sky130_fd_sc_hd__nand2_2 U17364 ( .A(n12684), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[4]), .Y(n17356) );
  sky130_fd_sc_hd__nand2_1 U17365 ( .A(n11557), .B(n11556), .Y(n17773) );
  sky130_fd_sc_hd__nand2_1 U17366 ( .A(n17767), .B(n17768), .Y(n11556) );
  sky130_fd_sc_hd__o21ai_1 U17367 ( .A1(n17767), .A2(n17768), .B1(n17766), .Y(
        n11557) );
  sky130_fd_sc_hd__xnor2_1 U17368 ( .A(n17766), .B(n11558), .Y(n17871) );
  sky130_fd_sc_hd__xnor2_1 U17369 ( .A(n17768), .B(n17767), .Y(n11558) );
  sky130_fd_sc_hd__nand3_2 U17370 ( .A(n11559), .B(n11929), .C(n11740), .Y(
        n23438) );
  sky130_fd_sc_hd__inv_2 U17371 ( .A(n12989), .Y(n11559) );
  sky130_fd_sc_hd__nand4_1 U17372 ( .A(n11000), .B(n23409), .C(n24583), .D(
        n24547), .Y(n12924) );
  sky130_fd_sc_hd__buf_6 U17373 ( .A(n18224), .X(n11561) );
  sky130_fd_sc_hd__nand2_1 U17374 ( .A(n12167), .B(n28047), .Y(n17446) );
  sky130_fd_sc_hd__inv_2 U17375 ( .A(n11562), .Y(n18224) );
  sky130_fd_sc_hd__o22ai_1 U17376 ( .A1(n22365), .A2(n22655), .B1(n19281), 
        .B2(n11561), .Y(n18252) );
  sky130_fd_sc_hd__nand2_1 U17377 ( .A(n21682), .B(n21683), .Y(n11565) );
  sky130_fd_sc_hd__nand2_1 U17378 ( .A(n24855), .B(n24452), .Y(n22415) );
  sky130_fd_sc_hd__nand2_1 U17379 ( .A(n29498), .B(n11853), .Y(n24432) );
  sky130_fd_sc_hd__nand2_1 U17380 ( .A(n11443), .B(n11566), .Y(n29498) );
  sky130_fd_sc_hd__inv_2 U17381 ( .A(n28130), .Y(n12815) );
  sky130_fd_sc_hd__inv_2 U17382 ( .A(n11929), .Y(n11687) );
  sky130_fd_sc_hd__nand2_1 U17383 ( .A(n11646), .B(n11567), .Y(n23441) );
  sky130_fd_sc_hd__o21ai_1 U17384 ( .A1(n12778), .A2(n23440), .B1(n11568), .Y(
        n11567) );
  sky130_fd_sc_hd__nand2_1 U17385 ( .A(n11929), .B(n28130), .Y(n11568) );
  sky130_fd_sc_hd__inv_2 U17386 ( .A(n11569), .Y(n13090) );
  sky130_fd_sc_hd__nand4_1 U17388 ( .A(n11577), .B(n11576), .C(n11575), .D(
        n11574), .Y(n11685) );
  sky130_fd_sc_hd__nand2_1 U17389 ( .A(j202_soc_core_memory0_ram_dout0[463]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11574) );
  sky130_fd_sc_hd__nand2_1 U17390 ( .A(j202_soc_core_memory0_ram_dout0[15]), 
        .B(n21639), .Y(n11575) );
  sky130_fd_sc_hd__nand2_1 U17391 ( .A(j202_soc_core_memory0_ram_dout0[431]), 
        .B(n12156), .Y(n11576) );
  sky130_fd_sc_hd__nand2_1 U17392 ( .A(j202_soc_core_memory0_ram_dout0[399]), 
        .B(n21496), .Y(n11577) );
  sky130_fd_sc_hd__nor2_1 U17393 ( .A(n12362), .B(n12278), .Y(n11581) );
  sky130_fd_sc_hd__inv_1 U17394 ( .A(n11582), .Y(n23451) );
  sky130_fd_sc_hd__nand2_1 U17395 ( .A(n23407), .B(n11582), .Y(n23950) );
  sky130_fd_sc_hd__nand3_1 U17396 ( .A(n24690), .B(n11582), .C(n24691), .Y(
        n24693) );
  sky130_fd_sc_hd__nand4_1 U17397 ( .A(n20259), .B(n20266), .C(n20262), .D(
        n20261), .Y(n11590) );
  sky130_fd_sc_hd__nor2_1 U17398 ( .A(n11590), .B(n11598), .Y(n11586) );
  sky130_fd_sc_hd__nor2_1 U17399 ( .A(n11590), .B(n11589), .Y(n20417) );
  sky130_fd_sc_hd__nand2_2 U17400 ( .A(n11583), .B(n11587), .Y(n20425) );
  sky130_fd_sc_hd__inv_1 U17402 ( .A(n11589), .Y(n11584) );
  sky130_fd_sc_hd__nand2_1 U17404 ( .A(n20440), .B(n21919), .Y(n11588) );
  sky130_fd_sc_hd__nand2_1 U17406 ( .A(n11593), .B(n11592), .Y(n10528) );
  sky130_fd_sc_hd__and3_1 U17407 ( .A(n28074), .B(n28394), .C(n24698), .X(
        n11592) );
  sky130_fd_sc_hd__nand2_1 U17408 ( .A(n11594), .B(n28417), .Y(n11593) );
  sky130_fd_sc_hd__nand3_1 U17409 ( .A(n28115), .B(n24594), .C(n24695), .Y(
        n11594) );
  sky130_fd_sc_hd__nand3_2 U17410 ( .A(n11595), .B(n23387), .C(n12316), .Y(
        n11660) );
  sky130_fd_sc_hd__nand2_1 U17411 ( .A(n21002), .B(n12110), .Y(n12920) );
  sky130_fd_sc_hd__nand3_2 U17412 ( .A(n11831), .B(n11830), .C(n19854), .Y(
        n22007) );
  sky130_fd_sc_hd__inv_1 U17413 ( .A(n10982), .Y(n11595) );
  sky130_fd_sc_hd__nand2_1 U17414 ( .A(n11608), .B(n11607), .Y(n23447) );
  sky130_fd_sc_hd__nor2_1 U17415 ( .A(n11596), .B(n11650), .Y(n11649) );
  sky130_fd_sc_hd__inv_2 U17416 ( .A(n11605), .Y(n12350) );
  sky130_fd_sc_hd__nand3_2 U17417 ( .A(n23393), .B(n24568), .C(n11597), .Y(
        n11605) );
  sky130_fd_sc_hd__nand2_1 U17419 ( .A(n11600), .B(n11599), .Y(n11598) );
  sky130_fd_sc_hd__nand2_1 U17420 ( .A(j202_soc_core_memory0_ram_dout0[35]), 
        .B(n21633), .Y(n11599) );
  sky130_fd_sc_hd__nand2_1 U17421 ( .A(j202_soc_core_memory0_ram_dout0[99]), 
        .B(n21488), .Y(n11600) );
  sky130_fd_sc_hd__nand2_1 U17423 ( .A(j202_soc_core_memory0_ram_dout0[259]), 
        .B(n21634), .Y(n11602) );
  sky130_fd_sc_hd__nand2_1 U17424 ( .A(j202_soc_core_memory0_ram_dout0[291]), 
        .B(n21503), .Y(n11603) );
  sky130_fd_sc_hd__nand2_1 U17425 ( .A(n23410), .B(n27983), .Y(n11606) );
  sky130_fd_sc_hd__nand2_2 U17426 ( .A(n12282), .B(n11607), .Y(n12362) );
  sky130_fd_sc_hd__nand2_1 U17428 ( .A(n29593), .B(n11610), .Y(n23389) );
  sky130_fd_sc_hd__nand2_1 U17429 ( .A(n29489), .B(n11610), .Y(n23602) );
  sky130_fd_sc_hd__nand3_1 U17430 ( .A(n24550), .B(n28409), .C(n11610), .Y(
        n24614) );
  sky130_fd_sc_hd__nand2_1 U17431 ( .A(n28091), .B(n11424), .Y(n28093) );
  sky130_fd_sc_hd__o21a_1 U17432 ( .A1(n24115), .A2(n27885), .B1(n11424), .X(
        n24422) );
  sky130_fd_sc_hd__nand2_1 U17434 ( .A(n27744), .B(n12716), .Y(n11609) );
  sky130_fd_sc_hd__inv_1 U17435 ( .A(n11611), .Y(n11618) );
  sky130_fd_sc_hd__nand4_1 U17436 ( .A(n11615), .B(n11614), .C(n11613), .D(
        n11612), .Y(n11611) );
  sky130_fd_sc_hd__nand2_1 U17437 ( .A(j202_soc_core_memory0_ram_dout0[368]), 
        .B(n21495), .Y(n11612) );
  sky130_fd_sc_hd__nand2_1 U17438 ( .A(j202_soc_core_memory0_ram_dout0[272]), 
        .B(n21634), .Y(n11613) );
  sky130_fd_sc_hd__nand2_1 U17439 ( .A(j202_soc_core_memory0_ram_dout0[400]), 
        .B(n21496), .Y(n11614) );
  sky130_fd_sc_hd__nand2_1 U17440 ( .A(j202_soc_core_memory0_ram_dout0[432]), 
        .B(n12156), .Y(n11615) );
  sky130_fd_sc_hd__nand3_2 U17441 ( .A(n11618), .B(n19849), .C(n11616), .Y(
        n19850) );
  sky130_fd_sc_hd__inv_1 U17442 ( .A(n11617), .Y(n11616) );
  sky130_fd_sc_hd__nand2_1 U17443 ( .A(n11619), .B(n11620), .Y(n11617) );
  sky130_fd_sc_hd__nand2_1 U17444 ( .A(j202_soc_core_memory0_ram_dout0[336]), 
        .B(n21490), .Y(n11619) );
  sky130_fd_sc_hd__nand2_1 U17445 ( .A(j202_soc_core_memory0_ram_dout0[464]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11620) );
  sky130_fd_sc_hd__inv_2 U17447 ( .A(n23403), .Y(n11621) );
  sky130_fd_sc_hd__nand4_1 U17451 ( .A(n12731), .B(n12732), .C(n19117), .D(
        n19118), .Y(n11623) );
  sky130_fd_sc_hd__nand2_1 U17452 ( .A(n11628), .B(n11627), .Y(n11626) );
  sky130_fd_sc_hd__nand2_1 U17453 ( .A(j202_soc_core_memory0_ram_dout0[10]), 
        .B(n21639), .Y(n11627) );
  sky130_fd_sc_hd__nand2_1 U17454 ( .A(j202_soc_core_memory0_ram_dout0[298]), 
        .B(n21503), .Y(n11628) );
  sky130_fd_sc_hd__nand2_1 U17455 ( .A(n12806), .B(n21650), .Y(n12627) );
  sky130_fd_sc_hd__nand2_1 U17456 ( .A(n12810), .B(n21650), .Y(n12626) );
  sky130_fd_sc_hd__a21boi_2 U17457 ( .A1(n12803), .A2(n21020), .B1_N(n21022), 
        .Y(n12629) );
  sky130_fd_sc_hd__inv_1 U17458 ( .A(n11907), .Y(n11635) );
  sky130_fd_sc_hd__nor2_1 U17459 ( .A(n11636), .B(n23457), .Y(n24115) );
  sky130_fd_sc_hd__nor2b_1 U17460 ( .B_N(n21917), .A(n11642), .Y(n11637) );
  sky130_fd_sc_hd__nand2_1 U17462 ( .A(n21025), .B(n11639), .Y(n11638) );
  sky130_fd_sc_hd__nand2_1 U17464 ( .A(n21021), .B(n11097), .Y(n11641) );
  sky130_fd_sc_hd__buf_6 U17465 ( .A(n11174), .X(n11646) );
  sky130_fd_sc_hd__nand2_1 U17467 ( .A(n23405), .B(n22009), .Y(n12238) );
  sky130_fd_sc_hd__nor2_2 U17468 ( .A(n27899), .B(n12989), .Y(n11648) );
  sky130_fd_sc_hd__nand2_1 U17469 ( .A(n11648), .B(n23406), .Y(n23407) );
  sky130_fd_sc_hd__nand2_1 U17470 ( .A(n11648), .B(n27979), .Y(n23445) );
  sky130_fd_sc_hd__nand2_1 U17471 ( .A(n11647), .B(n11176), .Y(n24683) );
  sky130_fd_sc_hd__nand2_1 U17472 ( .A(n23380), .B(n28130), .Y(n24551) );
  sky130_fd_sc_hd__nand2_1 U17473 ( .A(n12248), .B(n24592), .Y(n24610) );
  sky130_fd_sc_hd__nand2_1 U17474 ( .A(n11836), .B(n30078), .Y(n12248) );
  sky130_fd_sc_hd__nand4_1 U17475 ( .A(n11654), .B(n11653), .C(n11652), .D(
        n11651), .Y(n11940) );
  sky130_fd_sc_hd__nand2_1 U17476 ( .A(j202_soc_core_memory0_ram_dout0[189]), 
        .B(n21487), .Y(n11651) );
  sky130_fd_sc_hd__nand2_1 U17477 ( .A(j202_soc_core_memory0_ram_dout0[125]), 
        .B(n21488), .Y(n11652) );
  sky130_fd_sc_hd__nand2_1 U17478 ( .A(j202_soc_core_memory0_ram_dout0[413]), 
        .B(n21496), .Y(n11653) );
  sky130_fd_sc_hd__nand2_1 U17479 ( .A(j202_soc_core_memory0_ram_dout0[477]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11654) );
  sky130_fd_sc_hd__o21a_1 U17480 ( .A1(n11659), .A2(n11912), .B1(n11655), .X(
        n23605) );
  sky130_fd_sc_hd__nor2_1 U17481 ( .A(n11657), .B(n22009), .Y(n11656) );
  sky130_fd_sc_hd__inv_2 U17482 ( .A(n11184), .Y(n11657) );
  sky130_fd_sc_hd__inv_2 U17483 ( .A(n29488), .Y(n11658) );
  sky130_fd_sc_hd__nand2_2 U17484 ( .A(n11140), .B(n12717), .Y(n11912) );
  sky130_fd_sc_hd__nor2_2 U17486 ( .A(n11657), .B(n29488), .Y(n24127) );
  sky130_fd_sc_hd__inv_2 U17487 ( .A(n11912), .Y(n12716) );
  sky130_fd_sc_hd__inv_2 U17488 ( .A(n12321), .Y(n12717) );
  sky130_fd_sc_hd__nor2_1 U17489 ( .A(n12233), .B(n11660), .Y(n28038) );
  sky130_fd_sc_hd__nor2_1 U17490 ( .A(n23396), .B(n11660), .Y(n12212) );
  sky130_fd_sc_hd__nand2_1 U17491 ( .A(n12345), .B(n11665), .Y(n28114) );
  sky130_fd_sc_hd__inv_1 U17492 ( .A(n24964), .Y(n11665) );
  sky130_fd_sc_hd__nor2_1 U17493 ( .A(n24421), .B(n24700), .Y(n27910) );
  sky130_fd_sc_hd__inv_1 U17494 ( .A(n24964), .Y(n24594) );
  sky130_fd_sc_hd__nand2_1 U17495 ( .A(n25149), .B(n25147), .Y(n12060) );
  sky130_fd_sc_hd__nand2_1 U17498 ( .A(n11970), .B(n11192), .Y(n11667) );
  sky130_fd_sc_hd__clkinv_1 U17499 ( .A(n11668), .Y(n11970) );
  sky130_fd_sc_hd__nand3_1 U17500 ( .A(n12657), .B(n11971), .C(n11972), .Y(
        n11668) );
  sky130_fd_sc_hd__nand2_1 U17502 ( .A(j202_soc_core_memory0_ram_dout0[227]), 
        .B(n21641), .Y(n11670) );
  sky130_fd_sc_hd__nand2_1 U17504 ( .A(n11672), .B(n12251), .Y(n28197) );
  sky130_fd_sc_hd__nor2_1 U17506 ( .A(n11679), .B(n11674), .Y(n11673) );
  sky130_fd_sc_hd__nand4_1 U17507 ( .A(n11678), .B(n11677), .C(n11676), .D(
        n11675), .Y(n11674) );
  sky130_fd_sc_hd__nand2_1 U17508 ( .A(j202_soc_core_memory0_ram_dout0[335]), 
        .B(n21490), .Y(n11675) );
  sky130_fd_sc_hd__nand2_1 U17509 ( .A(j202_soc_core_memory0_ram_dout0[303]), 
        .B(n21503), .Y(n11676) );
  sky130_fd_sc_hd__nand2_1 U17510 ( .A(j202_soc_core_memory0_ram_dout0[47]), 
        .B(n21633), .Y(n11677) );
  sky130_fd_sc_hd__nand2_1 U17511 ( .A(j202_soc_core_memory0_ram_dout0[367]), 
        .B(n21495), .Y(n11678) );
  sky130_fd_sc_hd__nand4_1 U17512 ( .A(n11683), .B(n11682), .C(n11681), .D(
        n11680), .Y(n11679) );
  sky130_fd_sc_hd__nand2_1 U17513 ( .A(j202_soc_core_memory0_ram_dout0[79]), 
        .B(n21642), .Y(n11680) );
  sky130_fd_sc_hd__nand2_1 U17514 ( .A(j202_soc_core_memory0_ram_dout0[143]), 
        .B(n21489), .Y(n11681) );
  sky130_fd_sc_hd__nand2_1 U17515 ( .A(j202_soc_core_memory0_ram_dout0[207]), 
        .B(n21640), .Y(n11682) );
  sky130_fd_sc_hd__nand2_1 U17516 ( .A(j202_soc_core_memory0_ram_dout0[239]), 
        .B(n21641), .Y(n11683) );
  sky130_fd_sc_hd__nand4_1 U17517 ( .A(n11721), .B(n11722), .C(n11723), .D(
        n12454), .Y(n11686) );
  sky130_fd_sc_hd__inv_2 U17518 ( .A(n12316), .Y(n23955) );
  sky130_fd_sc_hd__nand2b_1 U17519 ( .A_N(n11912), .B(n12154), .Y(n28259) );
  sky130_fd_sc_hd__nand2_2 U17520 ( .A(n11687), .B(n28130), .Y(n24097) );
  sky130_fd_sc_hd__nand3_1 U17521 ( .A(n28266), .B(n28267), .C(n11687), .Y(
        n28268) );
  sky130_fd_sc_hd__nand2_1 U17522 ( .A(n11689), .B(n11688), .Y(n10536) );
  sky130_fd_sc_hd__nand2_1 U17523 ( .A(n24137), .B(n28417), .Y(n11688) );
  sky130_fd_sc_hd__inv_2 U17524 ( .A(n12060), .Y(n11689) );
  sky130_fd_sc_hd__nand2_1 U17525 ( .A(n11701), .B(n11690), .Y(n21336) );
  sky130_fd_sc_hd__nand4_1 U17526 ( .A(n11695), .B(n11694), .C(n11693), .D(
        n11692), .Y(n11691) );
  sky130_fd_sc_hd__nand2_1 U17527 ( .A(j202_soc_core_memory0_ram_dout0[425]), 
        .B(n12156), .Y(n11692) );
  sky130_fd_sc_hd__nand2_1 U17528 ( .A(j202_soc_core_memory0_ram_dout0[361]), 
        .B(n21495), .Y(n11693) );
  sky130_fd_sc_hd__nand2_1 U17529 ( .A(j202_soc_core_memory0_ram_dout0[457]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11694) );
  sky130_fd_sc_hd__nand2_1 U17530 ( .A(j202_soc_core_memory0_ram_dout0[297]), 
        .B(n21503), .Y(n11695) );
  sky130_fd_sc_hd__nand4_1 U17531 ( .A(n11700), .B(n11699), .C(n11698), .D(
        n11697), .Y(n11696) );
  sky130_fd_sc_hd__nand2_1 U17532 ( .A(j202_soc_core_memory0_ram_dout0[9]), 
        .B(n21639), .Y(n11697) );
  sky130_fd_sc_hd__nand2_1 U17533 ( .A(j202_soc_core_memory0_ram_dout0[169]), 
        .B(n21487), .Y(n11698) );
  sky130_fd_sc_hd__nand2_1 U17534 ( .A(j202_soc_core_memory0_ram_dout0[41]), 
        .B(n21633), .Y(n11699) );
  sky130_fd_sc_hd__nand2_1 U17535 ( .A(j202_soc_core_memory0_ram_dout0[233]), 
        .B(n21641), .Y(n11700) );
  sky130_fd_sc_hd__nand4_1 U17536 ( .A(n20591), .B(n20590), .C(n20592), .D(
        n11703), .Y(n11702) );
  sky130_fd_sc_hd__nand2_1 U17537 ( .A(j202_soc_core_memory0_ram_dout0[393]), 
        .B(n21496), .Y(n11703) );
  sky130_fd_sc_hd__nand4_1 U17538 ( .A(n20698), .B(n20699), .C(n20589), .D(
        n20697), .Y(n11704) );
  sky130_fd_sc_hd__nand2_1 U17539 ( .A(n12212), .B(n28133), .Y(n11784) );
  sky130_fd_sc_hd__inv_2 U17541 ( .A(n24578), .Y(n11706) );
  sky130_fd_sc_hd__nand2_1 U17542 ( .A(n12001), .B(n29587), .Y(n24660) );
  sky130_fd_sc_hd__nand3_2 U17543 ( .A(n30048), .B(n30086), .C(n13034), .Y(
        n12317) );
  sky130_fd_sc_hd__nand3_2 U17544 ( .A(n19850), .B(n11712), .C(n21650), .Y(
        n13034) );
  sky130_fd_sc_hd__inv_1 U17546 ( .A(n11763), .Y(n11708) );
  sky130_fd_sc_hd__inv_2 U17548 ( .A(n11713), .Y(n11712) );
  sky130_fd_sc_hd__nand2_1 U17549 ( .A(j202_soc_core_memory0_ram_dout0[114]), 
        .B(n20460), .Y(n11718) );
  sky130_fd_sc_hd__nand2_1 U17550 ( .A(n12628), .B(n20258), .Y(n11907) );
  sky130_fd_sc_hd__nand2_1 U17551 ( .A(n11714), .B(n21020), .Y(n12628) );
  sky130_fd_sc_hd__nand4_1 U17552 ( .A(n11717), .B(n11718), .C(n11715), .D(
        n11716), .Y(n11714) );
  sky130_fd_sc_hd__nand2_1 U17553 ( .A(j202_soc_core_memory0_ram_dout0[210]), 
        .B(n20455), .Y(n11715) );
  sky130_fd_sc_hd__nand2_1 U17554 ( .A(j202_soc_core_memory0_ram_dout0[242]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[7]), .Y(n11716) );
  sky130_fd_sc_hd__nand2_1 U17555 ( .A(j202_soc_core_memory0_ram_dout0[146]), 
        .B(n20456), .Y(n11717) );
  sky130_fd_sc_hd__nand4_1 U17557 ( .A(n12717), .B(n11140), .C(n23426), .D(
        n24593), .Y(n23429) );
  sky130_fd_sc_hd__nand3_1 U17558 ( .A(n11910), .B(n10981), .C(n23392), .Y(
        n28386) );
  sky130_fd_sc_hd__nand2_1 U17559 ( .A(n28386), .B(n11733), .Y(n28419) );
  sky130_fd_sc_hd__nand2_1 U17560 ( .A(j202_soc_core_memory0_ram_dout0[111]), 
        .B(n21488), .Y(n11721) );
  sky130_fd_sc_hd__nand2_1 U17561 ( .A(j202_soc_core_memory0_ram_dout0[175]), 
        .B(n21487), .Y(n11722) );
  sky130_fd_sc_hd__nand2_1 U17562 ( .A(j202_soc_core_memory0_ram_dout0[271]), 
        .B(n21634), .Y(n11723) );
  sky130_fd_sc_hd__nand3_1 U17564 ( .A(n11725), .B(n28356), .C(n28357), .Y(
        j202_soc_core_j22_cpu_id_idec_N937) );
  sky130_fd_sc_hd__clkbuf_2 U17567 ( .A(n27901), .X(n11729) );
  sky130_fd_sc_hd__nand2_1 U17568 ( .A(n11729), .B(n12844), .Y(n28415) );
  sky130_fd_sc_hd__nand2_1 U17569 ( .A(n11729), .B(n12326), .Y(n28262) );
  sky130_fd_sc_hd__nand2b_1 U17570 ( .A_N(n12844), .B(n11178), .Y(n11731) );
  sky130_fd_sc_hd__inv_2 U17571 ( .A(n11732), .Y(n23393) );
  sky130_fd_sc_hd__inv_2 U17572 ( .A(n28419), .Y(n24568) );
  sky130_fd_sc_hd__nand2_1 U17573 ( .A(n27901), .B(n24634), .Y(n11733) );
  sky130_fd_sc_hd__nand4_1 U17574 ( .A(n11735), .B(n27730), .C(n28387), .D(
        n28148), .Y(n24402) );
  sky130_fd_sc_hd__inv_2 U17577 ( .A(n12424), .Y(n28266) );
  sky130_fd_sc_hd__nor2_1 U17578 ( .A(n28264), .B(n24621), .Y(n27983) );
  sky130_fd_sc_hd__nand2_1 U17579 ( .A(n24684), .B(n27730), .Y(n24621) );
  sky130_fd_sc_hd__nand2_1 U17580 ( .A(j202_soc_core_memory0_ram_dout0[301]), 
        .B(n21503), .Y(n11736) );
  sky130_fd_sc_hd__nand2_1 U17581 ( .A(j202_soc_core_memory0_ram_dout0[269]), 
        .B(n21634), .Y(n11737) );
  sky130_fd_sc_hd__nand2_1 U17582 ( .A(j202_soc_core_memory0_ram_dout0[397]), 
        .B(n21496), .Y(n11738) );
  sky130_fd_sc_hd__inv_2 U17584 ( .A(n23610), .Y(n27901) );
  sky130_fd_sc_hd__nand3_2 U17585 ( .A(n23614), .B(n23436), .C(n23448), .Y(
        n23437) );
  sky130_fd_sc_hd__o21ai_1 U17586 ( .A1(n29560), .A2(n12417), .B1(n24563), .Y(
        n11740) );
  sky130_fd_sc_hd__nand2_1 U17587 ( .A(n12212), .B(n28027), .Y(n11741) );
  sky130_fd_sc_hd__nor2_2 U17588 ( .A(n23403), .B(n12524), .Y(n28027) );
  sky130_fd_sc_hd__nand2_1 U17589 ( .A(n23396), .B(n23397), .Y(n12232) );
  sky130_fd_sc_hd__nand2_1 U17590 ( .A(n11750), .B(n11749), .Y(n11742) );
  sky130_fd_sc_hd__nand3_2 U17591 ( .A(n11747), .B(n11750), .C(n11743), .Y(
        n12410) );
  sky130_fd_sc_hd__inv_2 U17592 ( .A(n11744), .Y(n11743) );
  sky130_fd_sc_hd__nand2_1 U17593 ( .A(n11749), .B(n11745), .Y(n11744) );
  sky130_fd_sc_hd__o21a_1 U17594 ( .A1(n23511), .A2(n19852), .B1(n23510), .X(
        n11745) );
  sky130_fd_sc_hd__nand2_1 U17595 ( .A(n11748), .B(
        j202_soc_core_j22_cpu_ma_M_address[1]), .Y(n11747) );
  sky130_fd_sc_hd__nand2_1 U17597 ( .A(n23508), .B(
        j202_soc_core_j22_cpu_ma_M_address[1]), .Y(n23503) );
  sky130_fd_sc_hd__nand2_1 U17598 ( .A(n19853), .B(n19852), .Y(n23508) );
  sky130_fd_sc_hd__nand4_1 U17599 ( .A(n11012), .B(n11887), .C(n11886), .D(
        n23511), .Y(n11750) );
  sky130_fd_sc_hd__nand3_2 U17600 ( .A(n11773), .B(n11751), .C(n11772), .Y(
        n24861) );
  sky130_fd_sc_hd__and3b_1 U17601 ( .B(n24857), .C(n24856), .A_N(n11752), .X(
        n11751) );
  sky130_fd_sc_hd__o21ai_1 U17602 ( .A1(n25658), .A2(n24851), .B1(n24850), .Y(
        n11752) );
  sky130_fd_sc_hd__nand2_1 U17603 ( .A(n19850), .B(n21650), .Y(n20975) );
  sky130_fd_sc_hd__nand4_1 U17604 ( .A(n11757), .B(n11756), .C(n11755), .D(
        n11754), .Y(n11753) );
  sky130_fd_sc_hd__nand2_1 U17605 ( .A(j202_soc_core_memory0_ram_dout0[0]), 
        .B(n21639), .Y(n11754) );
  sky130_fd_sc_hd__nand2_1 U17606 ( .A(j202_soc_core_memory0_ram_dout0[288]), 
        .B(n21503), .Y(n11755) );
  sky130_fd_sc_hd__nand2_1 U17607 ( .A(j202_soc_core_memory0_ram_dout0[160]), 
        .B(n21487), .Y(n11756) );
  sky130_fd_sc_hd__nand2_1 U17608 ( .A(j202_soc_core_memory0_ram_dout0[192]), 
        .B(n21640), .Y(n11757) );
  sky130_fd_sc_hd__nand4_1 U17609 ( .A(n12960), .B(n11761), .C(n11760), .D(
        n11759), .Y(n11758) );
  sky130_fd_sc_hd__nand2_1 U17610 ( .A(j202_soc_core_memory0_ram_dout0[96]), 
        .B(n21488), .Y(n11759) );
  sky130_fd_sc_hd__nand2_1 U17611 ( .A(j202_soc_core_memory0_ram_dout0[128]), 
        .B(n21489), .Y(n11760) );
  sky130_fd_sc_hd__nand2_1 U17612 ( .A(j202_soc_core_memory0_ram_dout0[64]), 
        .B(n21642), .Y(n11761) );
  sky130_fd_sc_hd__nand4_1 U17613 ( .A(n12963), .B(n12957), .C(n12958), .D(
        n12959), .Y(n11762) );
  sky130_fd_sc_hd__nand4_1 U17614 ( .A(n12956), .B(n12961), .C(n12962), .D(
        n12122), .Y(n11763) );
  sky130_fd_sc_hd__o211ai_2 U17615 ( .A1(n11771), .A2(n11770), .B1(n22266), 
        .C1(n11764), .Y(n22799) );
  sky130_fd_sc_hd__nand3_1 U17616 ( .A(n11765), .B(n21728), .C(n11766), .Y(
        n11764) );
  sky130_fd_sc_hd__nand3_2 U17617 ( .A(n11765), .B(n21728), .C(n11769), .Y(
        n11770) );
  sky130_fd_sc_hd__inv_1 U17618 ( .A(n12026), .Y(n11768) );
  sky130_fd_sc_hd__and2_0 U17619 ( .A(n11769), .B(n27355), .X(n11766) );
  sky130_fd_sc_hd__o21a_1 U17620 ( .A1(n26919), .A2(n11188), .B1(n21727), .X(
        n11769) );
  sky130_fd_sc_hd__nand2_1 U17621 ( .A(n22416), .B(n22415), .Y(n11771) );
  sky130_fd_sc_hd__nand2_1 U17622 ( .A(n24859), .B(n24849), .Y(n11772) );
  sky130_fd_sc_hd__nand2_1 U17624 ( .A(n11774), .B(n27111), .Y(n11773) );
  sky130_fd_sc_hd__nand2_1 U17625 ( .A(n11776), .B(n11775), .Y(n11774) );
  sky130_fd_sc_hd__nand2_1 U17626 ( .A(n28537), .B(n26916), .Y(n11776) );
  sky130_fd_sc_hd__nand2_1 U17627 ( .A(n17828), .B(n11777), .Y(n18684) );
  sky130_fd_sc_hd__nand2_1 U17628 ( .A(n11008), .B(n21650), .Y(n21024) );
  sky130_fd_sc_hd__inv_1 U17629 ( .A(n11779), .Y(n11778) );
  sky130_fd_sc_hd__nand2_1 U17630 ( .A(n12008), .B(n12009), .Y(n11779) );
  sky130_fd_sc_hd__inv_1 U17631 ( .A(n11781), .Y(n11780) );
  sky130_fd_sc_hd__nand2_1 U17632 ( .A(n12006), .B(n12007), .Y(n11781) );
  sky130_fd_sc_hd__inv_1 U17633 ( .A(n11783), .Y(n11782) );
  sky130_fd_sc_hd__nand2b_1 U17634 ( .A_N(n24637), .B(n11784), .Y(n24623) );
  sky130_fd_sc_hd__inv_1 U17635 ( .A(n11785), .Y(n12657) );
  sky130_fd_sc_hd__nand4_1 U17636 ( .A(n11789), .B(n11788), .C(n11787), .D(
        n11786), .Y(n11785) );
  sky130_fd_sc_hd__and2_0 U17637 ( .A(n21169), .B(n21161), .X(n11786) );
  sky130_fd_sc_hd__nand2_1 U17638 ( .A(j202_soc_core_memory0_ram_dout0[454]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11787) );
  sky130_fd_sc_hd__nand2_1 U17639 ( .A(j202_soc_core_memory0_ram_dout0[422]), 
        .B(n12156), .Y(n11788) );
  sky130_fd_sc_hd__nand2_1 U17640 ( .A(j202_soc_core_memory0_ram_dout0[358]), 
        .B(n21495), .Y(n11789) );
  sky130_fd_sc_hd__inv_2 U17641 ( .A(n11790), .Y(n22949) );
  sky130_fd_sc_hd__nand2_1 U17642 ( .A(n22868), .B(n22867), .Y(n11790) );
  sky130_fd_sc_hd__nand3_2 U17643 ( .A(n24789), .B(n22266), .C(n24790), .Y(
        n22868) );
  sky130_fd_sc_hd__nand2_1 U17644 ( .A(n21980), .B(n27355), .Y(n24789) );
  sky130_fd_sc_hd__nand2_1 U17646 ( .A(j202_soc_core_memory0_ram_dout0[219]), 
        .B(n21640), .Y(n11791) );
  sky130_fd_sc_hd__nand2_1 U17647 ( .A(j202_soc_core_memory0_ram_dout0[123]), 
        .B(n21488), .Y(n11792) );
  sky130_fd_sc_hd__nand2_1 U17648 ( .A(j202_soc_core_memory0_ram_dout0[379]), 
        .B(n21495), .Y(n11793) );
  sky130_fd_sc_hd__inv_2 U17649 ( .A(n11794), .Y(n23557) );
  sky130_fd_sc_hd__inv_2 U17651 ( .A(n10994), .Y(n24968) );
  sky130_fd_sc_hd__a22oi_2 U17653 ( .A1(n12495), .A2(n11795), .B1(n25349), 
        .B2(n22230), .Y(n12210) );
  sky130_fd_sc_hd__nand2_1 U17654 ( .A(n11796), .B(n22739), .Y(n21334) );
  sky130_fd_sc_hd__nand4_1 U17657 ( .A(n11802), .B(n11801), .C(n11800), .D(
        n11799), .Y(n11798) );
  sky130_fd_sc_hd__nand2_1 U17658 ( .A(j202_soc_core_memory0_ram_dout0[2]), 
        .B(n21639), .Y(n11799) );
  sky130_fd_sc_hd__nand2_1 U17659 ( .A(j202_soc_core_memory0_ram_dout0[194]), 
        .B(n21640), .Y(n11800) );
  sky130_fd_sc_hd__nand2_1 U17660 ( .A(j202_soc_core_memory0_ram_dout0[290]), 
        .B(n21503), .Y(n11801) );
  sky130_fd_sc_hd__nand2_1 U17661 ( .A(j202_soc_core_memory0_ram_dout0[34]), 
        .B(n21633), .Y(n11802) );
  sky130_fd_sc_hd__nand4_1 U17662 ( .A(n12664), .B(n11806), .C(n11805), .D(
        n11804), .Y(n11803) );
  sky130_fd_sc_hd__nand2_1 U17663 ( .A(j202_soc_core_memory0_ram_dout0[450]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11804) );
  sky130_fd_sc_hd__nand2_1 U17664 ( .A(j202_soc_core_memory0_ram_dout0[418]), 
        .B(n12156), .Y(n11805) );
  sky130_fd_sc_hd__nand2_1 U17665 ( .A(j202_soc_core_memory0_ram_dout0[386]), 
        .B(n21496), .Y(n11806) );
  sky130_fd_sc_hd__nor2_1 U17666 ( .A(n11809), .B(n11808), .Y(n11807) );
  sky130_fd_sc_hd__nand4_1 U17667 ( .A(n12750), .B(n12744), .C(n12745), .D(
        n12746), .Y(n11808) );
  sky130_fd_sc_hd__nand4_1 U17668 ( .A(n12747), .B(n12748), .C(n12749), .D(
        n12743), .Y(n11809) );
  sky130_fd_sc_hd__nand3_1 U17670 ( .A(n22688), .B(n22687), .C(n22686), .Y(
        n29514) );
  sky130_fd_sc_hd__nand2_1 U17671 ( .A(n30059), .B(n11205), .Y(n11825) );
  sky130_fd_sc_hd__nand2_1 U17672 ( .A(n11102), .B(n22232), .Y(n11823) );
  sky130_fd_sc_hd__a22oi_1 U17673 ( .A1(n30059), .A2(n11814), .B1(n11102), 
        .B2(n11812), .Y(n11811) );
  sky130_fd_sc_hd__nor2_1 U17674 ( .A(n25397), .B(n12557), .Y(n11812) );
  sky130_fd_sc_hd__nor2_1 U17675 ( .A(n25397), .B(n22229), .Y(n11814) );
  sky130_fd_sc_hd__nand3_1 U17676 ( .A(n11817), .B(n11829), .C(n11827), .Y(
        n11815) );
  sky130_fd_sc_hd__nand2_1 U17677 ( .A(n11185), .B(n22114), .Y(n11827) );
  sky130_fd_sc_hd__nand2_1 U17678 ( .A(n12023), .B(n22230), .Y(n11829) );
  sky130_fd_sc_hd__and2_0 U17679 ( .A(n11824), .B(n27786), .X(n11818) );
  sky130_fd_sc_hd__o21ai_0 U17680 ( .A1(n11824), .A2(n25397), .B1(n21935), .Y(
        n11821) );
  sky130_fd_sc_hd__nor2_1 U17681 ( .A(n25397), .B(n11149), .Y(n11822) );
  sky130_fd_sc_hd__nand2_1 U17682 ( .A(n22009), .B(n12278), .Y(n11911) );
  sky130_fd_sc_hd__nand2_1 U17683 ( .A(n19853), .B(n13083), .Y(n11830) );
  sky130_fd_sc_hd__nand2_1 U17684 ( .A(n12770), .B(n12124), .Y(n11831) );
  sky130_fd_sc_hd__nand3_1 U17685 ( .A(n12921), .B(n12920), .C(n20252), .Y(
        n23388) );
  sky130_fd_sc_hd__nand4_1 U17686 ( .A(n11835), .B(n11834), .C(n11833), .D(
        n11832), .Y(n11855) );
  sky130_fd_sc_hd__nand2_1 U17687 ( .A(j202_soc_core_memory0_ram_dout0[127]), 
        .B(n21488), .Y(n11832) );
  sky130_fd_sc_hd__nand2_1 U17688 ( .A(j202_soc_core_memory0_ram_dout0[31]), 
        .B(n21639), .Y(n11833) );
  sky130_fd_sc_hd__nand2_1 U17689 ( .A(j202_soc_core_memory0_ram_dout0[191]), 
        .B(n21487), .Y(n11834) );
  sky130_fd_sc_hd__nand2_1 U17690 ( .A(j202_soc_core_memory0_ram_dout0[351]), 
        .B(n21490), .Y(n11835) );
  sky130_fd_sc_hd__nor2_1 U17691 ( .A(n11837), .B(n23598), .Y(n23599) );
  sky130_fd_sc_hd__nand2_1 U17692 ( .A(n11839), .B(n11173), .Y(n11837) );
  sky130_fd_sc_hd__a21oi_1 U17693 ( .A1(n28134), .A2(n12716), .B1(n11838), .Y(
        n28136) );
  sky130_fd_sc_hd__inv_1 U17694 ( .A(n11839), .Y(n11838) );
  sky130_fd_sc_hd__nand2_1 U17695 ( .A(n12716), .B(n11840), .Y(n11839) );
  sky130_fd_sc_hd__nand2_1 U17696 ( .A(n11841), .B(n11179), .Y(n11840) );
  sky130_fd_sc_hd__nand3_1 U17697 ( .A(n11139), .B(n26162), .C(n11123), .Y(
        n11842) );
  sky130_fd_sc_hd__nand2_1 U17698 ( .A(n25941), .B(n25397), .Y(n11843) );
  sky130_fd_sc_hd__nand2_1 U17699 ( .A(n11844), .B(n25994), .Y(n25995) );
  sky130_fd_sc_hd__nand2_1 U17700 ( .A(n11846), .B(n11845), .Y(n21230) );
  sky130_fd_sc_hd__nand3_1 U17701 ( .A(n12184), .B(n26334), .C(n27785), .Y(
        n11845) );
  sky130_fd_sc_hd__nand3_1 U17702 ( .A(n11847), .B(n26376), .C(n26916), .Y(
        n11846) );
  sky130_fd_sc_hd__nand2_1 U17703 ( .A(n12184), .B(n26334), .Y(n26376) );
  sky130_fd_sc_hd__nand4_1 U17704 ( .A(n11851), .B(n11849), .C(n11850), .D(
        n11190), .Y(n11847) );
  sky130_fd_sc_hd__inv_2 U17706 ( .A(n26165), .Y(n11852) );
  sky130_fd_sc_hd__buf_6 U17707 ( .A(n11138), .X(n11853) );
  sky130_fd_sc_hd__clkbuf_1 U17708 ( .A(n21187), .X(n11854) );
  sky130_fd_sc_hd__nand2_1 U17709 ( .A(n29520), .B(n12214), .Y(n24503) );
  sky130_fd_sc_hd__inv_1 U17710 ( .A(j202_soc_core_j22_cpu_ml_bufa[9]), .Y(
        n12049) );
  sky130_fd_sc_hd__nand2_1 U17711 ( .A(n21195), .B(n11856), .Y(n19108) );
  sky130_fd_sc_hd__nand2_1 U17712 ( .A(n18660), .B(n18659), .Y(n11856) );
  sky130_fd_sc_hd__nand2_1 U17713 ( .A(n17906), .B(n17905), .Y(n17947) );
  sky130_fd_sc_hd__nand2_1 U17714 ( .A(n11858), .B(n11857), .Y(n18239) );
  sky130_fd_sc_hd__nand2_1 U17715 ( .A(n18235), .B(n11860), .Y(n11857) );
  sky130_fd_sc_hd__xnor2_1 U17717 ( .A(n18234), .B(n11859), .Y(n18243) );
  sky130_fd_sc_hd__xnor2_1 U17718 ( .A(n18235), .B(n11860), .Y(n11859) );
  sky130_fd_sc_hd__nand2_1 U17719 ( .A(n12214), .B(n29506), .Y(n24479) );
  sky130_fd_sc_hd__nand3_1 U17720 ( .A(n11862), .B(n22826), .C(n11861), .Y(
        n29506) );
  sky130_fd_sc_hd__nand2_1 U17721 ( .A(n11864), .B(n11863), .Y(n11862) );
  sky130_fd_sc_hd__a21boi_0 U17722 ( .A1(n25677), .A2(n27052), .B1_N(n27717), 
        .Y(n11863) );
  sky130_fd_sc_hd__nand2_1 U17723 ( .A(n25718), .B(n27828), .Y(n11864) );
  sky130_fd_sc_hd__o21ai_1 U17724 ( .A1(n22516), .A2(n11866), .B1(n22515), .Y(
        n22517) );
  sky130_fd_sc_hd__xor2_1 U17725 ( .A(n22565), .B(n11866), .X(n24458) );
  sky130_fd_sc_hd__o21ai_1 U17726 ( .A1(n11866), .A2(n22934), .B1(n22933), .Y(
        n22935) );
  sky130_fd_sc_hd__o21ai_1 U17728 ( .A1(n11866), .A2(n22609), .B1(n22608), .Y(
        n22610) );
  sky130_fd_sc_hd__o21ai_1 U17729 ( .A1(n11866), .A2(n22342), .B1(n22341), .Y(
        n22343) );
  sky130_fd_sc_hd__nand2_1 U17730 ( .A(n23037), .B(n11867), .Y(n23038) );
  sky130_fd_sc_hd__nand2_1 U17731 ( .A(n11099), .B(n11171), .Y(n11867) );
  sky130_fd_sc_hd__o21ai_1 U17732 ( .A1(n11866), .A2(n22182), .B1(n22181), .Y(
        n22183) );
  sky130_fd_sc_hd__nand2_1 U17733 ( .A(n11869), .B(n11868), .Y(n17946) );
  sky130_fd_sc_hd__nand2_1 U17734 ( .A(n17997), .B(n17998), .Y(n11868) );
  sky130_fd_sc_hd__nand2_1 U17735 ( .A(n17996), .B(n11870), .Y(n11869) );
  sky130_fd_sc_hd__inv_1 U17736 ( .A(n11871), .Y(n11870) );
  sky130_fd_sc_hd__nor2_1 U17737 ( .A(n17998), .B(n17997), .Y(n11871) );
  sky130_fd_sc_hd__xnor2_1 U17738 ( .A(n11872), .B(n17996), .Y(n18007) );
  sky130_fd_sc_hd__xnor2_1 U17739 ( .A(n17997), .B(n17998), .Y(n11872) );
  sky130_fd_sc_hd__nand2_1 U17740 ( .A(n18468), .B(n11876), .Y(n12506) );
  sky130_fd_sc_hd__nand2_1 U17741 ( .A(n11873), .B(n18467), .Y(n12507) );
  sky130_fd_sc_hd__nand2b_1 U17742 ( .A_N(n18468), .B(n11874), .Y(n11873) );
  sky130_fd_sc_hd__nand2_1 U17745 ( .A(n11878), .B(n11877), .Y(n18056) );
  sky130_fd_sc_hd__nand2_1 U17746 ( .A(n18045), .B(n18046), .Y(n11877) );
  sky130_fd_sc_hd__o21ai_1 U17747 ( .A1(n18046), .A2(n18045), .B1(n18044), .Y(
        n11878) );
  sky130_fd_sc_hd__xnor2_1 U17748 ( .A(n18045), .B(n11879), .Y(n18060) );
  sky130_fd_sc_hd__xnor2_1 U17749 ( .A(n18046), .B(n18044), .Y(n11879) );
  sky130_fd_sc_hd__nand2_1 U17750 ( .A(n11881), .B(n11880), .Y(n18562) );
  sky130_fd_sc_hd__nand2_1 U17751 ( .A(n18557), .B(n18556), .Y(n11880) );
  sky130_fd_sc_hd__xnor2_1 U17753 ( .A(n18555), .B(n11882), .Y(n18629) );
  sky130_fd_sc_hd__xnor2_1 U17754 ( .A(n18557), .B(n18556), .Y(n11882) );
  sky130_fd_sc_hd__nand2_1 U17755 ( .A(n12673), .B(n25679), .Y(n26448) );
  sky130_fd_sc_hd__nor2_1 U17756 ( .A(n11885), .B(n11883), .Y(n11891) );
  sky130_fd_sc_hd__nand2_1 U17758 ( .A(j202_soc_core_memory0_ram_dout0[287]), 
        .B(n21634), .Y(n11884) );
  sky130_fd_sc_hd__nand4_1 U17759 ( .A(n12581), .B(n12576), .C(n16385), .D(
        n12577), .Y(n11885) );
  sky130_fd_sc_hd__inv_1 U17760 ( .A(n11888), .Y(n11887) );
  sky130_fd_sc_hd__nand3_1 U17761 ( .A(n16386), .B(n11890), .C(n11889), .Y(
        n11888) );
  sky130_fd_sc_hd__nand2_1 U17762 ( .A(j202_soc_core_memory0_ram_dout0[383]), 
        .B(n21495), .Y(n11889) );
  sky130_fd_sc_hd__nand2_1 U17763 ( .A(j202_soc_core_memory0_ram_dout0[415]), 
        .B(n21496), .Y(n11890) );
  sky130_fd_sc_hd__nand3_1 U17764 ( .A(n11892), .B(n30021), .C(n28034), .Y(
        n11894) );
  sky130_fd_sc_hd__nand2_1 U17765 ( .A(n11923), .B(n11922), .Y(n11892) );
  sky130_fd_sc_hd__nand2_1 U17766 ( .A(n24123), .B(n11906), .Y(n11923) );
  sky130_fd_sc_hd__nor2_1 U17767 ( .A(n11895), .B(n11894), .Y(n28035) );
  sky130_fd_sc_hd__nand2_1 U17768 ( .A(n28083), .B(n11896), .Y(n11895) );
  sky130_fd_sc_hd__nand2_1 U17769 ( .A(n28152), .B(n28417), .Y(n11896) );
  sky130_fd_sc_hd__nand2_1 U17770 ( .A(n24125), .B(n11705), .Y(n28033) );
  sky130_fd_sc_hd__nor2_1 U17773 ( .A(n28032), .B(n11901), .Y(n11900) );
  sky130_fd_sc_hd__nor2_1 U17774 ( .A(n11903), .B(n11705), .Y(n11901) );
  sky130_fd_sc_hd__nand3b_1 U17775 ( .A_N(n12944), .B(n28028), .C(n24400), .Y(
        n28152) );
  sky130_fd_sc_hd__nor2_1 U17776 ( .A(n12926), .B(n24620), .Y(n12925) );
  sky130_fd_sc_hd__inv_1 U17777 ( .A(n11906), .Y(n24620) );
  sky130_fd_sc_hd__nand3_2 U17778 ( .A(n11908), .B(n11906), .C(n24958), .Y(
        n24133) );
  sky130_fd_sc_hd__nand4_1 U17779 ( .A(n11906), .B(n27729), .C(n24545), .D(
        n24546), .Y(n24549) );
  sky130_fd_sc_hd__nand2_1 U17780 ( .A(n28270), .B(n11904), .Y(n28271) );
  sky130_fd_sc_hd__clkinv_1 U17781 ( .A(n24133), .Y(n28121) );
  sky130_fd_sc_hd__nor2_1 U17782 ( .A(n11909), .B(n11669), .Y(n11908) );
  sky130_fd_sc_hd__nand2_1 U17783 ( .A(n11001), .B(n29481), .Y(n12321) );
  sky130_fd_sc_hd__inv_2 U17784 ( .A(n12317), .Y(n23382) );
  sky130_fd_sc_hd__nor2_1 U17785 ( .A(n11912), .B(n23609), .Y(n23612) );
  sky130_fd_sc_hd__nor2_1 U17787 ( .A(n11916), .B(n11915), .Y(n11914) );
  sky130_fd_sc_hd__nand4_1 U17789 ( .A(n11924), .B(n20905), .C(n20906), .D(
        n20907), .Y(n11918) );
  sky130_fd_sc_hd__nand2_1 U17790 ( .A(n11920), .B(n12716), .Y(n11921) );
  sky130_fd_sc_hd__nand4_1 U17791 ( .A(n23609), .B(n23385), .C(n11841), .D(
        n11179), .Y(n11920) );
  sky130_fd_sc_hd__nand2_1 U17792 ( .A(n23384), .B(n23604), .Y(n23609) );
  sky130_fd_sc_hd__nand2_1 U17793 ( .A(n24607), .B(n12716), .Y(n28260) );
  sky130_fd_sc_hd__nand2_1 U17794 ( .A(n11923), .B(n12417), .Y(n11946) );
  sky130_fd_sc_hd__nand2_1 U17795 ( .A(n11923), .B(n29491), .Y(n24131) );
  sky130_fd_sc_hd__nand2_1 U17796 ( .A(n11923), .B(n11384), .Y(n24609) );
  sky130_fd_sc_hd__nand4_1 U17797 ( .A(n11924), .B(n20906), .C(n20905), .D(
        n20907), .Y(n20908) );
  sky130_fd_sc_hd__nand2_1 U17798 ( .A(j202_soc_core_memory0_ram_dout0[108]), 
        .B(n21488), .Y(n11924) );
  sky130_fd_sc_hd__o21ba_1 U17799 ( .A1(n11925), .A2(n24401), .B1_N(n24960), 
        .X(n24961) );
  sky130_fd_sc_hd__clkinv_1 U17800 ( .A(n28417), .Y(n11925) );
  sky130_fd_sc_hd__nor2_1 U17801 ( .A(n11926), .B(n11945), .Y(n11944) );
  sky130_fd_sc_hd__nor2_1 U17802 ( .A(n12524), .B(n30072), .Y(n11927) );
  sky130_fd_sc_hd__nand4_1 U17803 ( .A(n11932), .B(n11933), .C(n11931), .D(
        n11930), .Y(n12457) );
  sky130_fd_sc_hd__nand2_1 U17804 ( .A(j202_soc_core_memory0_ram_dout0[60]), 
        .B(n21633), .Y(n11930) );
  sky130_fd_sc_hd__nand2_1 U17805 ( .A(j202_soc_core_memory0_ram_dout0[476]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11931) );
  sky130_fd_sc_hd__nand2_1 U17806 ( .A(j202_soc_core_memory0_ram_dout0[348]), 
        .B(n21490), .Y(n11932) );
  sky130_fd_sc_hd__nand2_1 U17807 ( .A(j202_soc_core_memory0_ram_dout0[188]), 
        .B(n21487), .Y(n11933) );
  sky130_fd_sc_hd__nand4_1 U17808 ( .A(n11937), .B(n11936), .C(n11934), .D(
        n11935), .Y(n12000) );
  sky130_fd_sc_hd__nand2_1 U17809 ( .A(j202_soc_core_memory0_ram_dout0[284]), 
        .B(n21634), .Y(n11934) );
  sky130_fd_sc_hd__nand2_1 U17810 ( .A(j202_soc_core_memory0_ram_dout0[220]), 
        .B(n21640), .Y(n11935) );
  sky130_fd_sc_hd__nand2_1 U17811 ( .A(j202_soc_core_memory0_ram_dout0[380]), 
        .B(n21495), .Y(n11936) );
  sky130_fd_sc_hd__nand2_1 U17812 ( .A(j202_soc_core_memory0_ram_dout0[444]), 
        .B(n12156), .Y(n11937) );
  sky130_fd_sc_hd__nand4_1 U17813 ( .A(n12448), .B(n15660), .C(n15663), .D(
        n12449), .Y(n11938) );
  sky130_fd_sc_hd__nand4_1 U17814 ( .A(n12447), .B(n15659), .C(n15661), .D(
        n13000), .Y(n11939) );
  sky130_fd_sc_hd__nand2_1 U17815 ( .A(n11941), .B(n24400), .Y(n28388) );
  sky130_fd_sc_hd__nand3_1 U17816 ( .A(n11942), .B(n28367), .C(n24597), .Y(
        n10540) );
  sky130_fd_sc_hd__nand2_1 U17817 ( .A(n11943), .B(n28417), .Y(n11942) );
  sky130_fd_sc_hd__nand4_1 U17818 ( .A(n11946), .B(n24595), .C(n24594), .D(
        n11944), .Y(n11943) );
  sky130_fd_sc_hd__nand2_1 U17820 ( .A(n11949), .B(n11948), .Y(n11947) );
  sky130_fd_sc_hd__and3_1 U17821 ( .A(n25852), .B(n25850), .C(n25851), .X(
        n11948) );
  sky130_fd_sc_hd__nand2_1 U17822 ( .A(n25855), .B(n25847), .Y(n11949) );
  sky130_fd_sc_hd__o21a_1 U17823 ( .A1(n11951), .A2(n25845), .B1(n25836), .X(
        n11950) );
  sky130_fd_sc_hd__or2_0 U17825 ( .A(n25838), .B(n25837), .X(n11951) );
  sky130_fd_sc_hd__nand2_1 U17826 ( .A(n12455), .B(n12456), .Y(n20090) );
  sky130_fd_sc_hd__inv_1 U17827 ( .A(n11952), .Y(n20586) );
  sky130_fd_sc_hd__nand3_1 U17828 ( .A(n12954), .B(n12969), .C(n12444), .Y(
        n12443) );
  sky130_fd_sc_hd__nand2_1 U17829 ( .A(n11952), .B(n21917), .Y(n12954) );
  sky130_fd_sc_hd__nand2_1 U17830 ( .A(n12756), .B(n16293), .Y(n11952) );
  sky130_fd_sc_hd__nand4_1 U17831 ( .A(n11956), .B(n11955), .C(n11954), .D(
        n11953), .Y(n12896) );
  sky130_fd_sc_hd__nand2_1 U17832 ( .A(j202_soc_core_memory0_ram_dout0[55]), 
        .B(n21633), .Y(n11953) );
  sky130_fd_sc_hd__nand2_1 U17833 ( .A(j202_soc_core_memory0_ram_dout0[247]), 
        .B(n21641), .Y(n11954) );
  sky130_fd_sc_hd__nand2_1 U17834 ( .A(j202_soc_core_memory0_ram_dout0[23]), 
        .B(n21639), .Y(n11955) );
  sky130_fd_sc_hd__nand2_1 U17835 ( .A(j202_soc_core_memory0_ram_dout0[183]), 
        .B(n21487), .Y(n11956) );
  sky130_fd_sc_hd__nand2_1 U17836 ( .A(n11960), .B(n11958), .Y(n17643) );
  sky130_fd_sc_hd__nand2_1 U17837 ( .A(n11959), .B(n11963), .Y(n11958) );
  sky130_fd_sc_hd__nand2_1 U17838 ( .A(n12224), .B(n11961), .Y(n11960) );
  sky130_fd_sc_hd__nand2_1 U17839 ( .A(n11964), .B(n11962), .Y(n17548) );
  sky130_fd_sc_hd__nand2b_1 U17840 ( .A_N(n17515), .B(n11963), .Y(n11962) );
  sky130_fd_sc_hd__inv_2 U17841 ( .A(n19002), .Y(n11963) );
  sky130_fd_sc_hd__nand2_1 U17842 ( .A(n12224), .B(n23567), .Y(n11964) );
  sky130_fd_sc_hd__nand2_1 U17843 ( .A(n11966), .B(n11965), .Y(n19025) );
  sky130_fd_sc_hd__nand2_1 U17844 ( .A(n11455), .B(n19002), .Y(n11965) );
  sky130_fd_sc_hd__o22ai_1 U17845 ( .A1(n19002), .A2(n18973), .B1(n17381), 
        .B2(n11967), .Y(n18959) );
  sky130_fd_sc_hd__o22ai_1 U17846 ( .A1(n19002), .A2(n18382), .B1(n18500), 
        .B2(n11967), .Y(n18501) );
  sky130_fd_sc_hd__o22ai_1 U17847 ( .A1(n19002), .A2(n18500), .B1(n18499), 
        .B2(n11967), .Y(n18582) );
  sky130_fd_sc_hd__o22ai_1 U17848 ( .A1(n19002), .A2(n17433), .B1(n18386), 
        .B2(n11967), .Y(n18351) );
  sky130_fd_sc_hd__o22ai_1 U17849 ( .A1(n19002), .A2(n17415), .B1(n17433), 
        .B2(n11967), .Y(n18417) );
  sky130_fd_sc_hd__o22ai_1 U17850 ( .A1(n19002), .A2(n18385), .B1(n18382), 
        .B2(n11455), .Y(n18464) );
  sky130_fd_sc_hd__o22ai_2 U17851 ( .A1(n19002), .A2(n17381), .B1(n17374), 
        .B2(n11967), .Y(n17378) );
  sky130_fd_sc_hd__o22ai_1 U17852 ( .A1(n17675), .A2(n11967), .B1(n18499), 
        .B2(n19002), .Y(n18552) );
  sky130_fd_sc_hd__o22ai_1 U17853 ( .A1(n19002), .A2(n18386), .B1(n18385), 
        .B2(n11967), .Y(n18396) );
  sky130_fd_sc_hd__o22ai_1 U17854 ( .A1(n19002), .A2(n17374), .B1(n17406), 
        .B2(n11455), .Y(n17404) );
  sky130_fd_sc_hd__o22ai_1 U17855 ( .A1(n19002), .A2(n19001), .B1(n18973), 
        .B2(n11455), .Y(n19004) );
  sky130_fd_sc_hd__o22ai_1 U17856 ( .A1(n19002), .A2(n17406), .B1(n17415), 
        .B2(n11455), .Y(n17436) );
  sky130_fd_sc_hd__inv_4 U17857 ( .A(n25246), .Y(n26451) );
  sky130_fd_sc_hd__nand2_2 U17858 ( .A(n11968), .B(n13101), .Y(n25246) );
  sky130_fd_sc_hd__nand2_1 U17859 ( .A(n11969), .B(n25225), .Y(n11968) );
  sky130_fd_sc_hd__nand2_1 U17860 ( .A(n25223), .B(n25222), .Y(n11969) );
  sky130_fd_sc_hd__nand2_1 U17861 ( .A(n11970), .B(n11192), .Y(n12495) );
  sky130_fd_sc_hd__inv_1 U17862 ( .A(n21064), .Y(n11971) );
  sky130_fd_sc_hd__nand3_1 U17863 ( .A(n23021), .B(n11187), .C(n22177), .Y(
        n11973) );
  sky130_fd_sc_hd__nand2_1 U17864 ( .A(n11973), .B(n11974), .Y(n22179) );
  sky130_fd_sc_hd__nand2_1 U17865 ( .A(n23021), .B(n22177), .Y(n11975) );
  sky130_fd_sc_hd__nand2_1 U17866 ( .A(n11975), .B(n22176), .Y(n22270) );
  sky130_fd_sc_hd__o21a_1 U17867 ( .A1(n22178), .A2(n22176), .B1(n22268), .X(
        n11974) );
  sky130_fd_sc_hd__nand3_1 U17868 ( .A(n13360), .B(n13358), .C(n13359), .Y(
        n15647) );
  sky130_fd_sc_hd__nand2_4 U17872 ( .A(n30062), .B(n18796), .Y(n23514) );
  sky130_fd_sc_hd__nand2_1 U17875 ( .A(n11988), .B(n12298), .Y(n11982) );
  sky130_fd_sc_hd__nand2_1 U17876 ( .A(n11987), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[6]), .Y(n11983) );
  sky130_fd_sc_hd__nand2_1 U17877 ( .A(n13347), .B(n11985), .Y(n11984) );
  sky130_fd_sc_hd__nand2b_1 U17878 ( .A_N(n11988), .B(n11987), .Y(n11986) );
  sky130_fd_sc_hd__nand2_1 U17879 ( .A(n24673), .B(n23498), .Y(n13304) );
  sky130_fd_sc_hd__mux2i_1 U17880 ( .A0(n13145), .A1(n13146), .S(n11989), .Y(
        n11988) );
  sky130_fd_sc_hd__nand4_1 U17881 ( .A(n11993), .B(n11992), .C(n11991), .D(
        n11990), .Y(n12653) );
  sky130_fd_sc_hd__nand2_1 U17882 ( .A(j202_soc_core_memory0_ram_dout0[326]), 
        .B(n21490), .Y(n11990) );
  sky130_fd_sc_hd__nand2_1 U17883 ( .A(j202_soc_core_memory0_ram_dout0[294]), 
        .B(n21503), .Y(n11991) );
  sky130_fd_sc_hd__nand2_1 U17884 ( .A(j202_soc_core_memory0_ram_dout0[262]), 
        .B(n21634), .Y(n11992) );
  sky130_fd_sc_hd__nand2_1 U17885 ( .A(j202_soc_core_memory0_ram_dout0[390]), 
        .B(n21496), .Y(n11993) );
  sky130_fd_sc_hd__inv_2 U17886 ( .A(j202_soc_core_rst), .Y(n28914) );
  sky130_fd_sc_hd__nor2_1 U17887 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .B(j202_soc_core_rst), 
        .Y(n23853) );
  sky130_fd_sc_hd__nand3_1 U17890 ( .A(n28416), .B(n28415), .C(n11994), .Y(
        n28418) );
  sky130_fd_sc_hd__nor2_1 U17891 ( .A(n11995), .B(n12000), .Y(n12455) );
  sky130_fd_sc_hd__nand4_1 U17892 ( .A(n11998), .B(n11999), .C(n11996), .D(
        n11997), .Y(n11995) );
  sky130_fd_sc_hd__nand2_1 U17893 ( .A(j202_soc_core_memory0_ram_dout0[28]), 
        .B(n21639), .Y(n11996) );
  sky130_fd_sc_hd__nand2_1 U17894 ( .A(j202_soc_core_memory0_ram_dout0[316]), 
        .B(n21503), .Y(n11997) );
  sky130_fd_sc_hd__nand2_1 U17895 ( .A(j202_soc_core_memory0_ram_dout0[412]), 
        .B(n21496), .Y(n11998) );
  sky130_fd_sc_hd__nand2_1 U17896 ( .A(j202_soc_core_memory0_ram_dout0[252]), 
        .B(n21641), .Y(n11999) );
  sky130_fd_sc_hd__nand2_1 U17899 ( .A(j202_soc_core_memory0_ram_dout0[56]), 
        .B(n21633), .Y(n12003) );
  sky130_fd_sc_hd__nand2_1 U17900 ( .A(j202_soc_core_memory0_ram_dout0[344]), 
        .B(n21490), .Y(n12004) );
  sky130_fd_sc_hd__nand2_1 U17901 ( .A(j202_soc_core_memory0_ram_dout0[280]), 
        .B(n21634), .Y(n12005) );
  sky130_fd_sc_hd__nand2_1 U17902 ( .A(j202_soc_core_memory0_ram_dout0[433]), 
        .B(n12156), .Y(n12006) );
  sky130_fd_sc_hd__nand2_1 U17903 ( .A(j202_soc_core_memory0_ram_dout0[465]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12007) );
  sky130_fd_sc_hd__nand2_1 U17904 ( .A(j202_soc_core_memory0_ram_dout0[401]), 
        .B(n21496), .Y(n12008) );
  sky130_fd_sc_hd__nand2_1 U17905 ( .A(j202_soc_core_memory0_ram_dout0[369]), 
        .B(n21495), .Y(n12009) );
  sky130_fd_sc_hd__nand4_1 U17906 ( .A(n12013), .B(n12012), .C(n12011), .D(
        n12010), .Y(n12528) );
  sky130_fd_sc_hd__nand2_1 U17907 ( .A(j202_soc_core_memory0_ram_dout0[307]), 
        .B(n21503), .Y(n12010) );
  sky130_fd_sc_hd__nand2_1 U17908 ( .A(j202_soc_core_memory0_ram_dout0[243]), 
        .B(n21641), .Y(n12011) );
  sky130_fd_sc_hd__nand2_1 U17909 ( .A(j202_soc_core_memory0_ram_dout0[19]), 
        .B(n21639), .Y(n12012) );
  sky130_fd_sc_hd__nand2_1 U17910 ( .A(j202_soc_core_memory0_ram_dout0[339]), 
        .B(n21490), .Y(n12013) );
  sky130_fd_sc_hd__inv_1 U17911 ( .A(n12015), .Y(n12014) );
  sky130_fd_sc_hd__nand3_1 U17912 ( .A(n12021), .B(n12649), .C(n12020), .Y(
        n12015) );
  sky130_fd_sc_hd__nand2_1 U17913 ( .A(n12940), .B(n12125), .Y(n12018) );
  sky130_fd_sc_hd__nand2_1 U17914 ( .A(n12654), .B(n21917), .Y(n12019) );
  sky130_fd_sc_hd__nand2_1 U17915 ( .A(n12828), .B(n12650), .Y(n12020) );
  sky130_fd_sc_hd__o21a_1 U17916 ( .A1(n11203), .A2(n15174), .B1(n21172), .X(
        n12021) );
  sky130_fd_sc_hd__nand2_1 U17917 ( .A(n21336), .B(n21335), .Y(n24074) );
  sky130_fd_sc_hd__nand2_1 U17918 ( .A(n12718), .B(n12721), .Y(n12751) );
  sky130_fd_sc_hd__inv_2 U17919 ( .A(n21932), .Y(n12023) );
  sky130_fd_sc_hd__nand2_1 U17920 ( .A(n12024), .B(n21025), .Y(n21932) );
  sky130_fd_sc_hd__nand3_1 U17921 ( .A(n21024), .B(n21022), .C(n21023), .Y(
        n12024) );
  sky130_fd_sc_hd__a21oi_2 U17922 ( .A1(n21936), .A2(n26375), .B1(n12025), .Y(
        n21980) );
  sky130_fd_sc_hd__nand2_1 U17923 ( .A(n21956), .B(n21955), .Y(n12025) );
  sky130_fd_sc_hd__o21ai_1 U17924 ( .A1(n12028), .A2(n12798), .B1(n12027), .Y(
        n12026) );
  sky130_fd_sc_hd__nand2_1 U17925 ( .A(n12798), .B(n25397), .Y(n12027) );
  sky130_fd_sc_hd__clkinv_1 U17926 ( .A(n11123), .Y(n12028) );
  sky130_fd_sc_hd__nand2_1 U17928 ( .A(n12029), .B(n15482), .Y(n12862) );
  sky130_fd_sc_hd__nand2_1 U17929 ( .A(n11388), .B(n21917), .Y(n20585) );
  sky130_fd_sc_hd__nand2_2 U17930 ( .A(n12560), .B(n10969), .Y(n12730) );
  sky130_fd_sc_hd__inv_2 U17931 ( .A(n12730), .Y(n27148) );
  sky130_fd_sc_hd__nand3_1 U17932 ( .A(n12210), .B(n22115), .C(n22116), .Y(
        n12039) );
  sky130_fd_sc_hd__inv_2 U17933 ( .A(n13444), .Y(n21925) );
  sky130_fd_sc_hd__inv_1 U17935 ( .A(n12052), .Y(n12053) );
  sky130_fd_sc_hd__nand2_2 U17937 ( .A(n29593), .B(n23549), .Y(n23448) );
  sky130_fd_sc_hd__buf_6 U17938 ( .A(n24480), .X(n12043) );
  sky130_fd_sc_hd__nand2_4 U17939 ( .A(n17340), .B(n18989), .Y(n12044) );
  sky130_fd_sc_hd__inv_2 U17940 ( .A(n24479), .Y(n24480) );
  sky130_fd_sc_hd__xnor2_2 U17941 ( .A(n22526), .B(n27767), .Y(n17340) );
  sky130_fd_sc_hd__a21o_1 U17942 ( .A1(n12044), .A2(n18989), .B1(n18927), .X(
        n18944) );
  sky130_fd_sc_hd__inv_1 U17943 ( .A(n28430), .Y(n12045) );
  sky130_fd_sc_hd__inv_2 U17944 ( .A(n24497), .Y(n24498) );
  sky130_fd_sc_hd__nand2_1 U17945 ( .A(n23551), .B(n24404), .Y(n12964) );
  sky130_fd_sc_hd__inv_2 U17946 ( .A(n18202), .Y(n12047) );
  sky130_fd_sc_hd__inv_4 U17947 ( .A(n12047), .Y(n12048) );
  sky130_fd_sc_hd__nand2_1 U17948 ( .A(n17494), .B(n17495), .Y(n18202) );
  sky130_fd_sc_hd__inv_2 U17949 ( .A(n12049), .Y(n12050) );
  sky130_fd_sc_hd__o21a_1 U17950 ( .A1(n26164), .A2(n12351), .B1(n26159), .X(
        n28518) );
  sky130_fd_sc_hd__nand2_1 U17951 ( .A(n23438), .B(n23437), .Y(n12051) );
  sky130_fd_sc_hd__inv_4 U17952 ( .A(n27896), .Y(n27857) );
  sky130_fd_sc_hd__nor2_1 U17953 ( .A(n12764), .B(n12759), .Y(n12055) );
  sky130_fd_sc_hd__inv_2 U17956 ( .A(n25630), .Y(n12058) );
  sky130_fd_sc_hd__inv_2 U17957 ( .A(n25630), .Y(n12059) );
  sky130_fd_sc_hd__inv_2 U17958 ( .A(n25630), .Y(n25604) );
  sky130_fd_sc_hd__nand2_1 U17959 ( .A(n23548), .B(n28417), .Y(n12061) );
  sky130_fd_sc_hd__nand2_1 U17960 ( .A(n11175), .B(n12239), .Y(n23606) );
  sky130_fd_sc_hd__inv_2 U17961 ( .A(n11177), .Y(n12239) );
  sky130_fd_sc_hd__inv_2 U17962 ( .A(n13839), .Y(n16514) );
  sky130_fd_sc_hd__nor2_1 U17963 ( .A(n24091), .B(n12360), .Y(n12065) );
  sky130_fd_sc_hd__nand2_4 U17964 ( .A(n23421), .B(n22003), .Y(n12524) );
  sky130_fd_sc_hd__nand2_1 U17965 ( .A(n23606), .B(n12598), .Y(n23948) );
  sky130_fd_sc_hd__nor2_2 U17966 ( .A(n24421), .B(n24700), .Y(n12345) );
  sky130_fd_sc_hd__nand2_2 U17967 ( .A(n22004), .B(n12239), .Y(n28095) );
  sky130_fd_sc_hd__nand2_1 U17968 ( .A(n12288), .B(n28417), .Y(n28349) );
  sky130_fd_sc_hd__inv_2 U17969 ( .A(n12220), .Y(n12066) );
  sky130_fd_sc_hd__buf_2 U17970 ( .A(n23610), .X(n12430) );
  sky130_fd_sc_hd__o21a_1 U17971 ( .A1(n28495), .A2(n26378), .B1(n26306), .X(
        n26247) );
  sky130_fd_sc_hd__o211ai_2 U17972 ( .A1(n23850), .A2(n23849), .B1(n23848), 
        .C1(n24712), .Y(n29749) );
  sky130_fd_sc_hd__inv_8 U17973 ( .A(n29760), .Y(n12070) );
  sky130_fd_sc_hd__inv_8 U17974 ( .A(n29760), .Y(n12071) );
  sky130_fd_sc_hd__inv_8 U17975 ( .A(n29758), .Y(n12072) );
  sky130_fd_sc_hd__inv_8 U17976 ( .A(n29758), .Y(n12073) );
  sky130_fd_sc_hd__inv_8 U17977 ( .A(n29757), .Y(n12074) );
  sky130_fd_sc_hd__inv_8 U17978 ( .A(n29757), .Y(n12075) );
  sky130_fd_sc_hd__inv_8 U17979 ( .A(n29759), .Y(n12076) );
  sky130_fd_sc_hd__inv_8 U17980 ( .A(n29759), .Y(n12077) );
  sky130_fd_sc_hd__inv_8 U17981 ( .A(n29756), .Y(n12078) );
  sky130_fd_sc_hd__inv_8 U17982 ( .A(n29756), .Y(n12079) );
  sky130_fd_sc_hd__inv_8 U17983 ( .A(n29755), .Y(n12080) );
  sky130_fd_sc_hd__inv_8 U17984 ( .A(n29755), .Y(n12081) );
  sky130_fd_sc_hd__nor2_1 U17985 ( .A(n26903), .B(n12085), .Y(n12083) );
  sky130_fd_sc_hd__inv_8 U17986 ( .A(n29760), .Y(n12311) );
  sky130_fd_sc_hd__inv_8 U17987 ( .A(n29760), .Y(n12310) );
  sky130_fd_sc_hd__inv_8 U17988 ( .A(n29758), .Y(n12301) );
  sky130_fd_sc_hd__inv_8 U17989 ( .A(n29758), .Y(n12300) );
  sky130_fd_sc_hd__inv_8 U17990 ( .A(n29758), .Y(n12377) );
  sky130_fd_sc_hd__inv_8 U17991 ( .A(n29757), .Y(n12307) );
  sky130_fd_sc_hd__inv_8 U17992 ( .A(n29757), .Y(n12306) );
  sky130_fd_sc_hd__inv_8 U17993 ( .A(n29757), .Y(n12383) );
  sky130_fd_sc_hd__inv_8 U17994 ( .A(n29755), .Y(n12303) );
  sky130_fd_sc_hd__inv_8 U17995 ( .A(n29755), .Y(n12302) );
  sky130_fd_sc_hd__inv_8 U17996 ( .A(n29755), .Y(n12379) );
  sky130_fd_sc_hd__nor2_2 U17997 ( .A(n13154), .B(n13162), .Y(n21634) );
  sky130_fd_sc_hd__nor2_2 U17999 ( .A(j202_soc_core_j22_cpu_regop_other__2_), 
        .B(n13337), .Y(n13436) );
  sky130_fd_sc_hd__nor2_1 U18000 ( .A(n12054), .B(n13426), .Y(n14378) );
  sky130_fd_sc_hd__clkinv_1 U18001 ( .A(j202_soc_core_j22_cpu_id_op2_v_), .Y(
        n19539) );
  sky130_fd_sc_hd__clkinv_1 U18002 ( .A(n13362), .Y(n23643) );
  sky130_fd_sc_hd__and2_0 U18003 ( .A(n16618), .B(n16617), .X(n16682) );
  sky130_fd_sc_hd__xor2_1 U18004 ( .A(n13026), .B(n22023), .X(n13027) );
  sky130_fd_sc_hd__clkinv_1 U18005 ( .A(j202_soc_core_j22_cpu_ml_bufa[31]), 
        .Y(n13026) );
  sky130_fd_sc_hd__buf_4 U18006 ( .A(n13027), .X(n13025) );
  sky130_fd_sc_hd__clkinv_1 U18007 ( .A(j202_soc_core_j22_cpu_regop_Ra__0_), 
        .Y(n13513) );
  sky130_fd_sc_hd__clkinv_1 U18008 ( .A(n19141), .Y(n20740) );
  sky130_fd_sc_hd__nand2b_1 U18009 ( .A_N(n20814), .B(n20485), .Y(n20742) );
  sky130_fd_sc_hd__o22ai_1 U18010 ( .A1(n18213), .A2(n18081), .B1(n18212), 
        .B2(n12538), .Y(n18231) );
  sky130_fd_sc_hd__clkinv_1 U18011 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .Y(n19119) );
  sky130_fd_sc_hd__clkinv_1 U18012 ( .A(n17007), .Y(n17099) );
  sky130_fd_sc_hd__clkinv_1 U18013 ( .A(n17009), .Y(n16992) );
  sky130_fd_sc_hd__clkinv_1 U18014 ( .A(n13167), .Y(n13172) );
  sky130_fd_sc_hd__inv_2 U18015 ( .A(n11093), .Y(n14477) );
  sky130_fd_sc_hd__o211ai_1 U18016 ( .A1(n12565), .A2(n12564), .B1(n12563), 
        .C1(n12561), .Y(n19237) );
  sky130_fd_sc_hd__nor2_1 U18017 ( .A(n12158), .B(n12562), .Y(n12561) );
  sky130_fd_sc_hd__nand2_1 U18018 ( .A(n14378), .B(
        j202_soc_core_j22_cpu_regop_imm__12_), .Y(n16524) );
  sky130_fd_sc_hd__clkinv_1 U18020 ( .A(n13860), .Y(n13861) );
  sky130_fd_sc_hd__nor2_1 U18021 ( .A(n13263), .B(n13272), .Y(n19605) );
  sky130_fd_sc_hd__nand3_1 U18022 ( .A(n11108), .B(n21841), .C(n12196), .Y(
        n12195) );
  sky130_fd_sc_hd__nand3_1 U18023 ( .A(n18818), .B(n18805), .C(n26340), .Y(
        n26048) );
  sky130_fd_sc_hd__clkinv_1 U18024 ( .A(n21517), .Y(n20786) );
  sky130_fd_sc_hd__clkinv_1 U18026 ( .A(n20456), .Y(n15195) );
  sky130_fd_sc_hd__clkinv_1 U18027 ( .A(n20458), .Y(n15196) );
  sky130_fd_sc_hd__nor2_1 U18028 ( .A(n15194), .B(n15198), .Y(n21487) );
  sky130_fd_sc_hd__clkinv_1 U18029 ( .A(n20459), .Y(n15194) );
  sky130_fd_sc_hd__nand3_2 U18030 ( .A(n13160), .B(n13163), .C(n13159), .Y(
        n15198) );
  sky130_fd_sc_hd__clkinv_1 U18031 ( .A(n13162), .Y(n13160) );
  sky130_fd_sc_hd__inv_2 U18032 ( .A(n11093), .Y(n14342) );
  sky130_fd_sc_hd__clkinv_1 U18033 ( .A(n20460), .Y(n15199) );
  sky130_fd_sc_hd__nor2_1 U18034 ( .A(n15197), .B(n15198), .Y(n21640) );
  sky130_fd_sc_hd__clkinv_1 U18035 ( .A(n20457), .Y(n15193) );
  sky130_fd_sc_hd__clkinv_1 U18036 ( .A(j202_soc_core_j22_cpu_opst[4]), .Y(
        n23413) );
  sky130_fd_sc_hd__nor2_1 U18037 ( .A(n20898), .B(n30066), .Y(n12269) );
  sky130_fd_sc_hd__a21oi_1 U18038 ( .A1(n21291), .A2(n16523), .B1(n14016), .Y(
        n27023) );
  sky130_fd_sc_hd__nor2_1 U18039 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[1]), .B(
        n18799), .Y(n26189) );
  sky130_fd_sc_hd__nand2b_1 U18040 ( .A_N(n26048), .B(n25822), .Y(n26939) );
  sky130_fd_sc_hd__nand2b_1 U18041 ( .A_N(n26048), .B(n25824), .Y(n26919) );
  sky130_fd_sc_hd__nor2_1 U18042 ( .A(n28264), .B(n24616), .Y(n24618) );
  sky130_fd_sc_hd__inv_2 U18043 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[0]), .Y(
        n28104) );
  sky130_fd_sc_hd__inv_2 U18044 ( .A(n12622), .Y(n12332) );
  sky130_fd_sc_hd__clkinv_1 U18045 ( .A(n23412), .Y(n28086) );
  sky130_fd_sc_hd__clkinv_1 U18046 ( .A(n26746), .Y(n28313) );
  sky130_fd_sc_hd__clkinv_1 U18047 ( .A(j202_soc_core_j22_cpu_opst[0]), .Y(
        n28355) );
  sky130_fd_sc_hd__clkinv_1 U18048 ( .A(n28103), .Y(n24302) );
  sky130_fd_sc_hd__nor2_1 U18049 ( .A(j202_soc_core_j22_cpu_opst[2]), .B(
        n28355), .Y(n28402) );
  sky130_fd_sc_hd__o22ai_1 U18050 ( .A1(n18486), .A2(n17478), .B1(n17496), 
        .B2(n18483), .Y(n17486) );
  sky130_fd_sc_hd__clkinv_1 U18051 ( .A(n18428), .Y(n13032) );
  sky130_fd_sc_hd__o22ai_1 U18052 ( .A1(n19023), .A2(n18910), .B1(n18934), 
        .B2(n19020), .Y(n18923) );
  sky130_fd_sc_hd__nor2_1 U18054 ( .A(n13025), .B(n17336), .Y(n17426) );
  sky130_fd_sc_hd__clkinv_1 U18055 ( .A(n18477), .Y(n18346) );
  sky130_fd_sc_hd__clkinv_1 U18056 ( .A(n18476), .Y(n18347) );
  sky130_fd_sc_hd__nand3_1 U18057 ( .A(n20673), .B(n14597), .C(n17251), .Y(
        n21571) );
  sky130_fd_sc_hd__nand3_1 U18058 ( .A(n17268), .B(n14597), .C(n20304), .Y(
        n21536) );
  sky130_fd_sc_hd__clkinv_1 U18059 ( .A(n20307), .Y(n17105) );
  sky130_fd_sc_hd__nor2_1 U18060 ( .A(n13025), .B(n18905), .Y(n22029) );
  sky130_fd_sc_hd__o22ai_1 U18061 ( .A1(n18211), .A2(n12538), .B1(n18213), 
        .B2(n18212), .Y(n18225) );
  sky130_fd_sc_hd__inv_2 U18062 ( .A(n22833), .Y(n22782) );
  sky130_fd_sc_hd__nor2_1 U18063 ( .A(n13025), .B(n22025), .Y(n22039) );
  sky130_fd_sc_hd__inv_2 U18064 ( .A(n22039), .Y(n22038) );
  sky130_fd_sc_hd__and2_0 U18065 ( .A(n21351), .B(n21364), .X(n21430) );
  sky130_fd_sc_hd__and2_0 U18066 ( .A(n21365), .B(n21421), .X(n21428) );
  sky130_fd_sc_hd__nor2_1 U18067 ( .A(n12841), .B(n12840), .Y(n12839) );
  sky130_fd_sc_hd__nor2_1 U18068 ( .A(n14597), .B(n20034), .Y(n12840) );
  sky130_fd_sc_hd__clkinv_1 U18069 ( .A(n20024), .Y(n20148) );
  sky130_fd_sc_hd__clkinv_1 U18070 ( .A(n17242), .Y(n18697) );
  sky130_fd_sc_hd__clkinv_1 U18071 ( .A(n16977), .Y(n16968) );
  sky130_fd_sc_hd__clkinv_1 U18072 ( .A(n16950), .Y(n16980) );
  sky130_fd_sc_hd__and2_0 U18074 ( .A(n20767), .B(n20675), .X(n19179) );
  sky130_fd_sc_hd__nor2_1 U18076 ( .A(n14597), .B(
        j202_soc_core_bootrom_00_address_w[4]), .Y(n20393) );
  sky130_fd_sc_hd__clkinv_1 U18077 ( .A(n18670), .Y(n12485) );
  sky130_fd_sc_hd__nand2_1 U18078 ( .A(n12368), .B(n22230), .Y(n21838) );
  sky130_fd_sc_hd__a2bb2oi_1 U18079 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[35]), .B2(n26730), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[38]), .A2_N(n26711), .Y(n23088) );
  sky130_fd_sc_hd__nor2_1 U18080 ( .A(n13199), .B(n17243), .Y(n20303) );
  sky130_fd_sc_hd__nor2_1 U18081 ( .A(n14597), .B(n19140), .Y(n20833) );
  sky130_fd_sc_hd__inv_2 U18082 ( .A(n20563), .Y(n20551) );
  sky130_fd_sc_hd__clkinv_1 U18083 ( .A(
        j202_soc_core_memory0_ram_dout0_sel[10]), .Y(n13157) );
  sky130_fd_sc_hd__clkinv_1 U18084 ( .A(n16206), .Y(n20385) );
  sky130_fd_sc_hd__nand2_1 U18085 ( .A(n24673), .B(n23755), .Y(n13300) );
  sky130_fd_sc_hd__inv_2 U18087 ( .A(n13631), .Y(n15958) );
  sky130_fd_sc_hd__clkinv_1 U18088 ( .A(j202_soc_core_memory0_ram_dout0_sel[9]), .Y(n13163) );
  sky130_fd_sc_hd__inv_2 U18089 ( .A(n14001), .Y(n15992) );
  sky130_fd_sc_hd__and2_0 U18090 ( .A(n25804), .B(n25803), .X(n13103) );
  sky130_fd_sc_hd__inv_2 U18091 ( .A(n11148), .Y(n16444) );
  sky130_fd_sc_hd__clkinv_1 U18093 ( .A(n13411), .Y(n13827) );
  sky130_fd_sc_hd__clkinv_1 U18095 ( .A(n13838), .Y(n13631) );
  sky130_fd_sc_hd__clkinv_1 U18096 ( .A(n13821), .Y(n13616) );
  sky130_fd_sc_hd__clkinv_1 U18097 ( .A(n12099), .Y(n12494) );
  sky130_fd_sc_hd__and2_0 U18098 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[1]), 
        .B(j202_soc_core_uart_TOP_rx_fifo_rp[0]), .X(n21505) );
  sky130_fd_sc_hd__o21ai_1 U18099 ( .A1(n16014), .A2(n16013), .B1(n16012), .Y(
        n16896) );
  sky130_fd_sc_hd__nand3_1 U18100 ( .A(n30085), .B(n21841), .C(n12198), .Y(
        n12197) );
  sky130_fd_sc_hd__nand2b_1 U18101 ( .A_N(n12367), .B(n11205), .Y(n21841) );
  sky130_fd_sc_hd__mux2_2 U18102 ( .A0(j202_soc_core_intc_core_00_rg_ipr[16]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[20]), .S(n27321), .X(n23224) );
  sky130_fd_sc_hd__mux2_2 U18103 ( .A0(n23233), .A1(n23232), .S(n27319), .X(
        n23260) );
  sky130_fd_sc_hd__nor2_1 U18104 ( .A(n11184), .B(n24128), .Y(n12599) );
  sky130_fd_sc_hd__nand4_1 U18105 ( .A(n26162), .B(n24788), .C(n27148), .D(
        n26161), .Y(n26163) );
  sky130_fd_sc_hd__clkinv_1 U18106 ( .A(n25088), .Y(n25063) );
  sky130_fd_sc_hd__nand2_1 U18107 ( .A(n26001), .B(n22850), .Y(n23004) );
  sky130_fd_sc_hd__clkinv_1 U18108 ( .A(n23120), .Y(n12701) );
  sky130_fd_sc_hd__inv_2 U18109 ( .A(n16551), .Y(n17034) );
  sky130_fd_sc_hd__nor2_1 U18110 ( .A(n22413), .B(n13273), .Y(n21513) );
  sky130_fd_sc_hd__clkinv_1 U18111 ( .A(n21512), .Y(n20759) );
  sky130_fd_sc_hd__nand2_1 U18112 ( .A(j202_soc_core_memory0_ram_dout0[313]), 
        .B(n21503), .Y(n12937) );
  sky130_fd_sc_hd__nor2_1 U18114 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[1]), 
        .B(n28104), .Y(n26295) );
  sky130_fd_sc_hd__clkinv_1 U18116 ( .A(n26939), .Y(n27791) );
  sky130_fd_sc_hd__nand2_1 U18117 ( .A(n17965), .B(n17964), .Y(n22365) );
  sky130_fd_sc_hd__inv_2 U18118 ( .A(n14052), .Y(n23776) );
  sky130_fd_sc_hd__inv_2 U18119 ( .A(n13616), .Y(n23754) );
  sky130_fd_sc_hd__nand3_1 U18120 ( .A(n12687), .B(n22126), .C(n12686), .Y(
        n12685) );
  sky130_fd_sc_hd__nand3_1 U18121 ( .A(n12688), .B(n22239), .C(n21843), .Y(
        n12687) );
  sky130_fd_sc_hd__clkbuf_1 U18122 ( .A(n29594), .X(n12669) );
  sky130_fd_sc_hd__nand2_1 U18123 ( .A(n23587), .B(n27052), .Y(n24463) );
  sky130_fd_sc_hd__and2_1 U18124 ( .A(n24764), .B(n27052), .X(n24461) );
  sky130_fd_sc_hd__clkinv_1 U18125 ( .A(j202_soc_core_j22_cpu_regop_Rs__1_), 
        .Y(n22996) );
  sky130_fd_sc_hd__nor2_1 U18126 ( .A(n12590), .B(n12585), .Y(n12584) );
  sky130_fd_sc_hd__nor2_1 U18127 ( .A(n12596), .B(n12595), .Y(n12594) );
  sky130_fd_sc_hd__a21oi_1 U18128 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__13_), .B1(n21173), .Y(n21174) );
  sky130_fd_sc_hd__clkinv_1 U18129 ( .A(n15094), .Y(n12651) );
  sky130_fd_sc_hd__inv_2 U18130 ( .A(n21650), .Y(n21816) );
  sky130_fd_sc_hd__nand3_1 U18131 ( .A(n17067), .B(n16738), .C(n17065), .Y(
        n12574) );
  sky130_fd_sc_hd__nand3_1 U18133 ( .A(n12522), .B(n12523), .C(n15375), .Y(
        n25633) );
  sky130_fd_sc_hd__nand4_1 U18134 ( .A(n20869), .B(n20868), .C(n20870), .D(
        n20865), .Y(n12977) );
  sky130_fd_sc_hd__clkbuf_1 U18135 ( .A(n23398), .X(n24591) );
  sky130_fd_sc_hd__nor2_1 U18136 ( .A(j202_soc_core_j22_cpu_regop_We__2_), .B(
        n23845), .Y(n24176) );
  sky130_fd_sc_hd__inv_2 U18137 ( .A(n28056), .Y(n24456) );
  sky130_fd_sc_hd__nand3_1 U18138 ( .A(n23443), .B(n12280), .C(n23441), .Y(
        n24964) );
  sky130_fd_sc_hd__nand3_2 U18139 ( .A(n13436), .B(
        j202_soc_core_j22_cpu_regop_other__0_), .C(n18859), .Y(n16487) );
  sky130_fd_sc_hd__nand2_2 U18140 ( .A(n13436), .B(n13302), .Y(n16488) );
  sky130_fd_sc_hd__and2_0 U18141 ( .A(n29270), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd), .X(n29262) );
  sky130_fd_sc_hd__clkinv_1 U18142 ( .A(n27484), .Y(n27477) );
  sky130_fd_sc_hd__clkinv_1 U18143 ( .A(n27656), .Y(n29080) );
  sky130_fd_sc_hd__clkinv_1 U18144 ( .A(n27658), .Y(n29082) );
  sky130_fd_sc_hd__nor2_1 U18145 ( .A(n29088), .B(n27658), .Y(n27656) );
  sky130_fd_sc_hd__clkinv_1 U18146 ( .A(n26744), .Y(n28311) );
  sky130_fd_sc_hd__nor2_1 U18147 ( .A(n29088), .B(n26746), .Y(n26744) );
  sky130_fd_sc_hd__clkinv_1 U18148 ( .A(n28233), .Y(n29074) );
  sky130_fd_sc_hd__clkinv_1 U18149 ( .A(n28235), .Y(n29076) );
  sky130_fd_sc_hd__clkinv_1 U18150 ( .A(n26702), .Y(n28308) );
  sky130_fd_sc_hd__clkinv_1 U18151 ( .A(n26704), .Y(n28310) );
  sky130_fd_sc_hd__nor2_1 U18152 ( .A(n29088), .B(n26704), .Y(n26702) );
  sky130_fd_sc_hd__and2_0 U18153 ( .A(n23560), .B(n23623), .X(n13056) );
  sky130_fd_sc_hd__clkinv_1 U18154 ( .A(n27023), .Y(n28467) );
  sky130_fd_sc_hd__a21boi_0 U18155 ( .A1(n25728), .A2(n27789), .B1_N(n25302), 
        .Y(n25306) );
  sky130_fd_sc_hd__clkinv_1 U18156 ( .A(n29196), .Y(n29263) );
  sky130_fd_sc_hd__clkinv_1 U18157 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .Y(n28647) );
  sky130_fd_sc_hd__clkinv_1 U18158 ( .A(n26467), .Y(n28651) );
  sky130_fd_sc_hd__clkbuf_1 U18159 ( .A(j202_soc_core_j22_cpu_ml_bufa[26]), 
        .X(n27767) );
  sky130_fd_sc_hd__clkinv_1 U18160 ( .A(n28425), .Y(n27388) );
  sky130_fd_sc_hd__o31ai_1 U18161 ( .A1(n24289), .A2(n24288), .A3(n24287), 
        .B1(n28428), .Y(n27764) );
  sky130_fd_sc_hd__inv_2 U18162 ( .A(j202_soc_core_intr_req_), .Y(n28376) );
  sky130_fd_sc_hd__nand2b_1 U18163 ( .A_N(n23838), .B(n23837), .Y(n27648) );
  sky130_fd_sc_hd__clkinv_1 U18164 ( .A(n27648), .Y(n27860) );
  sky130_fd_sc_hd__nand3_1 U18165 ( .A(n13442), .B(n13441), .C(n12101), .Y(
        n28519) );
  sky130_fd_sc_hd__clkinv_1 U18166 ( .A(n22845), .Y(n27768) );
  sky130_fd_sc_hd__inv_2 U18167 ( .A(j202_soc_core_j22_cpu_regop_We__0_), .Y(
        n24771) );
  sky130_fd_sc_hd__clkinv_1 U18168 ( .A(n29542), .Y(n29070) );
  sky130_fd_sc_hd__nand2b_1 U18169 ( .A_N(n28090), .B(n28267), .Y(n28097) );
  sky130_fd_sc_hd__nor2_1 U18170 ( .A(n12779), .B(n28094), .Y(n28096) );
  sky130_fd_sc_hd__o21a_1 U18171 ( .A1(n11002), .A2(n24112), .B1(n10981), .X(
        n24113) );
  sky130_fd_sc_hd__inv_1 U18172 ( .A(n23377), .Y(n12703) );
  sky130_fd_sc_hd__nor2_1 U18173 ( .A(n12708), .B(n24393), .Y(n12707) );
  sky130_fd_sc_hd__and2_0 U18174 ( .A(n12157), .B(n12710), .X(n12088) );
  sky130_fd_sc_hd__clkinv_1 U18175 ( .A(n23376), .Y(n12710) );
  sky130_fd_sc_hd__clkinv_1 U18176 ( .A(n27530), .Y(n27544) );
  sky130_fd_sc_hd__clkinv_1 U18177 ( .A(n27540), .Y(n26990) );
  sky130_fd_sc_hd__clkinv_1 U18178 ( .A(n27850), .Y(n26070) );
  sky130_fd_sc_hd__clkinv_1 U18179 ( .A(n27855), .Y(n25724) );
  sky130_fd_sc_hd__clkinv_1 U18180 ( .A(n28518), .Y(n27114) );
  sky130_fd_sc_hd__clkinv_1 U18182 ( .A(n12708), .Y(n12706) );
  sky130_fd_sc_hd__clkinv_1 U18183 ( .A(n23855), .Y(n28721) );
  sky130_fd_sc_hd__clkinv_1 U18184 ( .A(n28724), .Y(n28886) );
  sky130_fd_sc_hd__nor2_1 U18185 ( .A(j202_soc_core_wbqspiflash_00_state[3]), 
        .B(n23640), .Y(n28870) );
  sky130_fd_sc_hd__clkinv_1 U18186 ( .A(n21653), .Y(n20454) );
  sky130_fd_sc_hd__a21oi_1 U18187 ( .A1(n29581), .A2(n24302), .B1(n24301), .Y(
        n27091) );
  sky130_fd_sc_hd__o21a_1 U18188 ( .A1(n24040), .A2(n24039), .B1(n24038), .X(
        n27848) );
  sky130_fd_sc_hd__nand2b_1 U18189 ( .A_N(n24037), .B(n24033), .Y(n27850) );
  sky130_fd_sc_hd__clkinv_1 U18190 ( .A(n22309), .Y(n23044) );
  sky130_fd_sc_hd__nor2_1 U18191 ( .A(n24590), .B(n24303), .Y(n27717) );
  sky130_fd_sc_hd__nor2_1 U18192 ( .A(n20427), .B(n24613), .Y(n28360) );
  sky130_fd_sc_hd__nand2_1 U18193 ( .A(n28109), .B(n29745), .Y(n24613) );
  sky130_fd_sc_hd__nand3_1 U18194 ( .A(n13293), .B(n28402), .C(n28086), .Y(
        n28367) );
  sky130_fd_sc_hd__buf_2 U18195 ( .A(n28062), .X(n12842) );
  sky130_fd_sc_hd__nand2_1 U18196 ( .A(n28360), .B(n23419), .Y(n28394) );
  sky130_fd_sc_hd__clkinv_1 U18197 ( .A(n24489), .Y(n24490) );
  sky130_fd_sc_hd__inv_2 U18199 ( .A(gpio_en_o[3]), .Y(io_oeb[3]) );
  sky130_fd_sc_hd__inv_2 U18201 ( .A(gpio_en_o[11]), .Y(io_oeb[31]) );
  sky130_fd_sc_hd__nand3_1 U18202 ( .A(n20947), .B(n20946), .C(n20945), .Y(
        n29473) );
  sky130_fd_sc_hd__clkinv_1 U18206 ( .A(n17519), .Y(n12537) );
  sky130_fd_sc_hd__nor2_1 U18207 ( .A(n13025), .B(n17411), .Y(n18415) );
  sky130_fd_sc_hd__nor2_1 U18208 ( .A(n13025), .B(n17430), .Y(n18355) );
  sky130_fd_sc_hd__clkinv_1 U18209 ( .A(n15712), .Y(n15713) );
  sky130_fd_sc_hd__inv_2 U18210 ( .A(n15340), .Y(n15590) );
  sky130_fd_sc_hd__nor2_1 U18212 ( .A(n13025), .B(n17366), .Y(n17390) );
  sky130_fd_sc_hd__clkinv_1 U18213 ( .A(n18468), .Y(n12508) );
  sky130_fd_sc_hd__nor2_1 U18214 ( .A(n18358), .B(n18357), .Y(n12407) );
  sky130_fd_sc_hd__o22ai_1 U18215 ( .A1(n24854), .A2(n21745), .B1(n18179), 
        .B2(n18536), .Y(n17524) );
  sky130_fd_sc_hd__clkinv_1 U18216 ( .A(n17944), .Y(n17902) );
  sky130_fd_sc_hd__o22ai_1 U18217 ( .A1(n24854), .A2(n21687), .B1(n22764), 
        .B2(n18536), .Y(n17953) );
  sky130_fd_sc_hd__o22ai_1 U18218 ( .A1(n18492), .A2(n17798), .B1(n17885), 
        .B2(n18489), .Y(n12163) );
  sky130_fd_sc_hd__o22ai_1 U18219 ( .A1(n24854), .A2(n22112), .B1(n22148), 
        .B2(n11561), .Y(n17689) );
  sky130_fd_sc_hd__nor2_1 U18220 ( .A(n13025), .B(n17382), .Y(n18957) );
  sky130_fd_sc_hd__nor2_1 U18221 ( .A(n13025), .B(n17364), .Y(n17401) );
  sky130_fd_sc_hd__nor2_1 U18222 ( .A(n13025), .B(n18917), .Y(n18929) );
  sky130_fd_sc_hd__nor2_1 U18223 ( .A(n13025), .B(n18926), .Y(n18945) );
  sky130_fd_sc_hd__nor2_1 U18224 ( .A(n18509), .B(n18511), .Y(n12505) );
  sky130_fd_sc_hd__nor2_1 U18225 ( .A(n13025), .B(n18343), .Y(n18398) );
  sky130_fd_sc_hd__nor2_1 U18226 ( .A(n13025), .B(n18344), .Y(n18393) );
  sky130_fd_sc_hd__clkinv_1 U18227 ( .A(n16632), .Y(n16633) );
  sky130_fd_sc_hd__inv_2 U18228 ( .A(n15678), .Y(n17241) );
  sky130_fd_sc_hd__nand3_1 U18229 ( .A(n21074), .B(n14597), .C(n11150), .Y(
        n15683) );
  sky130_fd_sc_hd__nor2_1 U18230 ( .A(n15675), .B(n15676), .Y(n21146) );
  sky130_fd_sc_hd__clkinv_1 U18231 ( .A(n16776), .Y(n16140) );
  sky130_fd_sc_hd__and2_0 U18232 ( .A(n14656), .B(n16776), .X(n16784) );
  sky130_fd_sc_hd__inv_2 U18233 ( .A(n19521), .Y(n19771) );
  sky130_fd_sc_hd__nor2_1 U18235 ( .A(n13025), .B(n18943), .Y(n19035) );
  sky130_fd_sc_hd__nor2_1 U18236 ( .A(n13027), .B(n18965), .Y(n18984) );
  sky130_fd_sc_hd__nor2_1 U18237 ( .A(n13025), .B(n19000), .Y(n19026) );
  sky130_fd_sc_hd__clkinv_1 U18238 ( .A(n17948), .Y(n12475) );
  sky130_fd_sc_hd__and2_0 U18239 ( .A(n22541), .B(n22507), .X(n22509) );
  sky130_fd_sc_hd__o2bb2ai_1 U18240 ( .B1(n19002), .B2(n17593), .A1_N(n12481), 
        .A2_N(n12224), .Y(n12480) );
  sky130_fd_sc_hd__o22ai_1 U18241 ( .A1(n24854), .A2(n21893), .B1(n22630), 
        .B2(n18536), .Y(n17679) );
  sky130_fd_sc_hd__o22ai_1 U18242 ( .A1(n18474), .A2(n17633), .B1(n17586), 
        .B2(n18471), .Y(n12668) );
  sky130_fd_sc_hd__clkinv_1 U18243 ( .A(n17799), .Y(n12484) );
  sky130_fd_sc_hd__o22ai_1 U18244 ( .A1(n18209), .A2(n18029), .B1(n18074), 
        .B2(n18206), .Y(n18032) );
  sky130_fd_sc_hd__nor2_1 U18245 ( .A(n13025), .B(n18907), .Y(n18913) );
  sky130_fd_sc_hd__clkinv_1 U18246 ( .A(n18601), .Y(n12488) );
  sky130_fd_sc_hd__inv_2 U18247 ( .A(j202_soc_core_j22_cpu_regop_Rm__1_), .Y(
        n13381) );
  sky130_fd_sc_hd__clkinv_1 U18248 ( .A(n18592), .Y(n12672) );
  sky130_fd_sc_hd__nor2_1 U18249 ( .A(n13025), .B(n18909), .Y(n18922) );
  sky130_fd_sc_hd__nand2_1 U18250 ( .A(n13413), .B(
        j202_soc_core_j22_cpu_regop_Rm__2_), .Y(n13402) );
  sky130_fd_sc_hd__and2_0 U18251 ( .A(n21394), .B(n21575), .X(n21551) );
  sky130_fd_sc_hd__and2_0 U18252 ( .A(n21574), .B(n21536), .X(n21385) );
  sky130_fd_sc_hd__inv_2 U18253 ( .A(n22921), .Y(n21761) );
  sky130_fd_sc_hd__inv_2 U18254 ( .A(n22918), .Y(n21762) );
  sky130_fd_sc_hd__and2_0 U18255 ( .A(n19814), .B(n19781), .X(n19743) );
  sky130_fd_sc_hd__clkinv_1 U18256 ( .A(n19716), .Y(n19441) );
  sky130_fd_sc_hd__clkinv_1 U18257 ( .A(n28460), .Y(n26310) );
  sky130_fd_sc_hd__clkinv_1 U18258 ( .A(j202_soc_core_bootrom_00_address_w[10]), .Y(n18712) );
  sky130_fd_sc_hd__clkinv_1 U18259 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .Y(n13180) );
  sky130_fd_sc_hd__and2_0 U18260 ( .A(n21380), .B(n20058), .X(n21386) );
  sky130_fd_sc_hd__clkinv_1 U18261 ( .A(n19185), .Y(n15700) );
  sky130_fd_sc_hd__clkinv_1 U18262 ( .A(n20767), .Y(n20468) );
  sky130_fd_sc_hd__nand2b_1 U18263 ( .A_N(n20560), .B(n19119), .Y(n20837) );
  sky130_fd_sc_hd__inv_2 U18264 ( .A(n20634), .Y(n20680) );
  sky130_fd_sc_hd__nand4bb_1 U18265 ( .A_N(n20601), .B_N(n20600), .C(n20747), 
        .D(n20679), .Y(n20602) );
  sky130_fd_sc_hd__clkinv_1 U18266 ( .A(n20387), .Y(n19392) );
  sky130_fd_sc_hd__and2_0 U18267 ( .A(n19369), .B(n20348), .X(n19659) );
  sky130_fd_sc_hd__and2_0 U18268 ( .A(n20372), .B(n19369), .X(n20311) );
  sky130_fd_sc_hd__and2_0 U18269 ( .A(n20316), .B(n20390), .X(n19617) );
  sky130_fd_sc_hd__and2_0 U18270 ( .A(n19404), .B(n20380), .X(n19660) );
  sky130_fd_sc_hd__clkinv_1 U18271 ( .A(n20278), .Y(n20279) );
  sky130_fd_sc_hd__clkinv_1 U18272 ( .A(n20884), .Y(n12445) );
  sky130_fd_sc_hd__clkinv_1 U18273 ( .A(n17061), .Y(n16198) );
  sky130_fd_sc_hd__inv_2 U18275 ( .A(n13761), .Y(n15984) );
  sky130_fd_sc_hd__clkinv_1 U18276 ( .A(n26932), .Y(n24930) );
  sky130_fd_sc_hd__clkinv_1 U18277 ( .A(n27793), .Y(n26034) );
  sky130_fd_sc_hd__clkinv_1 U18278 ( .A(n18619), .Y(n18621) );
  sky130_fd_sc_hd__clkinv_1 U18279 ( .A(n17637), .Y(n12682) );
  sky130_fd_sc_hd__clkinv_1 U18280 ( .A(n17850), .Y(n17852) );
  sky130_fd_sc_hd__clkinv_1 U18281 ( .A(n13467), .Y(n14209) );
  sky130_fd_sc_hd__o2bb2ai_1 U18282 ( .B1(n17748), .B2(n17747), .A1_N(n17806), 
        .A2_N(n17807), .Y(n17811) );
  sky130_fd_sc_hd__clkinv_1 U18283 ( .A(n19010), .Y(n17395) );
  sky130_fd_sc_hd__clkinv_1 U18284 ( .A(n22105), .Y(n19062) );
  sky130_fd_sc_hd__inv_2 U18285 ( .A(n13385), .Y(n13408) );
  sky130_fd_sc_hd__nand2_1 U18286 ( .A(n23030), .B(n22923), .Y(n22925) );
  sky130_fd_sc_hd__nor2_1 U18287 ( .A(n22199), .B(n22190), .Y(n18668) );
  sky130_fd_sc_hd__and2_0 U18289 ( .A(n21392), .B(n21391), .X(n13044) );
  sky130_fd_sc_hd__clkinv_1 U18291 ( .A(n12202), .Y(n12200) );
  sky130_fd_sc_hd__clkinv_1 U18292 ( .A(n21862), .Y(n12196) );
  sky130_fd_sc_hd__inv_2 U18293 ( .A(n21193), .Y(n22202) );
  sky130_fd_sc_hd__inv_2 U18294 ( .A(n27115), .Y(n27800) );
  sky130_fd_sc_hd__inv_2 U18295 ( .A(n20175), .Y(n20130) );
  sky130_fd_sc_hd__clkinv_1 U18296 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .Y(n20485) );
  sky130_fd_sc_hd__mux2_2 U18297 ( .A0(n23135), .A1(n23134), .S(n27326), .X(
        n23256) );
  sky130_fd_sc_hd__o2bb2ai_1 U18298 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[12]), .B2(n25164), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[9]), .A2_N(n25162), .Y(n23151) );
  sky130_fd_sc_hd__and2_0 U18299 ( .A(n20533), .B(n20559), .X(n20534) );
  sky130_fd_sc_hd__clkinv_1 U18300 ( .A(
        j202_soc_core_memory0_ram_dout0_sel[12]), .Y(n13150) );
  sky130_fd_sc_hd__clkinv_1 U18301 ( .A(n19689), .Y(n19677) );
  sky130_fd_sc_hd__clkinv_1 U18302 ( .A(n20395), .Y(n19546) );
  sky130_fd_sc_hd__inv_2 U18303 ( .A(n16139), .Y(n20374) );
  sky130_fd_sc_hd__clkinv_1 U18304 ( .A(n16207), .Y(n20368) );
  sky130_fd_sc_hd__clkinv_1 U18307 ( .A(n16667), .Y(n20643) );
  sky130_fd_sc_hd__a21boi_0 U18308 ( .A1(n20406), .A2(n20757), .B1_N(n20405), 
        .Y(n20407) );
  sky130_fd_sc_hd__inv_2 U18309 ( .A(n18887), .Y(n17933) );
  sky130_fd_sc_hd__clkbuf_1 U18310 ( .A(n13587), .X(n16500) );
  sky130_fd_sc_hd__and2_0 U18311 ( .A(n24991), .B(n24990), .X(n24992) );
  sky130_fd_sc_hd__and2_0 U18312 ( .A(n24989), .B(n24988), .X(n24993) );
  sky130_fd_sc_hd__and2_0 U18313 ( .A(n24985), .B(n24984), .X(n24995) );
  sky130_fd_sc_hd__and2_0 U18314 ( .A(n24987), .B(n24986), .X(n24994) );
  sky130_fd_sc_hd__inv_2 U18315 ( .A(n13827), .Y(n16466) );
  sky130_fd_sc_hd__clkinv_1 U18316 ( .A(n27799), .Y(n26930) );
  sky130_fd_sc_hd__clkinv_1 U18317 ( .A(n27815), .Y(n25648) );
  sky130_fd_sc_hd__clkinv_1 U18318 ( .A(n22676), .Y(n12170) );
  sky130_fd_sc_hd__buf_2 U18319 ( .A(j202_soc_core_j22_cpu_ml_bufb[0]), .X(
        n18470) );
  sky130_fd_sc_hd__clkinv_1 U18320 ( .A(n13818), .Y(n13725) );
  sky130_fd_sc_hd__clkinv_1 U18321 ( .A(n24069), .Y(n25938) );
  sky130_fd_sc_hd__clkinv_1 U18322 ( .A(n25688), .Y(n27810) );
  sky130_fd_sc_hd__and2_0 U18323 ( .A(n27826), .B(n27052), .X(n27782) );
  sky130_fd_sc_hd__clkinv_1 U18324 ( .A(n25261), .Y(n25256) );
  sky130_fd_sc_hd__and2_0 U18325 ( .A(n23925), .B(n23924), .X(n23929) );
  sky130_fd_sc_hd__and2_0 U18326 ( .A(n23927), .B(n23926), .X(n23928) );
  sky130_fd_sc_hd__and2_0 U18327 ( .A(n23923), .B(n23922), .X(n23930) );
  sky130_fd_sc_hd__nor2_1 U18328 ( .A(n18846), .B(n18845), .Y(n27808) );
  sky130_fd_sc_hd__inv_2 U18329 ( .A(n25999), .Y(n18846) );
  sky130_fd_sc_hd__maj3_1 U18330 ( .A(n23315), .B(n23317), .C(n23304), .X(
        n23310) );
  sky130_fd_sc_hd__a21boi_0 U18331 ( .A1(n24044), .A2(n27789), .B1_N(n22254), 
        .Y(n22255) );
  sky130_fd_sc_hd__nand2_1 U18332 ( .A(n12393), .B(n29593), .Y(n23613) );
  sky130_fd_sc_hd__clkinv_1 U18334 ( .A(n26365), .Y(n26366) );
  sky130_fd_sc_hd__clkinv_1 U18335 ( .A(n26210), .Y(n26346) );
  sky130_fd_sc_hd__clkinv_1 U18336 ( .A(n26205), .Y(n26207) );
  sky130_fd_sc_hd__and2_0 U18337 ( .A(n21689), .B(n22230), .X(n12138) );
  sky130_fd_sc_hd__nand2_1 U18338 ( .A(n23427), .B(n11141), .Y(n12572) );
  sky130_fd_sc_hd__inv_1 U18339 ( .A(n22225), .Y(n12802) );
  sky130_fd_sc_hd__nor2_1 U18340 ( .A(n12115), .B(n20101), .Y(n19983) );
  sky130_fd_sc_hd__nand3_1 U18341 ( .A(n12829), .B(n12830), .C(n15092), .Y(
        n12828) );
  sky130_fd_sc_hd__clkinv_1 U18344 ( .A(n20200), .Y(n20179) );
  sky130_fd_sc_hd__nor2_1 U18345 ( .A(n13173), .B(n13172), .Y(n20460) );
  sky130_fd_sc_hd__a21oi_1 U18346 ( .A1(n23125), .A2(n23124), .B1(n12694), .Y(
        n12693) );
  sky130_fd_sc_hd__nor2_1 U18347 ( .A(n23124), .B(n23125), .Y(n12696) );
  sky130_fd_sc_hd__nand2_1 U18348 ( .A(j202_soc_core_memory0_ram_dout0[319]), 
        .B(n21503), .Y(n12577) );
  sky130_fd_sc_hd__o21a_1 U18349 ( .A1(n20863), .A2(n20862), .B1(n21629), .X(
        n20880) );
  sky130_fd_sc_hd__nor2_1 U18351 ( .A(n13277), .B(n13276), .Y(n21516) );
  sky130_fd_sc_hd__clkinv_1 U18352 ( .A(n21515), .Y(n20540) );
  sky130_fd_sc_hd__and3_1 U18353 ( .A(n21629), .B(n17264), .C(n21101), .X(
        n20784) );
  sky130_fd_sc_hd__and2_0 U18354 ( .A(n21629), .B(n16996), .X(n20757) );
  sky130_fd_sc_hd__clkinv_1 U18355 ( .A(n20684), .Y(n20856) );
  sky130_fd_sc_hd__and2_0 U18356 ( .A(n15256), .B(n21917), .X(n12125) );
  sky130_fd_sc_hd__and2_0 U18357 ( .A(n17333), .B(n21919), .X(n12109) );
  sky130_fd_sc_hd__clkinv_1 U18358 ( .A(n17205), .Y(n12743) );
  sky130_fd_sc_hd__clkinv_1 U18361 ( .A(n13072), .Y(n12776) );
  sky130_fd_sc_hd__nand2_1 U18362 ( .A(n11449), .B(n28394), .Y(n12926) );
  sky130_fd_sc_hd__clkinv_1 U18363 ( .A(j202_soc_core_gpio_core_00_reg_addr[1]), .Y(n26773) );
  sky130_fd_sc_hd__buf_4 U18364 ( .A(j202_soc_core_j22_cpu_ml_bufa[21]), .X(
        n22299) );
  sky130_fd_sc_hd__inv_2 U18365 ( .A(n24345), .Y(n17994) );
  sky130_fd_sc_hd__and2_0 U18366 ( .A(n28204), .B(n28202), .X(n25179) );
  sky130_fd_sc_hd__clkinv_1 U18367 ( .A(n25090), .Y(n29406) );
  sky130_fd_sc_hd__clkinv_1 U18368 ( .A(j202_soc_core_j22_cpu_rf_pr[12]), .Y(
        n21885) );
  sky130_fd_sc_hd__clkinv_1 U18369 ( .A(n18261), .Y(n12885) );
  sky130_fd_sc_hd__a21boi_0 U18370 ( .A1(n24947), .A2(n27789), .B1_N(n24946), 
        .Y(n24949) );
  sky130_fd_sc_hd__and2_0 U18371 ( .A(n24281), .B(n26189), .X(n24282) );
  sky130_fd_sc_hd__clkinv_1 U18372 ( .A(n28685), .Y(n26637) );
  sky130_fd_sc_hd__inv_2 U18373 ( .A(n18686), .Y(n22967) );
  sky130_fd_sc_hd__inv_1 U18374 ( .A(n22713), .Y(n22072) );
  sky130_fd_sc_hd__clkinv_1 U18375 ( .A(n27615), .Y(n24287) );
  sky130_fd_sc_hd__nand2_1 U18376 ( .A(n23485), .B(n24452), .Y(n22439) );
  sky130_fd_sc_hd__nand3_1 U18377 ( .A(n11171), .B(n12494), .C(n23030), .Y(
        n12490) );
  sky130_fd_sc_hd__o2bb2ai_1 U18378 ( .B1(n12494), .B2(n22106), .A1_N(n12493), 
        .A2_N(n22106), .Y(n12492) );
  sky130_fd_sc_hd__xnor2_1 U18379 ( .A(n23025), .B(n23024), .Y(n24439) );
  sky130_fd_sc_hd__and2_0 U18380 ( .A(n16096), .B(n16095), .X(n16302) );
  sky130_fd_sc_hd__nand3_1 U18381 ( .A(n20717), .B(n20716), .C(n22114), .Y(
        n12571) );
  sky130_fd_sc_hd__clkinv_1 U18382 ( .A(n27153), .Y(n12341) );
  sky130_fd_sc_hd__nor2_1 U18383 ( .A(n12819), .B(n12220), .Y(n12818) );
  sky130_fd_sc_hd__inv_2 U18384 ( .A(n26341), .Y(n24910) );
  sky130_fd_sc_hd__nand3_1 U18385 ( .A(n27572), .B(n26916), .C(n26064), .Y(
        n26065) );
  sky130_fd_sc_hd__nand2_1 U18386 ( .A(n23577), .B(n24452), .Y(n25993) );
  sky130_fd_sc_hd__clkinv_1 U18387 ( .A(n21519), .Y(n21446) );
  sky130_fd_sc_hd__clkinv_1 U18388 ( .A(n27807), .Y(n26323) );
  sky130_fd_sc_hd__clkinv_1 U18389 ( .A(n18818), .Y(n27789) );
  sky130_fd_sc_hd__clkinv_1 U18390 ( .A(n24758), .Y(n24732) );
  sky130_fd_sc_hd__and2_0 U18391 ( .A(n10971), .B(n26189), .X(n25214) );
  sky130_fd_sc_hd__nand2_1 U18392 ( .A(n23469), .B(n24452), .Y(n22405) );
  sky130_fd_sc_hd__and2_0 U18394 ( .A(j202_soc_core_intc_core_00_bs_addr[2]), 
        .B(j202_soc_core_intc_core_00_bs_addr[8]), .X(n25062) );
  sky130_fd_sc_hd__clkinv_1 U18395 ( .A(n28326), .Y(n28238) );
  sky130_fd_sc_hd__clkinv_1 U18396 ( .A(n22084), .Y(n22986) );
  sky130_fd_sc_hd__clkinv_1 U18398 ( .A(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n21768) );
  sky130_fd_sc_hd__clkinv_1 U18399 ( .A(n15527), .Y(n20196) );
  sky130_fd_sc_hd__nand3_1 U18400 ( .A(n20461), .B(n12608), .C(n12607), .Y(
        n12606) );
  sky130_fd_sc_hd__inv_1 U18401 ( .A(n23273), .Y(n23366) );
  sky130_fd_sc_hd__clkinv_1 U18402 ( .A(n23076), .Y(n27328) );
  sky130_fd_sc_hd__a21oi_1 U18403 ( .A1(n23297), .A2(n23296), .B1(n23295), .Y(
        n27339) );
  sky130_fd_sc_hd__nand2_1 U18404 ( .A(n23171), .B(n23170), .Y(n27316) );
  sky130_fd_sc_hd__clkinv_1 U18405 ( .A(n24757), .Y(n24738) );
  sky130_fd_sc_hd__clkinv_1 U18406 ( .A(n28676), .Y(n27195) );
  sky130_fd_sc_hd__clkinv_1 U18407 ( .A(n27193), .Y(n27196) );
  sky130_fd_sc_hd__and2_0 U18408 ( .A(n28837), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .X(n28655) );
  sky130_fd_sc_hd__clkinv_1 U18409 ( .A(n27288), .Y(n27291) );
  sky130_fd_sc_hd__clkinv_1 U18410 ( .A(n27289), .Y(n27290) );
  sky130_fd_sc_hd__and2_0 U18411 ( .A(n27430), .B(n26534), .X(n26538) );
  sky130_fd_sc_hd__clkinv_1 U18412 ( .A(n28729), .Y(n26535) );
  sky130_fd_sc_hd__clkinv_1 U18413 ( .A(n27240), .Y(n28828) );
  sky130_fd_sc_hd__and2_0 U18415 ( .A(n21817), .B(n21815), .X(n19926) );
  sky130_fd_sc_hd__nor2_1 U18416 ( .A(n11203), .B(n16294), .Y(n12879) );
  sky130_fd_sc_hd__nand2_1 U18417 ( .A(j202_soc_core_memory0_ram_dout0[345]), 
        .B(n21490), .Y(n12939) );
  sky130_fd_sc_hd__clkinv_1 U18418 ( .A(n19857), .Y(n21916) );
  sky130_fd_sc_hd__nand3_1 U18419 ( .A(n12805), .B(n13177), .C(n12804), .Y(
        n12803) );
  sky130_fd_sc_hd__inv_2 U18420 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[5]), .Y(
        n26142) );
  sky130_fd_sc_hd__clkinv_1 U18421 ( .A(n24852), .Y(n24452) );
  sky130_fd_sc_hd__inv_2 U18422 ( .A(j202_soc_core_intc_core_00_rg_ipr[8]), 
        .Y(n25164) );
  sky130_fd_sc_hd__clkinv_1 U18423 ( .A(j202_soc_core_intc_core_00_rg_ipr[53]), 
        .Y(n25576) );
  sky130_fd_sc_hd__clkinv_1 U18424 ( .A(j202_soc_core_intc_core_00_bs_addr[0]), 
        .Y(n25050) );
  sky130_fd_sc_hd__clkinv_1 U18425 ( .A(j202_soc_core_intc_core_00_bs_addr[1]), 
        .Y(n25046) );
  sky130_fd_sc_hd__clkinv_1 U18426 ( .A(n28817), .Y(n28888) );
  sky130_fd_sc_hd__and2_0 U18428 ( .A(n29270), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[2]), .X(n29648) );
  sky130_fd_sc_hd__nand3_2 U18429 ( .A(n14295), .B(n14294), .C(n14293), .Y(
        n28489) );
  sky130_fd_sc_hd__and2_0 U18430 ( .A(n28837), .B(n26485), .X(n28864) );
  sky130_fd_sc_hd__clkinv_1 U18431 ( .A(n25594), .Y(n12222) );
  sky130_fd_sc_hd__clkinv_1 U18432 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[4]), .Y(n28930) );
  sky130_fd_sc_hd__clkinv_1 U18433 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[8]), .Y(n28958) );
  sky130_fd_sc_hd__clkinv_1 U18434 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[16]), .Y(n29015) );
  sky130_fd_sc_hd__clkinv_1 U18435 ( .A(gpio_en_o[24]), .Y(n29052) );
  sky130_fd_sc_hd__clkinv_1 U18436 ( .A(gpio_en_o[28]), .Y(n29059) );
  sky130_fd_sc_hd__clkinv_1 U18437 ( .A(n29061), .Y(n29039) );
  sky130_fd_sc_hd__clkinv_1 U18438 ( .A(n28595), .Y(n29300) );
  sky130_fd_sc_hd__and2_0 U18439 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[0]), 
        .B(j202_soc_core_uart_TOP_tx_fifo_rp[1]), .X(n29302) );
  sky130_fd_sc_hd__a21oi_1 U18440 ( .A1(n22997), .A2(n16523), .B1(n14182), .Y(
        n25451) );
  sky130_fd_sc_hd__inv_1 U18441 ( .A(n28535), .Y(n28437) );
  sky130_fd_sc_hd__clkinv_1 U18442 ( .A(n26311), .Y(n28443) );
  sky130_fd_sc_hd__and2_0 U18443 ( .A(j202_soc_core_cmt_core_00_cnt0[0]), .B(
        j202_soc_core_cmt_core_00_cnt0[1]), .X(n27472) );
  sky130_fd_sc_hd__clkinv_1 U18444 ( .A(n28219), .Y(n28220) );
  sky130_fd_sc_hd__clkinv_1 U18445 ( .A(n25083), .Y(n28317) );
  sky130_fd_sc_hd__nor2_1 U18446 ( .A(n12429), .B(n25887), .Y(n12428) );
  sky130_fd_sc_hd__a21boi_0 U18447 ( .A1(n22848), .A2(n24764), .B1_N(n22847), 
        .Y(n25307) );
  sky130_fd_sc_hd__nand3_2 U18448 ( .A(n14433), .B(n12096), .C(n14432), .Y(
        n26051) );
  sky130_fd_sc_hd__nor2_1 U18449 ( .A(n25098), .B(n25097), .Y(n28330) );
  sky130_fd_sc_hd__clkinv_1 U18450 ( .A(j202_soc_core_intc_core_00_rg_ipr[50]), 
        .Y(n26736) );
  sky130_fd_sc_hd__clkinv_1 U18452 ( .A(j202_soc_core_intc_core_00_rg_ipr[32]), 
        .Y(n26727) );
  sky130_fd_sc_hd__nand2_1 U18453 ( .A(n25069), .B(n25068), .Y(n26760) );
  sky130_fd_sc_hd__nand2_1 U18454 ( .A(n28316), .B(n29827), .Y(n28314) );
  sky130_fd_sc_hd__inv_2 U18456 ( .A(j202_soc_core_intc_core_00_rg_ipr[10]), 
        .Y(n25071) );
  sky130_fd_sc_hd__nand2_1 U18457 ( .A(n29143), .B(n25084), .Y(n28064) );
  sky130_fd_sc_hd__inv_2 U18458 ( .A(n29565), .Y(n27090) );
  sky130_fd_sc_hd__inv_2 U18459 ( .A(n28466), .Y(n28113) );
  sky130_fd_sc_hd__clkinv_1 U18460 ( .A(n28459), .Y(n26670) );
  sky130_fd_sc_hd__inv_2 U18461 ( .A(n26961), .Y(n26965) );
  sky130_fd_sc_hd__inv_2 U18462 ( .A(n28483), .Y(n26975) );
  sky130_fd_sc_hd__clkinv_1 U18463 ( .A(n26416), .Y(n28429) );
  sky130_fd_sc_hd__clkinv_1 U18464 ( .A(n27271), .Y(n27234) );
  sky130_fd_sc_hd__clkinv_1 U18465 ( .A(n27119), .Y(n25776) );
  sky130_fd_sc_hd__buf_4 U18466 ( .A(j202_soc_core_j22_cpu_ml_bufa[29]), .X(
        n25389) );
  sky130_fd_sc_hd__a21boi_1 U18467 ( .A1(n22525), .A2(n24764), .B1_N(n22524), 
        .Y(n27021) );
  sky130_fd_sc_hd__clkbuf_1 U18468 ( .A(j202_soc_core_j22_cpu_ml_bufa[22]), 
        .X(n25627) );
  sky130_fd_sc_hd__buf_4 U18469 ( .A(j202_soc_core_j22_cpu_ml_bufa[15]), .X(
        n18887) );
  sky130_fd_sc_hd__and2_1 U18470 ( .A(n21706), .B(n21705), .X(n24353) );
  sky130_fd_sc_hd__a21oi_1 U18471 ( .A1(n22908), .A2(n16523), .B1(n15894), .Y(
        n26276) );
  sky130_fd_sc_hd__clkinv_1 U18472 ( .A(n29483), .Y(n28910) );
  sky130_fd_sc_hd__nand2_1 U18473 ( .A(n23847), .B(n23846), .Y(n27841) );
  sky130_fd_sc_hd__inv_2 U18474 ( .A(n27841), .Y(n24712) );
  sky130_fd_sc_hd__inv_2 U18475 ( .A(n25981), .Y(n27836) );
  sky130_fd_sc_hd__nand2_1 U18477 ( .A(n22415), .B(n22416), .Y(n27645) );
  sky130_fd_sc_hd__inv_1 U18478 ( .A(n27775), .Y(n27862) );
  sky130_fd_sc_hd__clkinv_1 U18479 ( .A(n27774), .Y(n27861) );
  sky130_fd_sc_hd__clkinv_1 U18480 ( .A(n28512), .Y(n28533) );
  sky130_fd_sc_hd__clkinv_1 U18481 ( .A(n28491), .Y(n28539) );
  sky130_fd_sc_hd__nand2_1 U18482 ( .A(n13328), .B(n13075), .Y(n28538) );
  sky130_fd_sc_hd__clkinv_1 U18483 ( .A(n12690), .Y(n18814) );
  sky130_fd_sc_hd__nand2_1 U18484 ( .A(n22394), .B(n22393), .Y(n27462) );
  sky130_fd_sc_hd__inv_2 U18485 ( .A(n28453), .Y(n25556) );
  sky130_fd_sc_hd__clkinv_1 U18487 ( .A(n27858), .Y(n25963) );
  sky130_fd_sc_hd__nand3_1 U18488 ( .A(n24176), .B(
        j202_soc_core_j22_cpu_regop_We__3_), .C(n24771), .Y(n27858) );
  sky130_fd_sc_hd__buf_4 U18489 ( .A(n24770), .X(n24778) );
  sky130_fd_sc_hd__buf_2 U18490 ( .A(n12822), .X(n12821) );
  sky130_fd_sc_hd__clkinv_1 U18491 ( .A(n25555), .Y(n25420) );
  sky130_fd_sc_hd__inv_2 U18493 ( .A(n28501), .Y(n27433) );
  sky130_fd_sc_hd__clkbuf_1 U18494 ( .A(n27896), .X(n12181) );
  sky130_fd_sc_hd__clkinv_1 U18495 ( .A(n25468), .Y(n25461) );
  sky130_fd_sc_hd__nand2_1 U18497 ( .A(n22405), .B(n22404), .Y(n27153) );
  sky130_fd_sc_hd__inv_2 U18498 ( .A(j202_soc_core_intc_core_00_rg_ipr[13]), 
        .Y(n25162) );
  sky130_fd_sc_hd__clkinv_1 U18499 ( .A(n27848), .Y(n26071) );
  sky130_fd_sc_hd__nor2_1 U18500 ( .A(n25094), .B(n25095), .Y(n28320) );
  sky130_fd_sc_hd__nor2_1 U18501 ( .A(n25098), .B(n25095), .Y(n28331) );
  sky130_fd_sc_hd__nor2_1 U18502 ( .A(n29088), .B(n28231), .Y(n28321) );
  sky130_fd_sc_hd__nor2_1 U18503 ( .A(n25094), .B(n25097), .Y(n28329) );
  sky130_fd_sc_hd__nor2_1 U18504 ( .A(n29088), .B(n25096), .Y(n28323) );
  sky130_fd_sc_hd__clkinv_1 U18505 ( .A(n28861), .Y(n28731) );
  sky130_fd_sc_hd__inv_2 U18506 ( .A(n24695), .Y(n24700) );
  sky130_fd_sc_hd__clkinv_1 U18507 ( .A(n29550), .Y(n23623) );
  sky130_fd_sc_hd__nand3_1 U18508 ( .A(n12461), .B(n21043), .C(n21044), .Y(
        n21046) );
  sky130_fd_sc_hd__inv_1 U18509 ( .A(n29441), .Y(n21044) );
  sky130_fd_sc_hd__clkinv_1 U18510 ( .A(n28734), .Y(n28887) );
  sky130_fd_sc_hd__clkinv_1 U18511 ( .A(n28865), .Y(n28843) );
  sky130_fd_sc_hd__and2_0 U18512 ( .A(n21175), .B(n21919), .X(n12111) );
  sky130_fd_sc_hd__and2_0 U18513 ( .A(n20719), .B(n21917), .X(n12123) );
  sky130_fd_sc_hd__and2_0 U18514 ( .A(n21335), .B(n21919), .X(n12112) );
  sky130_fd_sc_hd__clkinv_1 U18515 ( .A(n23949), .Y(n12327) );
  sky130_fd_sc_hd__nand3_2 U18516 ( .A(n13723), .B(n13722), .C(n12091), .Y(
        n28515) );
  sky130_fd_sc_hd__nand2_1 U18517 ( .A(n21242), .B(n16523), .Y(n13723) );
  sky130_fd_sc_hd__clkinv_1 U18518 ( .A(n11144), .Y(n12354) );
  sky130_fd_sc_hd__clkinv_1 U18520 ( .A(n27717), .Y(n24467) );
  sky130_fd_sc_hd__nand2_1 U18521 ( .A(n19311), .B(n19310), .Y(n27773) );
  sky130_fd_sc_hd__nor2b_1 U18523 ( .B_N(n26911), .A(n26904), .Y(n29390) );
  sky130_fd_sc_hd__clkinv_1 U18524 ( .A(n28257), .Y(n29394) );
  sky130_fd_sc_hd__clkinv_1 U18525 ( .A(n29311), .Y(n29392) );
  sky130_fd_sc_hd__clkinv_1 U18526 ( .A(n28254), .Y(n29389) );
  sky130_fd_sc_hd__clkinv_1 U18527 ( .A(n29310), .Y(n29393) );
  sky130_fd_sc_hd__nor2_1 U18528 ( .A(n26906), .B(n26905), .Y(n29391) );
  sky130_fd_sc_hd__inv_2 U18529 ( .A(n28360), .Y(n28405) );
  sky130_fd_sc_hd__clkinv_1 U18530 ( .A(n24513), .Y(n24514) );
  sky130_fd_sc_hd__clkinv_1 U18532 ( .A(n24507), .Y(n24508) );
  sky130_fd_sc_hd__clkinv_1 U18533 ( .A(n24500), .Y(n24501) );
  sky130_fd_sc_hd__clkinv_1 U18534 ( .A(n12467), .Y(n24499) );
  sky130_fd_sc_hd__clkinv_1 U18536 ( .A(n24483), .Y(n24484) );
  sky130_fd_sc_hd__clkinv_1 U18537 ( .A(n24481), .Y(n24482) );
  sky130_fd_sc_hd__clkinv_1 U18538 ( .A(n24477), .Y(n24478) );
  sky130_fd_sc_hd__and2_0 U18540 ( .A(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[0]), .B(n23898), .X(io_out[10]) );
  sky130_fd_sc_hd__and2_0 U18541 ( .A(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[1]), .B(n23898), .X(io_out[11]) );
  sky130_fd_sc_hd__and2_1 U18542 ( .A(n28078), .B(n28394), .X(n12151) );
  sky130_fd_sc_hd__and2_0 U18543 ( .A(n24277), .B(n24276), .X(n29744) );
  sky130_fd_sc_hd__inv_1 U18544 ( .A(n24384), .Y(n29497) );
  sky130_fd_sc_hd__buf_2 U18545 ( .A(n10714), .X(n29824) );
  sky130_fd_sc_hd__and2_0 U18546 ( .A(n26900), .B(n24274), .X(n29743) );
  sky130_fd_sc_hd__clkinv_1 U18547 ( .A(j202_soc_core_intc_core_00_rg_ie[29]), 
        .Y(n25489) );
  sky130_fd_sc_hd__and2_0 U18548 ( .A(j202_soc_core_uart_TOP_hold_reg[1]), .B(
        n29300), .X(j202_soc_core_uart_TOP_N25) );
  sky130_fd_sc_hd__and2_0 U18549 ( .A(j202_soc_core_uart_TOP_tx_bit_cnt[0]), 
        .B(j202_soc_core_uart_TOP_tx_bit_cnt[1]), .X(n24263) );
  sky130_fd_sc_hd__nand4bb_1 U18550 ( .A_N(
        j202_soc_core_uart_TOP_tx_bit_cnt[1]), .B_N(
        j202_soc_core_uart_TOP_tx_bit_cnt[2]), .C(
        j202_soc_core_uart_TOP_tx_bit_cnt[0]), .D(
        j202_soc_core_uart_TOP_tx_bit_cnt[3]), .Y(j202_soc_core_uart_TOP_N123)
         );
  sky130_fd_sc_hd__clkinv_1 U18551 ( .A(j202_soc_core_uart_TOP_tx_fifo_gb), 
        .Y(n28585) );
  sky130_fd_sc_hd__and2_0 U18552 ( .A(n28589), .B(n29173), .X(n10949) );
  sky130_fd_sc_hd__and2_0 U18553 ( .A(n24273), .B(n29172), .X(n29742) );
  sky130_fd_sc_hd__o21a_1 U18554 ( .A1(n23018), .A2(n25391), .B1(n23017), .X(
        n23046) );
  sky130_fd_sc_hd__clkinv_1 U18555 ( .A(j202_soc_core_intc_core_00_rg_ipr[41]), 
        .Y(n26733) );
  sky130_fd_sc_hd__clkinv_1 U18556 ( .A(j202_soc_core_intc_core_00_rg_ipr[105]), .Y(n27935) );
  sky130_fd_sc_hd__clkinv_1 U18557 ( .A(j202_soc_core_intc_core_00_rg_ie[25]), 
        .Y(n27168) );
  sky130_fd_sc_hd__clkinv_1 U18558 ( .A(j202_soc_core_intc_core_00_rg_ipr[113]), .Y(n25744) );
  sky130_fd_sc_hd__clkinv_1 U18559 ( .A(j202_soc_core_intc_core_00_rg_ipr[115]), .Y(n25322) );
  sky130_fd_sc_hd__clkinv_1 U18560 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[100]), .Y(n25320) );
  sky130_fd_sc_hd__clkinv_1 U18561 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[108]), .Y(n25321) );
  sky130_fd_sc_hd__clkinv_1 U18562 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[116]), .Y(n25326) );
  sky130_fd_sc_hd__clkinv_1 U18563 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[124]), .Y(n25327) );
  sky130_fd_sc_hd__clkinv_1 U18564 ( .A(j202_soc_core_intc_core_00_rg_ipr[112]), .Y(n27097) );
  sky130_fd_sc_hd__clkinv_1 U18565 ( .A(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_), .Y(n27699) );
  sky130_fd_sc_hd__clkinv_1 U18566 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[119]), .Y(n27599) );
  sky130_fd_sc_hd__clkinv_1 U18567 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[118]), .Y(n27076) );
  sky130_fd_sc_hd__clkinv_1 U18568 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[115]), .Y(n26125) );
  sky130_fd_sc_hd__clkinv_1 U18569 ( .A(j202_soc_core_intc_core_00_rg_itgt[83]), .Y(n26884) );
  sky130_fd_sc_hd__clkinv_1 U18570 ( .A(j202_soc_core_intc_core_00_rg_itgt[51]), .Y(n25792) );
  sky130_fd_sc_hd__clkinv_1 U18571 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[114]), .Y(n27004) );
  sky130_fd_sc_hd__clkinv_1 U18572 ( .A(j202_soc_core_intc_core_00_rg_itgt[82]), .Y(n25078) );
  sky130_fd_sc_hd__clkinv_1 U18573 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[113]), .Y(n27562) );
  sky130_fd_sc_hd__clkinv_1 U18574 ( .A(j202_soc_core_intc_core_00_rg_itgt[81]), .Y(n27449) );
  sky130_fd_sc_hd__clkinv_1 U18575 ( .A(j202_soc_core_intc_core_00_rg_itgt[49]), .Y(n27413) );
  sky130_fd_sc_hd__clkinv_1 U18576 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[112]), .Y(n27685) );
  sky130_fd_sc_hd__clkinv_1 U18577 ( .A(j202_soc_core_intc_core_00_rg_itgt[48]), .Y(n29081) );
  sky130_fd_sc_hd__clkinv_1 U18578 ( .A(j202_soc_core_intc_core_00_rg_itgt[23]), .Y(n27396) );
  sky130_fd_sc_hd__clkinv_1 U18579 ( .A(j202_soc_core_intc_core_00_rg_itgt[22]), .Y(n27657) );
  sky130_fd_sc_hd__clkinv_1 U18580 ( .A(j202_soc_core_intc_core_00_rg_itgt[21]), .Y(n27370) );
  sky130_fd_sc_hd__clkinv_1 U18581 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[111]), .Y(n27595) );
  sky130_fd_sc_hd__clkinv_1 U18582 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[110]), .Y(n27072) );
  sky130_fd_sc_hd__clkinv_1 U18583 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[107]), .Y(n26120) );
  sky130_fd_sc_hd__clkinv_1 U18584 ( .A(j202_soc_core_intc_core_00_rg_itgt[75]), .Y(n26881) );
  sky130_fd_sc_hd__clkinv_1 U18585 ( .A(j202_soc_core_intc_core_00_rg_itgt[43]), .Y(n25788) );
  sky130_fd_sc_hd__clkinv_1 U18586 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[106]), .Y(n27002) );
  sky130_fd_sc_hd__clkinv_1 U18587 ( .A(j202_soc_core_intc_core_00_rg_itgt[74]), .Y(n25065) );
  sky130_fd_sc_hd__clkinv_1 U18588 ( .A(j202_soc_core_intc_core_00_rg_itgt[73]), .Y(n27447) );
  sky130_fd_sc_hd__clkinv_1 U18589 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[104]), .Y(n27682) );
  sky130_fd_sc_hd__clkinv_1 U18590 ( .A(j202_soc_core_intc_core_00_rg_itgt[40]), .Y(n28312) );
  sky130_fd_sc_hd__clkinv_1 U18591 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[127]), .Y(n27600) );
  sky130_fd_sc_hd__clkinv_1 U18592 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[126]), .Y(n27077) );
  sky130_fd_sc_hd__clkinv_1 U18593 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[123]), .Y(n26126) );
  sky130_fd_sc_hd__clkinv_1 U18594 ( .A(j202_soc_core_intc_core_00_rg_itgt[91]), .Y(n26885) );
  sky130_fd_sc_hd__clkinv_1 U18595 ( .A(j202_soc_core_intc_core_00_rg_itgt[59]), .Y(n25793) );
  sky130_fd_sc_hd__clkinv_1 U18596 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[122]), .Y(n27005) );
  sky130_fd_sc_hd__clkinv_1 U18597 ( .A(j202_soc_core_intc_core_00_rg_itgt[90]), .Y(n25080) );
  sky130_fd_sc_hd__clkinv_1 U18598 ( .A(j202_soc_core_intc_core_00_rg_itgt[89]), .Y(n27451) );
  sky130_fd_sc_hd__clkinv_1 U18599 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[120]), .Y(n27687) );
  sky130_fd_sc_hd__clkinv_1 U18600 ( .A(j202_soc_core_intc_core_00_rg_itgt[56]), .Y(n29075) );
  sky130_fd_sc_hd__clkinv_1 U18601 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[103]), .Y(n27594) );
  sky130_fd_sc_hd__clkinv_1 U18602 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[102]), .Y(n27071) );
  sky130_fd_sc_hd__clkinv_1 U18603 ( .A(j202_soc_core_intc_core_00_rg_itgt[99]), .Y(n26119) );
  sky130_fd_sc_hd__clkinv_1 U18604 ( .A(j202_soc_core_intc_core_00_rg_itgt[67]), .Y(n26880) );
  sky130_fd_sc_hd__clkinv_1 U18605 ( .A(j202_soc_core_intc_core_00_rg_itgt[35]), .Y(n25787) );
  sky130_fd_sc_hd__clkinv_1 U18606 ( .A(j202_soc_core_intc_core_00_rg_itgt[98]), .Y(n27001) );
  sky130_fd_sc_hd__clkinv_1 U18607 ( .A(j202_soc_core_intc_core_00_rg_itgt[66]), .Y(n25060) );
  sky130_fd_sc_hd__clkinv_1 U18608 ( .A(j202_soc_core_intc_core_00_rg_itgt[97]), .Y(n27559) );
  sky130_fd_sc_hd__clkinv_1 U18609 ( .A(j202_soc_core_intc_core_00_rg_itgt[65]), .Y(n27446) );
  sky130_fd_sc_hd__clkinv_1 U18610 ( .A(j202_soc_core_intc_core_00_rg_itgt[33]), .Y(n27410) );
  sky130_fd_sc_hd__clkinv_1 U18611 ( .A(j202_soc_core_intc_core_00_rg_itgt[96]), .Y(n27681) );
  sky130_fd_sc_hd__clkinv_1 U18612 ( .A(j202_soc_core_intc_core_00_rg_itgt[32]), .Y(n28309) );
  sky130_fd_sc_hd__clkinv_1 U18613 ( .A(j202_soc_core_intc_core_00_rg_ipr[62]), 
        .Y(n26741) );
  sky130_fd_sc_hd__clkinv_1 U18614 ( .A(j202_soc_core_intc_core_00_rg_ipr[46]), 
        .Y(n26731) );
  sky130_fd_sc_hd__clkinv_1 U18615 ( .A(j202_soc_core_intc_core_00_rg_ipr[33]), 
        .Y(n26725) );
  sky130_fd_sc_hd__clkinv_1 U18616 ( .A(j202_soc_core_intc_core_00_rg_ipr[127]), .Y(n27596) );
  sky130_fd_sc_hd__clkinv_1 U18617 ( .A(j202_soc_core_intc_core_00_rg_ipr[126]), .Y(n27997) );
  sky130_fd_sc_hd__clkinv_1 U18618 ( .A(j202_soc_core_intc_core_00_rg_ipr[123]), .Y(n27073) );
  sky130_fd_sc_hd__clkinv_1 U18619 ( .A(j202_soc_core_intc_core_00_rg_ipr[120]), .Y(n27652) );
  sky130_fd_sc_hd__clkinv_1 U18620 ( .A(j202_soc_core_intc_core_00_rg_ipr[119]), .Y(n27628) );
  sky130_fd_sc_hd__clkinv_1 U18621 ( .A(j202_soc_core_intc_core_00_rg_ipr[116]), .Y(n27368) );
  sky130_fd_sc_hd__clkinv_1 U18622 ( .A(j202_soc_core_intc_core_00_rg_ipr[114]), .Y(n27131) );
  sky130_fd_sc_hd__clkinv_1 U18623 ( .A(j202_soc_core_intc_core_00_rg_ipr[111]), .Y(n26121) );
  sky130_fd_sc_hd__clkinv_1 U18624 ( .A(j202_soc_core_intc_core_00_rg_ipr[110]), .Y(n26882) );
  sky130_fd_sc_hd__clkinv_1 U18625 ( .A(j202_soc_core_intc_core_00_rg_ipr[109]), .Y(n25789) );
  sky130_fd_sc_hd__clkinv_1 U18626 ( .A(j202_soc_core_intc_core_00_rg_ipr[107]), .Y(n27003) );
  sky130_fd_sc_hd__clkinv_1 U18627 ( .A(j202_soc_core_intc_core_00_rg_ipr[106]), .Y(n25067) );
  sky130_fd_sc_hd__clkinv_1 U18628 ( .A(j202_soc_core_intc_core_00_rg_ipr[104]), .Y(n27969) );
  sky130_fd_sc_hd__clkinv_1 U18629 ( .A(j202_soc_core_intc_core_00_rg_ipr[102]), .Y(n27448) );
  sky130_fd_sc_hd__clkinv_1 U18630 ( .A(j202_soc_core_intc_core_00_rg_ipr[100]), .Y(n27496) );
  sky130_fd_sc_hd__clkinv_1 U18631 ( .A(j202_soc_core_intc_core_00_rg_ipr[99]), 
        .Y(n27683) );
  sky130_fd_sc_hd__clkinv_1 U18632 ( .A(j202_soc_core_intc_core_00_rg_ipr[97]), 
        .Y(n28315) );
  sky130_fd_sc_hd__clkinv_1 U18633 ( .A(j202_soc_core_intc_core_00_rg_ipr[96]), 
        .Y(n28229) );
  sky130_fd_sc_hd__clkinv_1 U18634 ( .A(j202_soc_core_intc_core_00_rg_ie[31]), 
        .Y(n27597) );
  sky130_fd_sc_hd__clkinv_1 U18635 ( .A(j202_soc_core_intc_core_00_rg_ie[30]), 
        .Y(n27998) );
  sky130_fd_sc_hd__clkinv_1 U18636 ( .A(j202_soc_core_intc_core_00_rg_ie[28]), 
        .Y(n27393) );
  sky130_fd_sc_hd__clkinv_1 U18637 ( .A(j202_soc_core_intc_core_00_rg_ie[27]), 
        .Y(n27074) );
  sky130_fd_sc_hd__clkinv_1 U18638 ( .A(j202_soc_core_intc_core_00_rg_ie[24]), 
        .Y(n27653) );
  sky130_fd_sc_hd__clkinv_1 U18639 ( .A(j202_soc_core_intc_core_00_rg_ie[23]), 
        .Y(n27629) );
  sky130_fd_sc_hd__clkinv_1 U18640 ( .A(j202_soc_core_intc_core_00_rg_ie[22]), 
        .Y(n25609) );
  sky130_fd_sc_hd__clkinv_1 U18641 ( .A(j202_soc_core_intc_core_00_rg_ie[21]), 
        .Y(n25577) );
  sky130_fd_sc_hd__clkinv_1 U18642 ( .A(j202_soc_core_intc_core_00_rg_eimk[2]), 
        .Y(n28184) );
  sky130_fd_sc_hd__clkinv_1 U18643 ( .A(n27091), .Y(n12532) );
  sky130_fd_sc_hd__nand3_1 U18644 ( .A(n21186), .B(n21185), .C(n21184), .Y(
        n29549) );
  sky130_fd_sc_hd__and2_0 U18645 ( .A(n28026), .B(
        j202_soc_core_wbqspiflash_00_spi_out[26]), .X(n29683) );
  sky130_fd_sc_hd__and2_0 U18646 ( .A(n28026), .B(
        j202_soc_core_wbqspiflash_00_spi_out[25]), .X(n29684) );
  sky130_fd_sc_hd__and2_0 U18647 ( .A(n28026), .B(
        j202_soc_core_wbqspiflash_00_spi_out[24]), .X(n29685) );
  sky130_fd_sc_hd__and2_0 U18648 ( .A(n28026), .B(
        j202_soc_core_wbqspiflash_00_spi_out[23]), .X(n29686) );
  sky130_fd_sc_hd__and2_0 U18649 ( .A(n28026), .B(
        j202_soc_core_wbqspiflash_00_spi_out[22]), .X(n29687) );
  sky130_fd_sc_hd__and2_0 U18650 ( .A(n28026), .B(
        j202_soc_core_wbqspiflash_00_spi_out[13]), .X(n29688) );
  sky130_fd_sc_hd__and2_0 U18651 ( .A(n28026), .B(
        j202_soc_core_wbqspiflash_00_spi_out[12]), .X(n29689) );
  sky130_fd_sc_hd__and2_0 U18652 ( .A(n28026), .B(
        j202_soc_core_wbqspiflash_00_spi_out[11]), .X(n29690) );
  sky130_fd_sc_hd__and2_0 U18653 ( .A(n28026), .B(
        j202_soc_core_wbqspiflash_00_spi_out[10]), .X(n29691) );
  sky130_fd_sc_hd__and2_0 U18654 ( .A(n28026), .B(
        j202_soc_core_wbqspiflash_00_spi_out[9]), .X(n29692) );
  sky130_fd_sc_hd__and2_0 U18655 ( .A(n28026), .B(
        j202_soc_core_wbqspiflash_00_spi_out[8]), .X(n29693) );
  sky130_fd_sc_hd__and2_1 U18658 ( .A(n27119), .B(n23572), .X(n13079) );
  sky130_fd_sc_hd__and2_1 U18659 ( .A(n27119), .B(n23564), .X(n13081) );
  sky130_fd_sc_hd__and2_1 U18661 ( .A(n27119), .B(n23575), .X(n13095) );
  sky130_fd_sc_hd__nand3_1 U18662 ( .A(n12204), .B(n27118), .C(n27119), .Y(
        n29844) );
  sky130_fd_sc_hd__and2_0 U18663 ( .A(n29169), .B(n24267), .X(n29732) );
  sky130_fd_sc_hd__and2_0 U18664 ( .A(n29169), .B(n24270), .X(n29733) );
  sky130_fd_sc_hd__o22ai_1 U18665 ( .A1(n25982), .A2(n27897), .B1(n27837), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N3040) );
  sky130_fd_sc_hd__and2_1 U18666 ( .A(j202_soc_core_j22_cpu_ml_N428), .B(
        n28441), .X(n29650) );
  sky130_fd_sc_hd__clkinv_1 U18668 ( .A(n12035), .Y(n12340) );
  sky130_fd_sc_hd__nor3_1 U18669 ( .A(n23643), .B(n24651), .C(n23642), .Y(
        n29879) );
  sky130_fd_sc_hd__clkinv_1 U18670 ( .A(n12037), .Y(n12339) );
  sky130_fd_sc_hd__a21oi_1 U18671 ( .A1(n27344), .A2(n12088), .B1(n29583), .Y(
        n12709) );
  sky130_fd_sc_hd__nand3_1 U18672 ( .A(n12703), .B(n27344), .C(n12157), .Y(
        n12705) );
  sky130_fd_sc_hd__a21boi_1 U18674 ( .A1(n21290), .A2(n27717), .B1_N(n21304), 
        .Y(n12408) );
  sky130_fd_sc_hd__nand3_1 U18675 ( .A(n21018), .B(n21017), .C(n21016), .Y(
        n29547) );
  sky130_fd_sc_hd__nand3_1 U18676 ( .A(n24594), .B(n24600), .C(n24599), .Y(
        n24601) );
  sky130_fd_sc_hd__and2_0 U18677 ( .A(n25340), .B(n26548), .X(n23636) );
  sky130_fd_sc_hd__clkinv_1 U18679 ( .A(n13033), .Y(n29444) );
  sky130_fd_sc_hd__clkbuf_1 U18680 ( .A(n21056), .X(n29747) );
  sky130_fd_sc_hd__and2_0 U18681 ( .A(n24259), .B(
        j202_soc_core_intc_core_00_rg_ie[16]), .X(n29722) );
  sky130_fd_sc_hd__clkinv_1 U18682 ( .A(n24726), .Y(n24727) );
  sky130_fd_sc_hd__clkinv_1 U18683 ( .A(n26502), .Y(n23880) );
  sky130_fd_sc_hd__clkinv_1 U18684 ( .A(n12877), .Y(n12876) );
  sky130_fd_sc_hd__nand2_1 U18685 ( .A(n24039), .B(n23893), .Y(n29748) );
  sky130_fd_sc_hd__clkbuf_1 U18686 ( .A(n10711), .X(n29826) );
  sky130_fd_sc_hd__nor2_1 U18688 ( .A(j202_soc_core_aquc_WE_), .B(n25033), .Y(
        n29435) );
  sky130_fd_sc_hd__clkinv_1 U18689 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[6]), .Y(n12298) );
  sky130_fd_sc_hd__and2_0 U18690 ( .A(n24201), .B(n24520), .X(n29694) );
  sky130_fd_sc_hd__and2_0 U18691 ( .A(n29745), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]), .X(n29728) );
  sky130_fd_sc_hd__clkinv_1 U18692 ( .A(la_oenb[31]), .Y(n24184) );
  sky130_fd_sc_hd__clkinv_1 U18693 ( .A(la_oenb[30]), .Y(n24185) );
  sky130_fd_sc_hd__clkinv_1 U18694 ( .A(la_oenb[29]), .Y(n24186) );
  sky130_fd_sc_hd__clkinv_1 U18695 ( .A(la_oenb[28]), .Y(n24187) );
  sky130_fd_sc_hd__clkinv_1 U18696 ( .A(la_oenb[27]), .Y(n24188) );
  sky130_fd_sc_hd__clkinv_1 U18697 ( .A(la_oenb[26]), .Y(n24189) );
  sky130_fd_sc_hd__clkinv_1 U18698 ( .A(la_oenb[25]), .Y(n24190) );
  sky130_fd_sc_hd__clkinv_1 U18699 ( .A(la_oenb[24]), .Y(n24191) );
  sky130_fd_sc_hd__clkinv_1 U18700 ( .A(la_oenb[23]), .Y(n24192) );
  sky130_fd_sc_hd__clkinv_1 U18701 ( .A(la_oenb[22]), .Y(n24193) );
  sky130_fd_sc_hd__clkinv_1 U18702 ( .A(la_oenb[21]), .Y(n24194) );
  sky130_fd_sc_hd__clkinv_1 U18703 ( .A(la_oenb[20]), .Y(n24195) );
  sky130_fd_sc_hd__clkinv_1 U18704 ( .A(la_oenb[19]), .Y(n24196) );
  sky130_fd_sc_hd__clkinv_1 U18705 ( .A(la_oenb[18]), .Y(n24197) );
  sky130_fd_sc_hd__clkinv_1 U18706 ( .A(la_oenb[17]), .Y(n24198) );
  sky130_fd_sc_hd__and2_0 U18707 ( .A(io_in[35]), .B(n29830), .X(n29668) );
  sky130_fd_sc_hd__and2_0 U18708 ( .A(io_in[31]), .B(n29830), .X(n29632) );
  sky130_fd_sc_hd__and2_0 U18709 ( .A(io_in[2]), .B(n29745), .X(n29680) );
  sky130_fd_sc_hd__and2_0 U18710 ( .A(n29610), .B(wbs_dat_i[1]), .X(n13) );
  sky130_fd_sc_hd__and2_0 U18711 ( .A(n29610), .B(wbs_dat_i[2]), .X(n14) );
  sky130_fd_sc_hd__and2_0 U18712 ( .A(n29610), .B(wbs_dat_i[3]), .X(n15) );
  sky130_fd_sc_hd__and2_0 U18713 ( .A(n29610), .B(wbs_dat_i[4]), .X(n16) );
  sky130_fd_sc_hd__and2_0 U18714 ( .A(n29610), .B(wbs_dat_i[5]), .X(n17) );
  sky130_fd_sc_hd__and2_0 U18715 ( .A(n29610), .B(wbs_dat_i[6]), .X(n18) );
  sky130_fd_sc_hd__and2_0 U18716 ( .A(n29610), .B(wbs_dat_i[7]), .X(n19) );
  sky130_fd_sc_hd__and2_0 U18717 ( .A(n29610), .B(wbs_dat_i[8]), .X(n21) );
  sky130_fd_sc_hd__and2_0 U18718 ( .A(n24025), .B(wbs_dat_i[9]), .X(n220) );
  sky130_fd_sc_hd__and2_0 U18719 ( .A(n24025), .B(wbs_dat_i[10]), .X(n230) );
  sky130_fd_sc_hd__and2_0 U18720 ( .A(n24025), .B(wbs_dat_i[11]), .X(n240) );
  sky130_fd_sc_hd__and2_0 U18721 ( .A(n24025), .B(wbs_dat_i[12]), .X(n250) );
  sky130_fd_sc_hd__and2_0 U18722 ( .A(n24025), .B(wbs_dat_i[13]), .X(n260) );
  sky130_fd_sc_hd__and2_0 U18723 ( .A(n24025), .B(wbs_dat_i[14]), .X(n270) );
  sky130_fd_sc_hd__a31o_1 U18724 ( .A1(n29610), .A2(wbs_we_i), .A3(
        wbs_sel_i[1]), .B1(wb_rst_i), .X(n20) );
  sky130_fd_sc_hd__and2_0 U18725 ( .A(n24025), .B(wbs_dat_i[15]), .X(n280) );
  sky130_fd_sc_hd__and2_0 U18726 ( .A(n24025), .B(wbs_dat_i[16]), .X(n300) );
  sky130_fd_sc_hd__and2_0 U18727 ( .A(n24025), .B(wbs_dat_i[17]), .X(n310) );
  sky130_fd_sc_hd__and2_0 U18728 ( .A(n24025), .B(wbs_dat_i[18]), .X(n320) );
  sky130_fd_sc_hd__and2_0 U18729 ( .A(n24025), .B(wbs_dat_i[19]), .X(n330) );
  sky130_fd_sc_hd__and2_0 U18730 ( .A(n24025), .B(wbs_dat_i[20]), .X(n340) );
  sky130_fd_sc_hd__and2_0 U18731 ( .A(n29610), .B(wbs_dat_i[21]), .X(n350) );
  sky130_fd_sc_hd__and2_0 U18732 ( .A(n29610), .B(wbs_dat_i[22]), .X(n360) );
  sky130_fd_sc_hd__a31o_1 U18733 ( .A1(n29610), .A2(wbs_we_i), .A3(
        wbs_sel_i[2]), .B1(wb_rst_i), .X(n290) );
  sky130_fd_sc_hd__and2_0 U18734 ( .A(n29610), .B(wbs_dat_i[23]), .X(n370) );
  sky130_fd_sc_hd__and2_0 U18735 ( .A(n29610), .B(wbs_dat_i[24]), .X(n390) );
  sky130_fd_sc_hd__and2_0 U18736 ( .A(n24025), .B(wbs_dat_i[25]), .X(n400) );
  sky130_fd_sc_hd__and2_0 U18737 ( .A(n29610), .B(wbs_dat_i[26]), .X(n410) );
  sky130_fd_sc_hd__and2_0 U18738 ( .A(n29610), .B(wbs_dat_i[27]), .X(n420) );
  sky130_fd_sc_hd__and2_0 U18739 ( .A(n29610), .B(wbs_dat_i[28]), .X(n430) );
  sky130_fd_sc_hd__and2_0 U18740 ( .A(n29610), .B(wbs_dat_i[29]), .X(n440) );
  sky130_fd_sc_hd__and2_0 U18741 ( .A(n29610), .B(wbs_dat_i[30]), .X(n450) );
  sky130_fd_sc_hd__a31o_1 U18742 ( .A1(n29610), .A2(wbs_we_i), .A3(
        wbs_sel_i[3]), .B1(wb_rst_i), .X(n380) );
  sky130_fd_sc_hd__and2_0 U18743 ( .A(n29610), .B(wbs_dat_i[31]), .X(n460) );
  sky130_fd_sc_hd__clkbuf_1 U18744 ( .A(n24025), .X(n29610) );
  sky130_fd_sc_hd__inv_8 U18745 ( .A(n29760), .Y(n12387) );
  sky130_fd_sc_hd__inv_8 U18746 ( .A(n29758), .Y(n12376) );
  sky130_fd_sc_hd__inv_8 U18747 ( .A(n29757), .Y(n12382) );
  sky130_fd_sc_hd__inv_8 U18748 ( .A(n29755), .Y(n12378) );
  sky130_fd_sc_hd__inv_8 U18749 ( .A(n29759), .Y(n12309) );
  sky130_fd_sc_hd__inv_8 U18750 ( .A(n29756), .Y(n12305) );
  sky130_fd_sc_hd__inv_8 U18751 ( .A(n29759), .Y(n12308) );
  sky130_fd_sc_hd__inv_8 U18752 ( .A(n29756), .Y(n12304) );
  sky130_fd_sc_hd__inv_8 U18753 ( .A(n29760), .Y(n12388) );
  sky130_fd_sc_hd__inv_8 U18754 ( .A(n29759), .Y(n12385) );
  sky130_fd_sc_hd__inv_8 U18755 ( .A(n29756), .Y(n12381) );
  sky130_fd_sc_hd__clkinv_1 U18756 ( .A(n18805), .Y(n26414) );
  sky130_fd_sc_hd__inv_2 U18757 ( .A(n13796), .Y(n14985) );
  sky130_fd_sc_hd__inv_2 U18758 ( .A(n13796), .Y(n16447) );
  sky130_fd_sc_hd__inv_2 U18760 ( .A(j202_soc_core_intc_core_00_rg_ipr[48]), 
        .Y(n26739) );
  sky130_fd_sc_hd__clkinv_1 U18761 ( .A(n26414), .Y(n26926) );
  sky130_fd_sc_hd__clkinv_1 U18762 ( .A(n22678), .Y(n22929) );
  sky130_fd_sc_hd__o21ai_2 U18763 ( .A1(n24717), .A2(n23839), .B1(n27861), .Y(
        j202_soc_core_j22_cpu_rf_N3371) );
  sky130_fd_sc_hd__inv_4 U18764 ( .A(n19726), .Y(n19816) );
  sky130_fd_sc_hd__inv_2 U18765 ( .A(n24854), .Y(n22940) );
  sky130_fd_sc_hd__nor2_2 U18766 ( .A(n30011), .B(n14312), .Y(n14743) );
  sky130_fd_sc_hd__inv_2 U18767 ( .A(n13448), .Y(n14107) );
  sky130_fd_sc_hd__inv_2 U18768 ( .A(n14107), .Y(n15937) );
  sky130_fd_sc_hd__nand2_4 U18769 ( .A(n13364), .B(n13363), .Y(n13365) );
  sky130_fd_sc_hd__or2_2 U18770 ( .A(n14597), .B(n21088), .X(n12089) );
  sky130_fd_sc_hd__inv_2 U18772 ( .A(n14209), .Y(n16398) );
  sky130_fd_sc_hd__inv_2 U18773 ( .A(n14209), .Y(n15783) );
  sky130_fd_sc_hd__inv_2 U18774 ( .A(n13946), .Y(n16410) );
  sky130_fd_sc_hd__inv_2 U18775 ( .A(n13951), .Y(n16433) );
  sky130_fd_sc_hd__inv_2 U18776 ( .A(n13951), .Y(n15907) );
  sky130_fd_sc_hd__and4_1 U18778 ( .A(n13721), .B(n13720), .C(n13719), .D(
        n13718), .X(n12091) );
  sky130_fd_sc_hd__and4_1 U18779 ( .A(n13806), .B(n13805), .C(n13804), .D(
        n13803), .X(n12092) );
  sky130_fd_sc_hd__inv_2 U18780 ( .A(n13952), .Y(n16446) );
  sky130_fd_sc_hd__inv_2 U18781 ( .A(n14082), .Y(n16432) );
  sky130_fd_sc_hd__inv_2 U18782 ( .A(n14082), .Y(n14828) );
  sky130_fd_sc_hd__inv_2 U18783 ( .A(n14033), .Y(n16425) );
  sky130_fd_sc_hd__inv_2 U18784 ( .A(n14033), .Y(n14986) );
  sky130_fd_sc_hd__inv_2 U18785 ( .A(n13546), .Y(n13796) );
  sky130_fd_sc_hd__inv_2 U18786 ( .A(n14220), .Y(n15925) );
  sky130_fd_sc_hd__inv_2 U18787 ( .A(n14220), .Y(n16448) );
  sky130_fd_sc_hd__inv_2 U18788 ( .A(n29588), .Y(n12861) );
  sky130_fd_sc_hd__clkinv_1 U18789 ( .A(n20139), .Y(n12841) );
  sky130_fd_sc_hd__a21o_1 U18790 ( .A1(n25473), .A2(n17225), .B1(n16099), .X(
        n12094) );
  sky130_fd_sc_hd__and4_1 U18791 ( .A(n14086), .B(n14085), .C(n14084), .D(
        n14083), .X(n12095) );
  sky130_fd_sc_hd__and4_1 U18792 ( .A(n14425), .B(n14424), .C(n14423), .D(
        n14422), .X(n12096) );
  sky130_fd_sc_hd__and4_1 U18793 ( .A(n13473), .B(n13472), .C(n13471), .D(
        n13470), .X(n12097) );
  sky130_fd_sc_hd__and4_1 U18794 ( .A(n14925), .B(n14924), .C(n14923), .D(
        n14922), .X(n12100) );
  sky130_fd_sc_hd__and4_1 U18795 ( .A(n13440), .B(n13439), .C(n13438), .D(
        n13437), .X(n12101) );
  sky130_fd_sc_hd__o211a_2 U18796 ( .A1(n13512), .A2(n16444), .B1(n13511), 
        .C1(n13510), .X(n12102) );
  sky130_fd_sc_hd__and4_1 U18797 ( .A(n14997), .B(n14996), .C(n14995), .D(
        n14994), .X(n12103) );
  sky130_fd_sc_hd__and4_1 U18798 ( .A(n14942), .B(n14941), .C(n14940), .D(
        n14939), .X(n12104) );
  sky130_fd_sc_hd__and4_1 U18799 ( .A(n14447), .B(n14446), .C(n14445), .D(
        n14444), .X(n12105) );
  sky130_fd_sc_hd__and4_1 U18800 ( .A(n14502), .B(n14501), .C(n14500), .D(
        n14499), .X(n12106) );
  sky130_fd_sc_hd__clkinv_1 U18801 ( .A(n13054), .Y(n24791) );
  sky130_fd_sc_hd__clkinv_1 U18802 ( .A(n29553), .Y(n24818) );
  sky130_fd_sc_hd__clkinv_1 U18803 ( .A(n29557), .Y(n24817) );
  sky130_fd_sc_hd__clkinv_1 U18804 ( .A(n29556), .Y(n25035) );
  sky130_fd_sc_hd__clkinv_1 U18805 ( .A(n29545), .Y(n25053) );
  sky130_fd_sc_hd__clkinv_1 U18806 ( .A(n29554), .Y(n25054) );
  sky130_fd_sc_hd__clkinv_1 U18807 ( .A(n29555), .Y(n25036) );
  sky130_fd_sc_hd__clkinv_1 U18808 ( .A(n29552), .Y(n27951) );
  sky130_fd_sc_hd__clkinv_1 U18809 ( .A(n29548), .Y(n25051) );
  sky130_fd_sc_hd__o211a_1 U18810 ( .A1(n26926), .A2(n26866), .B1(n25960), 
        .C1(n25959), .X(n12113) );
  sky130_fd_sc_hd__and4_1 U18811 ( .A(n14068), .B(n14067), .C(n14066), .D(
        n14065), .X(n12114) );
  sky130_fd_sc_hd__and4_1 U18812 ( .A(n15911), .B(n15910), .C(n15909), .D(
        n15908), .X(n12119) );
  sky130_fd_sc_hd__and4_1 U18813 ( .A(n13881), .B(n13880), .C(n13879), .D(
        n13878), .X(n12120) );
  sky130_fd_sc_hd__o211a_2 U18814 ( .A1(n27027), .A2(n11186), .B1(n15486), 
        .C1(n15485), .X(n12121) );
  sky130_fd_sc_hd__and4_1 U18815 ( .A(n19687), .B(n19677), .C(n19676), .D(
        n19685), .X(n12122) );
  sky130_fd_sc_hd__and2_1 U18816 ( .A(n19851), .B(n21917), .X(n12124) );
  sky130_fd_sc_hd__and4_1 U18817 ( .A(n19229), .B(n19228), .C(n19215), .D(
        n19226), .X(n12126) );
  sky130_fd_sc_hd__and4_1 U18818 ( .A(n19413), .B(n19412), .C(n19421), .D(
        n19423), .X(n12137) );
  sky130_fd_sc_hd__a21boi_1 U18819 ( .A1(n27362), .A2(n27361), .B1_N(n27360), 
        .Y(n27363) );
  sky130_fd_sc_hd__and2_1 U18821 ( .A(n27093), .B(n29553), .X(n12144) );
  sky130_fd_sc_hd__and2_1 U18822 ( .A(n27093), .B(n29557), .X(n12145) );
  sky130_fd_sc_hd__and2_1 U18823 ( .A(n27093), .B(n29545), .X(n12146) );
  sky130_fd_sc_hd__and2_1 U18824 ( .A(n27093), .B(n29554), .X(n12147) );
  sky130_fd_sc_hd__and2_1 U18826 ( .A(n27093), .B(n29555), .X(n12149) );
  sky130_fd_sc_hd__nand2_1 U18827 ( .A(n30025), .B(n21915), .Y(n29501) );
  sky130_fd_sc_hd__nand3_2 U18828 ( .A(n27721), .B(n23046), .C(n23045), .Y(
        n29517) );
  sky130_fd_sc_hd__or2b_4 U18829 ( .A(n29603), .B_N(n29745), .X(n23851) );
  sky130_fd_sc_hd__clkinv_1 U18830 ( .A(n27847), .Y(n25964) );
  sky130_fd_sc_hd__clkinv_1 U18831 ( .A(j202_soc_core_j22_cpu_macop_MAC_[0]), 
        .Y(n27828) );
  sky130_fd_sc_hd__clkinv_1 U18832 ( .A(n27828), .Y(n27052) );
  sky130_fd_sc_hd__nand2_1 U18834 ( .A(n27858), .B(n24681), .Y(n27859) );
  sky130_fd_sc_hd__nand2b_1 U18836 ( .A_N(n24613), .B(n20427), .Y(n28379) );
  sky130_fd_sc_hd__buf_4 U18839 ( .A(j202_soc_core_j22_cpu_ml_bufa[19]), .X(
        n22811) );
  sky130_fd_sc_hd__clkinv_1 U18840 ( .A(n27355), .Y(n27152) );
  sky130_fd_sc_hd__clkinv_1 U18841 ( .A(n27711), .Y(n29583) );
  sky130_fd_sc_hd__clkinv_1 U18842 ( .A(j202_soc_core_intc_core_00_rg_ipr[54]), 
        .Y(n12697) );
  sky130_fd_sc_hd__clkinv_1 U18843 ( .A(j202_soc_core_intc_core_00_rg_ipr[52]), 
        .Y(n12695) );
  sky130_fd_sc_hd__nand2_1 U18844 ( .A(n12161), .B(n12160), .Y(n17886) );
  sky130_fd_sc_hd__nand2_1 U18845 ( .A(n17917), .B(n17916), .Y(n12160) );
  sky130_fd_sc_hd__o21ai_1 U18846 ( .A1(n17916), .A2(n17917), .B1(n12163), .Y(
        n12161) );
  sky130_fd_sc_hd__xnor2_1 U18847 ( .A(n17917), .B(n12162), .Y(n17971) );
  sky130_fd_sc_hd__xnor2_1 U18848 ( .A(n12163), .B(n17916), .Y(n12162) );
  sky130_fd_sc_hd__nand2_1 U18849 ( .A(n12165), .B(n12164), .Y(n18006) );
  sky130_fd_sc_hd__nand2_1 U18850 ( .A(n18001), .B(n18000), .Y(n12164) );
  sky130_fd_sc_hd__o21ai_1 U18851 ( .A1(n18000), .A2(n18001), .B1(n17999), .Y(
        n12165) );
  sky130_fd_sc_hd__xnor2_1 U18853 ( .A(n18000), .B(n18001), .Y(n12166) );
  sky130_fd_sc_hd__nor2_2 U18854 ( .A(n18284), .B(n18285), .Y(n22976) );
  sky130_fd_sc_hd__nand3_1 U18855 ( .A(n22677), .B(n22929), .C(n22789), .Y(
        n12168) );
  sky130_fd_sc_hd__nand2_1 U18856 ( .A(n22677), .B(n23021), .Y(n12171) );
  sky130_fd_sc_hd__nand3_1 U18857 ( .A(n12169), .B(n22928), .C(n12168), .Y(
        n22679) );
  sky130_fd_sc_hd__nand2_1 U18858 ( .A(n22676), .B(n22929), .Y(n12169) );
  sky130_fd_sc_hd__nand2_1 U18859 ( .A(n12171), .B(n12170), .Y(n22931) );
  sky130_fd_sc_hd__nand2_1 U18860 ( .A(n12173), .B(n12172), .Y(n19067) );
  sky130_fd_sc_hd__nand2_1 U18861 ( .A(n19018), .B(n19019), .Y(n12172) );
  sky130_fd_sc_hd__o21ai_1 U18862 ( .A1(n19019), .A2(n19018), .B1(n19017), .Y(
        n12173) );
  sky130_fd_sc_hd__xnor2_1 U18863 ( .A(n19018), .B(n12174), .Y(n19066) );
  sky130_fd_sc_hd__xnor2_1 U18864 ( .A(n19019), .B(n19017), .Y(n12174) );
  sky130_fd_sc_hd__nand2_1 U18865 ( .A(n12176), .B(n12175), .Y(n18282) );
  sky130_fd_sc_hd__nand2_1 U18866 ( .A(n18276), .B(n18277), .Y(n12175) );
  sky130_fd_sc_hd__nand2_1 U18867 ( .A(n18275), .B(n12177), .Y(n12176) );
  sky130_fd_sc_hd__nand2_1 U18868 ( .A(n12179), .B(n12178), .Y(n12177) );
  sky130_fd_sc_hd__xnor2_1 U18869 ( .A(n18275), .B(n12180), .Y(n18278) );
  sky130_fd_sc_hd__xnor2_1 U18870 ( .A(n18277), .B(n18276), .Y(n12180) );
  sky130_fd_sc_hd__nand3_2 U18871 ( .A(n12182), .B(n12183), .C(n27824), .Y(
        n27896) );
  sky130_fd_sc_hd__and2_1 U18872 ( .A(n27833), .B(n27832), .X(n12183) );
  sky130_fd_sc_hd__nand2_1 U18874 ( .A(n12184), .B(n21696), .Y(n21212) );
  sky130_fd_sc_hd__nand2_1 U18875 ( .A(n12184), .B(n25724), .Y(n24085) );
  sky130_fd_sc_hd__nand2_1 U18876 ( .A(n12184), .B(n28539), .Y(n28517) );
  sky130_fd_sc_hd__a22oi_1 U18877 ( .A1(n24773), .A2(n27862), .B1(n12184), 
        .B2(n27861), .Y(n24776) );
  sky130_fd_sc_hd__nor2_1 U18878 ( .A(n12184), .B(n26188), .Y(n26199) );
  sky130_fd_sc_hd__o21ai_1 U18879 ( .A1(n12190), .A2(n12185), .B1(n20454), .Y(
        n12523) );
  sky130_fd_sc_hd__nand4_1 U18880 ( .A(n12189), .B(n12188), .C(n12187), .D(
        n12186), .Y(n12185) );
  sky130_fd_sc_hd__nand2_1 U18881 ( .A(j202_soc_core_memory0_ram_dout0[52]), 
        .B(n21633), .Y(n12186) );
  sky130_fd_sc_hd__nand2_1 U18882 ( .A(j202_soc_core_memory0_ram_dout0[308]), 
        .B(n21503), .Y(n12187) );
  sky130_fd_sc_hd__nand2_1 U18883 ( .A(j202_soc_core_memory0_ram_dout0[436]), 
        .B(n12156), .Y(n12188) );
  sky130_fd_sc_hd__nand2_1 U18884 ( .A(j202_soc_core_memory0_ram_dout0[468]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12189) );
  sky130_fd_sc_hd__nand2_1 U18885 ( .A(j202_soc_core_memory0_ram_dout0[372]), 
        .B(n21495), .Y(n12191) );
  sky130_fd_sc_hd__nand2_1 U18886 ( .A(j202_soc_core_memory0_ram_dout0[276]), 
        .B(n21634), .Y(n12192) );
  sky130_fd_sc_hd__nand2_1 U18887 ( .A(j202_soc_core_memory0_ram_dout0[340]), 
        .B(n21490), .Y(n12193) );
  sky130_fd_sc_hd__nand2_1 U18888 ( .A(n30085), .B(n21841), .Y(n28508) );
  sky130_fd_sc_hd__nand2_1 U18889 ( .A(n12195), .B(n12194), .Y(n21864) );
  sky130_fd_sc_hd__or2_0 U18890 ( .A(n21862), .B(n21863), .X(n12194) );
  sky130_fd_sc_hd__and2_0 U18891 ( .A(n21842), .B(n26411), .X(n12198) );
  sky130_fd_sc_hd__nand2b_1 U18892 ( .A_N(n11108), .B(n12200), .Y(n12199) );
  sky130_fd_sc_hd__o21a_1 U18893 ( .A1(n12202), .A2(n21841), .B1(n22136), .X(
        n12201) );
  sky130_fd_sc_hd__nand2b_1 U18894 ( .A_N(n27785), .B(n21842), .Y(n12202) );
  sky130_fd_sc_hd__nand2_1 U18895 ( .A(n21865), .B(n21864), .Y(n27359) );
  sky130_fd_sc_hd__buf_6 U18896 ( .A(n25381), .X(n12203) );
  sky130_fd_sc_hd__inv_2 U18897 ( .A(n25381), .Y(n25779) );
  sky130_fd_sc_hd__nand2_1 U18898 ( .A(n25381), .B(n27117), .Y(n12204) );
  sky130_fd_sc_hd__o21a_2 U18899 ( .A1(n24695), .A2(n28379), .B1(n24420), .X(
        n24426) );
  sky130_fd_sc_hd__nand3_1 U18900 ( .A(n30083), .B(n24683), .C(n12780), .Y(
        n24688) );
  sky130_fd_sc_hd__nand3_1 U18901 ( .A(n28097), .B(n28096), .C(n28095), .Y(
        n28393) );
  sky130_fd_sc_hd__nand3_1 U18902 ( .A(n18856), .B(n18857), .C(n22266), .Y(
        n12206) );
  sky130_fd_sc_hd__buf_4 U18903 ( .A(n24472), .X(n12207) );
  sky130_fd_sc_hd__a21oi_1 U18904 ( .A1(n22147), .A2(n26426), .B1(n22146), .Y(
        n12209) );
  sky130_fd_sc_hd__nand2_1 U18906 ( .A(n11175), .B(n27728), .Y(n28261) );
  sky130_fd_sc_hd__buf_2 U18907 ( .A(n11138), .X(n12213) );
  sky130_fd_sc_hd__buf_6 U18908 ( .A(n11138), .X(n12214) );
  sky130_fd_sc_hd__nand2_1 U18910 ( .A(n12216), .B(n12217), .Y(n12219) );
  sky130_fd_sc_hd__inv_2 U18911 ( .A(n23509), .Y(n24179) );
  sky130_fd_sc_hd__nand2_1 U18912 ( .A(n28430), .B(n27785), .Y(n26409) );
  sky130_fd_sc_hd__a21o_1 U18914 ( .A1(n18189), .A2(n18192), .B1(n17508), .X(
        n17475) );
  sky130_fd_sc_hd__nor2b_1 U18915 ( .B_N(n18470), .A(n18192), .Y(n18114) );
  sky130_fd_sc_hd__a21oi_1 U18917 ( .A1(n23955), .A2(n24423), .B1(n23607), .Y(
        n23618) );
  sky130_fd_sc_hd__clkbuf_1 U18918 ( .A(n25633), .X(n12368) );
  sky130_fd_sc_hd__nand2_8 U18919 ( .A(n18213), .B(n17462), .Y(n12538) );
  sky130_fd_sc_hd__nand2_1 U18920 ( .A(n21872), .B(n27355), .Y(n12223) );
  sky130_fd_sc_hd__inv_1 U18921 ( .A(n12352), .Y(n21872) );
  sky130_fd_sc_hd__and2_4 U18922 ( .A(n17369), .B(n17368), .X(n12224) );
  sky130_fd_sc_hd__inv_2 U18923 ( .A(n24915), .Y(n12225) );
  sky130_fd_sc_hd__nand2_1 U18924 ( .A(n23408), .B(n11176), .Y(n23395) );
  sky130_fd_sc_hd__and2_4 U18925 ( .A(n29501), .B(n12214), .X(n12231) );
  sky130_fd_sc_hd__inv_8 U18926 ( .A(n29759), .Y(n12384) );
  sky130_fd_sc_hd__buf_2 U18927 ( .A(n28378), .X(n12235) );
  sky130_fd_sc_hd__nand4_1 U18928 ( .A(n23619), .B(n12350), .C(n23617), .D(
        n23618), .Y(n12237) );
  sky130_fd_sc_hd__fah_1 U18929 ( .A(n19027), .B(n19026), .CI(n19025), .COUT(
        n19043), .SUM(n19030) );
  sky130_fd_sc_hd__o21ai_1 U18930 ( .A1(n23023), .A2(n12349), .B1(n23022), .Y(
        n23024) );
  sky130_fd_sc_hd__o21ai_1 U18931 ( .A1(n21911), .A2(n12349), .B1(n21910), .Y(
        n21912) );
  sky130_fd_sc_hd__nor2_1 U18933 ( .A(n24421), .B(n22010), .Y(n12240) );
  sky130_fd_sc_hd__nor2_1 U18934 ( .A(n24421), .B(n22010), .Y(n12847) );
  sky130_fd_sc_hd__nand3_2 U18935 ( .A(n22267), .B(n22265), .C(n22266), .Y(
        n12241) );
  sky130_fd_sc_hd__and2_4 U18936 ( .A(n29517), .B(n11853), .X(n12242) );
  sky130_fd_sc_hd__and2_4 U18937 ( .A(n29517), .B(n11853), .X(n12243) );
  sky130_fd_sc_hd__and2_4 U18938 ( .A(n29552), .B(n12271), .X(n23982) );
  sky130_fd_sc_hd__inv_1 U18939 ( .A(n22004), .Y(n12244) );
  sky130_fd_sc_hd__clkbuf_1 U18940 ( .A(n12781), .X(n12779) );
  sky130_fd_sc_hd__inv_2 U18941 ( .A(n25856), .Y(n12246) );
  sky130_fd_sc_hd__inv_2 U18942 ( .A(n25856), .Y(n27386) );
  sky130_fd_sc_hd__clkbuf_1 U18943 ( .A(n27884), .X(n12249) );
  sky130_fd_sc_hd__buf_8 U18944 ( .A(n12371), .X(n12312) );
  sky130_fd_sc_hd__a2bb2oi_2 U18945 ( .B1(n25392), .B2(n29487), .A1_N(n12367), 
        .A2_N(n24069), .Y(n26162) );
  sky130_fd_sc_hd__inv_1 U18946 ( .A(n23379), .Y(n12453) );
  sky130_fd_sc_hd__nor2_1 U18949 ( .A(n12220), .B(n27739), .Y(n24112) );
  sky130_fd_sc_hd__nand2_1 U18950 ( .A(n22450), .B(n21871), .Y(n21874) );
  sky130_fd_sc_hd__inv_2 U18951 ( .A(n29822), .Y(n12372) );
  sky130_fd_sc_hd__inv_1 U18952 ( .A(n23408), .Y(n12253) );
  sky130_fd_sc_hd__inv_2 U18953 ( .A(n29761), .Y(n12386) );
  sky130_fd_sc_hd__inv_2 U18955 ( .A(n29822), .Y(n12373) );
  sky130_fd_sc_hd__nand2_1 U18957 ( .A(n23408), .B(n12220), .Y(n12434) );
  sky130_fd_sc_hd__mux2i_1 U18958 ( .A0(n26670), .A1(n26669), .S(n24832), .Y(
        j202_soc_core_j22_cpu_rf_N3283) );
  sky130_fd_sc_hd__inv_2 U18959 ( .A(n24861), .Y(n12256) );
  sky130_fd_sc_hd__inv_2 U18960 ( .A(n24861), .Y(n28060) );
  sky130_fd_sc_hd__inv_2 U18964 ( .A(n12259), .Y(n12260) );
  sky130_fd_sc_hd__inv_8 U18965 ( .A(n29756), .Y(n12380) );
  sky130_fd_sc_hd__a21oi_1 U18966 ( .A1(n21777), .A2(n21451), .B1(n11204), .Y(
        n21484) );
  sky130_fd_sc_hd__nand3_1 U18967 ( .A(n21439), .B(n21438), .C(n21437), .Y(
        n21440) );
  sky130_fd_sc_hd__inv_1 U18968 ( .A(n26160), .Y(n12542) );
  sky130_fd_sc_hd__nor2_1 U18971 ( .A(n20898), .B(n20897), .Y(n12270) );
  sky130_fd_sc_hd__o21a_1 U18972 ( .A1(n25696), .A2(n25701), .B1(n25700), .X(
        n12261) );
  sky130_fd_sc_hd__nand2_1 U18973 ( .A(n12261), .B(n25699), .Y(n25702) );
  sky130_fd_sc_hd__nand2_1 U18974 ( .A(n25961), .B(n26009), .Y(n12263) );
  sky130_fd_sc_hd__and2_4 U18975 ( .A(n12263), .B(n12113), .X(n25968) );
  sky130_fd_sc_hd__nand3_1 U18976 ( .A(n25943), .B(n26919), .C(n25942), .Y(
        n25961) );
  sky130_fd_sc_hd__inv_2 U18977 ( .A(n28442), .Y(n27572) );
  sky130_fd_sc_hd__nor2_1 U18978 ( .A(n24403), .B(n24402), .Y(n28123) );
  sky130_fd_sc_hd__inv_2 U18979 ( .A(n25383), .Y(n12266) );
  sky130_fd_sc_hd__inv_2 U18980 ( .A(n25383), .Y(n12267) );
  sky130_fd_sc_hd__nor2_1 U18983 ( .A(n20898), .B(n20897), .Y(n23999) );
  sky130_fd_sc_hd__inv_2 U18984 ( .A(n12271), .Y(n12272) );
  sky130_fd_sc_hd__nand2_1 U18985 ( .A(n23614), .B(n12393), .Y(n12335) );
  sky130_fd_sc_hd__nand3b_1 U18987 ( .A_N(n12923), .B(n24407), .C(n12922), .Y(
        n27884) );
  sky130_fd_sc_hd__buf_6 U18988 ( .A(n12534), .X(n12533) );
  sky130_fd_sc_hd__inv_2 U18989 ( .A(n23434), .Y(n23551) );
  sky130_fd_sc_hd__nor2_1 U18992 ( .A(n23439), .B(n12051), .Y(n12280) );
  sky130_fd_sc_hd__a21bo_2 U18993 ( .A1(n27645), .A2(n27152), .B1_N(n27649), 
        .X(n12281) );
  sky130_fd_sc_hd__nand2_1 U18994 ( .A(n12393), .B(n29593), .Y(n12285) );
  sky130_fd_sc_hd__inv_4 U18995 ( .A(n29760), .Y(n12289) );
  sky130_fd_sc_hd__o21a_1 U18996 ( .A1(n29593), .A2(n12235), .B1(n28345), .X(
        n13048) );
  sky130_fd_sc_hd__inv_4 U18997 ( .A(n29760), .Y(n12290) );
  sky130_fd_sc_hd__inv_1 U18998 ( .A(n30058), .Y(n12291) );
  sky130_fd_sc_hd__a21oi_1 U18999 ( .A1(n13012), .A2(n13001), .B1(n15630), .Y(
        n22226) );
  sky130_fd_sc_hd__nand2_1 U19000 ( .A(n16739), .B(n20454), .Y(n12846) );
  sky130_fd_sc_hd__and2_1 U19001 ( .A(n15494), .B(n12121), .X(n12728) );
  sky130_fd_sc_hd__nand2b_1 U19002 ( .A_N(n29746), .B(n29745), .Y(n10600) );
  sky130_fd_sc_hd__nor2_1 U19003 ( .A(n13403), .B(n13402), .Y(n13821) );
  sky130_fd_sc_hd__nor2_1 U19004 ( .A(n21042), .B(n12574), .Y(n21043) );
  sky130_fd_sc_hd__nor2_1 U19008 ( .A(n14575), .B(n14576), .Y(n20984) );
  sky130_fd_sc_hd__buf_8 U19009 ( .A(n12371), .X(n12313) );
  sky130_fd_sc_hd__buf_8 U19010 ( .A(n12371), .X(n12314) );
  sky130_fd_sc_hd__inv_12 U19011 ( .A(n23982), .Y(n29760) );
  sky130_fd_sc_hd__and2b_4 U19012 ( .B(n29557), .A_N(n30070), .X(n23988) );
  sky130_fd_sc_hd__o21ai_1 U19013 ( .A1(n28133), .A2(n23547), .B1(n12064), .Y(
        n24545) );
  sky130_fd_sc_hd__and2_4 U19014 ( .A(n29501), .B(n12214), .X(n12319) );
  sky130_fd_sc_hd__nand3_4 U19016 ( .A(n24427), .B(n24425), .C(n24426), .Y(
        n12364) );
  sky130_fd_sc_hd__nand2_1 U19017 ( .A(n24632), .B(n12151), .Y(n10641) );
  sky130_fd_sc_hd__o22ai_2 U19018 ( .A1(n23252), .A2(n23237), .B1(n23236), 
        .B2(n23235), .Y(n23245) );
  sky130_fd_sc_hd__nand2_2 U19019 ( .A(n27345), .B(n29480), .Y(n24384) );
  sky130_fd_sc_hd__nor2_2 U19021 ( .A(n24387), .B(n27336), .Y(n24391) );
  sky130_fd_sc_hd__a22oi_2 U19022 ( .A1(j202_soc_core_memory0_ram_dout0[103]), 
        .A2(n21488), .B1(n21487), .B2(j202_soc_core_memory0_ram_dout0[167]), 
        .Y(n17233) );
  sky130_fd_sc_hd__nor2_2 U19023 ( .A(n19063), .B(n19064), .Y(n22920) );
  sky130_fd_sc_hd__fah_1 U19025 ( .A(n18466), .B(n18465), .CI(n18464), .COUT(
        n18424), .SUM(n18539) );
  sky130_fd_sc_hd__nand3_1 U19026 ( .A(n21922), .B(n21921), .C(n21923), .Y(
        n12323) );
  sky130_fd_sc_hd__nand3_1 U19027 ( .A(n12240), .B(n24116), .C(n28150), .Y(
        n24117) );
  sky130_fd_sc_hd__a21o_1 U19029 ( .A1(n25381), .A2(n25380), .B1(n25776), .X(
        j202_soc_core_j22_cpu_ml_machj[21]) );
  sky130_fd_sc_hd__nand2_1 U19030 ( .A(n12594), .B(n12584), .Y(n21002) );
  sky130_fd_sc_hd__nand3_1 U19034 ( .A(n12140), .B(n12728), .C(n12726), .Y(
        n12725) );
  sky130_fd_sc_hd__o22a_1 U19035 ( .A1(n26276), .A2(n22745), .B1(n22705), .B2(
        n25286), .X(n16305) );
  sky130_fd_sc_hd__nand2_1 U19036 ( .A(n12526), .B(n12159), .Y(n22261) );
  sky130_fd_sc_hd__nor2_1 U19037 ( .A(n12094), .B(n12535), .Y(n24144) );
  sky130_fd_sc_hd__inv_2 U19038 ( .A(n26968), .Y(n12330) );
  sky130_fd_sc_hd__inv_2 U19039 ( .A(n26968), .Y(n24363) );
  sky130_fd_sc_hd__nor2_1 U19040 ( .A(n19303), .B(n21268), .Y(n22956) );
  sky130_fd_sc_hd__a22oi_2 U19041 ( .A1(j202_soc_core_memory0_ram_dout0[48]), 
        .A2(n21633), .B1(n21503), .B2(j202_soc_core_memory0_ram_dout0[304]), 
        .Y(n19849) );
  sky130_fd_sc_hd__fah_1 U19042 ( .A(n18413), .B(n18412), .CI(n18411), .COUT(
        n18438), .SUM(n18436) );
  sky130_fd_sc_hd__nor2_1 U19043 ( .A(n12458), .B(n12457), .Y(n12456) );
  sky130_fd_sc_hd__fah_1 U19045 ( .A(n17648), .B(n17647), .CI(n17646), .COUT(
        n18567), .SUM(n17671) );
  sky130_fd_sc_hd__and2b_4 U19046 ( .B(n29553), .A_N(n30070), .X(n23987) );
  sky130_fd_sc_hd__inv_1 U19047 ( .A(n23553), .Y(n12337) );
  sky130_fd_sc_hd__and3_1 U19048 ( .A(n28148), .B(n28147), .C(n28387), .X(
        n28149) );
  sky130_fd_sc_hd__nand4_1 U19049 ( .A(n24103), .B(n27909), .C(n27905), .D(
        n28148), .Y(n12338) );
  sky130_fd_sc_hd__nand2_2 U19050 ( .A(n12241), .B(n22952), .Y(n24447) );
  sky130_fd_sc_hd__and2b_4 U19051 ( .B(n29556), .A_N(n30070), .X(n23983) );
  sky130_fd_sc_hd__buf_6 U19053 ( .A(n27363), .X(n12344) );
  sky130_fd_sc_hd__and2b_4 U19054 ( .B(n29554), .A_N(n30070), .X(n23985) );
  sky130_fd_sc_hd__inv_2 U19055 ( .A(n17870), .Y(n18338) );
  sky130_fd_sc_hd__and2b_4 U19056 ( .B(n29555), .A_N(n30070), .X(n23984) );
  sky130_fd_sc_hd__nand3_1 U19057 ( .A(n12646), .B(n19848), .C(n12645), .Y(
        n12644) );
  sky130_fd_sc_hd__nand2_2 U19059 ( .A(n23375), .B(n23374), .Y(n23377) );
  sky130_fd_sc_hd__nand3_2 U19060 ( .A(n14752), .B(n14751), .C(n14750), .Y(
        n27807) );
  sky130_fd_sc_hd__nand2_1 U19061 ( .A(n16543), .B(n11144), .Y(n12355) );
  sky130_fd_sc_hd__nand2_1 U19062 ( .A(n16088), .B(n28529), .Y(n12356) );
  sky130_fd_sc_hd__nand2_1 U19063 ( .A(n21993), .B(n16523), .Y(n13786) );
  sky130_fd_sc_hd__nand4_1 U19064 ( .A(n13776), .B(n13775), .C(n13774), .D(
        n30023), .Y(n21993) );
  sky130_fd_sc_hd__inv_2 U19065 ( .A(n16541), .Y(n16088) );
  sky130_fd_sc_hd__nor2_2 U19067 ( .A(n19069), .B(n19070), .Y(n21907) );
  sky130_fd_sc_hd__inv_1 U19068 ( .A(n24626), .Y(n24640) );
  sky130_fd_sc_hd__nand3_1 U19069 ( .A(n20417), .B(n30200), .C(n11107), .Y(
        n20441) );
  sky130_fd_sc_hd__nand3_1 U19070 ( .A(n12820), .B(n12332), .C(n23421), .Y(
        n24409) );
  sky130_fd_sc_hd__o211ai_1 U19071 ( .A1(j202_soc_core_intc_core_00_rg_ipr[17]), .A2(n25578), .B1(n23186), .C1(n23185), .Y(n23188) );
  sky130_fd_sc_hd__nand3_1 U19072 ( .A(n18797), .B(n23505), .C(n23514), .Y(
        n25941) );
  sky130_fd_sc_hd__o21a_1 U19073 ( .A1(n27648), .A2(n25968), .B1(n25967), .X(
        n25969) );
  sky130_fd_sc_hd__buf_6 U19074 ( .A(n17334), .X(n18474) );
  sky130_fd_sc_hd__inv_1 U19077 ( .A(n23395), .Y(n23380) );
  sky130_fd_sc_hd__nand3_1 U19078 ( .A(n21874), .B(n12223), .C(n22266), .Y(
        n12365) );
  sky130_fd_sc_hd__inv_2 U19079 ( .A(n25271), .Y(n26431) );
  sky130_fd_sc_hd__buf_2 U19080 ( .A(n26166), .X(n12367) );
  sky130_fd_sc_hd__nor2_1 U19081 ( .A(n12908), .B(n12903), .Y(n12902) );
  sky130_fd_sc_hd__nand3_1 U19082 ( .A(n13638), .B(n13637), .C(n13636), .Y(
        n22282) );
  sky130_fd_sc_hd__nand2_1 U19083 ( .A(n10959), .B(n29436), .Y(n21045) );
  sky130_fd_sc_hd__inv_1 U19084 ( .A(n18815), .Y(n22752) );
  sky130_fd_sc_hd__nand3_1 U19085 ( .A(n24143), .B(n12334), .C(n12574), .Y(
        n17080) );
  sky130_fd_sc_hd__nand2_1 U19087 ( .A(n25282), .B(n12391), .Y(n12390) );
  sky130_fd_sc_hd__or2_0 U19088 ( .A(n25682), .B(n25265), .X(n12391) );
  sky130_fd_sc_hd__and2_0 U19089 ( .A(n25277), .B(n25278), .X(n12392) );
  sky130_fd_sc_hd__a22oi_2 U19090 ( .A1(j202_soc_core_memory0_ram_dout0[135]), 
        .A2(n21489), .B1(n21642), .B2(j202_soc_core_memory0_ram_dout0[71]), 
        .Y(n17232) );
  sky130_fd_sc_hd__a22oi_2 U19091 ( .A1(j202_soc_core_memory0_ram_dout0[116]), 
        .A2(n20460), .B1(n20459), .B2(j202_soc_core_memory0_ram_dout0[180]), 
        .Y(n15370) );
  sky130_fd_sc_hd__inv_1 U19092 ( .A(n17321), .Y(n12768) );
  sky130_fd_sc_hd__buf_2 U19093 ( .A(n24404), .X(n12393) );
  sky130_fd_sc_hd__o21ai_1 U19094 ( .A1(n12394), .A2(n12793), .B1(n20454), .Y(
        n12792) );
  sky130_fd_sc_hd__nand3_1 U19095 ( .A(n14726), .B(n12791), .C(n12790), .Y(
        n12789) );
  sky130_fd_sc_hd__buf_2 U19096 ( .A(n12816), .X(n12621) );
  sky130_fd_sc_hd__clkbuf_1 U19097 ( .A(n28492), .X(n12396) );
  sky130_fd_sc_hd__nand2_2 U19098 ( .A(n12397), .B(n25373), .Y(n25630) );
  sky130_fd_sc_hd__or2_0 U19099 ( .A(n25658), .B(n25371), .X(n12398) );
  sky130_fd_sc_hd__clkbuf_1 U19100 ( .A(n28089), .X(n12399) );
  sky130_fd_sc_hd__inv_1 U19102 ( .A(n23600), .Y(n23619) );
  sky130_fd_sc_hd__nand3_1 U19103 ( .A(n25145), .B(n22394), .C(n22393), .Y(
        n12510) );
  sky130_fd_sc_hd__nand2_1 U19104 ( .A(n12404), .B(n12403), .Y(n18408) );
  sky130_fd_sc_hd__nand2b_1 U19105 ( .A_N(n12407), .B(n18362), .Y(n12403) );
  sky130_fd_sc_hd__nand2_1 U19106 ( .A(n18361), .B(n12405), .Y(n12404) );
  sky130_fd_sc_hd__nand2b_1 U19107 ( .A_N(n18362), .B(n12407), .Y(n12405) );
  sky130_fd_sc_hd__xor2_1 U19108 ( .A(n12406), .B(n18361), .X(n18523) );
  sky130_fd_sc_hd__xnor2_1 U19109 ( .A(n18362), .B(n12407), .Y(n12406) );
  sky130_fd_sc_hd__nand3_1 U19110 ( .A(n17332), .B(n17331), .C(n17330), .Y(
        n17333) );
  sky130_fd_sc_hd__nand3_2 U19111 ( .A(n21241), .B(n21240), .C(n22266), .Y(
        n22826) );
  sky130_fd_sc_hd__nand3_1 U19112 ( .A(n27991), .B(n24968), .C(n25148), .Y(
        n23401) );
  sky130_fd_sc_hd__clkbuf_1 U19113 ( .A(n24068), .X(n12409) );
  sky130_fd_sc_hd__o22ai_1 U19115 ( .A1(n18486), .A2(n17447), .B1(n17478), 
        .B2(n18483), .Y(n17477) );
  sky130_fd_sc_hd__nand2_4 U19116 ( .A(n18486), .B(n17444), .Y(n18483) );
  sky130_fd_sc_hd__xnor2_1 U19117 ( .A(n17572), .B(n12411), .Y(n17860) );
  sky130_fd_sc_hd__xnor2_1 U19118 ( .A(n17574), .B(n17573), .Y(n12411) );
  sky130_fd_sc_hd__nand2_1 U19119 ( .A(n12413), .B(n12412), .Y(n17861) );
  sky130_fd_sc_hd__nand2_1 U19120 ( .A(n17573), .B(n17574), .Y(n12412) );
  sky130_fd_sc_hd__nor2_1 U19123 ( .A(n12531), .B(n12530), .Y(n12529) );
  sky130_fd_sc_hd__o21ai_1 U19124 ( .A1(n27355), .A2(n25866), .B1(n25891), .Y(
        n12429) );
  sky130_fd_sc_hd__nand2_1 U19125 ( .A(n12415), .B(n12414), .Y(n17570) );
  sky130_fd_sc_hd__nand2_1 U19126 ( .A(n17532), .B(n17531), .Y(n12414) );
  sky130_fd_sc_hd__o21ai_1 U19127 ( .A1(n17531), .A2(n17532), .B1(n17530), .Y(
        n12415) );
  sky130_fd_sc_hd__xnor2_1 U19128 ( .A(n17532), .B(n12416), .Y(n17834) );
  sky130_fd_sc_hd__xnor2_1 U19129 ( .A(n17530), .B(n17531), .Y(n12416) );
  sky130_fd_sc_hd__a21oi_2 U19130 ( .A1(n23507), .A2(n23506), .B1(n26189), .Y(
        n23515) );
  sky130_fd_sc_hd__nand2_1 U19131 ( .A(n25563), .B(n12420), .Y(n12419) );
  sky130_fd_sc_hd__nor2b_1 U19132 ( .B_N(n25558), .A(n25557), .Y(n12420) );
  sky130_fd_sc_hd__clkbuf_1 U19133 ( .A(n24144), .X(n12421) );
  sky130_fd_sc_hd__inv_2 U19134 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]), 
        .Y(n12684) );
  sky130_fd_sc_hd__and2_4 U19135 ( .A(n27152), .B(n27016), .X(n12426) );
  sky130_fd_sc_hd__clkbuf_1 U19136 ( .A(n26165), .X(n12423) );
  sky130_fd_sc_hd__nand3_1 U19137 ( .A(n11174), .B(n23604), .C(n24593), .Y(
        n12424) );
  sky130_fd_sc_hd__clkbuf_1 U19138 ( .A(j202_soc_core_j22_cpu_ml_bufa[30]), 
        .X(n12425) );
  sky130_fd_sc_hd__nor2_8 U19139 ( .A(n12426), .B(n25935), .Y(n28111) );
  sky130_fd_sc_hd__nor2_4 U19140 ( .A(n23403), .B(n24564), .Y(n28133) );
  sky130_fd_sc_hd__nand3_1 U19141 ( .A(n12441), .B(n12442), .C(n12440), .Y(
        n12758) );
  sky130_fd_sc_hd__nand2_1 U19142 ( .A(n25888), .B(n27115), .Y(n12427) );
  sky130_fd_sc_hd__o21ai_1 U19144 ( .A1(n27919), .A2(n27918), .B1(n12155), .Y(
        j202_soc_core_ahb2aqu_00_N161) );
  sky130_fd_sc_hd__a21oi_2 U19146 ( .A1(n21880), .A2(n12432), .B1(n18288), .Y(
        n18881) );
  sky130_fd_sc_hd__nor2_1 U19147 ( .A(n22976), .B(n22971), .Y(n12432) );
  sky130_fd_sc_hd__nand2_1 U19148 ( .A(n23486), .B(n23487), .Y(n12433) );
  sky130_fd_sc_hd__buf_6 U19149 ( .A(n18224), .X(n18536) );
  sky130_fd_sc_hd__clkbuf_1 U19150 ( .A(n22211), .X(n12435) );
  sky130_fd_sc_hd__clkbuf_1 U19151 ( .A(j202_soc_core_j22_cpu_ml_bufa[2]), .X(
        n12436) );
  sky130_fd_sc_hd__nand2_1 U19152 ( .A(n12438), .B(n12437), .Y(n18092) );
  sky130_fd_sc_hd__nand2_1 U19153 ( .A(n18090), .B(n18089), .Y(n12437) );
  sky130_fd_sc_hd__o21ai_1 U19154 ( .A1(n18089), .A2(n18090), .B1(n18088), .Y(
        n12438) );
  sky130_fd_sc_hd__xnor2_1 U19155 ( .A(n18088), .B(n12439), .Y(n18281) );
  sky130_fd_sc_hd__xnor2_1 U19156 ( .A(n18090), .B(n18089), .Y(n12439) );
  sky130_fd_sc_hd__nand2_1 U19157 ( .A(j202_soc_core_memory0_ram_dout0[89]), 
        .B(n20458), .Y(n12440) );
  sky130_fd_sc_hd__nand2_1 U19158 ( .A(j202_soc_core_memory0_ram_dout0[25]), 
        .B(n20457), .Y(n12441) );
  sky130_fd_sc_hd__nand2_1 U19159 ( .A(j202_soc_core_memory0_ram_dout0[217]), 
        .B(n20455), .Y(n12442) );
  sky130_fd_sc_hd__nor2_1 U19160 ( .A(n12445), .B(n12952), .Y(n12444) );
  sky130_fd_sc_hd__nand2_1 U19161 ( .A(n12970), .B(n12111), .Y(n12969) );
  sky130_fd_sc_hd__nand2_1 U19162 ( .A(n12968), .B(n12953), .Y(n12446) );
  sky130_fd_sc_hd__nand2_1 U19163 ( .A(n21336), .B(n12112), .Y(n12953) );
  sky130_fd_sc_hd__nand2_1 U19166 ( .A(j202_soc_core_memory0_ram_dout0[381]), 
        .B(n21495), .Y(n12448) );
  sky130_fd_sc_hd__nand2_1 U19167 ( .A(j202_soc_core_memory0_ram_dout0[349]), 
        .B(n21490), .Y(n12449) );
  sky130_fd_sc_hd__nand2_1 U19168 ( .A(j202_soc_core_memory0_ram_dout0[285]), 
        .B(n21634), .Y(n12450) );
  sky130_fd_sc_hd__nand2_1 U19169 ( .A(j202_soc_core_memory0_ram_dout0[221]), 
        .B(n21640), .Y(n12451) );
  sky130_fd_sc_hd__o21bai_1 U19170 ( .A1(n12235), .A2(n28380), .B1_N(n12211), 
        .Y(n28358) );
  sky130_fd_sc_hd__nand2b_1 U19171 ( .A_N(n23379), .B(n12452), .Y(n28348) );
  sky130_fd_sc_hd__and3_1 U19173 ( .A(n18784), .B(n18788), .C(n18791), .X(
        n12454) );
  sky130_fd_sc_hd__inv_1 U19174 ( .A(n12252), .Y(n23459) );
  sky130_fd_sc_hd__nand4_1 U19175 ( .A(n16936), .B(n16937), .C(n16935), .D(
        n17017), .Y(n12458) );
  sky130_fd_sc_hd__nand2_1 U19177 ( .A(n25633), .B(n22739), .Y(n12462) );
  sky130_fd_sc_hd__nand2_1 U19178 ( .A(n15374), .B(n20462), .Y(n12522) );
  sky130_fd_sc_hd__nand3_1 U19180 ( .A(n22653), .B(n22316), .C(n12464), .Y(
        n29516) );
  sky130_fd_sc_hd__and2_0 U19181 ( .A(n12465), .B(n22651), .X(n12464) );
  sky130_fd_sc_hd__or2_0 U19182 ( .A(n22330), .B(
        j202_soc_core_j22_cpu_memop_MEM__0_), .X(n12465) );
  sky130_fd_sc_hd__nand2_1 U19183 ( .A(n29516), .B(n11853), .Y(n12467) );
  sky130_fd_sc_hd__nand2_1 U19184 ( .A(n12469), .B(n12468), .Y(n18511) );
  sky130_fd_sc_hd__nand2_1 U19185 ( .A(n18424), .B(n18425), .Y(n12468) );
  sky130_fd_sc_hd__o21ai_1 U19186 ( .A1(n18424), .A2(n18425), .B1(n18423), .Y(
        n12469) );
  sky130_fd_sc_hd__xnor2_1 U19187 ( .A(n18423), .B(n12470), .Y(n18521) );
  sky130_fd_sc_hd__xnor2_1 U19188 ( .A(n18424), .B(n18425), .Y(n12470) );
  sky130_fd_sc_hd__nand2b_1 U19189 ( .A_N(n27460), .B(n27576), .Y(n26862) );
  sky130_fd_sc_hd__nand2_1 U19190 ( .A(n12473), .B(n12472), .Y(n18326) );
  sky130_fd_sc_hd__nand2b_1 U19191 ( .A_N(n12476), .B(n17948), .Y(n12472) );
  sky130_fd_sc_hd__nand2_1 U19192 ( .A(n12474), .B(n17947), .Y(n12473) );
  sky130_fd_sc_hd__nand2_1 U19193 ( .A(n12476), .B(n12475), .Y(n12474) );
  sky130_fd_sc_hd__xor2_1 U19194 ( .A(n17877), .B(n17876), .X(n12476) );
  sky130_fd_sc_hd__nand2_1 U19195 ( .A(n12478), .B(n12477), .Y(n17618) );
  sky130_fd_sc_hd__nand2_1 U19196 ( .A(n17582), .B(n12480), .Y(n12477) );
  sky130_fd_sc_hd__o21ai_1 U19197 ( .A1(n12480), .A2(n17582), .B1(n17581), .Y(
        n12478) );
  sky130_fd_sc_hd__xnor2_1 U19198 ( .A(n17582), .B(n12479), .Y(n17590) );
  sky130_fd_sc_hd__xnor2_1 U19199 ( .A(n12480), .B(n17581), .Y(n12479) );
  sky130_fd_sc_hd__nand2_1 U19200 ( .A(n12483), .B(n12482), .Y(n17872) );
  sky130_fd_sc_hd__nand2_1 U19201 ( .A(n17801), .B(n17800), .Y(n12482) );
  sky130_fd_sc_hd__o21ai_1 U19202 ( .A1(n17800), .A2(n17801), .B1(n17799), .Y(
        n12483) );
  sky130_fd_sc_hd__nand2b_4 U19204 ( .A_N(n21192), .B(n12485), .Y(n22107) );
  sky130_fd_sc_hd__nor2_2 U19206 ( .A(n21189), .B(n19105), .Y(n22193) );
  sky130_fd_sc_hd__nand2_1 U19207 ( .A(n12487), .B(n12486), .Y(n18626) );
  sky130_fd_sc_hd__nand2_1 U19208 ( .A(n18600), .B(n18601), .Y(n12486) );
  sky130_fd_sc_hd__o21ai_1 U19209 ( .A1(n18601), .A2(n18600), .B1(n18599), .Y(
        n12487) );
  sky130_fd_sc_hd__xnor3_1 U19210 ( .A(n12488), .B(n18600), .C(n18599), .X(
        n18634) );
  sky130_fd_sc_hd__nand3_1 U19212 ( .A(n22106), .B(n11866), .C(n12099), .Y(
        n12491) );
  sky130_fd_sc_hd__nand2_1 U19213 ( .A(n22107), .B(n12099), .Y(n12493) );
  sky130_fd_sc_hd__nand2_1 U19214 ( .A(n23477), .B(n24452), .Y(n22394) );
  sky130_fd_sc_hd__nand2_1 U19215 ( .A(n12834), .B(n20454), .Y(n12496) );
  sky130_fd_sc_hd__nand2_1 U19216 ( .A(n12656), .B(n12655), .Y(n12654) );
  sky130_fd_sc_hd__xnor2_1 U19217 ( .A(n18561), .B(n18562), .Y(n12499) );
  sky130_fd_sc_hd__xnor2_1 U19218 ( .A(n18560), .B(n12499), .Y(n18660) );
  sky130_fd_sc_hd__nand2_1 U19219 ( .A(n12500), .B(n18429), .Y(n12504) );
  sky130_fd_sc_hd__nand2b_1 U19220 ( .A_N(n12505), .B(n18508), .Y(n12500) );
  sky130_fd_sc_hd__xnor2_1 U19221 ( .A(n12504), .B(n12501), .Y(n18517) );
  sky130_fd_sc_hd__xnor2_1 U19222 ( .A(n18433), .B(n18432), .Y(n12501) );
  sky130_fd_sc_hd__nand2_1 U19223 ( .A(n12503), .B(n12502), .Y(n18448) );
  sky130_fd_sc_hd__nand2_1 U19224 ( .A(n18432), .B(n18433), .Y(n12502) );
  sky130_fd_sc_hd__xor2_1 U19226 ( .A(n13032), .B(n13031), .X(n18508) );
  sky130_fd_sc_hd__nand2_1 U19227 ( .A(n12507), .B(n12506), .Y(n18425) );
  sky130_fd_sc_hd__nand2_1 U19228 ( .A(n12209), .B(n27355), .Y(n12509) );
  sky130_fd_sc_hd__nand2_1 U19229 ( .A(n12990), .B(n20454), .Y(n12512) );
  sky130_fd_sc_hd__nand4_1 U19230 ( .A(n12994), .B(n12993), .C(n12992), .D(
        n12991), .Y(n12990) );
  sky130_fd_sc_hd__nand2_1 U19231 ( .A(n12848), .B(n12851), .Y(n12515) );
  sky130_fd_sc_hd__inv_1 U19232 ( .A(n12517), .Y(n12516) );
  sky130_fd_sc_hd__nand2_1 U19233 ( .A(n12766), .B(n12849), .Y(n12517) );
  sky130_fd_sc_hd__nand2_1 U19234 ( .A(n12519), .B(n21485), .Y(n22002) );
  sky130_fd_sc_hd__nand2_1 U19235 ( .A(n12521), .B(n12520), .Y(n12519) );
  sky130_fd_sc_hd__nand2_1 U19236 ( .A(n21486), .B(n11203), .Y(n12520) );
  sky130_fd_sc_hd__nand2_1 U19238 ( .A(n22258), .B(n11123), .Y(n12525) );
  sky130_fd_sc_hd__nand2_1 U19239 ( .A(n22257), .B(n22258), .Y(n12526) );
  sky130_fd_sc_hd__inv_1 U19240 ( .A(n22257), .Y(n26381) );
  sky130_fd_sc_hd__nand4_1 U19241 ( .A(n12870), .B(n12871), .C(n12872), .D(
        n12873), .Y(n12527) );
  sky130_fd_sc_hd__nand4_1 U19242 ( .A(n12869), .B(n12863), .C(n12864), .D(
        n12865), .Y(n12530) );
  sky130_fd_sc_hd__nor2b_1 U19243 ( .B_N(n12532), .A(n12533), .Y(
        j202_soc_core_ahb2apb_01_N56) );
  sky130_fd_sc_hd__nor2_1 U19244 ( .A(n24719), .B(n12533), .Y(
        j202_soc_core_ahb2apb_01_N32) );
  sky130_fd_sc_hd__nor2_1 U19245 ( .A(n27919), .B(n12533), .Y(
        j202_soc_core_ahb2apb_01_N24) );
  sky130_fd_sc_hd__nor2_1 U19246 ( .A(n27090), .B(n12533), .Y(
        j202_soc_core_ahb2apb_01_N23) );
  sky130_fd_sc_hd__nor2_1 U19247 ( .A(n24817), .B(n12533), .Y(
        j202_soc_core_ahb2apb_01_N25) );
  sky130_fd_sc_hd__nor2_1 U19248 ( .A(n24818), .B(n12533), .Y(
        j202_soc_core_ahb2apb_01_N26) );
  sky130_fd_sc_hd__nor2_1 U19249 ( .A(n27951), .B(n12533), .Y(
        j202_soc_core_ahb2apb_01_N31) );
  sky130_fd_sc_hd__nor2_1 U19250 ( .A(n25035), .B(n12533), .Y(
        j202_soc_core_ahb2apb_01_N30) );
  sky130_fd_sc_hd__nor2_1 U19251 ( .A(n25036), .B(n12533), .Y(
        j202_soc_core_ahb2apb_01_N29) );
  sky130_fd_sc_hd__nor2_1 U19252 ( .A(n25476), .B(n12533), .Y(
        j202_soc_core_ahb2apb_01_N57) );
  sky130_fd_sc_hd__nor2_1 U19253 ( .A(n25051), .B(n12533), .Y(
        j202_soc_core_ahb2apb_01_N33) );
  sky130_fd_sc_hd__nor2_1 U19254 ( .A(n25052), .B(n12533), .Y(
        j202_soc_core_ahb2apb_01_N34) );
  sky130_fd_sc_hd__nor2_1 U19255 ( .A(n25053), .B(n12533), .Y(
        j202_soc_core_ahb2apb_01_N27) );
  sky130_fd_sc_hd__nor2_1 U19256 ( .A(n25054), .B(n12533), .Y(
        j202_soc_core_ahb2apb_01_N28) );
  sky130_fd_sc_hd__nor2_1 U19257 ( .A(n25040), .B(n12533), .Y(
        j202_soc_core_ahb2apb_01_N89) );
  sky130_fd_sc_hd__nor2_1 U19258 ( .A(n12533), .B(n12842), .Y(
        j202_soc_core_ahb2apb_01_N55) );
  sky130_fd_sc_hd__nor2_1 U19259 ( .A(n12725), .B(n12535), .Y(n12724) );
  sky130_fd_sc_hd__nor2_1 U19260 ( .A(n17053), .B(n12816), .Y(n12535) );
  sky130_fd_sc_hd__nand2_2 U19261 ( .A(n13024), .B(n23561), .Y(n25381) );
  sky130_fd_sc_hd__nand2_1 U19262 ( .A(n12537), .B(n12536), .Y(n17541) );
  sky130_fd_sc_hd__nand2_1 U19263 ( .A(n12538), .B(n18213), .Y(n12536) );
  sky130_fd_sc_hd__o22ai_1 U19264 ( .A1(n18213), .A2(n17883), .B1(n17935), 
        .B2(n12538), .Y(n17973) );
  sky130_fd_sc_hd__o22ai_1 U19265 ( .A1(n18213), .A2(n17987), .B1(n17986), 
        .B2(n12538), .Y(n18014) );
  sky130_fd_sc_hd__o22ai_1 U19266 ( .A1(n18213), .A2(n17694), .B1(n17743), 
        .B2(n12538), .Y(n17707) );
  sky130_fd_sc_hd__o22ai_1 U19267 ( .A1(n18213), .A2(n17742), .B1(n17793), 
        .B2(n12538), .Y(n17895) );
  sky130_fd_sc_hd__o22ai_1 U19268 ( .A1(n18213), .A2(n17519), .B1(n17465), 
        .B2(n12538), .Y(n17482) );
  sky130_fd_sc_hd__o22ai_1 U19269 ( .A1(n18213), .A2(n17465), .B1(n17500), 
        .B2(n12538), .Y(n17472) );
  sky130_fd_sc_hd__o22ai_1 U19270 ( .A1(n18213), .A2(n17499), .B1(n17694), 
        .B2(n12538), .Y(n17711) );
  sky130_fd_sc_hd__o22ai_1 U19271 ( .A1(n18213), .A2(n17500), .B1(n17499), 
        .B2(n12538), .Y(n17756) );
  sky130_fd_sc_hd__o22ai_1 U19272 ( .A1(n18213), .A2(n17935), .B1(n17987), 
        .B2(n12538), .Y(n17959) );
  sky130_fd_sc_hd__o22ai_1 U19273 ( .A1(n18213), .A2(n17986), .B1(n18020), 
        .B2(n12538), .Y(n18055) );
  sky130_fd_sc_hd__o22ai_1 U19274 ( .A1(n18213), .A2(n17793), .B1(n17883), 
        .B2(n12538), .Y(n17920) );
  sky130_fd_sc_hd__o22ai_1 U19275 ( .A1(n18213), .A2(n17743), .B1(n17742), 
        .B2(n12538), .Y(n17780) );
  sky130_fd_sc_hd__o22ai_1 U19276 ( .A1(n18213), .A2(n18020), .B1(n18021), 
        .B2(n12538), .Y(n18087) );
  sky130_fd_sc_hd__nand2b_1 U19277 ( .A_N(n12541), .B(n17857), .Y(n22870) );
  sky130_fd_sc_hd__inv_2 U19278 ( .A(n12539), .Y(n22869) );
  sky130_fd_sc_hd__nand2_1 U19279 ( .A(n12541), .B(n12540), .Y(n12539) );
  sky130_fd_sc_hd__xnor2_1 U19280 ( .A(n17854), .B(n17853), .Y(n12541) );
  sky130_fd_sc_hd__nand2_1 U19281 ( .A(n12542), .B(n26181), .Y(n24833) );
  sky130_fd_sc_hd__nand3_2 U19282 ( .A(n12551), .B(n12547), .C(n12543), .Y(
        n16739) );
  sky130_fd_sc_hd__inv_2 U19283 ( .A(n12544), .Y(n12543) );
  sky130_fd_sc_hd__nand2_1 U19284 ( .A(n12546), .B(n12545), .Y(n12544) );
  sky130_fd_sc_hd__nand2_1 U19285 ( .A(j202_soc_core_memory0_ram_dout0[58]), 
        .B(n21633), .Y(n12545) );
  sky130_fd_sc_hd__nand2_1 U19286 ( .A(j202_soc_core_memory0_ram_dout0[314]), 
        .B(n21503), .Y(n12546) );
  sky130_fd_sc_hd__inv_2 U19287 ( .A(n12548), .Y(n12547) );
  sky130_fd_sc_hd__nand2_1 U19288 ( .A(n12550), .B(n12549), .Y(n12548) );
  sky130_fd_sc_hd__nand2_1 U19289 ( .A(j202_soc_core_memory0_ram_dout0[282]), 
        .B(n21634), .Y(n12549) );
  sky130_fd_sc_hd__nand2_1 U19290 ( .A(j202_soc_core_memory0_ram_dout0[346]), 
        .B(n21490), .Y(n12550) );
  sky130_fd_sc_hd__nand2_1 U19291 ( .A(j202_soc_core_memory0_ram_dout0[410]), 
        .B(n21496), .Y(n12552) );
  sky130_fd_sc_hd__nand2_1 U19292 ( .A(j202_soc_core_memory0_ram_dout0[378]), 
        .B(n21495), .Y(n12553) );
  sky130_fd_sc_hd__nand2_1 U19293 ( .A(j202_soc_core_memory0_ram_dout0[442]), 
        .B(n12156), .Y(n12554) );
  sky130_fd_sc_hd__nand2_1 U19294 ( .A(j202_soc_core_memory0_ram_dout0[474]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12555) );
  sky130_fd_sc_hd__nand2_1 U19296 ( .A(n20255), .B(n22232), .Y(n12558) );
  sky130_fd_sc_hd__nand2_1 U19297 ( .A(n12569), .B(n12568), .Y(n12559) );
  sky130_fd_sc_hd__nor2_1 U19298 ( .A(n25397), .B(n12566), .Y(n12562) );
  sky130_fd_sc_hd__nand2_1 U19299 ( .A(n12565), .B(n27785), .Y(n12563) );
  sky130_fd_sc_hd__nand2_1 U19300 ( .A(n12566), .B(n27786), .Y(n12564) );
  sky130_fd_sc_hd__nand3_1 U19301 ( .A(n12846), .B(n12845), .C(n12143), .Y(
        n12569) );
  sky130_fd_sc_hd__nand2b_1 U19302 ( .A_N(n11205), .B(n12570), .Y(n12568) );
  sky130_fd_sc_hd__nand2_1 U19303 ( .A(n20717), .B(n20716), .Y(n24090) );
  sky130_fd_sc_hd__or2_0 U19304 ( .A(n21934), .B(n20257), .X(n12570) );
  sky130_fd_sc_hd__nand2_1 U19305 ( .A(n20254), .B(n20253), .Y(n19236) );
  sky130_fd_sc_hd__nand2_1 U19306 ( .A(n11002), .B(n12332), .Y(n27886) );
  sky130_fd_sc_hd__nand2_1 U19307 ( .A(j202_soc_core_memory0_ram_dout0[63]), 
        .B(n21633), .Y(n12576) );
  sky130_fd_sc_hd__nand2_1 U19308 ( .A(j202_soc_core_memory0_ram_dout0[255]), 
        .B(n21641), .Y(n12578) );
  sky130_fd_sc_hd__nand2_1 U19309 ( .A(j202_soc_core_memory0_ram_dout0[223]), 
        .B(n21640), .Y(n12579) );
  sky130_fd_sc_hd__nand2_1 U19311 ( .A(n12583), .B(n23555), .Y(n25146) );
  sky130_fd_sc_hd__nand4_1 U19312 ( .A(n12589), .B(n12588), .C(n12587), .D(
        n12586), .Y(n12585) );
  sky130_fd_sc_hd__nand2_1 U19313 ( .A(j202_soc_core_memory0_ram_dout0[238]), 
        .B(n21641), .Y(n12586) );
  sky130_fd_sc_hd__nand2_1 U19314 ( .A(j202_soc_core_memory0_ram_dout0[14]), 
        .B(n21639), .Y(n12587) );
  sky130_fd_sc_hd__nand2_1 U19315 ( .A(j202_soc_core_memory0_ram_dout0[206]), 
        .B(n21640), .Y(n12588) );
  sky130_fd_sc_hd__nand2_1 U19316 ( .A(j202_soc_core_memory0_ram_dout0[334]), 
        .B(n21490), .Y(n12589) );
  sky130_fd_sc_hd__nand4_1 U19317 ( .A(n20094), .B(n12593), .C(n12592), .D(
        n12591), .Y(n12590) );
  sky130_fd_sc_hd__nand2_1 U19318 ( .A(j202_soc_core_memory0_ram_dout0[142]), 
        .B(n21489), .Y(n12591) );
  sky130_fd_sc_hd__nand2_1 U19319 ( .A(j202_soc_core_memory0_ram_dout0[398]), 
        .B(n21496), .Y(n12592) );
  sky130_fd_sc_hd__nand2_1 U19320 ( .A(j202_soc_core_memory0_ram_dout0[270]), 
        .B(n21634), .Y(n12593) );
  sky130_fd_sc_hd__nand4_1 U19321 ( .A(n12948), .B(n12949), .C(n20096), .D(
        n20095), .Y(n12595) );
  sky130_fd_sc_hd__nand4_1 U19322 ( .A(n20097), .B(n12946), .C(n12947), .D(
        n12950), .Y(n12596) );
  sky130_fd_sc_hd__nand2_1 U19323 ( .A(n12597), .B(n29488), .Y(n25904) );
  sky130_fd_sc_hd__nand2_1 U19324 ( .A(n12597), .B(n24127), .Y(n24111) );
  sky130_fd_sc_hd__o21ai_1 U19326 ( .A1(n12606), .A2(n12601), .B1(n20462), .Y(
        n12600) );
  sky130_fd_sc_hd__nand4_1 U19327 ( .A(n12605), .B(n12604), .C(n12603), .D(
        n12602), .Y(n12601) );
  sky130_fd_sc_hd__nand2_1 U19328 ( .A(j202_soc_core_memory0_ram_dout0[136]), 
        .B(n20456), .Y(n12602) );
  sky130_fd_sc_hd__nand2_1 U19329 ( .A(j202_soc_core_memory0_ram_dout0[232]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[7]), .Y(n12603) );
  sky130_fd_sc_hd__nand2_1 U19330 ( .A(j202_soc_core_memory0_ram_dout0[200]), 
        .B(n20455), .Y(n12604) );
  sky130_fd_sc_hd__nand2_1 U19331 ( .A(j202_soc_core_memory0_ram_dout0[104]), 
        .B(n20460), .Y(n12605) );
  sky130_fd_sc_hd__nand2_1 U19332 ( .A(j202_soc_core_memory0_ram_dout0[168]), 
        .B(n20459), .Y(n12607) );
  sky130_fd_sc_hd__nand2_1 U19333 ( .A(j202_soc_core_memory0_ram_dout0[8]), 
        .B(n20457), .Y(n12608) );
  sky130_fd_sc_hd__o21ai_1 U19334 ( .A1(n12615), .A2(n12610), .B1(n20454), .Y(
        n12609) );
  sky130_fd_sc_hd__nand4_1 U19335 ( .A(n12614), .B(n12613), .C(n12612), .D(
        n12611), .Y(n12610) );
  sky130_fd_sc_hd__nand2_1 U19336 ( .A(j202_soc_core_memory0_ram_dout0[392]), 
        .B(n21496), .Y(n12611) );
  sky130_fd_sc_hd__nand2_1 U19337 ( .A(j202_soc_core_memory0_ram_dout0[360]), 
        .B(n21495), .Y(n12612) );
  sky130_fd_sc_hd__nand2_1 U19338 ( .A(j202_soc_core_memory0_ram_dout0[424]), 
        .B(n12156), .Y(n12613) );
  sky130_fd_sc_hd__nand2_1 U19339 ( .A(j202_soc_core_memory0_ram_dout0[456]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12614) );
  sky130_fd_sc_hd__nand4_1 U19340 ( .A(n12619), .B(n12618), .C(n12617), .D(
        n12616), .Y(n12615) );
  sky130_fd_sc_hd__nand2_1 U19341 ( .A(j202_soc_core_memory0_ram_dout0[40]), 
        .B(n21633), .Y(n12616) );
  sky130_fd_sc_hd__nand2_1 U19342 ( .A(j202_soc_core_memory0_ram_dout0[296]), 
        .B(n21503), .Y(n12617) );
  sky130_fd_sc_hd__nand2_1 U19343 ( .A(j202_soc_core_memory0_ram_dout0[264]), 
        .B(n21634), .Y(n12618) );
  sky130_fd_sc_hd__nand2_1 U19344 ( .A(j202_soc_core_memory0_ram_dout0[328]), 
        .B(n21490), .Y(n12619) );
  sky130_fd_sc_hd__nor2_1 U19345 ( .A(n24574), .B(n27726), .Y(n12620) );
  sky130_fd_sc_hd__nand4_1 U19346 ( .A(n12150), .B(n28124), .C(n11005), .D(
        n28115), .Y(n28126) );
  sky130_fd_sc_hd__nand2_1 U19347 ( .A(n11536), .B(n26189), .Y(n26185) );
  sky130_fd_sc_hd__nand2_1 U19348 ( .A(n11536), .B(n25938), .Y(n25393) );
  sky130_fd_sc_hd__inv_1 U19349 ( .A(n27743), .Y(n12622) );
  sky130_fd_sc_hd__nand4_1 U19350 ( .A(n12629), .B(n12627), .C(n12626), .D(
        n12628), .Y(n20254) );
  sky130_fd_sc_hd__nand2_1 U19351 ( .A(n12625), .B(n20258), .Y(n12624) );
  sky130_fd_sc_hd__nand2_1 U19352 ( .A(n20253), .B(n21917), .Y(n12625) );
  sky130_fd_sc_hd__nand2_1 U19353 ( .A(n12742), .B(n17218), .Y(n12631) );
  sky130_fd_sc_hd__inv_1 U19355 ( .A(n12636), .Y(n12635) );
  sky130_fd_sc_hd__nand2_1 U19356 ( .A(n12638), .B(n12637), .Y(n12636) );
  sky130_fd_sc_hd__nand2_1 U19357 ( .A(j202_soc_core_memory0_ram_dout0[144]), 
        .B(n20456), .Y(n12637) );
  sky130_fd_sc_hd__nand2_1 U19358 ( .A(j202_soc_core_memory0_ram_dout0[240]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[7]), .Y(n12638) );
  sky130_fd_sc_hd__inv_1 U19359 ( .A(n12640), .Y(n12639) );
  sky130_fd_sc_hd__nand2_1 U19360 ( .A(n12642), .B(n12641), .Y(n12640) );
  sky130_fd_sc_hd__nand2_1 U19361 ( .A(j202_soc_core_memory0_ram_dout0[208]), 
        .B(n20455), .Y(n12641) );
  sky130_fd_sc_hd__nand2_1 U19362 ( .A(j202_soc_core_memory0_ram_dout0[112]), 
        .B(n20460), .Y(n12642) );
  sky130_fd_sc_hd__nand2_1 U19363 ( .A(j202_soc_core_memory0_ram_dout0[176]), 
        .B(n20459), .Y(n12645) );
  sky130_fd_sc_hd__nand2_1 U19364 ( .A(j202_soc_core_memory0_ram_dout0[16]), 
        .B(n20457), .Y(n12646) );
  sky130_fd_sc_hd__nand3_1 U19365 ( .A(n12834), .B(n20454), .C(n21917), .Y(
        n12649) );
  sky130_fd_sc_hd__nand2_1 U19366 ( .A(n12648), .B(n15174), .Y(n12647) );
  sky130_fd_sc_hd__nand2_1 U19367 ( .A(n12828), .B(n15094), .Y(n12648) );
  sky130_fd_sc_hd__nor2_1 U19368 ( .A(n11203), .B(n12651), .Y(n12650) );
  sky130_fd_sc_hd__nand2_1 U19369 ( .A(n12823), .B(n15094), .Y(n12655) );
  sky130_fd_sc_hd__inv_1 U19370 ( .A(n12658), .Y(n24410) );
  sky130_fd_sc_hd__nand2_1 U19371 ( .A(j202_soc_core_memory0_ram_dout0[443]), 
        .B(n12156), .Y(n12660) );
  sky130_fd_sc_hd__nand2_1 U19372 ( .A(j202_soc_core_memory0_ram_dout0[155]), 
        .B(n21489), .Y(n12661) );
  sky130_fd_sc_hd__nand2_1 U19373 ( .A(j202_soc_core_memory0_ram_dout0[187]), 
        .B(n21487), .Y(n12662) );
  sky130_fd_sc_hd__nand2_1 U19374 ( .A(j202_soc_core_memory0_ram_dout0[91]), 
        .B(n21642), .Y(n12663) );
  sky130_fd_sc_hd__nand2_1 U19375 ( .A(j202_soc_core_memory0_ram_dout0[354]), 
        .B(n21495), .Y(n12664) );
  sky130_fd_sc_hd__nand2_1 U19376 ( .A(n12666), .B(n12665), .Y(n17653) );
  sky130_fd_sc_hd__nand2_1 U19377 ( .A(n17612), .B(n12668), .Y(n12665) );
  sky130_fd_sc_hd__xnor3_1 U19379 ( .A(n12667), .B(n17611), .C(n17612), .X(
        n17616) );
  sky130_fd_sc_hd__inv_2 U19380 ( .A(n12964), .Y(n23553) );
  sky130_fd_sc_hd__xnor2_1 U19381 ( .A(n18614), .B(n12670), .Y(n17866) );
  sky130_fd_sc_hd__xnor2_1 U19382 ( .A(n18615), .B(n12678), .Y(n12670) );
  sky130_fd_sc_hd__xor2_1 U19383 ( .A(n18593), .B(n12671), .X(n18615) );
  sky130_fd_sc_hd__xnor2_1 U19384 ( .A(n12672), .B(n18591), .Y(n12671) );
  sky130_fd_sc_hd__nor2_1 U19385 ( .A(n24439), .B(n12673), .Y(n23487) );
  sky130_fd_sc_hd__nand2_1 U19386 ( .A(n12673), .B(n24452), .Y(n19095) );
  sky130_fd_sc_hd__nand4_1 U19387 ( .A(n24439), .B(n12673), .C(n23483), .D(
        n24453), .Y(n23461) );
  sky130_fd_sc_hd__nand2_1 U19388 ( .A(n12675), .B(n12674), .Y(n18649) );
  sky130_fd_sc_hd__nand2_1 U19389 ( .A(n12678), .B(n18615), .Y(n12674) );
  sky130_fd_sc_hd__nand2_1 U19390 ( .A(n18614), .B(n12676), .Y(n12675) );
  sky130_fd_sc_hd__nand2b_1 U19391 ( .A_N(n12678), .B(n12677), .Y(n12676) );
  sky130_fd_sc_hd__nand2_1 U19392 ( .A(n12679), .B(n17663), .Y(n12678) );
  sky130_fd_sc_hd__nand2_1 U19393 ( .A(n12681), .B(n12680), .Y(n17669) );
  sky130_fd_sc_hd__nand2_1 U19394 ( .A(n17637), .B(n17638), .Y(n12680) );
  sky130_fd_sc_hd__o21ai_1 U19395 ( .A1(n17638), .A2(n17637), .B1(n12683), .Y(
        n12681) );
  sky130_fd_sc_hd__xnor3_1 U19396 ( .A(n17638), .B(n12683), .C(n12682), .X(
        n17641) );
  sky130_fd_sc_hd__nand2_1 U19397 ( .A(n12685), .B(n22125), .Y(n12690) );
  sky130_fd_sc_hd__nand2_1 U19398 ( .A(n22238), .B(n22239), .Y(n12686) );
  sky130_fd_sc_hd__nand2_1 U19399 ( .A(n21846), .B(n21844), .Y(n12688) );
  sky130_fd_sc_hd__nand2_1 U19400 ( .A(n22240), .B(n12692), .Y(n12691) );
  sky130_fd_sc_hd__nand2_1 U19401 ( .A(n12688), .B(n21843), .Y(n12692) );
  sky130_fd_sc_hd__nand2_1 U19402 ( .A(n12689), .B(n18812), .Y(n21730) );
  sky130_fd_sc_hd__nand2_1 U19403 ( .A(n12690), .B(n12141), .Y(n12689) );
  sky130_fd_sc_hd__nand2_1 U19404 ( .A(n12691), .B(n22239), .Y(n22124) );
  sky130_fd_sc_hd__o22ai_1 U19405 ( .A1(n23077), .A2(n23085), .B1(n12696), 
        .B2(n12693), .Y(n23079) );
  sky130_fd_sc_hd__nand2_1 U19406 ( .A(n23133), .B(n23134), .Y(n12694) );
  sky130_fd_sc_hd__mux2i_1 U19407 ( .A0(n26739), .A1(n12695), .S(n27328), .Y(
        n23133) );
  sky130_fd_sc_hd__mux2i_1 U19408 ( .A0(n26736), .A1(n12697), .S(n27328), .Y(
        n23085) );
  sky130_fd_sc_hd__o21ai_1 U19409 ( .A1(n23136), .A2(n23259), .B1(n12702), .Y(
        n12699) );
  sky130_fd_sc_hd__nand3_1 U19410 ( .A(n12699), .B(n12700), .C(n12698), .Y(
        n23140) );
  sky130_fd_sc_hd__nand2_1 U19411 ( .A(n23259), .B(n23136), .Y(n12698) );
  sky130_fd_sc_hd__nand2_1 U19412 ( .A(n23150), .B(n23137), .Y(n12700) );
  sky130_fd_sc_hd__mux2i_1 U19413 ( .A0(n12701), .A1(n23113), .S(n27330), .Y(
        n23137) );
  sky130_fd_sc_hd__nand2_2 U19414 ( .A(n27331), .B(n23119), .Y(n27330) );
  sky130_fd_sc_hd__nand2_1 U19415 ( .A(n23256), .B(n23254), .Y(n12702) );
  sky130_fd_sc_hd__inv_2 U19416 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[0]), 
        .Y(n24677) );
  sky130_fd_sc_hd__nand3_1 U19417 ( .A(n12705), .B(n12709), .C(n12704), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N4) );
  sky130_fd_sc_hd__nand2_1 U19418 ( .A(n23377), .B(n12707), .Y(n12704) );
  sky130_fd_sc_hd__nand2_1 U19419 ( .A(n23377), .B(n12706), .Y(n27712) );
  sky130_fd_sc_hd__nand2_1 U19420 ( .A(n23376), .B(n12069), .Y(n12708) );
  sky130_fd_sc_hd__nand2_1 U19421 ( .A(n12711), .B(n23277), .Y(n23279) );
  sky130_fd_sc_hd__nand2_1 U19422 ( .A(n12712), .B(n23271), .Y(n12711) );
  sky130_fd_sc_hd__nand3_1 U19423 ( .A(n12715), .B(n12714), .C(n12713), .Y(
        n12712) );
  sky130_fd_sc_hd__nand2_1 U19424 ( .A(n23270), .B(n23281), .Y(n12713) );
  sky130_fd_sc_hd__nand2_1 U19425 ( .A(n23263), .B(n23349), .Y(n12714) );
  sky130_fd_sc_hd__o21ai_1 U19426 ( .A1(n23349), .A2(n23263), .B1(n23350), .Y(
        n12715) );
  sky130_fd_sc_hd__nand2_1 U19427 ( .A(n23394), .B(n12716), .Y(n27736) );
  sky130_fd_sc_hd__nand4_1 U19428 ( .A(n12987), .B(n12978), .C(n12983), .D(
        n12981), .Y(n12720) );
  sky130_fd_sc_hd__nor2_1 U19429 ( .A(n12720), .B(n12719), .Y(n12718) );
  sky130_fd_sc_hd__nand4_1 U19430 ( .A(n12739), .B(n12741), .C(n12979), .D(
        n12982), .Y(n12719) );
  sky130_fd_sc_hd__nor2_1 U19431 ( .A(n12723), .B(n12722), .Y(n12721) );
  sky130_fd_sc_hd__nand4_1 U19432 ( .A(n12986), .B(n12984), .C(n12985), .D(
        n12988), .Y(n12722) );
  sky130_fd_sc_hd__nand4_1 U19433 ( .A(n12738), .B(n12740), .C(n12980), .D(
        n12137), .Y(n12723) );
  sky130_fd_sc_hd__nand2_1 U19436 ( .A(n12730), .B(n25724), .Y(n24051) );
  sky130_fd_sc_hd__nand2_1 U19437 ( .A(n12730), .B(n28539), .Y(n28523) );
  sky130_fd_sc_hd__a22oi_1 U19438 ( .A1(n27125), .A2(n27862), .B1(n12730), 
        .B2(n27861), .Y(n27126) );
  sky130_fd_sc_hd__a22oi_1 U19439 ( .A1(n12730), .A2(n26929), .B1(n11442), 
        .B2(n26377), .Y(n26379) );
  sky130_fd_sc_hd__nand4_1 U19440 ( .A(n12882), .B(n12884), .C(n12883), .D(
        n19220), .Y(n20717) );
  sky130_fd_sc_hd__nand2_1 U19441 ( .A(j202_soc_core_memory0_ram_dout0[458]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12731) );
  sky130_fd_sc_hd__nand2_1 U19442 ( .A(j202_soc_core_memory0_ram_dout0[362]), 
        .B(n21495), .Y(n12732) );
  sky130_fd_sc_hd__nand2_1 U19443 ( .A(j202_soc_core_memory0_ram_dout0[202]), 
        .B(n21640), .Y(n12733) );
  sky130_fd_sc_hd__nand2_1 U19444 ( .A(j202_soc_core_memory0_ram_dout0[394]), 
        .B(n21496), .Y(n12734) );
  sky130_fd_sc_hd__nand2_1 U19445 ( .A(j202_soc_core_memory0_ram_dout0[266]), 
        .B(n21634), .Y(n12735) );
  sky130_fd_sc_hd__nand2_1 U19446 ( .A(j202_soc_core_memory0_ram_dout0[234]), 
        .B(n21641), .Y(n12736) );
  sky130_fd_sc_hd__nand2_1 U19447 ( .A(j202_soc_core_memory0_ram_dout0[106]), 
        .B(n21488), .Y(n12737) );
  sky130_fd_sc_hd__nand2_1 U19448 ( .A(j202_soc_core_memory0_ram_dout0[225]), 
        .B(n21641), .Y(n12738) );
  sky130_fd_sc_hd__nand2_1 U19449 ( .A(j202_soc_core_memory0_ram_dout0[385]), 
        .B(n21496), .Y(n12739) );
  sky130_fd_sc_hd__nand2_1 U19450 ( .A(j202_soc_core_memory0_ram_dout0[33]), 
        .B(n21633), .Y(n12740) );
  sky130_fd_sc_hd__nand2_1 U19451 ( .A(j202_soc_core_memory0_ram_dout0[449]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12741) );
  sky130_fd_sc_hd__nand2_1 U19452 ( .A(j202_soc_core_memory0_ram_dout0[226]), 
        .B(n21641), .Y(n12744) );
  sky130_fd_sc_hd__nand2_1 U19453 ( .A(j202_soc_core_memory0_ram_dout0[66]), 
        .B(n21642), .Y(n12745) );
  sky130_fd_sc_hd__nand2_1 U19454 ( .A(j202_soc_core_memory0_ram_dout0[258]), 
        .B(n21634), .Y(n12746) );
  sky130_fd_sc_hd__nand2_1 U19455 ( .A(j202_soc_core_memory0_ram_dout0[130]), 
        .B(n21489), .Y(n12747) );
  sky130_fd_sc_hd__nand2_1 U19456 ( .A(j202_soc_core_memory0_ram_dout0[322]), 
        .B(n21490), .Y(n12748) );
  sky130_fd_sc_hd__nand2_1 U19457 ( .A(j202_soc_core_memory0_ram_dout0[162]), 
        .B(n21487), .Y(n12749) );
  sky130_fd_sc_hd__nand2_1 U19458 ( .A(j202_soc_core_memory0_ram_dout0[98]), 
        .B(n21488), .Y(n12750) );
  sky130_fd_sc_hd__nand2_1 U19459 ( .A(j202_soc_core_memory0_ram_dout0[13]), 
        .B(n21639), .Y(n12752) );
  sky130_fd_sc_hd__nand2_1 U19460 ( .A(j202_soc_core_memory0_ram_dout0[141]), 
        .B(n21489), .Y(n12753) );
  sky130_fd_sc_hd__nand2_1 U19461 ( .A(j202_soc_core_memory0_ram_dout0[237]), 
        .B(n21641), .Y(n12754) );
  sky130_fd_sc_hd__nand2_1 U19462 ( .A(j202_soc_core_memory0_ram_dout0[77]), 
        .B(n21642), .Y(n12755) );
  sky130_fd_sc_hd__o21ai_1 U19463 ( .A1(n12758), .A2(n12757), .B1(n20462), .Y(
        n12756) );
  sky130_fd_sc_hd__nand4_1 U19464 ( .A(n16202), .B(n16201), .C(n16200), .D(
        n16203), .Y(n12757) );
  sky130_fd_sc_hd__nand2_1 U19465 ( .A(j202_soc_core_memory0_ram_dout0[205]), 
        .B(n21640), .Y(n12760) );
  sky130_fd_sc_hd__nand2_1 U19466 ( .A(j202_soc_core_memory0_ram_dout0[45]), 
        .B(n21633), .Y(n12761) );
  sky130_fd_sc_hd__nand2_1 U19467 ( .A(j202_soc_core_memory0_ram_dout0[173]), 
        .B(n21487), .Y(n12762) );
  sky130_fd_sc_hd__nand2_1 U19468 ( .A(j202_soc_core_memory0_ram_dout0[109]), 
        .B(n21488), .Y(n12763) );
  sky130_fd_sc_hd__nand2_1 U19469 ( .A(j202_soc_core_memory0_ram_dout0[94]), 
        .B(n20458), .Y(n12765) );
  sky130_fd_sc_hd__nand2_1 U19470 ( .A(j202_soc_core_memory0_ram_dout0[222]), 
        .B(n20455), .Y(n12766) );
  sky130_fd_sc_hd__nand2_1 U19471 ( .A(j202_soc_core_memory0_ram_dout0[190]), 
        .B(n20459), .Y(n12767) );
  sky130_fd_sc_hd__nand3_1 U19472 ( .A(n11092), .B(n12945), .C(n24622), .Y(
        n24626) );
  sky130_fd_sc_hd__and2_0 U19473 ( .A(n21917), .B(n21650), .X(n12771) );
  sky130_fd_sc_hd__nand2_1 U19474 ( .A(j202_soc_core_memory0_ram_dout0[49]), 
        .B(n21633), .Y(n12772) );
  sky130_fd_sc_hd__nand2_1 U19475 ( .A(j202_soc_core_memory0_ram_dout0[305]), 
        .B(n21503), .Y(n12773) );
  sky130_fd_sc_hd__nand2_1 U19476 ( .A(j202_soc_core_memory0_ram_dout0[273]), 
        .B(n21634), .Y(n12774) );
  sky130_fd_sc_hd__nand2_1 U19477 ( .A(j202_soc_core_memory0_ram_dout0[337]), 
        .B(n21490), .Y(n12775) );
  sky130_fd_sc_hd__inv_1 U19478 ( .A(n12778), .Y(n23603) );
  sky130_fd_sc_hd__inv_1 U19479 ( .A(n12779), .Y(n12780) );
  sky130_fd_sc_hd__o21ai_1 U19480 ( .A1(n12789), .A2(n12784), .B1(n20462), .Y(
        n12783) );
  sky130_fd_sc_hd__nand4_1 U19481 ( .A(n12788), .B(n12787), .C(n12786), .D(
        n12785), .Y(n12784) );
  sky130_fd_sc_hd__nand2_1 U19482 ( .A(j202_soc_core_memory0_ram_dout0[152]), 
        .B(n20456), .Y(n12785) );
  sky130_fd_sc_hd__nand2_1 U19483 ( .A(j202_soc_core_memory0_ram_dout0[248]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[7]), .Y(n12786) );
  sky130_fd_sc_hd__nand2_1 U19484 ( .A(j202_soc_core_memory0_ram_dout0[216]), 
        .B(n20455), .Y(n12787) );
  sky130_fd_sc_hd__nand2_1 U19485 ( .A(j202_soc_core_memory0_ram_dout0[120]), 
        .B(n20460), .Y(n12788) );
  sky130_fd_sc_hd__nand2_1 U19486 ( .A(j202_soc_core_memory0_ram_dout0[184]), 
        .B(n20459), .Y(n12790) );
  sky130_fd_sc_hd__nand2_1 U19487 ( .A(j202_soc_core_memory0_ram_dout0[24]), 
        .B(n20457), .Y(n12791) );
  sky130_fd_sc_hd__nand4_1 U19488 ( .A(n12797), .B(n12796), .C(n12795), .D(
        n12794), .Y(n12793) );
  sky130_fd_sc_hd__nand2_1 U19489 ( .A(j202_soc_core_memory0_ram_dout0[408]), 
        .B(n21496), .Y(n12794) );
  sky130_fd_sc_hd__nand2_1 U19490 ( .A(j202_soc_core_memory0_ram_dout0[376]), 
        .B(n21495), .Y(n12795) );
  sky130_fd_sc_hd__nand2_1 U19491 ( .A(j202_soc_core_memory0_ram_dout0[440]), 
        .B(n12156), .Y(n12796) );
  sky130_fd_sc_hd__nand2_1 U19492 ( .A(j202_soc_core_memory0_ram_dout0[472]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12797) );
  sky130_fd_sc_hd__nand2_1 U19493 ( .A(n21690), .B(n12138), .Y(n12799) );
  sky130_fd_sc_hd__nand2_1 U19494 ( .A(n12800), .B(n12801), .Y(n20948) );
  sky130_fd_sc_hd__nand2_1 U19495 ( .A(j202_soc_core_memory0_ram_dout0[178]), 
        .B(n20459), .Y(n12804) );
  sky130_fd_sc_hd__nand2_1 U19496 ( .A(j202_soc_core_memory0_ram_dout0[18]), 
        .B(n20457), .Y(n12805) );
  sky130_fd_sc_hd__nand2_1 U19497 ( .A(j202_soc_core_memory0_ram_dout0[402]), 
        .B(n21496), .Y(n12807) );
  sky130_fd_sc_hd__nand2_1 U19498 ( .A(j202_soc_core_memory0_ram_dout0[434]), 
        .B(n12156), .Y(n12808) );
  sky130_fd_sc_hd__nand2_1 U19499 ( .A(j202_soc_core_memory0_ram_dout0[466]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12809) );
  sky130_fd_sc_hd__nand4_1 U19500 ( .A(n12814), .B(n12813), .C(n12812), .D(
        n12811), .Y(n12810) );
  sky130_fd_sc_hd__nand2_1 U19501 ( .A(j202_soc_core_memory0_ram_dout0[50]), 
        .B(n21633), .Y(n12811) );
  sky130_fd_sc_hd__nand2_1 U19502 ( .A(j202_soc_core_memory0_ram_dout0[306]), 
        .B(n21503), .Y(n12812) );
  sky130_fd_sc_hd__nand2_1 U19503 ( .A(j202_soc_core_memory0_ram_dout0[274]), 
        .B(n21634), .Y(n12813) );
  sky130_fd_sc_hd__nand2_1 U19504 ( .A(j202_soc_core_memory0_ram_dout0[338]), 
        .B(n21490), .Y(n12814) );
  sky130_fd_sc_hd__inv_2 U19505 ( .A(n24564), .Y(n23604) );
  sky130_fd_sc_hd__nand3_1 U19506 ( .A(n12055), .B(n30198), .C(n20949), .Y(
        n22224) );
  sky130_fd_sc_hd__nand2_1 U19507 ( .A(n12820), .B(n12818), .Y(n24592) );
  sky130_fd_sc_hd__nand2_1 U19508 ( .A(n11395), .B(n27743), .Y(n12819) );
  sky130_fd_sc_hd__nand2_1 U19509 ( .A(n24575), .B(n12821), .Y(n24577) );
  sky130_fd_sc_hd__nand2_1 U19510 ( .A(n28142), .B(n12128), .Y(n23960) );
  sky130_fd_sc_hd__nand4_1 U19511 ( .A(n12827), .B(n12826), .C(n12825), .D(
        n12824), .Y(n12823) );
  sky130_fd_sc_hd__nand2_1 U19512 ( .A(j202_soc_core_memory0_ram_dout0[150]), 
        .B(n20456), .Y(n12824) );
  sky130_fd_sc_hd__nand2_1 U19513 ( .A(j202_soc_core_memory0_ram_dout0[246]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[7]), .Y(n12825) );
  sky130_fd_sc_hd__nand2_1 U19514 ( .A(j202_soc_core_memory0_ram_dout0[214]), 
        .B(n20455), .Y(n12826) );
  sky130_fd_sc_hd__nand2_1 U19515 ( .A(j202_soc_core_memory0_ram_dout0[118]), 
        .B(n20460), .Y(n12827) );
  sky130_fd_sc_hd__nand2_1 U19516 ( .A(j202_soc_core_memory0_ram_dout0[182]), 
        .B(n20459), .Y(n12829) );
  sky130_fd_sc_hd__nand2_1 U19517 ( .A(j202_soc_core_memory0_ram_dout0[22]), 
        .B(n20457), .Y(n12830) );
  sky130_fd_sc_hd__nand2_1 U19518 ( .A(j202_soc_core_memory0_ram_dout0[374]), 
        .B(n21495), .Y(n12831) );
  sky130_fd_sc_hd__nand2_1 U19519 ( .A(j202_soc_core_memory0_ram_dout0[438]), 
        .B(n12156), .Y(n12832) );
  sky130_fd_sc_hd__nand2_1 U19520 ( .A(j202_soc_core_memory0_ram_dout0[470]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12833) );
  sky130_fd_sc_hd__nand4_1 U19521 ( .A(n12838), .B(n12837), .C(n12836), .D(
        n12835), .Y(n12834) );
  sky130_fd_sc_hd__nand2_1 U19522 ( .A(j202_soc_core_memory0_ram_dout0[54]), 
        .B(n21633), .Y(n12835) );
  sky130_fd_sc_hd__nand2_1 U19523 ( .A(j202_soc_core_memory0_ram_dout0[310]), 
        .B(n21503), .Y(n12836) );
  sky130_fd_sc_hd__nand2_1 U19524 ( .A(j202_soc_core_memory0_ram_dout0[278]), 
        .B(n21634), .Y(n12837) );
  sky130_fd_sc_hd__nand2_1 U19525 ( .A(j202_soc_core_memory0_ram_dout0[342]), 
        .B(n21490), .Y(n12838) );
  sky130_fd_sc_hd__nand3_1 U19526 ( .A(n16959), .B(n16963), .C(n12118), .Y(
        n16942) );
  sky130_fd_sc_hd__nand2b_1 U19527 ( .A_N(n16356), .B(n19129), .Y(n16677) );
  sky130_fd_sc_hd__nand2_1 U19528 ( .A(n19816), .B(n17250), .Y(n16356) );
  sky130_fd_sc_hd__nand2_1 U19529 ( .A(n21146), .B(n19119), .Y(n16959) );
  sky130_fd_sc_hd__nand2_1 U19530 ( .A(n18752), .B(n21088), .Y(n15676) );
  sky130_fd_sc_hd__nand2_1 U19531 ( .A(n19119), .B(n14597), .Y(n16206) );
  sky130_fd_sc_hd__nand2_1 U19532 ( .A(n18764), .B(n14597), .Y(n18700) );
  sky130_fd_sc_hd__nand2_1 U19533 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .B(n14597), .Y(n16207) );
  sky130_fd_sc_hd__nand2_1 U19534 ( .A(n13179), .B(n14597), .Y(n18730) );
  sky130_fd_sc_hd__nand2_1 U19535 ( .A(n19124), .B(n14597), .Y(n15759) );
  sky130_fd_sc_hd__nand2_1 U19536 ( .A(n17271), .B(n14597), .Y(n21593) );
  sky130_fd_sc_hd__nand2_1 U19537 ( .A(n17285), .B(n14597), .Y(n21354) );
  sky130_fd_sc_hd__nand2_1 U19538 ( .A(n17272), .B(n14597), .Y(n21554) );
  sky130_fd_sc_hd__nand2_1 U19539 ( .A(n21613), .B(n14597), .Y(n21521) );
  sky130_fd_sc_hd__nand2_1 U19540 ( .A(n21142), .B(n14597), .Y(n21399) );
  sky130_fd_sc_hd__nand2_1 U19541 ( .A(n16634), .B(n14597), .Y(n16689) );
  sky130_fd_sc_hd__nand2_1 U19542 ( .A(n20033), .B(n12839), .Y(n20035) );
  sky130_fd_sc_hd__nor2_1 U19543 ( .A(n12843), .B(n12842), .Y(n29644) );
  sky130_fd_sc_hd__nand2_1 U19544 ( .A(n26158), .B(n22739), .Y(n16907) );
  sky130_fd_sc_hd__nand2_1 U19545 ( .A(n16886), .B(n20462), .Y(n12845) );
  sky130_fd_sc_hd__nand2_1 U19546 ( .A(n12240), .B(n24547), .Y(n23391) );
  sky130_fd_sc_hd__nand3_1 U19547 ( .A(n12240), .B(n24544), .C(n28029), .Y(
        n24557) );
  sky130_fd_sc_hd__nand2_1 U19548 ( .A(j202_soc_core_memory0_ram_dout0[126]), 
        .B(n20460), .Y(n12848) );
  sky130_fd_sc_hd__nand2_1 U19549 ( .A(j202_soc_core_memory0_ram_dout0[158]), 
        .B(n20456), .Y(n12849) );
  sky130_fd_sc_hd__nand2_1 U19550 ( .A(j202_soc_core_memory0_ram_dout0[30]), 
        .B(n20457), .Y(n12850) );
  sky130_fd_sc_hd__nand2_1 U19551 ( .A(j202_soc_core_memory0_ram_dout0[254]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[7]), .Y(n12851) );
  sky130_fd_sc_hd__nand2_1 U19553 ( .A(j202_soc_core_memory0_ram_dout0[145]), 
        .B(n20456), .Y(n12853) );
  sky130_fd_sc_hd__nand2_1 U19554 ( .A(j202_soc_core_memory0_ram_dout0[241]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[7]), .Y(n12854) );
  sky130_fd_sc_hd__nand2_1 U19556 ( .A(j202_soc_core_memory0_ram_dout0[209]), 
        .B(n20455), .Y(n12856) );
  sky130_fd_sc_hd__nand2_1 U19557 ( .A(j202_soc_core_memory0_ram_dout0[113]), 
        .B(n20460), .Y(n12857) );
  sky130_fd_sc_hd__nand3_1 U19558 ( .A(n19431), .B(n12860), .C(n12859), .Y(
        n12858) );
  sky130_fd_sc_hd__nand2_1 U19559 ( .A(j202_soc_core_memory0_ram_dout0[177]), 
        .B(n20459), .Y(n12859) );
  sky130_fd_sc_hd__nand2_1 U19560 ( .A(j202_soc_core_memory0_ram_dout0[17]), 
        .B(n20457), .Y(n12860) );
  sky130_fd_sc_hd__nand2_1 U19561 ( .A(j202_soc_core_memory0_ram_dout0[275]), 
        .B(n21634), .Y(n12863) );
  sky130_fd_sc_hd__nand2_1 U19562 ( .A(j202_soc_core_memory0_ram_dout0[467]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12864) );
  sky130_fd_sc_hd__nand2_1 U19563 ( .A(j202_soc_core_memory0_ram_dout0[211]), 
        .B(n21640), .Y(n12865) );
  sky130_fd_sc_hd__nand2_1 U19564 ( .A(j202_soc_core_memory0_ram_dout0[435]), 
        .B(n12156), .Y(n12866) );
  sky130_fd_sc_hd__nand2_1 U19565 ( .A(j202_soc_core_memory0_ram_dout0[115]), 
        .B(n21488), .Y(n12867) );
  sky130_fd_sc_hd__nand2_1 U19566 ( .A(j202_soc_core_memory0_ram_dout0[51]), 
        .B(n21633), .Y(n12868) );
  sky130_fd_sc_hd__nand2_1 U19567 ( .A(j202_soc_core_memory0_ram_dout0[371]), 
        .B(n21495), .Y(n12869) );
  sky130_fd_sc_hd__nand2_1 U19568 ( .A(j202_soc_core_memory0_ram_dout0[403]), 
        .B(n21496), .Y(n12870) );
  sky130_fd_sc_hd__nand2_1 U19569 ( .A(j202_soc_core_memory0_ram_dout0[83]), 
        .B(n21642), .Y(n12871) );
  sky130_fd_sc_hd__nand2_1 U19570 ( .A(j202_soc_core_memory0_ram_dout0[147]), 
        .B(n21489), .Y(n12872) );
  sky130_fd_sc_hd__nand2_1 U19571 ( .A(j202_soc_core_memory0_ram_dout0[179]), 
        .B(n21487), .Y(n12873) );
  sky130_fd_sc_hd__nand3_4 U19572 ( .A(n12880), .B(n12876), .C(n12875), .Y(
        n29587) );
  sky130_fd_sc_hd__nand2_1 U19573 ( .A(n12878), .B(n12881), .Y(n12877) );
  sky130_fd_sc_hd__nand2_1 U19574 ( .A(n16886), .B(n12879), .Y(n12878) );
  sky130_fd_sc_hd__o21a_1 U19575 ( .A1(n11203), .A2(n16887), .B1(n20718), .X(
        n12881) );
  sky130_fd_sc_hd__nand4_1 U19576 ( .A(n23484), .B(n23485), .C(n27362), .D(
        n25890), .Y(n23462) );
  sky130_fd_sc_hd__nand2_1 U19578 ( .A(n12889), .B(n12888), .Y(n18267) );
  sky130_fd_sc_hd__nand2_1 U19579 ( .A(n18243), .B(n18244), .Y(n12888) );
  sky130_fd_sc_hd__xnor2_1 U19580 ( .A(n18242), .B(n12890), .Y(n18256) );
  sky130_fd_sc_hd__xnor2_1 U19581 ( .A(n18244), .B(n18243), .Y(n12890) );
  sky130_fd_sc_hd__xor2_1 U19582 ( .A(n12891), .B(n18223), .X(n18237) );
  sky130_fd_sc_hd__nand2_1 U19583 ( .A(n23036), .B(n19086), .Y(n12892) );
  sky130_fd_sc_hd__nand2_1 U19584 ( .A(n25775), .B(n23044), .Y(n12894) );
  sky130_fd_sc_hd__and2_0 U19585 ( .A(n19096), .B(n19097), .X(n12895) );
  sky130_fd_sc_hd__nand4_1 U19586 ( .A(n12901), .B(n12900), .C(n12899), .D(
        n12898), .Y(n12897) );
  sky130_fd_sc_hd__nand2_1 U19587 ( .A(j202_soc_core_memory0_ram_dout0[215]), 
        .B(n21640), .Y(n12898) );
  sky130_fd_sc_hd__nand2_1 U19588 ( .A(j202_soc_core_memory0_ram_dout0[119]), 
        .B(n21488), .Y(n12899) );
  sky130_fd_sc_hd__nand2_1 U19589 ( .A(j202_soc_core_memory0_ram_dout0[151]), 
        .B(n21489), .Y(n12900) );
  sky130_fd_sc_hd__nand2_1 U19590 ( .A(j202_soc_core_memory0_ram_dout0[87]), 
        .B(n21642), .Y(n12901) );
  sky130_fd_sc_hd__nand4_1 U19591 ( .A(n12907), .B(n12906), .C(n12904), .D(
        n12905), .Y(n12903) );
  sky130_fd_sc_hd__nand2_1 U19592 ( .A(j202_soc_core_memory0_ram_dout0[279]), 
        .B(n21634), .Y(n12904) );
  sky130_fd_sc_hd__nand2_1 U19593 ( .A(j202_soc_core_memory0_ram_dout0[407]), 
        .B(n21496), .Y(n12905) );
  sky130_fd_sc_hd__nand2_1 U19594 ( .A(j202_soc_core_memory0_ram_dout0[439]), 
        .B(n12156), .Y(n12906) );
  sky130_fd_sc_hd__nand2_1 U19595 ( .A(j202_soc_core_memory0_ram_dout0[471]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12907) );
  sky130_fd_sc_hd__nand4_1 U19596 ( .A(n12910), .B(n12912), .C(n12911), .D(
        n30028), .Y(n12908) );
  sky130_fd_sc_hd__nand2_1 U19597 ( .A(j202_soc_core_memory0_ram_dout0[343]), 
        .B(n21490), .Y(n12910) );
  sky130_fd_sc_hd__nand2_1 U19598 ( .A(j202_soc_core_memory0_ram_dout0[311]), 
        .B(n21503), .Y(n12911) );
  sky130_fd_sc_hd__nand2_1 U19599 ( .A(j202_soc_core_memory0_ram_dout0[375]), 
        .B(n21495), .Y(n12912) );
  sky130_fd_sc_hd__and2_0 U19600 ( .A(n22381), .B(n22380), .X(n12913) );
  sky130_fd_sc_hd__inv_2 U19601 ( .A(n12914), .Y(n24682) );
  sky130_fd_sc_hd__nand3_1 U19602 ( .A(n12916), .B(n18854), .C(n12915), .Y(
        n12914) );
  sky130_fd_sc_hd__nand2_1 U19603 ( .A(n12360), .B(n18853), .Y(n12915) );
  sky130_fd_sc_hd__nand2_1 U19604 ( .A(n12917), .B(n18807), .Y(n12916) );
  sky130_fd_sc_hd__nor2_1 U19605 ( .A(n12918), .B(n12361), .Y(n12917) );
  sky130_fd_sc_hd__nand2_1 U19606 ( .A(n24879), .B(n27786), .Y(n12918) );
  sky130_fd_sc_hd__nand2_1 U19607 ( .A(n30057), .B(n20454), .Y(n12919) );
  sky130_fd_sc_hd__nand2_1 U19608 ( .A(n12922), .B(n27745), .Y(n24581) );
  sky130_fd_sc_hd__o21ai_1 U19610 ( .A1(n12930), .A2(n12935), .B1(n20454), .Y(
        n20588) );
  sky130_fd_sc_hd__nand3_1 U19611 ( .A(n12928), .B(n20587), .C(n12927), .Y(
        n12952) );
  sky130_fd_sc_hd__nand2_1 U19612 ( .A(n12930), .B(n12929), .Y(n12927) );
  sky130_fd_sc_hd__nand2_1 U19613 ( .A(n12935), .B(n12929), .Y(n12928) );
  sky130_fd_sc_hd__and2_0 U19614 ( .A(n20454), .B(n21917), .X(n12929) );
  sky130_fd_sc_hd__nand4_1 U19615 ( .A(n12934), .B(n12933), .C(n12932), .D(
        n12931), .Y(n12930) );
  sky130_fd_sc_hd__nand2_1 U19616 ( .A(j202_soc_core_memory0_ram_dout0[409]), 
        .B(n21496), .Y(n12931) );
  sky130_fd_sc_hd__nand2_1 U19617 ( .A(j202_soc_core_memory0_ram_dout0[377]), 
        .B(n21495), .Y(n12932) );
  sky130_fd_sc_hd__nand2_1 U19618 ( .A(j202_soc_core_memory0_ram_dout0[441]), 
        .B(n12156), .Y(n12933) );
  sky130_fd_sc_hd__nand2_1 U19619 ( .A(j202_soc_core_memory0_ram_dout0[473]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12934) );
  sky130_fd_sc_hd__nand4_1 U19620 ( .A(n12939), .B(n12938), .C(n12937), .D(
        n12936), .Y(n12935) );
  sky130_fd_sc_hd__nand2_1 U19621 ( .A(j202_soc_core_memory0_ram_dout0[57]), 
        .B(n21633), .Y(n12936) );
  sky130_fd_sc_hd__nand2_1 U19622 ( .A(j202_soc_core_memory0_ram_dout0[281]), 
        .B(n21634), .Y(n12938) );
  sky130_fd_sc_hd__nand2_1 U19623 ( .A(n23435), .B(n30132), .Y(n23436) );
  sky130_fd_sc_hd__nand2_1 U19624 ( .A(n28091), .B(n30132), .Y(n27745) );
  sky130_fd_sc_hd__nand2_1 U19625 ( .A(n27980), .B(n12942), .Y(n24566) );
  sky130_fd_sc_hd__inv_2 U19626 ( .A(n24106), .Y(n12942) );
  sky130_fd_sc_hd__inv_1 U19627 ( .A(n24617), .Y(n12944) );
  sky130_fd_sc_hd__nand2_1 U19628 ( .A(j202_soc_core_memory0_ram_dout0[462]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12946) );
  sky130_fd_sc_hd__nand2_1 U19629 ( .A(j202_soc_core_memory0_ram_dout0[366]), 
        .B(n21495), .Y(n12947) );
  sky130_fd_sc_hd__nand2_1 U19630 ( .A(j202_soc_core_memory0_ram_dout0[430]), 
        .B(n12156), .Y(n12948) );
  sky130_fd_sc_hd__nand2_1 U19631 ( .A(j202_soc_core_memory0_ram_dout0[110]), 
        .B(n21488), .Y(n12949) );
  sky130_fd_sc_hd__and3_1 U19632 ( .A(n20241), .B(n20246), .C(n20249), .X(
        n12950) );
  sky130_fd_sc_hd__o21a_1 U19633 ( .A1(n12557), .A2(n13033), .B1(n21692), .X(
        n12955) );
  sky130_fd_sc_hd__nand2_1 U19634 ( .A(j202_soc_core_memory0_ram_dout0[32]), 
        .B(n21633), .Y(n12956) );
  sky130_fd_sc_hd__nand2_1 U19635 ( .A(j202_soc_core_memory0_ram_dout0[320]), 
        .B(n21490), .Y(n12957) );
  sky130_fd_sc_hd__nand2_1 U19636 ( .A(j202_soc_core_memory0_ram_dout0[256]), 
        .B(n21634), .Y(n12958) );
  sky130_fd_sc_hd__nand2_1 U19637 ( .A(j202_soc_core_memory0_ram_dout0[384]), 
        .B(n21496), .Y(n12959) );
  sky130_fd_sc_hd__nand2_1 U19638 ( .A(j202_soc_core_memory0_ram_dout0[224]), 
        .B(n21641), .Y(n12960) );
  sky130_fd_sc_hd__nand2_1 U19639 ( .A(j202_soc_core_memory0_ram_dout0[416]), 
        .B(n12156), .Y(n12961) );
  sky130_fd_sc_hd__nand2_1 U19640 ( .A(j202_soc_core_memory0_ram_dout0[352]), 
        .B(n21495), .Y(n12962) );
  sky130_fd_sc_hd__nand2_1 U19641 ( .A(j202_soc_core_memory0_ram_dout0[448]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12963) );
  sky130_fd_sc_hd__nand2_1 U19642 ( .A(n12965), .B(n12327), .Y(n27747) );
  sky130_fd_sc_hd__a21oi_1 U19643 ( .A1(n11423), .A2(n11175), .B1(n12966), .Y(
        n12965) );
  sky130_fd_sc_hd__nand3_1 U19644 ( .A(n12297), .B(n12972), .C(n12973), .Y(
        n12967) );
  sky130_fd_sc_hd__nand3_1 U19646 ( .A(n12971), .B(n30194), .C(n30020), .Y(
        n21176) );
  sky130_fd_sc_hd__nand3_1 U19647 ( .A(n12974), .B(n12973), .C(n12972), .Y(
        n20720) );
  sky130_fd_sc_hd__inv_1 U19648 ( .A(n16109), .Y(n12972) );
  sky130_fd_sc_hd__nand2_1 U19651 ( .A(j202_soc_core_memory0_ram_dout0[65]), 
        .B(n21642), .Y(n12978) );
  sky130_fd_sc_hd__nand2_1 U19652 ( .A(j202_soc_core_memory0_ram_dout0[193]), 
        .B(n21640), .Y(n12979) );
  sky130_fd_sc_hd__nand2_1 U19653 ( .A(j202_soc_core_memory0_ram_dout0[97]), 
        .B(n21488), .Y(n12980) );
  sky130_fd_sc_hd__nand2_1 U19654 ( .A(j202_soc_core_memory0_ram_dout0[321]), 
        .B(n21490), .Y(n12981) );
  sky130_fd_sc_hd__nand2_1 U19655 ( .A(j202_soc_core_memory0_ram_dout0[257]), 
        .B(n21634), .Y(n12982) );
  sky130_fd_sc_hd__nand2_1 U19656 ( .A(j202_soc_core_memory0_ram_dout0[417]), 
        .B(n12156), .Y(n12983) );
  sky130_fd_sc_hd__nand2_1 U19657 ( .A(j202_soc_core_memory0_ram_dout0[353]), 
        .B(n21495), .Y(n12984) );
  sky130_fd_sc_hd__nand2_1 U19658 ( .A(j202_soc_core_memory0_ram_dout0[161]), 
        .B(n21487), .Y(n12985) );
  sky130_fd_sc_hd__nand2_1 U19659 ( .A(j202_soc_core_memory0_ram_dout0[1]), 
        .B(n21639), .Y(n12986) );
  sky130_fd_sc_hd__nand2_1 U19660 ( .A(j202_soc_core_memory0_ram_dout0[289]), 
        .B(n21503), .Y(n12987) );
  sky130_fd_sc_hd__nand2_1 U19661 ( .A(j202_soc_core_memory0_ram_dout0[129]), 
        .B(n21489), .Y(n12988) );
  sky130_fd_sc_hd__nand3_2 U19662 ( .A(n24560), .B(n23426), .C(n23955), .Y(
        n12989) );
  sky130_fd_sc_hd__nand2_1 U19663 ( .A(j202_soc_core_memory0_ram_dout0[414]), 
        .B(n21496), .Y(n12991) );
  sky130_fd_sc_hd__nand2_1 U19664 ( .A(j202_soc_core_memory0_ram_dout0[382]), 
        .B(n21495), .Y(n12992) );
  sky130_fd_sc_hd__nand2_1 U19665 ( .A(j202_soc_core_memory0_ram_dout0[446]), 
        .B(n12156), .Y(n12993) );
  sky130_fd_sc_hd__nand2_1 U19666 ( .A(j202_soc_core_memory0_ram_dout0[478]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12994) );
  sky130_fd_sc_hd__nand2_1 U19667 ( .A(j202_soc_core_memory0_ram_dout0[62]), 
        .B(n21633), .Y(n12996) );
  sky130_fd_sc_hd__nand2_1 U19668 ( .A(j202_soc_core_memory0_ram_dout0[318]), 
        .B(n21503), .Y(n12997) );
  sky130_fd_sc_hd__nand2_1 U19669 ( .A(j202_soc_core_memory0_ram_dout0[286]), 
        .B(n21634), .Y(n12998) );
  sky130_fd_sc_hd__nand2_1 U19670 ( .A(j202_soc_core_memory0_ram_dout0[350]), 
        .B(n21490), .Y(n12999) );
  sky130_fd_sc_hd__and3_1 U19671 ( .A(n15770), .B(n15778), .C(n15780), .X(
        n13000) );
  sky130_fd_sc_hd__nand4_1 U19672 ( .A(n13004), .B(n13005), .C(n13006), .D(
        n13003), .Y(n13002) );
  sky130_fd_sc_hd__nand2_1 U19673 ( .A(j202_soc_core_memory0_ram_dout0[373]), 
        .B(n21495), .Y(n13003) );
  sky130_fd_sc_hd__nand2_1 U19674 ( .A(j202_soc_core_memory0_ram_dout0[469]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n13004) );
  sky130_fd_sc_hd__nand2_1 U19675 ( .A(j202_soc_core_memory0_ram_dout0[341]), 
        .B(n21490), .Y(n13005) );
  sky130_fd_sc_hd__nand2_1 U19676 ( .A(j202_soc_core_memory0_ram_dout0[277]), 
        .B(n21634), .Y(n13006) );
  sky130_fd_sc_hd__nand4_1 U19677 ( .A(n13009), .B(n13011), .C(n13010), .D(
        n13008), .Y(n13007) );
  sky130_fd_sc_hd__nand2_1 U19678 ( .A(j202_soc_core_memory0_ram_dout0[405]), 
        .B(n21496), .Y(n13009) );
  sky130_fd_sc_hd__nand2_1 U19679 ( .A(j202_soc_core_memory0_ram_dout0[21]), 
        .B(n21639), .Y(n13010) );
  sky130_fd_sc_hd__nand2_1 U19680 ( .A(j202_soc_core_memory0_ram_dout0[437]), 
        .B(n12156), .Y(n13011) );
  sky130_fd_sc_hd__nand4_1 U19681 ( .A(n13017), .B(n13016), .C(n13014), .D(
        n13015), .Y(n13013) );
  sky130_fd_sc_hd__nand2_1 U19682 ( .A(j202_soc_core_memory0_ram_dout0[53]), 
        .B(n21633), .Y(n13014) );
  sky130_fd_sc_hd__nand2_1 U19683 ( .A(j202_soc_core_memory0_ram_dout0[181]), 
        .B(n21487), .Y(n13015) );
  sky130_fd_sc_hd__nand2_1 U19684 ( .A(j202_soc_core_memory0_ram_dout0[245]), 
        .B(n21641), .Y(n13016) );
  sky130_fd_sc_hd__nand2_1 U19685 ( .A(j202_soc_core_memory0_ram_dout0[309]), 
        .B(n21503), .Y(n13017) );
  sky130_fd_sc_hd__nand4_1 U19686 ( .A(n13022), .B(n13021), .C(n13020), .D(
        n13019), .Y(n13018) );
  sky130_fd_sc_hd__nand2_1 U19687 ( .A(j202_soc_core_memory0_ram_dout0[149]), 
        .B(n21489), .Y(n13019) );
  sky130_fd_sc_hd__nand2_1 U19688 ( .A(j202_soc_core_memory0_ram_dout0[85]), 
        .B(n21642), .Y(n13020) );
  sky130_fd_sc_hd__nand2_1 U19689 ( .A(j202_soc_core_memory0_ram_dout0[213]), 
        .B(n21640), .Y(n13021) );
  sky130_fd_sc_hd__nand2_1 U19690 ( .A(j202_soc_core_memory0_ram_dout0[117]), 
        .B(n21488), .Y(n13022) );
  sky130_fd_sc_hd__nand2_1 U19691 ( .A(n29488), .B(n11141), .Y(n28129) );
  sky130_fd_sc_hd__nand2_4 U19692 ( .A(n13023), .B(n24764), .Y(n24312) );
  sky130_fd_sc_hd__nand2_4 U19693 ( .A(n24360), .B(n13023), .Y(n27770) );
  sky130_fd_sc_hd__nand3_1 U19694 ( .A(n24811), .B(n12203), .C(n13023), .Y(
        j202_soc_core_j22_cpu_ml_machj[0]) );
  sky130_fd_sc_hd__nand2_4 U19695 ( .A(n13024), .B(n23493), .Y(n13023) );
  sky130_fd_sc_hd__nor2b_1 U19696 ( .B_N(n18470), .A(n13025), .Y(n18358) );
  sky130_fd_sc_hd__nand2_1 U19697 ( .A(n13030), .B(n13029), .Y(n18442) );
  sky130_fd_sc_hd__nand2_1 U19698 ( .A(n18428), .B(n18427), .Y(n13029) );
  sky130_fd_sc_hd__o21ai_1 U19699 ( .A1(n18427), .A2(n18428), .B1(n18426), .Y(
        n13030) );
  sky130_fd_sc_hd__nand2_1 U19701 ( .A(n13037), .B(n19692), .Y(n13033) );
  sky130_fd_sc_hd__nand2_1 U19702 ( .A(n25965), .B(n27152), .Y(n25970) );
  sky130_fd_sc_hd__nand2_1 U19703 ( .A(n25421), .B(n27152), .Y(n25427) );
  sky130_fd_sc_hd__fah_1 U19704 ( .A(n18419), .B(n18418), .CI(n18417), .COUT(
        n18439), .SUM(n18434) );
  sky130_fd_sc_hd__a21oi_1 U19705 ( .A1(n22595), .A2(n18671), .B1(n22594), .Y(
        n22596) );
  sky130_fd_sc_hd__nand3_1 U19706 ( .A(n25676), .B(n25680), .C(n25681), .Y(
        n22812) );
  sky130_fd_sc_hd__buf_4 U19707 ( .A(n24470), .X(n29771) );
  sky130_fd_sc_hd__buf_4 U19708 ( .A(n24470), .X(n29770) );
  sky130_fd_sc_hd__a21o_1 U19709 ( .A1(n21993), .A2(n22996), .B1(n21992), .X(
        n22866) );
  sky130_fd_sc_hd__inv_2 U19710 ( .A(n17239), .Y(n21104) );
  sky130_fd_sc_hd__nor2_1 U19711 ( .A(j202_soc_core_j22_cpu_regop_other__0_), 
        .B(n18861), .Y(n22987) );
  sky130_fd_sc_hd__a21o_1 U19712 ( .A1(n25806), .A2(n25805), .B1(n13103), .X(
        n26271) );
  sky130_fd_sc_hd__inv_2 U19713 ( .A(n27809), .Y(n27026) );
  sky130_fd_sc_hd__o22a_1 U19714 ( .A1(n15887), .A2(n15886), .B1(n15885), .B2(
        n14342), .X(n15893) );
  sky130_fd_sc_hd__o22a_1 U19715 ( .A1(n14344), .A2(n15886), .B1(n14343), .B2(
        n14342), .X(n14351) );
  sky130_fd_sc_hd__o22a_1 U19716 ( .A1(n21738), .A2(n15886), .B1(n16487), .B2(
        n22741), .X(n14261) );
  sky130_fd_sc_hd__o22a_1 U19717 ( .A1(n14174), .A2(n15886), .B1(n14173), .B2(
        n14342), .X(n14181) );
  sky130_fd_sc_hd__o22a_1 U19718 ( .A1(n14973), .A2(n15886), .B1(n14972), .B2(
        n14477), .X(n14979) );
  sky130_fd_sc_hd__o22a_1 U19719 ( .A1(n14479), .A2(n15886), .B1(n14478), .B2(
        n14477), .X(n14486) );
  sky130_fd_sc_hd__nand2b_1 U19720 ( .A_N(n20002), .B(n21101), .Y(n20172) );
  sky130_fd_sc_hd__nand2b_1 U19721 ( .A_N(n17288), .B(n21101), .Y(n17293) );
  sky130_fd_sc_hd__nand2b_1 U19722 ( .A_N(n19707), .B(n21101), .Y(n19701) );
  sky130_fd_sc_hd__inv_2 U19723 ( .A(n13450), .Y(n13957) );
  sky130_fd_sc_hd__nand2_2 U19724 ( .A(n30127), .B(n27355), .Y(n27123) );
  sky130_fd_sc_hd__nand2b_1 U19726 ( .A_N(n20560), .B(n20464), .Y(n20830) );
  sky130_fd_sc_hd__nand2b_1 U19727 ( .A_N(n20560), .B(n18744), .Y(n20344) );
  sky130_fd_sc_hd__nand2b_1 U19728 ( .A_N(n20560), .B(n19140), .Y(n20349) );
  sky130_fd_sc_hd__nand3_2 U19729 ( .A(n15006), .B(n12103), .C(n15005), .Y(
        n26329) );
  sky130_fd_sc_hd__inv_2 U19730 ( .A(n25845), .Y(n25855) );
  sky130_fd_sc_hd__nand2_4 U19731 ( .A(n22705), .B(n13365), .Y(n22747) );
  sky130_fd_sc_hd__inv_1 U19732 ( .A(n19129), .Y(n15150) );
  sky130_fd_sc_hd__o22a_1 U19733 ( .A1(n13365), .A2(n25933), .B1(n27025), .B2(
        n11186), .X(n21178) );
  sky130_fd_sc_hd__o22a_1 U19734 ( .A1(n13365), .A2(n17226), .B1(n27147), .B2(
        n11186), .X(n17228) );
  sky130_fd_sc_hd__o22a_1 U19735 ( .A1(n13365), .A2(n25428), .B1(n26321), .B2(
        n11186), .X(n20961) );
  sky130_fd_sc_hd__nand3_1 U19736 ( .A(n13365), .B(
        j202_soc_core_j22_cpu_memop_Ma__0_), .C(
        j202_soc_core_j22_cpu_memop_Ma__1_), .Y(n17053) );
  sky130_fd_sc_hd__nand3_2 U19737 ( .A(n13365), .B(
        j202_soc_core_j22_cpu_memop_Ma__1_), .C(n13379), .Y(n22743) );
  sky130_fd_sc_hd__nand3_2 U19738 ( .A(n14950), .B(n12104), .C(n14949), .Y(
        n26331) );
  sky130_fd_sc_hd__buf_2 U19739 ( .A(n11091), .X(n16506) );
  sky130_fd_sc_hd__inv_2 U19740 ( .A(n19158), .Y(n20664) );
  sky130_fd_sc_hd__a21oi_2 U19741 ( .A1(n18815), .A2(n14411), .B1(n14410), .Y(
        n16557) );
  sky130_fd_sc_hd__nand2b_1 U19742 ( .A_N(n20814), .B(n19148), .Y(n16321) );
  sky130_fd_sc_hd__fah_1 U19745 ( .A(n18175), .B(n18174), .CI(n18173), .COUT(
        n18183), .SUM(n18166) );
  sky130_fd_sc_hd__nor2_2 U19746 ( .A(n18764), .B(n18699), .Y(n20199) );
  sky130_fd_sc_hd__o22ai_1 U19747 ( .A1(n18492), .A2(n17731), .B1(n17730), 
        .B2(n18489), .Y(n17740) );
  sky130_fd_sc_hd__nand3_1 U19749 ( .A(n25460), .B(n25459), .C(n25458), .Y(
        n25468) );
  sky130_fd_sc_hd__nand3_2 U19750 ( .A(n13696), .B(n13051), .C(n13695), .Y(
        n26929) );
  sky130_fd_sc_hd__nand3_1 U19752 ( .A(n26920), .B(n26919), .C(n26918), .Y(
        n26921) );
  sky130_fd_sc_hd__inv_4 U19753 ( .A(n28498), .Y(n25594) );
  sky130_fd_sc_hd__a31oi_2 U19754 ( .A1(n23880), .A2(n26583), .A3(n26649), 
        .B1(n29088), .Y(n29877) );
  sky130_fd_sc_hd__nand3_2 U19756 ( .A(n14070), .B(n14069), .C(n12114), .Y(
        n28460) );
  sky130_fd_sc_hd__nand2_1 U19757 ( .A(n22439), .B(n22438), .Y(n24772) );
  sky130_fd_sc_hd__nand2_1 U19758 ( .A(n19295), .B(n19078), .Y(n19080) );
  sky130_fd_sc_hd__nand2_1 U19759 ( .A(n22161), .B(n16523), .Y(n13584) );
  sky130_fd_sc_hd__nor2_1 U19760 ( .A(n21260), .B(n19076), .Y(n19078) );
  sky130_fd_sc_hd__a22oi_1 U19761 ( .A1(j202_soc_core_j22_cpu_ml_mach[29]), 
        .A2(n23041), .B1(n23040), .B2(n24452), .Y(n23042) );
  sky130_fd_sc_hd__a2bb2oi_1 U19762 ( .B1(n14378), .B2(
        j202_soc_core_j22_cpu_regop_imm__7_), .A1_N(n18871), .A2_N(n16525), 
        .Y(n14288) );
  sky130_fd_sc_hd__o2bb2ai_1 U19763 ( .B1(n25556), .B2(n25986), .A1_N(n25555), 
        .A2_N(n25986), .Y(j202_soc_core_j22_cpu_rf_N2988) );
  sky130_fd_sc_hd__o2bb2ai_1 U19764 ( .B1(n25556), .B2(n25989), .A1_N(n25555), 
        .A2_N(n25989), .Y(j202_soc_core_j22_cpu_rf_N2766) );
  sky130_fd_sc_hd__o2bb2ai_1 U19765 ( .B1(n25556), .B2(n25979), .A1_N(n25555), 
        .A2_N(n25979), .Y(j202_soc_core_j22_cpu_rf_N3210) );
  sky130_fd_sc_hd__o2bb2ai_1 U19766 ( .B1(n25556), .B2(n25987), .A1_N(n25555), 
        .A2_N(n25987), .Y(j202_soc_core_j22_cpu_rf_N3136) );
  sky130_fd_sc_hd__o2bb2ai_1 U19767 ( .B1(n25556), .B2(n25983), .A1_N(n25555), 
        .A2_N(n25983), .Y(j202_soc_core_j22_cpu_rf_N3062) );
  sky130_fd_sc_hd__o2bb2ai_1 U19768 ( .B1(n25556), .B2(n25980), .A1_N(n25555), 
        .A2_N(n25980), .Y(j202_soc_core_j22_cpu_rf_N2803) );
  sky130_fd_sc_hd__o2bb2ai_1 U19769 ( .B1(n25556), .B2(n25977), .A1_N(n25555), 
        .A2_N(n25977), .Y(j202_soc_core_j22_cpu_rf_N2877) );
  sky130_fd_sc_hd__fah_1 U19770 ( .A(n17526), .B(n17525), .CI(n17524), .COUT(
        n17557), .SUM(n17836) );
  sky130_fd_sc_hd__fah_1 U19771 ( .A(n19048), .B(n19047), .CI(n19046), .COUT(
        n19052), .SUM(n19056) );
  sky130_fd_sc_hd__fah_1 U19772 ( .A(n18391), .B(n18390), .CI(n18389), .COUT(
        n18446), .SUM(n18440) );
  sky130_fd_sc_hd__a21boi_1 U19773 ( .A1(n23036), .A2(n21909), .B1_N(n21908), 
        .Y(n21910) );
  sky130_fd_sc_hd__a21oi_1 U19774 ( .A1(n23036), .A2(n13086), .B1(n19062), .Y(
        n18674) );
  sky130_fd_sc_hd__nand2_1 U19776 ( .A(n18858), .B(n16523), .Y(n14295) );
  sky130_fd_sc_hd__nand3_1 U19777 ( .A(n13912), .B(n13911), .C(n13910), .Y(
        n19264) );
  sky130_fd_sc_hd__nand3_2 U19778 ( .A(n22236), .B(n22235), .C(n22234), .Y(
        n28501) );
  sky130_fd_sc_hd__nand2b_1 U19779 ( .A_N(n25763), .B(n27152), .Y(n25310) );
  sky130_fd_sc_hd__nand2b_1 U19780 ( .A_N(n25763), .B(n23044), .Y(n22865) );
  sky130_fd_sc_hd__nand2_1 U19781 ( .A(n25128), .B(n27152), .Y(n25131) );
  sky130_fd_sc_hd__fah_1 U19782 ( .A(n17546), .B(n17545), .CI(n17544), .COUT(
        n17579), .SUM(n17538) );
  sky130_fd_sc_hd__fah_1 U19783 ( .A(n17888), .B(n17887), .CI(n17886), .COUT(
        n17910), .SUM(n17996) );
  sky130_fd_sc_hd__nor2b_1 U19784 ( .B_N(n18470), .A(n18213), .Y(n18201) );
  sky130_fd_sc_hd__o211ai_1 U19785 ( .A1(n28430), .A2(n26411), .B1(n26410), 
        .C1(n26409), .Y(n26412) );
  sky130_fd_sc_hd__a21o_1 U19786 ( .A1(n12260), .A2(n25724), .B1(n24182), .X(
        n29646) );
  sky130_fd_sc_hd__inv_2 U19788 ( .A(n27588), .Y(n26450) );
  sky130_fd_sc_hd__fah_1 U19789 ( .A(n17960), .B(n17959), .CI(n17958), .COUT(
        n17957), .SUM(n18058) );
  sky130_fd_sc_hd__nand3_1 U19790 ( .A(n22316), .B(n22461), .C(n22460), .Y(
        n29522) );
  sky130_fd_sc_hd__fah_1 U19791 ( .A(n18019), .B(n18018), .CI(n18017), .COUT(
        n18068), .SUM(n18065) );
  sky130_fd_sc_hd__nand2_8 U19792 ( .A(n17338), .B(n18533), .Y(n18530) );
  sky130_fd_sc_hd__fah_1 U19793 ( .A(n18400), .B(n18399), .CI(n18398), .COUT(
        n18426), .SUM(n18476) );
  sky130_fd_sc_hd__nor2_1 U19795 ( .A(n13802), .B(n13801), .Y(n13817) );
  sky130_fd_sc_hd__inv_6 U19796 ( .A(n23588), .Y(n27766) );
  sky130_fd_sc_hd__a21oi_2 U19797 ( .A1(n22855), .A2(n16523), .B1(n14487), .Y(
        n26285) );
  sky130_fd_sc_hd__o21ai_1 U19798 ( .A1(n22625), .A2(n11866), .B1(n22624), .Y(
        n22626) );
  sky130_fd_sc_hd__o21a_1 U19799 ( .A1(n23018), .A2(n25144), .B1(n22591), .X(
        n22617) );
  sky130_fd_sc_hd__nand3_1 U19800 ( .A(n24153), .B(n25679), .C(n24173), .Y(
        n24174) );
  sky130_fd_sc_hd__fah_1 U19801 ( .A(n18055), .B(n18054), .CI(n18053), .COUT(
        n18045), .SUM(n18071) );
  sky130_fd_sc_hd__fah_1 U19802 ( .A(n17481), .B(n17480), .CI(n17479), .COUT(
        n17539), .SUM(n17514) );
  sky130_fd_sc_hd__nand2b_4 U19803 ( .A_N(n14588), .B(n24033), .Y(n22745) );
  sky130_fd_sc_hd__nand2b_1 U19804 ( .A_N(n24673), .B(n24672), .Y(n27760) );
  sky130_fd_sc_hd__fah_1 U19805 ( .A(n17894), .B(n17893), .CI(n17892), .COUT(
        n17801), .SUM(n17923) );
  sky130_fd_sc_hd__nor2_1 U19807 ( .A(n22215), .B(n22211), .Y(n18329) );
  sky130_fd_sc_hd__fah_1 U19808 ( .A(n17474), .B(n17473), .CI(n17472), .COUT(
        n17530), .SUM(n17821) );
  sky130_fd_sc_hd__nand2_2 U19809 ( .A(n13479), .B(n13513), .Y(n14312) );
  sky130_fd_sc_hd__nand2_1 U19810 ( .A(n13477), .B(n28376), .Y(n13479) );
  sky130_fd_sc_hd__inv_2 U19811 ( .A(n16086), .Y(n16543) );
  sky130_fd_sc_hd__nand2_1 U19812 ( .A(n13555), .B(n13792), .Y(n16086) );
  sky130_fd_sc_hd__xnor2_1 U19813 ( .A(n17533), .B(n17552), .Y(n17851) );
  sky130_fd_sc_hd__o21a_1 U19814 ( .A1(n24469), .A2(n24468), .B1(n12213), .X(
        n24470) );
  sky130_fd_sc_hd__nand2_1 U19815 ( .A(n29513), .B(n12213), .Y(n24493) );
  sky130_fd_sc_hd__o21ai_1 U19816 ( .A1(n22807), .A2(n12349), .B1(n22806), .Y(
        n22808) );
  sky130_fd_sc_hd__a21oi_1 U19817 ( .A1(n18830), .A2(n18834), .B1(n28056), .Y(
        n22980) );
  sky130_fd_sc_hd__fah_1 U19818 ( .A(n18016), .B(n18015), .CI(n18014), .COUT(
        n18069), .SUM(n18066) );
  sky130_fd_sc_hd__buf_6 U19819 ( .A(n17461), .X(n18213) );
  sky130_fd_sc_hd__o21bai_1 U19820 ( .A1(n27648), .A2(n25766), .B1_N(n25285), 
        .Y(j202_soc_core_j22_cpu_rf_N3373) );
  sky130_fd_sc_hd__fah_1 U19821 ( .A(n17716), .B(n17714), .CI(n17715), .COUT(
        n17703), .SUM(n17750) );
  sky130_fd_sc_hd__fah_1 U19822 ( .A(n17700), .B(n17699), .CI(n17698), .COUT(
        n17702), .SUM(n17769) );
  sky130_fd_sc_hd__fah_1 U19823 ( .A(n18551), .B(n18550), .CI(n18549), .COUT(
        n18564), .SUM(n18566) );
  sky130_fd_sc_hd__a2bb2oi_2 U19824 ( .B1(n23516), .B2(n22230), .A1_N(n22229), 
        .A2_N(n12621), .Y(n22236) );
  sky130_fd_sc_hd__fah_1 U19825 ( .A(n17691), .B(n17690), .CI(n17689), .COUT(
        n17819), .SUM(n17824) );
  sky130_fd_sc_hd__a22oi_2 U19826 ( .A1(j202_soc_core_memory0_ram_dout0[26]), 
        .A2(n20457), .B1(n20456), .B2(j202_soc_core_memory0_ram_dout0[154]), 
        .Y(n16884) );
  sky130_fd_sc_hd__buf_4 U19828 ( .A(n17724), .X(n18209) );
  sky130_fd_sc_hd__a22oi_2 U19829 ( .A1(j202_soc_core_memory0_ram_dout0[122]), 
        .A2(n20460), .B1(n20459), .B2(j202_soc_core_memory0_ram_dout0[186]), 
        .Y(n16882) );
  sky130_fd_sc_hd__nor2_2 U19831 ( .A(n18661), .B(n18662), .Y(n21189) );
  sky130_fd_sc_hd__fah_1 U19832 ( .A(n18946), .B(n18945), .CI(n18944), .COUT(
        n18939), .SUM(n19047) );
  sky130_fd_sc_hd__fah_1 U19833 ( .A(n17741), .B(n17740), .CI(n17739), .COUT(
        n17767), .SUM(n17799) );
  sky130_fd_sc_hd__o2bb2ai_1 U19834 ( .B1(n26896), .B2(n27859), .A1_N(n25963), 
        .A2_N(n30051), .Y(j202_soc_core_j22_cpu_rf_N3325) );
  sky130_fd_sc_hd__o2bb2ai_1 U19835 ( .B1(n26896), .B2(n27841), .A1_N(n30051), 
        .A2_N(n27841), .Y(j202_soc_core_j22_cpu_rf_N3249) );
  sky130_fd_sc_hd__o2bb2ai_1 U19836 ( .B1(n26896), .B2(n25964), .A1_N(n25964), 
        .A2_N(n30050), .Y(j202_soc_core_j22_cpu_rf_N2694) );
  sky130_fd_sc_hd__o2bb2ai_1 U19837 ( .B1(n26896), .B2(n26894), .A1_N(n26895), 
        .A2_N(n26894), .Y(j202_soc_core_j22_cpu_rf_N2916) );
  sky130_fd_sc_hd__o2bb2ai_1 U19838 ( .B1(n26896), .B2(n25982), .A1_N(n26895), 
        .A2_N(n25982), .Y(j202_soc_core_j22_cpu_rf_N3027) );
  sky130_fd_sc_hd__o2bb2ai_1 U19839 ( .B1(n26896), .B2(n25981), .A1_N(n26895), 
        .A2_N(n25981), .Y(j202_soc_core_j22_cpu_rf_N3175) );
  sky130_fd_sc_hd__o2bb2ai_1 U19840 ( .B1(n26896), .B2(n25986), .A1_N(n30050), 
        .A2_N(n25986), .Y(j202_soc_core_j22_cpu_rf_N2990) );
  sky130_fd_sc_hd__o2bb2ai_1 U19841 ( .B1(n26896), .B2(n25988), .A1_N(n26895), 
        .A2_N(n25988), .Y(j202_soc_core_j22_cpu_rf_N2842) );
  sky130_fd_sc_hd__o2bb2ai_1 U19842 ( .B1(n26896), .B2(n25985), .A1_N(n30050), 
        .A2_N(n25985), .Y(j202_soc_core_j22_cpu_rf_N3101) );
  sky130_fd_sc_hd__o2bb2ai_1 U19843 ( .B1(n26896), .B2(n25984), .A1_N(n30051), 
        .A2_N(n25984), .Y(j202_soc_core_j22_cpu_rf_N2731) );
  sky130_fd_sc_hd__o2bb2ai_1 U19844 ( .B1(n26896), .B2(n25978), .A1_N(n30051), 
        .A2_N(n25978), .Y(j202_soc_core_j22_cpu_rf_N2953) );
  sky130_fd_sc_hd__o2bb2ai_1 U19845 ( .B1(n26896), .B2(n25987), .A1_N(n30050), 
        .A2_N(n25987), .Y(j202_soc_core_j22_cpu_rf_N3138) );
  sky130_fd_sc_hd__o2bb2ai_1 U19846 ( .B1(n26896), .B2(n25983), .A1_N(n30051), 
        .A2_N(n25983), .Y(j202_soc_core_j22_cpu_rf_N3064) );
  sky130_fd_sc_hd__o2bb2ai_1 U19847 ( .B1(n26896), .B2(n25980), .A1_N(n30050), 
        .A2_N(n25980), .Y(j202_soc_core_j22_cpu_rf_N2805) );
  sky130_fd_sc_hd__o2bb2ai_1 U19848 ( .B1(n26896), .B2(n25979), .A1_N(n26895), 
        .A2_N(n25979), .Y(j202_soc_core_j22_cpu_rf_N3212) );
  sky130_fd_sc_hd__o2bb2ai_1 U19849 ( .B1(n26896), .B2(n25977), .A1_N(n30051), 
        .A2_N(n25977), .Y(j202_soc_core_j22_cpu_rf_N2879) );
  sky130_fd_sc_hd__fah_1 U19850 ( .A(n17706), .B(n17705), .CI(n17704), .COUT(
        n17770), .SUM(n17777) );
  sky130_fd_sc_hd__fah_1 U19851 ( .A(n18198), .B(n18197), .CI(n18196), .COUT(
        n18254), .SUM(n18182) );
  sky130_fd_sc_hd__fah_1 U19852 ( .A(n18584), .B(n18583), .CI(n18582), .COUT(
        n18544), .SUM(n18604) );
  sky130_fd_sc_hd__inv_1 U19853 ( .A(n28118), .Y(n23452) );
  sky130_fd_sc_hd__a21oi_2 U19854 ( .A1(n21730), .A2(n18222), .B1(n18221), .Y(
        n19279) );
  sky130_fd_sc_hd__a21oi_4 U19855 ( .A1(n23160), .A2(n23159), .B1(n23158), .Y(
        n27315) );
  sky130_fd_sc_hd__fah_1 U19856 ( .A(n18958), .B(n18957), .CI(n18956), .COUT(
        n19008), .SUM(n18978) );
  sky130_fd_sc_hd__nand2_1 U19857 ( .A(n23483), .B(n25679), .Y(n25260) );
  sky130_fd_sc_hd__fah_1 U19859 ( .A(n17780), .B(n17779), .CI(n17778), .COUT(
        n17766), .SUM(n17891) );
  sky130_fd_sc_hd__nor2_1 U19860 ( .A(n18217), .B(n18218), .Y(n22885) );
  sky130_fd_sc_hd__fah_1 U19861 ( .A(n18043), .B(n18042), .CI(n18041), .COUT(
        n18061), .SUM(n18089) );
  sky130_fd_sc_hd__nand2b_1 U19862 ( .A_N(n26001), .B(n12436), .Y(n22429) );
  sky130_fd_sc_hd__a22oi_2 U19863 ( .A1(j202_soc_core_memory0_ram_dout0[327]), 
        .A2(n21490), .B1(n21634), .B2(j202_soc_core_memory0_ram_dout0[263]), 
        .Y(n17319) );
  sky130_fd_sc_hd__a22oi_2 U19864 ( .A1(j202_soc_core_memory0_ram_dout0[391]), 
        .A2(n21496), .B1(n21641), .B2(j202_soc_core_memory0_ram_dout0[231]), 
        .Y(n17317) );
  sky130_fd_sc_hd__nand2_2 U19865 ( .A(n23547), .B(n12064), .Y(n28387) );
  sky130_fd_sc_hd__nor2_2 U19866 ( .A(n18322), .B(n18323), .Y(n21235) );
  sky130_fd_sc_hd__and4_1 U19867 ( .A(n13977), .B(n13976), .C(n13975), .D(
        n13974), .X(n13038) );
  sky130_fd_sc_hd__and4_1 U19868 ( .A(n14031), .B(n14030), .C(n14029), .D(
        n14028), .X(n13039) );
  sky130_fd_sc_hd__and4_1 U19869 ( .A(n13956), .B(n13955), .C(n13954), .D(
        n13953), .X(n13040) );
  sky130_fd_sc_hd__and4_1 U19870 ( .A(n13950), .B(n13949), .C(n13948), .D(
        n13947), .X(n13041) );
  sky130_fd_sc_hd__and4_1 U19871 ( .A(n13962), .B(n13961), .C(n13960), .D(
        n13959), .X(n13042) );
  sky130_fd_sc_hd__xor2_1 U19873 ( .A(n28697), .B(n28698), .X(n13045) );
  sky130_fd_sc_hd__xnor2_1 U19874 ( .A(n15631), .B(n22298), .Y(n13047) );
  sky130_fd_sc_hd__and4_1 U19875 ( .A(n15935), .B(n15934), .C(n15933), .D(
        n15932), .X(n13049) );
  sky130_fd_sc_hd__and4_1 U19876 ( .A(n13810), .B(n13809), .C(n13808), .D(
        n13807), .X(n13050) );
  sky130_fd_sc_hd__o211a_2 U19877 ( .A1(n13914), .A2(n16444), .B1(n13684), 
        .C1(n13683), .X(n13051) );
  sky130_fd_sc_hd__xor2_1 U19878 ( .A(j202_soc_core_qspi_wb_addr[12]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[12]), .X(n13052) );
  sky130_fd_sc_hd__o211a_2 U19879 ( .A1(n27849), .A2(n22705), .B1(n16891), 
        .C1(n16890), .X(n13055) );
  sky130_fd_sc_hd__and4_1 U19880 ( .A(n11180), .B(n26381), .C(n26380), .D(
        n26385), .X(n13057) );
  sky130_fd_sc_hd__and4_1 U19881 ( .A(n15996), .B(n15995), .C(n15994), .D(
        n15993), .X(n13058) );
  sky130_fd_sc_hd__a22o_1 U19882 ( .A1(n18454), .A2(n18453), .B1(n18456), .B2(
        n17437), .X(n13059) );
  sky130_fd_sc_hd__and4_1 U19883 ( .A(n14870), .B(n14869), .C(n14868), .D(
        n14867), .X(n13060) );
  sky130_fd_sc_hd__o211a_2 U19884 ( .A1(n13660), .A2(n16444), .B1(n13659), 
        .C1(n13658), .X(n13061) );
  sky130_fd_sc_hd__o211a_2 U19885 ( .A1(n14259), .A2(n16444), .B1(n14195), 
        .C1(n14194), .X(n13062) );
  sky130_fd_sc_hd__and4_1 U19886 ( .A(n16443), .B(n16442), .C(n16441), .D(
        n16440), .X(n13063) );
  sky130_fd_sc_hd__and4_1 U19887 ( .A(n14309), .B(n14308), .C(n14307), .D(
        n14306), .X(n13064) );
  sky130_fd_sc_hd__inv_2 U19888 ( .A(n13826), .Y(n13761) );
  sky130_fd_sc_hd__inv_2 U19889 ( .A(n13761), .Y(n16507) );
  sky130_fd_sc_hd__inv_2 U19890 ( .A(n13456), .Y(n14106) );
  sky130_fd_sc_hd__inv_2 U19891 ( .A(n14106), .Y(n16399) );
  sky130_fd_sc_hd__o211a_2 U19892 ( .A1(n13047), .A2(n22705), .B1(n15634), 
        .C1(n15633), .X(n13065) );
  sky130_fd_sc_hd__xor2_1 U19893 ( .A(j202_soc_core_qspi_wb_addr[15]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[15]), .X(n13066) );
  sky130_fd_sc_hd__and4_1 U19894 ( .A(n15962), .B(n15961), .C(n15960), .D(
        n15959), .X(n13067) );
  sky130_fd_sc_hd__xor2_1 U19895 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]), .B(
        j202_soc_core_qspi_wb_addr[16]), .X(n13068) );
  sky130_fd_sc_hd__xor2_1 U19896 ( .A(j202_soc_core_qspi_wb_addr[9]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[9]), .X(n13069) );
  sky130_fd_sc_hd__xor2_1 U19897 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .B(
        j202_soc_core_qspi_wb_addr[22]), .X(n13070) );
  sky130_fd_sc_hd__or3_1 U19898 ( .A(n29088), .B(n24681), .C(n25963), .X(
        n13071) );
  sky130_fd_sc_hd__inv_2 U19899 ( .A(n15410), .Y(n17237) );
  sky130_fd_sc_hd__nor2_1 U19900 ( .A(n24030), .B(n28895), .Y(n29603) );
  sky130_fd_sc_hd__clkinv_1 U19901 ( .A(n29603), .Y(n28898) );
  sky130_fd_sc_hd__xor2_1 U19902 ( .A(j202_soc_core_qspi_wb_addr[10]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[10]), .X(n13073) );
  sky130_fd_sc_hd__inv_2 U19903 ( .A(n15886), .Y(n14775) );
  sky130_fd_sc_hd__inv_2 U19904 ( .A(n14095), .Y(n16426) );
  sky130_fd_sc_hd__inv_2 U19905 ( .A(n14095), .Y(n16043) );
  sky130_fd_sc_hd__inv_2 U19906 ( .A(n13952), .Y(n16044) );
  sky130_fd_sc_hd__inv_2 U19907 ( .A(n13538), .Y(n13946) );
  sky130_fd_sc_hd__inv_2 U19908 ( .A(n13526), .Y(n14220) );
  sky130_fd_sc_hd__inv_2 U19909 ( .A(n12086), .Y(n15788) );
  sky130_fd_sc_hd__inv_2 U19910 ( .A(n12086), .Y(n14821) );
  sky130_fd_sc_hd__inv_2 U19911 ( .A(n14200), .Y(n16427) );
  sky130_fd_sc_hd__inv_2 U19912 ( .A(n14200), .Y(n15796) );
  sky130_fd_sc_hd__clkinv_1 U19914 ( .A(n22364), .Y(n23593) );
  sky130_fd_sc_hd__clkinv_1 U19915 ( .A(n22317), .Y(n23589) );
  sky130_fd_sc_hd__or2_1 U19916 ( .A(n18259), .B(n18260), .X(n13076) );
  sky130_fd_sc_hd__clkinv_1 U19917 ( .A(n21121), .Y(n21126) );
  sky130_fd_sc_hd__clkinv_1 U19918 ( .A(j202_soc_core_j22_cpu_pc[11]), .Y(
        n14009) );
  sky130_fd_sc_hd__clkinv_1 U19919 ( .A(j202_soc_core_j22_cpu_pc[2]), .Y(
        n13913) );
  sky130_fd_sc_hd__clkinv_1 U19920 ( .A(j202_soc_core_j22_cpu_pc[24]), .Y(
        n22725) );
  sky130_fd_sc_hd__clkinv_1 U19921 ( .A(j202_soc_core_j22_cpu_pc[10]), .Y(
        n14345) );
  sky130_fd_sc_hd__clkinv_1 U19922 ( .A(j202_soc_core_j22_cpu_pc[20]), .Y(
        n22322) );
  sky130_fd_sc_hd__clkinv_1 U19923 ( .A(j202_soc_core_j22_cpu_pc[18]), .Y(
        n13377) );
  sky130_fd_sc_hd__clkinv_1 U19924 ( .A(j202_soc_core_j22_cpu_pc[21]), .Y(
        n22298) );
  sky130_fd_sc_hd__clkinv_1 U19925 ( .A(j202_soc_core_j22_cpu_pc[15]), .Y(
        n14563) );
  sky130_fd_sc_hd__clkinv_1 U19926 ( .A(j202_soc_core_j22_cpu_pc[23]), .Y(
        n15260) );
  sky130_fd_sc_hd__clkinv_1 U19927 ( .A(j202_soc_core_j22_cpu_pc[19]), .Y(
        n15484) );
  sky130_fd_sc_hd__nor2_1 U19928 ( .A(n24034), .B(n24037), .Y(n26068) );
  sky130_fd_sc_hd__clkinv_1 U19929 ( .A(j202_soc_core_j22_cpu_pc[9]), .Y(
        n14375) );
  sky130_fd_sc_hd__clkinv_1 U19930 ( .A(j202_soc_core_j22_cpu_pc[5]), .Y(
        n13640) );
  sky130_fd_sc_hd__and4_1 U19931 ( .A(n15034), .B(n15033), .C(n15032), .D(
        n15031), .X(n13084) );
  sky130_fd_sc_hd__clkinv_1 U19932 ( .A(j202_soc_core_j22_cpu_pc[22]), .Y(
        n22164) );
  sky130_fd_sc_hd__clkinv_1 U19933 ( .A(j202_soc_core_j22_cpu_pc[17]), .Y(
        n22849) );
  sky130_fd_sc_hd__nor2_1 U19935 ( .A(n24282), .B(n26160), .Y(n25696) );
  sky130_fd_sc_hd__clkinv_1 U19936 ( .A(j202_soc_core_j22_cpu_pc[8]), .Y(
        n22741) );
  sky130_fd_sc_hd__and4_1 U19937 ( .A(n14224), .B(n14223), .C(n14222), .D(
        n14221), .X(n13085) );
  sky130_fd_sc_hd__clkinv_1 U19938 ( .A(j202_soc_core_j22_cpu_pc[7]), .Y(
        n14285) );
  sky130_fd_sc_hd__or2_1 U19939 ( .A(n18672), .B(n18673), .X(n13086) );
  sky130_fd_sc_hd__and2_1 U19940 ( .A(n27093), .B(n29581), .X(n13088) );
  sky130_fd_sc_hd__clkinv_1 U19941 ( .A(j202_soc_core_j22_cpu_pc[16]), .Y(
        n22769) );
  sky130_fd_sc_hd__inv_2 U19942 ( .A(n13827), .Y(n15950) );
  sky130_fd_sc_hd__inv_2 U19943 ( .A(n14053), .Y(n15017) );
  sky130_fd_sc_hd__inv_2 U19944 ( .A(n14053), .Y(n16064) );
  sky130_fd_sc_hd__and4_1 U19945 ( .A(n13844), .B(n13843), .C(n13842), .D(
        n13841), .X(n13089) );
  sky130_fd_sc_hd__inv_2 U19946 ( .A(n13835), .Y(n13392) );
  sky130_fd_sc_hd__and4_1 U19947 ( .A(n15974), .B(n15973), .C(n15972), .D(
        n15971), .X(n13091) );
  sky130_fd_sc_hd__clkinv_1 U19948 ( .A(j202_soc_core_j22_cpu_pc[14]), .Y(
        n14143) );
  sky130_fd_sc_hd__and4_1 U19949 ( .A(n14111), .B(n14110), .C(n14109), .D(
        n14108), .X(n13093) );
  sky130_fd_sc_hd__clkinv_1 U19950 ( .A(j202_soc_core_j22_cpu_pc[13]), .Y(
        n14175) );
  sky130_fd_sc_hd__and4_1 U19951 ( .A(n14783), .B(n14782), .C(n14781), .D(
        n14780), .X(n13094) );
  sky130_fd_sc_hd__and4_1 U19952 ( .A(n15064), .B(n15063), .C(n15062), .D(
        n15061), .X(n13096) );
  sky130_fd_sc_hd__and4_1 U19953 ( .A(n16008), .B(n16007), .C(n16006), .D(
        n16005), .X(n13099) );
  sky130_fd_sc_hd__and2_1 U19954 ( .A(n25243), .B(n25242), .X(n13101) );
  sky130_fd_sc_hd__clkinv_1 U19955 ( .A(j202_soc_core_j22_cpu_pc[6]), .Y(
        n13576) );
  sky130_fd_sc_hd__clkinv_1 U19956 ( .A(j202_soc_core_j22_cpu_pc[4]), .Y(
        n13750) );
  sky130_fd_sc_hd__and4_1 U19957 ( .A(n15860), .B(n15859), .C(n15858), .D(
        n15857), .X(n13107) );
  sky130_fd_sc_hd__and4_1 U19958 ( .A(n16538), .B(n16537), .C(n16536), .D(
        n16535), .X(n13108) );
  sky130_fd_sc_hd__and4_1 U19959 ( .A(n13582), .B(n13581), .C(n13580), .D(
        n13579), .X(n13110) );
  sky130_fd_sc_hd__nor2_2 U19960 ( .A(n29088), .B(n25336), .Y(n29752) );
  sky130_fd_sc_hd__clkinv_1 U19961 ( .A(n18576), .Y(n18573) );
  sky130_fd_sc_hd__clkinv_1 U19963 ( .A(n22498), .Y(n22493) );
  sky130_fd_sc_hd__nand2_1 U19964 ( .A(n13860), .B(n13787), .Y(n16541) );
  sky130_fd_sc_hd__a21oi_1 U19965 ( .A1(n23036), .A2(n22923), .B1(n22922), .Y(
        n22924) );
  sky130_fd_sc_hd__inv_2 U19966 ( .A(n27042), .Y(n27804) );
  sky130_fd_sc_hd__inv_2 U19967 ( .A(n21272), .Y(n22965) );
  sky130_fd_sc_hd__clkinv_1 U19968 ( .A(n18151), .Y(n18149) );
  sky130_fd_sc_hd__nor2_1 U19969 ( .A(n18806), .B(n26048), .Y(n27786) );
  sky130_fd_sc_hd__inv_2 U19970 ( .A(n26329), .Y(n26280) );
  sky130_fd_sc_hd__nand2_1 U19971 ( .A(n13155), .B(n13157), .Y(n13162) );
  sky130_fd_sc_hd__nand3_2 U19972 ( .A(n13436), .B(n18869), .C(n18859), .Y(
        n16490) );
  sky130_fd_sc_hd__nand3_1 U19973 ( .A(n17354), .B(n17353), .C(n17352), .Y(
        n18830) );
  sky130_fd_sc_hd__inv_2 U19974 ( .A(n14525), .Y(n14001) );
  sky130_fd_sc_hd__nand3_1 U19975 ( .A(n25436), .B(n25435), .C(n25434), .Y(
        n25437) );
  sky130_fd_sc_hd__nand3_1 U19976 ( .A(n28204), .B(n19605), .C(n19598), .Y(
        n21517) );
  sky130_fd_sc_hd__nand2_1 U19977 ( .A(n21650), .B(n21768), .Y(n21653) );
  sky130_fd_sc_hd__a21oi_2 U19978 ( .A1(n21744), .A2(n16523), .B1(n14264), .Y(
        n24931) );
  sky130_fd_sc_hd__nand2_1 U19979 ( .A(n24453), .B(n24452), .Y(n24460) );
  sky130_fd_sc_hd__clkinv_1 U19980 ( .A(n13815), .Y(n13816) );
  sky130_fd_sc_hd__nand2_1 U19981 ( .A(n23483), .B(n24452), .Y(n24798) );
  sky130_fd_sc_hd__a21oi_1 U19982 ( .A1(n17040), .A2(n16193), .B1(n16192), .Y(
        n16196) );
  sky130_fd_sc_hd__nor2_1 U19983 ( .A(n24122), .B(n24121), .Y(n24123) );
  sky130_fd_sc_hd__clkinv_1 U19984 ( .A(n20580), .Y(n21629) );
  sky130_fd_sc_hd__nor2_1 U19985 ( .A(n13368), .B(n28102), .Y(n24034) );
  sky130_fd_sc_hd__nor2_1 U19986 ( .A(j202_soc_core_j22_cpu_ma_M_area[1]), .B(
        j202_soc_core_j22_cpu_ma_M_area[0]), .Y(n21650) );
  sky130_fd_sc_hd__buf_2 U19987 ( .A(n13426), .X(n16523) );
  sky130_fd_sc_hd__clkinv_1 U19988 ( .A(n29261), .Y(n29264) );
  sky130_fd_sc_hd__nand2_1 U19989 ( .A(n27514), .B(n29170), .Y(n27540) );
  sky130_fd_sc_hd__clkbuf_1 U19990 ( .A(n27398), .X(n28328) );
  sky130_fd_sc_hd__nor2_1 U19991 ( .A(n25084), .B(n25083), .Y(n28326) );
  sky130_fd_sc_hd__nand3_1 U19992 ( .A(n24798), .B(n24797), .C(n24796), .Y(
        n24904) );
  sky130_fd_sc_hd__nand3_1 U19993 ( .A(n24176), .B(
        j202_soc_core_j22_cpu_regop_We__0_), .C(n23888), .Y(n27775) );
  sky130_fd_sc_hd__nand2_1 U19994 ( .A(n23314), .B(n23313), .Y(n24392) );
  sky130_fd_sc_hd__nor2_1 U19995 ( .A(n13075), .B(n24283), .Y(n28425) );
  sky130_fd_sc_hd__nor2_1 U19996 ( .A(n28211), .B(n24756), .Y(n28295) );
  sky130_fd_sc_hd__clkinv_1 U19997 ( .A(n26397), .Y(n26393) );
  sky130_fd_sc_hd__o31a_1 U19998 ( .A1(n26904), .A2(n26783), .A3(n26903), .B1(
        n29745), .X(n29061) );
  sky130_fd_sc_hd__inv_2 U20000 ( .A(j202_soc_core_intc_core_00_rg_ipr[21]), 
        .Y(n25578) );
  sky130_fd_sc_hd__nor2_1 U20001 ( .A(n24755), .B(n28210), .Y(n27486) );
  sky130_fd_sc_hd__clkinv_1 U20002 ( .A(n28177), .Y(n28545) );
  sky130_fd_sc_hd__nor2_1 U20003 ( .A(n29088), .B(n28235), .Y(n28233) );
  sky130_fd_sc_hd__nand2_1 U20006 ( .A(n23828), .B(n23827), .Y(n25981) );
  sky130_fd_sc_hd__nor2_1 U20007 ( .A(n13325), .B(n28512), .Y(n28540) );
  sky130_fd_sc_hd__nand2_1 U20008 ( .A(n24732), .B(n24736), .Y(n28289) );
  sky130_fd_sc_hd__a2bb2oi_1 U20009 ( .B1(n28870), .B2(n27231), .A1_N(n26564), 
        .A2_N(n27224), .Y(n26565) );
  sky130_fd_sc_hd__nand2_1 U20010 ( .A(n23887), .B(n29745), .Y(n27855) );
  sky130_fd_sc_hd__clkinv_1 U20011 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[22]), .Y(n26831) );
  sky130_fd_sc_hd__buf_4 U20012 ( .A(j202_soc_core_rst), .X(n29088) );
  sky130_fd_sc_hd__nor3_1 U20013 ( .A(wb_rst_i), .B(wbs_ack_o), .C(n13111), 
        .Y(n24025) );
  sky130_fd_sc_hd__nand3_1 U20015 ( .A(n22865), .B(n22864), .C(n22868), .Y(
        n29504) );
  sky130_fd_sc_hd__o2bb2ai_1 U20016 ( .B1(n26896), .B2(n25989), .A1_N(n26895), 
        .A2_N(n25989), .Y(j202_soc_core_j22_cpu_rf_N2768) );
  sky130_fd_sc_hd__and3_1 U20017 ( .A(n26479), .B(n26467), .C(n29830), .X(
        n29631) );
  sky130_fd_sc_hd__o2bb2ai_1 U20018 ( .B1(n25556), .B2(n27841), .A1_N(n25555), 
        .A2_N(n27841), .Y(j202_soc_core_j22_cpu_rf_N3247) );
  sky130_fd_sc_hd__o2bb2ai_1 U20019 ( .B1(n25556), .B2(n25981), .A1_N(n25555), 
        .A2_N(n25981), .Y(j202_soc_core_j22_cpu_rf_N3173) );
  sky130_fd_sc_hd__o2bb2ai_1 U20020 ( .B1(n25556), .B2(n25985), .A1_N(n25555), 
        .A2_N(n25985), .Y(j202_soc_core_j22_cpu_rf_N3099) );
  sky130_fd_sc_hd__o2bb2ai_1 U20021 ( .B1(n25556), .B2(n25982), .A1_N(n25555), 
        .A2_N(n25982), .Y(j202_soc_core_j22_cpu_rf_N3025) );
  sky130_fd_sc_hd__o2bb2ai_1 U20022 ( .B1(n25556), .B2(n25978), .A1_N(n25555), 
        .A2_N(n25978), .Y(j202_soc_core_j22_cpu_rf_N2951) );
  sky130_fd_sc_hd__o2bb2ai_1 U20023 ( .B1(n25556), .B2(n26894), .A1_N(n25555), 
        .A2_N(n26894), .Y(j202_soc_core_j22_cpu_rf_N2914) );
  sky130_fd_sc_hd__o2bb2ai_1 U20024 ( .B1(n25556), .B2(n25988), .A1_N(n25555), 
        .A2_N(n25988), .Y(j202_soc_core_j22_cpu_rf_N2840) );
  sky130_fd_sc_hd__o2bb2ai_1 U20025 ( .B1(n25556), .B2(n25984), .A1_N(n25555), 
        .A2_N(n25984), .Y(j202_soc_core_j22_cpu_rf_N2729) );
  sky130_fd_sc_hd__o2bb2ai_1 U20026 ( .B1(n25556), .B2(n25964), .A1_N(n25555), 
        .A2_N(n25964), .Y(j202_soc_core_j22_cpu_rf_N2692) );
  sky130_fd_sc_hd__nand2b_1 U20027 ( .A_N(n27062), .B(n27061), .Y(
        j202_soc_core_j22_cpu_rf_N3375) );
  sky130_fd_sc_hd__nand2_1 U20028 ( .A(n28540), .B(n24430), .Y(
        j202_soc_core_j22_cpu_ml_N428) );
  sky130_fd_sc_hd__o2bb2ai_1 U20029 ( .B1(n25556), .B2(n27859), .A1_N(n25555), 
        .A2_N(n25963), .Y(j202_soc_core_j22_cpu_rf_N3324) );
  sky130_fd_sc_hd__a21oi_1 U20030 ( .A1(n23637), .A2(n23636), .B1(n29088), .Y(
        n29876) );
  sky130_fd_sc_hd__clkbuf_1 U20031 ( .A(n29876), .X(n29754) );
  sky130_fd_sc_hd__clkbuf_1 U20032 ( .A(io_oeb[12]), .X(io_oeb[13]) );
  sky130_fd_sc_hd__clkbuf_1 U20033 ( .A(la_data_out[2]), .X(io_out[2]) );
  sky130_fd_sc_hd__clkbuf_1 U20034 ( .A(la_data_out[11]), .X(io_out[31]) );
  sky130_fd_sc_hd__nand3_1 U20035 ( .A(start_n_reg[1]), .B(wbs_cyc_i), .C(
        wbs_stb_i), .Y(n13111) );
  sky130_fd_sc_hd__nor2_1 U20036 ( .A(n29088), .B(n28258), .Y(n29598) );
  sky130_fd_sc_hd__nor2_1 U20037 ( .A(n29088), .B(n26831), .Y(n29579) );
  sky130_fd_sc_hd__nor2_1 U20038 ( .A(n29088), .B(n29051), .Y(n29605) );
  sky130_fd_sc_hd__nor2_1 U20039 ( .A(j202_soc_core_rst), .B(n26809), .Y(
        n29578) );
  sky130_fd_sc_hd__nor2_1 U20040 ( .A(n29088), .B(n29058), .Y(n29606) );
  sky130_fd_sc_hd__nor2_1 U20041 ( .A(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[0]), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[1]), .Y(n13114) );
  sky130_fd_sc_hd__xnor2_1 U20042 ( .A(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[0]), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[0]), .Y(n13113) );
  sky130_fd_sc_hd__xnor2_1 U20043 ( .A(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[1]), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[1]), .Y(n13112) );
  sky130_fd_sc_hd__nand2_1 U20044 ( .A(n13113), .B(n13112), .Y(n13115) );
  sky130_fd_sc_hd__or4_1 U20045 ( .A(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[2]), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[2]), .C(n13114), 
        .D(n13115), .X(n28157) );
  sky130_fd_sc_hd__nand3_1 U20046 ( .A(n13116), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[2]), .C(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[2]), .Y(n28160) );
  sky130_fd_sc_hd__nand2_1 U20047 ( .A(n28157), .B(n28160), .Y(n29599) );
  sky130_fd_sc_hd__xnor2_1 U20048 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .B(
        j202_soc_core_bldc_core_00_pwm_period[0]), .Y(n13118) );
  sky130_fd_sc_hd__xnor2_1 U20049 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .B(
        j202_soc_core_bldc_core_00_pwm_period[10]), .Y(n13117) );
  sky130_fd_sc_hd__nand2_1 U20050 ( .A(n13118), .B(n13117), .Y(n13135) );
  sky130_fd_sc_hd__xor2_1 U20051 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[11]), .B(
        j202_soc_core_bldc_core_00_pwm_period[11]), .X(n13120) );
  sky130_fd_sc_hd__xor2_1 U20052 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]), .B(
        j202_soc_core_bldc_core_00_pwm_period[5]), .X(n13119) );
  sky130_fd_sc_hd__nor2_1 U20053 ( .A(n13120), .B(n13119), .Y(n13130) );
  sky130_fd_sc_hd__xnor2_1 U20054 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .B(n27445), .Y(
        n13122) );
  sky130_fd_sc_hd__xor2_1 U20055 ( .A(j202_soc_core_bldc_core_00_pwm_period[2]), .B(j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[2]), .X(n13121) );
  sky130_fd_sc_hd__nor2_1 U20056 ( .A(n13122), .B(n13121), .Y(n13129) );
  sky130_fd_sc_hd__xnor2_1 U20057 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .B(n27968), .Y(
        n13124) );
  sky130_fd_sc_hd__xnor2_1 U20058 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[7]), .B(n24531), .Y(n13123) );
  sky130_fd_sc_hd__nor2_1 U20059 ( .A(n13124), .B(n13123), .Y(n13128) );
  sky130_fd_sc_hd__xnor2_1 U20060 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[3]), .B(n24521), .Y(n13126) );
  sky130_fd_sc_hd__xnor2_1 U20061 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .B(n28307), .Y(
        n13125) );
  sky130_fd_sc_hd__nor2_1 U20062 ( .A(n13126), .B(n13125), .Y(n13127) );
  sky130_fd_sc_hd__nand4_1 U20063 ( .A(n13130), .B(n13129), .C(n13128), .D(
        n13127), .Y(n13133) );
  sky130_fd_sc_hd__xnor2_1 U20064 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]), .B(
        j202_soc_core_bldc_core_00_pwm_period[9]), .Y(n13132) );
  sky130_fd_sc_hd__xnor2_1 U20065 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[4]), .B(
        j202_soc_core_bldc_core_00_pwm_period[4]), .Y(n13131) );
  sky130_fd_sc_hd__nand3b_1 U20066 ( .A_N(n13133), .B(n13132), .C(n13131), .Y(
        n13134) );
  sky130_fd_sc_hd__nor2_1 U20067 ( .A(n13135), .B(n13134), .Y(n29115) );
  sky130_fd_sc_hd__nand2b_1 U20068 ( .A_N(n29115), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .Y(n29493) );
  sky130_fd_sc_hd__nor2_1 U20069 ( .A(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[1]), .B(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[0]), .Y(n13136) );
  sky130_fd_sc_hd__nand3_1 U20070 ( .A(n13136), .B(j202_soc_core_aquc_STB_), 
        .C(j202_soc_core_aquc_CE__0_), .Y(n25033) );
  sky130_fd_sc_hd__nand2_1 U20071 ( .A(n21049), .B(n24724), .Y(n24177) );
  sky130_fd_sc_hd__nand2_1 U20072 ( .A(n24177), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[0]), .Y(n13138) );
  sky130_fd_sc_hd__nor2_1 U20073 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[2]), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[1]), .Y(n13137) );
  sky130_fd_sc_hd__nand2_1 U20074 ( .A(n13138), .B(n13137), .Y(n13140) );
  sky130_fd_sc_hd__nor2_1 U20075 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[3]), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[4]), .Y(n13139) );
  sky130_fd_sc_hd__nand2_1 U20076 ( .A(n13140), .B(n13139), .Y(n13144) );
  sky130_fd_sc_hd__nor2_1 U20077 ( .A(j202_soc_core_ahb2apb_01_state[0]), .B(
        j202_soc_core_ahb2apb_01_state[1]), .Y(n25039) );
  sky130_fd_sc_hd__nand2_1 U20078 ( .A(n25039), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[1]), .Y(n13142) );
  sky130_fd_sc_hd__inv_2 U20079 ( .A(j202_soc_core_ahb2apb_02_state[1]), .Y(
        n24296) );
  sky130_fd_sc_hd__nand2_1 U20080 ( .A(n24296), .B(n24260), .Y(n13141) );
  sky130_fd_sc_hd__mux2i_1 U20081 ( .A0(n13142), .A1(n13141), .S(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[2]), .Y(n13143) );
  sky130_fd_sc_hd__nor2_1 U20082 ( .A(n13144), .B(n13143), .Y(n13146) );
  sky130_fd_sc_hd__nor2_1 U20083 ( .A(j202_soc_core_memory0_ram_dout0_sel[14]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[13]), .Y(n13151) );
  sky130_fd_sc_hd__nand2_1 U20084 ( .A(n13151), .B(n13150), .Y(n13153) );
  sky130_fd_sc_hd__nand2_1 U20085 ( .A(n13163), .B(
        j202_soc_core_memory0_ram_dout0_sel[8]), .Y(n13154) );
  sky130_fd_sc_hd__nor2_1 U20086 ( .A(j202_soc_core_memory0_ram_dout0_sel[7]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[6]), .Y(n13174) );
  sky130_fd_sc_hd__nand2_1 U20087 ( .A(n13174), .B(n13176), .Y(n13169) );
  sky130_fd_sc_hd__nor2_1 U20088 ( .A(j202_soc_core_memory0_ram_dout0_sel[4]), 
        .B(n13169), .Y(n13167) );
  sky130_fd_sc_hd__nor2_1 U20089 ( .A(j202_soc_core_memory0_ram_dout0_sel[2]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[3]), .Y(n13158) );
  sky130_fd_sc_hd__nand3_1 U20090 ( .A(n13167), .B(
        j202_soc_core_memory0_ram_dout0_sel[1]), .C(n13158), .Y(n13161) );
  sky130_fd_sc_hd__nor2_1 U20091 ( .A(j202_soc_core_memory0_ram_dout0_sel[7]), 
        .B(n13164), .Y(n20455) );
  sky130_fd_sc_hd__nand4_1 U20092 ( .A(n13166), .B(n13173), .C(
        j202_soc_core_memory0_ram_dout0_sel[0]), .D(n13165), .Y(n13168) );
  sky130_fd_sc_hd__nand2_1 U20093 ( .A(n13173), .B(
        j202_soc_core_memory0_ram_dout0_sel[2]), .Y(n13171) );
  sky130_fd_sc_hd__nand2_1 U20094 ( .A(j202_soc_core_memory0_ram_dout0[82]), 
        .B(n20458), .Y(n13177) );
  sky130_fd_sc_hd__nand2_1 U20096 ( .A(n21650), .B(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n21022) );
  sky130_fd_sc_hd__nand2_1 U20097 ( .A(n13178), .B(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n20253) );
  sky130_fd_sc_hd__inv_2 U20098 ( .A(n13180), .Y(n20464) );
  sky130_fd_sc_hd__nand2_1 U20099 ( .A(n18712), .B(n11150), .Y(n15678) );
  sky130_fd_sc_hd__nor2_1 U20100 ( .A(n15685), .B(n15678), .Y(n19712) );
  sky130_fd_sc_hd__nand2_1 U20101 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .B(n13199), .Y(n15527) );
  sky130_fd_sc_hd__nand2_1 U20102 ( .A(n19712), .B(n20196), .Y(n15535) );
  sky130_fd_sc_hd__inv_2 U20103 ( .A(n21145), .Y(n21101) );
  sky130_fd_sc_hd__inv_4 U20104 ( .A(n19130), .Y(n21088) );
  sky130_fd_sc_hd__nor2_1 U20105 ( .A(n21101), .B(n19726), .Y(n13201) );
  sky130_fd_sc_hd__nor2_2 U20106 ( .A(j202_soc_core_bootrom_00_address_w[11]), 
        .B(n18712), .Y(n17250) );
  sky130_fd_sc_hd__nand2_1 U20107 ( .A(n17250), .B(n20464), .Y(n16985) );
  sky130_fd_sc_hd__nor2_1 U20108 ( .A(n21145), .B(n18744), .Y(n15610) );
  sky130_fd_sc_hd__nand2_1 U20109 ( .A(n19124), .B(n15610), .Y(n19777) );
  sky130_fd_sc_hd__nor2_1 U20110 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n20464), .Y(n19129) );
  sky130_fd_sc_hd__nor2_1 U20111 ( .A(n18712), .B(n15150), .Y(n15394) );
  sky130_fd_sc_hd__inv_4 U20112 ( .A(n18744), .Y(n19140) );
  sky130_fd_sc_hd__nand2_1 U20113 ( .A(n13182), .B(n21145), .Y(n13203) );
  sky130_fd_sc_hd__nor2_1 U20114 ( .A(n19140), .B(n13203), .Y(n19866) );
  sky130_fd_sc_hd__nand2_1 U20115 ( .A(n15394), .B(n19866), .Y(n19753) );
  sky130_fd_sc_hd__nor2_1 U20116 ( .A(n19140), .B(n21145), .Y(n15516) );
  sky130_fd_sc_hd__nand2_1 U20117 ( .A(n17250), .B(n15516), .Y(n20034) );
  sky130_fd_sc_hd__nand2b_1 U20118 ( .A_N(n20034), .B(n16338), .Y(n19763) );
  sky130_fd_sc_hd__nand3_1 U20119 ( .A(n19777), .B(n19753), .C(n19763), .Y(
        n13184) );
  sky130_fd_sc_hd__nand2_1 U20120 ( .A(n11150), .B(n19140), .Y(n18713) );
  sky130_fd_sc_hd__nand2_1 U20121 ( .A(n18727), .B(n21101), .Y(n13181) );
  sky130_fd_sc_hd__nor2_1 U20122 ( .A(n20464), .B(n13179), .Y(n15684) );
  sky130_fd_sc_hd__nand2_1 U20123 ( .A(n15684), .B(n18712), .Y(n13190) );
  sky130_fd_sc_hd__nor2_1 U20124 ( .A(n13181), .B(n13190), .Y(n19507) );
  sky130_fd_sc_hd__nand2_1 U20125 ( .A(n17241), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n17100) );
  sky130_fd_sc_hd__nor2_1 U20126 ( .A(n19119), .B(n17100), .Y(n15303) );
  sky130_fd_sc_hd__nor2_1 U20127 ( .A(n19140), .B(n21101), .Y(n16205) );
  sky130_fd_sc_hd__nand2_1 U20128 ( .A(n15303), .B(n16205), .Y(n19523) );
  sky130_fd_sc_hd__nand2_1 U20129 ( .A(n11150), .B(n21145), .Y(n17265) );
  sky130_fd_sc_hd__nor2_1 U20130 ( .A(n19140), .B(n18764), .Y(n16160) );
  sky130_fd_sc_hd__nand2_1 U20131 ( .A(n18742), .B(n16160), .Y(n18704) );
  sky130_fd_sc_hd__nor2_1 U20132 ( .A(n15150), .B(n18704), .Y(n15435) );
  sky130_fd_sc_hd__nand3_1 U20133 ( .A(n19738), .B(n19523), .C(n19770), .Y(
        n15393) );
  sky130_fd_sc_hd__nor2_1 U20135 ( .A(n13183), .B(n19120), .Y(n15409) );
  sky130_fd_sc_hd__nand2_1 U20136 ( .A(n21145), .B(n19140), .Y(n15106) );
  sky130_fd_sc_hd__nand2_1 U20137 ( .A(n19124), .B(n15577), .Y(n19813) );
  sky130_fd_sc_hd__nand2b_1 U20138 ( .A_N(n20034), .B(n19129), .Y(n13234) );
  sky130_fd_sc_hd__nand2_1 U20139 ( .A(n15303), .B(n15610), .Y(n19764) );
  sky130_fd_sc_hd__nand4_1 U20140 ( .A(n19728), .B(n19813), .C(n13234), .D(
        n19764), .Y(n19779) );
  sky130_fd_sc_hd__nor3_1 U20141 ( .A(n13184), .B(n15393), .C(n19779), .Y(
        n13185) );
  sky130_fd_sc_hd__nand2_1 U20142 ( .A(n15303), .B(n15577), .Y(n19714) );
  sky130_fd_sc_hd__nand2_1 U20143 ( .A(n19712), .B(n16205), .Y(n19490) );
  sky130_fd_sc_hd__nand2_1 U20144 ( .A(n19714), .B(n19490), .Y(n15424) );
  sky130_fd_sc_hd__nand2_1 U20145 ( .A(n19712), .B(n15577), .Y(n15431) );
  sky130_fd_sc_hd__nand2_1 U20146 ( .A(n20464), .B(n21359), .Y(n15747) );
  sky130_fd_sc_hd__nor2_1 U20147 ( .A(n18712), .B(n15747), .Y(n19504) );
  sky130_fd_sc_hd__nand2_1 U20148 ( .A(n19866), .B(n19504), .Y(n15396) );
  sky130_fd_sc_hd__nand2_1 U20149 ( .A(n15431), .B(n15396), .Y(n19465) );
  sky130_fd_sc_hd__nor2_1 U20150 ( .A(n17265), .B(n13190), .Y(n19827) );
  sky130_fd_sc_hd__nand2_1 U20151 ( .A(n19827), .B(n19140), .Y(n19814) );
  sky130_fd_sc_hd__nand2b_1 U20152 ( .A_N(n19465), .B(n19814), .Y(n15422) );
  sky130_fd_sc_hd__nor2_1 U20153 ( .A(n15424), .B(n15422), .Y(n19711) );
  sky130_fd_sc_hd__nand2_1 U20154 ( .A(n13185), .B(n19711), .Y(n13186) );
  sky130_fd_sc_hd__nand2_1 U20155 ( .A(n19148), .B(n21088), .Y(n15410) );
  sky130_fd_sc_hd__nand2_1 U20156 ( .A(n13186), .B(n17237), .Y(n13198) );
  sky130_fd_sc_hd__nand2_1 U20157 ( .A(n15684), .B(n18764), .Y(n15155) );
  sky130_fd_sc_hd__nor2_1 U20158 ( .A(n19140), .B(n13182), .Y(n18706) );
  sky130_fd_sc_hd__nand2_1 U20159 ( .A(n18706), .B(n21101), .Y(n18699) );
  sky130_fd_sc_hd__nor2_1 U20160 ( .A(n15155), .B(n18699), .Y(n13187) );
  sky130_fd_sc_hd__nand2_1 U20161 ( .A(n19124), .B(n19866), .Y(n19755) );
  sky130_fd_sc_hd__nand3_1 U20162 ( .A(n15394), .B(n19140), .C(n21360), .Y(
        n19810) );
  sky130_fd_sc_hd__nand3_1 U20163 ( .A(n19755), .B(n19764), .C(n19810), .Y(
        n19483) );
  sky130_fd_sc_hd__nor2_1 U20164 ( .A(n13187), .B(n19483), .Y(n19775) );
  sky130_fd_sc_hd__nand3_1 U20165 ( .A(n19738), .B(n19523), .C(n13234), .Y(
        n19516) );
  sky130_fd_sc_hd__nand2_1 U20166 ( .A(n19712), .B(n15516), .Y(n19432) );
  sky130_fd_sc_hd__nand4_1 U20167 ( .A(n19775), .B(n19739), .C(n13188), .D(
        n19432), .Y(n13189) );
  sky130_fd_sc_hd__nand2_1 U20168 ( .A(n13189), .B(n21103), .Y(n13197) );
  sky130_fd_sc_hd__nand3_1 U20169 ( .A(n19755), .B(n19523), .C(n13234), .Y(
        n13243) );
  sky130_fd_sc_hd__nor2_1 U20170 ( .A(n13235), .B(n15409), .Y(n19801) );
  sky130_fd_sc_hd__nand2_1 U20171 ( .A(n19505), .B(n13191), .Y(n19706) );
  sky130_fd_sc_hd__nand2_1 U20172 ( .A(n19712), .B(n15106), .Y(n19522) );
  sky130_fd_sc_hd__and3_1 U20173 ( .A(n19706), .B(n15396), .C(n19522), .X(
        n13192) );
  sky130_fd_sc_hd__nand4_1 U20174 ( .A(n19801), .B(n13192), .C(n19764), .D(
        n19777), .Y(n13193) );
  sky130_fd_sc_hd__inv_2 U20175 ( .A(n12089), .Y(n19804) );
  sky130_fd_sc_hd__o21ai_1 U20176 ( .A1(n13243), .A2(n13193), .B1(n19804), .Y(
        n13196) );
  sky130_fd_sc_hd__nor2_1 U20177 ( .A(n11150), .B(n18744), .Y(n18695) );
  sky130_fd_sc_hd__nand3_1 U20178 ( .A(n15394), .B(n18695), .C(n21101), .Y(
        n19782) );
  sky130_fd_sc_hd__nand2_1 U20179 ( .A(n19523), .B(n19782), .Y(n13205) );
  sky130_fd_sc_hd__a21oi_1 U20180 ( .A1(n19712), .A2(n19140), .B1(n15435), .Y(
        n13229) );
  sky130_fd_sc_hd__o31ai_1 U20181 ( .A1(n18712), .A2(n13179), .A3(n18699), 
        .B1(n13229), .Y(n13194) );
  sky130_fd_sc_hd__o21ai_1 U20182 ( .A1(n13205), .A2(n13194), .B1(n19816), .Y(
        n13195) );
  sky130_fd_sc_hd__nand4_1 U20183 ( .A(n13198), .B(n13197), .C(n13196), .D(
        n13195), .Y(n13200) );
  sky130_fd_sc_hd__nor2_1 U20184 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(j202_soc_core_bootrom_00_address_w[8]), .Y(n20126) );
  sky130_fd_sc_hd__a22oi_1 U20185 ( .A1(n15605), .A2(n13201), .B1(n13200), 
        .B2(n20126), .Y(n13254) );
  sky130_fd_sc_hd__nand2_1 U20186 ( .A(n19712), .B(n15610), .Y(n19811) );
  sky130_fd_sc_hd__nand2_1 U20187 ( .A(n18712), .B(n21101), .Y(n13202) );
  sky130_fd_sc_hd__nor2_1 U20188 ( .A(n18713), .B(n13202), .Y(n18703) );
  sky130_fd_sc_hd__nand2_1 U20189 ( .A(n18703), .B(n19129), .Y(n19781) );
  sky130_fd_sc_hd__nand2_1 U20190 ( .A(n19811), .B(n19781), .Y(n19509) );
  sky130_fd_sc_hd__nor2_1 U20191 ( .A(n13220), .B(n19509), .Y(n19767) );
  sky130_fd_sc_hd__nand2_1 U20192 ( .A(n19767), .B(n15396), .Y(n13204) );
  sky130_fd_sc_hd__nor2_1 U20193 ( .A(n15747), .B(n20034), .Y(n19521) );
  sky130_fd_sc_hd__nand2_1 U20194 ( .A(n19523), .B(n15431), .Y(n19511) );
  sky130_fd_sc_hd__nor2_1 U20195 ( .A(n19521), .B(n19511), .Y(n19437) );
  sky130_fd_sc_hd__nor2_1 U20196 ( .A(n18712), .B(n13203), .Y(n18715) );
  sky130_fd_sc_hd__nand2_1 U20197 ( .A(n18715), .B(n15684), .Y(n19694) );
  sky130_fd_sc_hd__nand2b_1 U20198 ( .A_N(n19694), .B(n18744), .Y(n19715) );
  sky130_fd_sc_hd__nand2_1 U20199 ( .A(n19715), .B(n19755), .Y(n19795) );
  sky130_fd_sc_hd__nand2_1 U20200 ( .A(n19437), .B(n19825), .Y(n15426) );
  sky130_fd_sc_hd__o21ai_1 U20201 ( .A1(n13204), .A2(n15426), .B1(n21103), .Y(
        n13214) );
  sky130_fd_sc_hd__nand2_1 U20202 ( .A(n20199), .B(n20531), .Y(n19783) );
  sky130_fd_sc_hd__nand2_1 U20203 ( .A(n19783), .B(n19490), .Y(n19434) );
  sky130_fd_sc_hd__nand2_1 U20204 ( .A(n19827), .B(n18744), .Y(n19765) );
  sky130_fd_sc_hd__nand4_1 U20205 ( .A(n19480), .B(n19512), .C(n19517), .D(
        n19765), .Y(n13208) );
  sky130_fd_sc_hd__nand2b_1 U20206 ( .A_N(n19694), .B(n19140), .Y(n19812) );
  sky130_fd_sc_hd__nand2_1 U20207 ( .A(n19812), .B(n19810), .Y(n19796) );
  sky130_fd_sc_hd__nand2_1 U20208 ( .A(n20199), .B(n19129), .Y(n19729) );
  sky130_fd_sc_hd__nand4b_1 U20209 ( .A_N(n19509), .B(n19814), .C(n19729), .D(
        n19763), .Y(n13206) );
  sky130_fd_sc_hd__o31a_1 U20210 ( .A1(n15424), .A2(n19796), .A3(n13206), .B1(
        n17237), .X(n13207) );
  sky130_fd_sc_hd__a21oi_1 U20211 ( .A1(n13208), .A2(n19804), .B1(n13207), .Y(
        n13213) );
  sky130_fd_sc_hd__nand2_1 U20212 ( .A(n18712), .B(n19140), .Y(n13209) );
  sky130_fd_sc_hd__nor2_1 U20213 ( .A(n17265), .B(n13209), .Y(n18753) );
  sky130_fd_sc_hd__nand2_1 U20214 ( .A(n18753), .B(n19129), .Y(n19809) );
  sky130_fd_sc_hd__nand4_1 U20215 ( .A(n19771), .B(n19783), .C(n19809), .D(
        n19770), .Y(n13210) );
  sky130_fd_sc_hd__nand2_1 U20216 ( .A(n19814), .B(n19706), .Y(n19797) );
  sky130_fd_sc_hd__nand2_1 U20218 ( .A(n19813), .B(n19729), .Y(n13233) );
  sky130_fd_sc_hd__nand2_1 U20219 ( .A(n19726), .B(n12089), .Y(n19486) );
  sky130_fd_sc_hd__nand2_1 U20220 ( .A(n13233), .B(n19486), .Y(n13211) );
  sky130_fd_sc_hd__nand4_1 U20221 ( .A(n13214), .B(n13213), .C(n13212), .D(
        n13211), .Y(n13215) );
  sky130_fd_sc_hd__nand2_1 U20222 ( .A(n13215), .B(n20196), .Y(n13253) );
  sky130_fd_sc_hd__and3_1 U20223 ( .A(n19755), .B(n19783), .C(n19753), .X(
        n19467) );
  sky130_fd_sc_hd__nand2_1 U20224 ( .A(n19504), .B(n18695), .Y(n19707) );
  sky130_fd_sc_hd__nand2b_1 U20225 ( .A_N(n19707), .B(n21145), .Y(n19754) );
  sky130_fd_sc_hd__nand2_1 U20226 ( .A(n19729), .B(n19754), .Y(n19698) );
  sky130_fd_sc_hd__nand4_1 U20227 ( .A(n19467), .B(n19720), .C(n19432), .D(
        n19809), .Y(n13219) );
  sky130_fd_sc_hd__nand2_1 U20228 ( .A(n19714), .B(n19706), .Y(n15438) );
  sky130_fd_sc_hd__o21ai_1 U20229 ( .A1(n15438), .A2(n19511), .B1(n19486), .Y(
        n13217) );
  sky130_fd_sc_hd__nand2b_1 U20230 ( .A_N(n15435), .B(n19522), .Y(n19470) );
  sky130_fd_sc_hd__nand2_1 U20232 ( .A(n13217), .B(n13216), .Y(n13218) );
  sky130_fd_sc_hd__a21oi_1 U20233 ( .A1(n13219), .A2(n19804), .B1(n13218), .Y(
        n13226) );
  sky130_fd_sc_hd__nor2_1 U20234 ( .A(n19708), .B(n19483), .Y(n19481) );
  sky130_fd_sc_hd__nor2_1 U20235 ( .A(n19521), .B(n13220), .Y(n13221) );
  sky130_fd_sc_hd__nand4_1 U20236 ( .A(n19481), .B(n19512), .C(n13221), .D(
        n19754), .Y(n13222) );
  sky130_fd_sc_hd__nand2_1 U20237 ( .A(n13222), .B(n17237), .Y(n13225) );
  sky130_fd_sc_hd__nand2b_1 U20238 ( .A_N(n19509), .B(n19753), .Y(n19716) );
  sky130_fd_sc_hd__nand2b_1 U20239 ( .A_N(n20034), .B(n20810), .Y(n19463) );
  sky130_fd_sc_hd__nand2_1 U20240 ( .A(n19463), .B(n19809), .Y(n19733) );
  sky130_fd_sc_hd__nor2_1 U20241 ( .A(n19733), .B(n13240), .Y(n19518) );
  sky130_fd_sc_hd__nand4_1 U20242 ( .A(n19711), .B(n19441), .C(n19720), .D(
        n19518), .Y(n13223) );
  sky130_fd_sc_hd__nand2_1 U20243 ( .A(n13223), .B(n21103), .Y(n13224) );
  sky130_fd_sc_hd__nand3_1 U20244 ( .A(n13226), .B(n13225), .C(n13224), .Y(
        n13227) );
  sky130_fd_sc_hd__nor2_1 U20245 ( .A(n13199), .B(n17264), .Y(n20194) );
  sky130_fd_sc_hd__nand2_1 U20246 ( .A(n13227), .B(n20194), .Y(n13252) );
  sky130_fd_sc_hd__nand2_1 U20247 ( .A(n19432), .B(n19810), .Y(n13228) );
  sky130_fd_sc_hd__nand2_1 U20248 ( .A(n19765), .B(n19701), .Y(n13239) );
  sky130_fd_sc_hd__nor2_1 U20249 ( .A(n13228), .B(n13239), .Y(n19759) );
  sky130_fd_sc_hd__nand2b_1 U20250 ( .A_N(n19507), .B(n19729), .Y(n19821) );
  sky130_fd_sc_hd__nor3_1 U20251 ( .A(n13235), .B(n13230), .C(n19821), .Y(
        n13231) );
  sky130_fd_sc_hd__nand4_1 U20252 ( .A(n19759), .B(n13231), .C(n19467), .D(
        n19513), .Y(n13232) );
  sky130_fd_sc_hd__nand2_1 U20253 ( .A(n13232), .B(n19804), .Y(n13249) );
  sky130_fd_sc_hd__nor2_1 U20254 ( .A(n13241), .B(n13233), .Y(n15425) );
  sky130_fd_sc_hd__nand2_1 U20255 ( .A(n19765), .B(n13234), .Y(n19807) );
  sky130_fd_sc_hd__nor2_1 U20256 ( .A(n19509), .B(n19807), .Y(n15430) );
  sky130_fd_sc_hd__nor2_1 U20257 ( .A(n13236), .B(n13235), .Y(n13237) );
  sky130_fd_sc_hd__nand4_1 U20258 ( .A(n15425), .B(n19480), .C(n19823), .D(
        n13237), .Y(n13238) );
  sky130_fd_sc_hd__nand2_1 U20259 ( .A(n13238), .B(n19816), .Y(n13248) );
  sky130_fd_sc_hd__nor2_1 U20260 ( .A(n13241), .B(n13240), .Y(n19695) );
  sky130_fd_sc_hd__and3_1 U20261 ( .A(n19783), .B(n19771), .C(n19753), .X(
        n19446) );
  sky130_fd_sc_hd__nand4_1 U20262 ( .A(n19773), .B(n19823), .C(n19695), .D(
        n19446), .Y(n13242) );
  sky130_fd_sc_hd__nand2_1 U20263 ( .A(n13242), .B(n17237), .Y(n13247) );
  sky130_fd_sc_hd__nand2_1 U20264 ( .A(n19763), .B(n15396), .Y(n15455) );
  sky130_fd_sc_hd__nor2_1 U20265 ( .A(n15455), .B(n15438), .Y(n19440) );
  sky130_fd_sc_hd__nand2_1 U20266 ( .A(n19812), .B(n19701), .Y(n15413) );
  sky130_fd_sc_hd__nand4_1 U20267 ( .A(n19440), .B(n13244), .C(n19719), .D(
        n19754), .Y(n13245) );
  sky130_fd_sc_hd__nand2_1 U20268 ( .A(n13245), .B(n21103), .Y(n13246) );
  sky130_fd_sc_hd__nand4_1 U20269 ( .A(n13249), .B(n13248), .C(n13247), .D(
        n13246), .Y(n13250) );
  sky130_fd_sc_hd__nor2_1 U20270 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .B(n20485), .Y(n20235) );
  sky130_fd_sc_hd__nand2_1 U20271 ( .A(n13250), .B(n20235), .Y(n13251) );
  sky130_fd_sc_hd__nand4_1 U20272 ( .A(n13254), .B(n13253), .C(n13252), .D(
        n13251), .Y(n13285) );
  sky130_fd_sc_hd__nor2_1 U20273 ( .A(j202_soc_core_bootrom_00_address_w[14]), 
        .B(j202_soc_core_bootrom_00_address_w[12]), .Y(n13256) );
  sky130_fd_sc_hd__nor2_1 U20274 ( .A(j202_soc_core_bootrom_00_address_w[15]), 
        .B(j202_soc_core_bootrom_00_address_w[13]), .Y(n13255) );
  sky130_fd_sc_hd__nand2_1 U20275 ( .A(n13256), .B(n13255), .Y(n13259) );
  sky130_fd_sc_hd__nor2_1 U20276 ( .A(j202_soc_core_bootrom_00_address_w[17]), 
        .B(j202_soc_core_bootrom_00_address_w[16]), .Y(n13257) );
  sky130_fd_sc_hd__nand4_1 U20277 ( .A(n13274), .B(n13257), .C(
        j202_soc_core_j22_cpu_ma_M_area[1]), .D(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[6]), .Y(n13258) );
  sky130_fd_sc_hd__mux2_2 U20278 ( .A0(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[4]), .A1(
        j202_soc_core_aquc_ADR__4_), .S(n29435), .X(n19593) );
  sky130_fd_sc_hd__mux2_2 U20279 ( .A0(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[3]), .A1(
        j202_soc_core_aquc_ADR__3_), .S(n29435), .X(n22760) );
  sky130_fd_sc_hd__nor2_1 U20280 ( .A(n19593), .B(n22760), .Y(n28204) );
  sky130_fd_sc_hd__nor2_1 U20281 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[6]), .B(n13260), .Y(n13275) );
  sky130_fd_sc_hd__nor2_1 U20282 ( .A(j202_soc_core_j22_cpu_ma_M_area[0]), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[5]), .Y(n13262) );
  sky130_fd_sc_hd__nand3_1 U20283 ( .A(n13275), .B(n13262), .C(n13261), .Y(
        n13272) );
  sky130_fd_sc_hd__nor2_1 U20284 ( .A(j202_soc_core_aquc_ADR__7_), .B(
        j202_soc_core_aquc_ADR__6_), .Y(n13265) );
  sky130_fd_sc_hd__nand3_1 U20285 ( .A(n29435), .B(n13265), .C(n13264), .Y(
        n17200) );
  sky130_fd_sc_hd__nand2b_1 U20286 ( .A_N(n17200), .B(n13266), .Y(n13271) );
  sky130_fd_sc_hd__nand2_1 U20287 ( .A(n13268), .B(n13267), .Y(n13269) );
  sky130_fd_sc_hd__mux2_2 U20288 ( .A0(n13270), .A1(n13269), .S(n29435), .X(
        n17198) );
  sky130_fd_sc_hd__nor2_1 U20289 ( .A(n13271), .B(n17198), .Y(n19598) );
  sky130_fd_sc_hd__nor2_1 U20290 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[3]), .B(n13272), .Y(n17192) );
  sky130_fd_sc_hd__nand2_1 U20291 ( .A(n17192), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[2]), .Y(n21515) );
  sky130_fd_sc_hd__nand2_1 U20292 ( .A(n20540), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[50]), .Y(n13282) );
  sky130_fd_sc_hd__nand2_1 U20293 ( .A(n21513), .B(j202_soc_core_uart_div1[2]), 
        .Y(n13281) );
  sky130_fd_sc_hd__nand2_1 U20294 ( .A(n13274), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[5]), .Y(n13277) );
  sky130_fd_sc_hd__nand2_1 U20295 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[18]), .Y(n13280) );
  sky130_fd_sc_hd__nand3_1 U20296 ( .A(n17192), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[1]), .C(n13278), .Y(n21512) );
  sky130_fd_sc_hd__nand2_1 U20297 ( .A(n20759), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[82]), .Y(n13279) );
  sky130_fd_sc_hd__nand4_1 U20298 ( .A(n13282), .B(n13281), .C(n13280), .D(
        n13279), .Y(n13283) );
  sky130_fd_sc_hd__a21oi_1 U20299 ( .A1(n20786), .A2(
        j202_soc_core_bldc_core_00_pwm_duty[6]), .B1(n13283), .Y(n13284) );
  sky130_fd_sc_hd__a21boi_1 U20300 ( .A1(n13285), .A2(n21629), .B1_N(n13284), 
        .Y(n20257) );
  sky130_fd_sc_hd__nand2_1 U20301 ( .A(n19236), .B(n20257), .Y(n26164) );
  sky130_fd_sc_hd__nand2_1 U20302 ( .A(n24673), .B(
        j202_soc_core_j22_cpu_ifetchl), .Y(n23883) );
  sky130_fd_sc_hd__nand2_1 U20303 ( .A(n24771), .B(
        j202_soc_core_j22_cpu_regop_We__2_), .Y(n13288) );
  sky130_fd_sc_hd__nor2_1 U20304 ( .A(n23888), .B(n13288), .Y(n13290) );
  sky130_fd_sc_hd__nor2_1 U20305 ( .A(j202_soc_core_j22_cpu_regop_We__3_), .B(
        n13305), .Y(n23836) );
  sky130_fd_sc_hd__nor2_1 U20306 ( .A(j202_soc_core_j22_cpu_regop_We__0_), .B(
        n23842), .Y(n13289) );
  sky130_fd_sc_hd__mux2i_1 U20307 ( .A0(n13290), .A1(n13289), .S(n12347), .Y(
        n13292) );
  sky130_fd_sc_hd__nor2_1 U20308 ( .A(n12040), .B(
        j202_soc_core_j22_cpu_memop_MEM__1_), .Y(n15656) );
  sky130_fd_sc_hd__nand2_1 U20309 ( .A(n15656), .B(n24647), .Y(n16933) );
  sky130_fd_sc_hd__nand2b_1 U20310 ( .A_N(n16933), .B(
        j202_soc_core_j22_cpu_memop_MEM__0_), .Y(n28103) );
  sky130_fd_sc_hd__nor2_1 U20311 ( .A(j202_soc_core_j22_cpu_memop_MEM__0_), 
        .B(j202_soc_core_j22_cpu_memop_MEM__3_), .Y(n15654) );
  sky130_fd_sc_hd__nand3_1 U20312 ( .A(n15654), .B(
        j202_soc_core_j22_cpu_memop_MEM__1_), .C(n12041), .Y(n13291) );
  sky130_fd_sc_hd__nand3_1 U20313 ( .A(n13292), .B(n28103), .C(n13291), .Y(
        n13293) );
  sky130_fd_sc_hd__nand3_1 U20314 ( .A(n23413), .B(n28373), .C(n20428), .Y(
        n23412) );
  sky130_fd_sc_hd__nand2_1 U20315 ( .A(n23836), .B(
        j202_soc_core_j22_cpu_regop_We__0_), .Y(n13351) );
  sky130_fd_sc_hd__nor2_1 U20316 ( .A(n12348), .B(n13351), .Y(n23755) );
  sky130_fd_sc_hd__xnor2_1 U20318 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__2_), 
        .B(n12032), .Y(n13298) );
  sky130_fd_sc_hd__xnor2_1 U20319 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__1_), 
        .B(n12030), .Y(n13297) );
  sky130_fd_sc_hd__xnor2_1 U20320 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__3_), 
        .B(n12340), .Y(n13296) );
  sky130_fd_sc_hd__xnor2_1 U20321 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__0_), 
        .B(n12339), .Y(n13295) );
  sky130_fd_sc_hd__nand4_1 U20322 ( .A(n13298), .B(n13297), .C(n13296), .D(
        n13295), .Y(n13299) );
  sky130_fd_sc_hd__a21o_1 U20323 ( .A1(n13300), .A2(n13294), .B1(n13299), .X(
        n13316) );
  sky130_fd_sc_hd__nor2_1 U20324 ( .A(n12347), .B(n13351), .Y(n23498) );
  sky130_fd_sc_hd__nand2_1 U20325 ( .A(j202_soc_core_j22_cpu_regop_other__1_), 
        .B(j202_soc_core_j22_cpu_regop_other__0_), .Y(n13428) );
  sky130_fd_sc_hd__nand2_1 U20327 ( .A(n13301), .B(
        j202_soc_core_j22_cpu_regop_Rs__1_), .Y(n22084) );
  sky130_fd_sc_hd__nand2_1 U20328 ( .A(j202_soc_core_j22_cpu_regop_Ra__0_), 
        .B(j202_soc_core_j22_cpu_regop_Ra__1_), .Y(n13303) );
  sky130_fd_sc_hd__nand2_1 U20329 ( .A(n12054), .B(
        j202_soc_core_j22_cpu_regop_Rb__1_), .Y(n13337) );
  sky130_fd_sc_hd__nand4_1 U20330 ( .A(n13304), .B(n22084), .C(n13303), .D(
        n16488), .Y(n13350) );
  sky130_fd_sc_hd__nor2_1 U20331 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__1_), 
        .B(j202_soc_core_j22_cpu_regop_M_Rn__0_), .Y(n23807) );
  sky130_fd_sc_hd__nor2_1 U20332 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__2_), 
        .B(j202_soc_core_j22_cpu_regop_M_Rn__3_), .Y(n23760) );
  sky130_fd_sc_hd__nand3_1 U20333 ( .A(n13350), .B(n23807), .C(n23760), .Y(
        n13315) );
  sky130_fd_sc_hd__nor2_1 U20334 ( .A(n12347), .B(n23888), .Y(n23889) );
  sky130_fd_sc_hd__nand2_1 U20335 ( .A(n23889), .B(n13305), .Y(n24715) );
  sky130_fd_sc_hd__nor2_1 U20336 ( .A(j202_soc_core_j22_cpu_regop_We__0_), .B(
        n24715), .Y(n23753) );
  sky130_fd_sc_hd__nand2_1 U20337 ( .A(n12054), .B(n16523), .Y(n13307) );
  sky130_fd_sc_hd__nand2_1 U20338 ( .A(n22996), .B(
        j202_soc_core_j22_cpu_regop_Rs__0_), .Y(n13306) );
  sky130_fd_sc_hd__nand3_1 U20339 ( .A(n13308), .B(n13307), .C(n13306), .Y(
        n13353) );
  sky130_fd_sc_hd__xor2_1 U20340 ( .A(j202_soc_core_j22_cpu_regop_Rm__0_), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__0_), .X(n13310) );
  sky130_fd_sc_hd__xor2_1 U20341 ( .A(j202_soc_core_j22_cpu_regop_Rm__1_), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__1_), .X(n13309) );
  sky130_fd_sc_hd__nor2_1 U20342 ( .A(n13310), .B(n13309), .Y(n13313) );
  sky130_fd_sc_hd__xnor2_1 U20343 ( .A(j202_soc_core_j22_cpu_regop_Rm__3_), 
        .B(j202_soc_core_j22_cpu_regop_M_Rn__3_), .Y(n13312) );
  sky130_fd_sc_hd__xnor2_1 U20344 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__2_), 
        .B(j202_soc_core_j22_cpu_regop_Rm__2_), .Y(n13311) );
  sky130_fd_sc_hd__nand4_1 U20345 ( .A(n13353), .B(n13313), .C(n13312), .D(
        n13311), .Y(n13314) );
  sky130_fd_sc_hd__nand3_1 U20346 ( .A(n13316), .B(n13315), .C(n13314), .Y(
        n13317) );
  sky130_fd_sc_hd__nand3_1 U20347 ( .A(n13341), .B(n23831), .C(
        j202_soc_core_j22_cpu_regop_M_Wm__1_), .Y(n13336) );
  sky130_fd_sc_hd__nor2_1 U20348 ( .A(n24718), .B(n13336), .Y(n23750) );
  sky130_fd_sc_hd__nand2_1 U20349 ( .A(n13317), .B(n23750), .Y(n13360) );
  sky130_fd_sc_hd__nor2_1 U20350 ( .A(j202_soc_core_j22_cpu_macop_MAC_[3]), 
        .B(j202_soc_core_j22_cpu_macop_MAC_[2]), .Y(n24289) );
  sky130_fd_sc_hd__nand4_1 U20351 ( .A(n24289), .B(n28053), .C(n27763), .D(
        n27828), .Y(n13335) );
  sky130_fd_sc_hd__nand3_1 U20352 ( .A(n13322), .B(n28044), .C(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[4]), .Y(n24285) );
  sky130_fd_sc_hd__nand2_1 U20353 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]), .B(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .Y(n13318) );
  sky130_fd_sc_hd__nand2_1 U20354 ( .A(n13319), .B(n13318), .Y(n23625) );
  sky130_fd_sc_hd__nand2_1 U20355 ( .A(n13321), .B(n13320), .Y(n24284) );
  sky130_fd_sc_hd__nor2_1 U20356 ( .A(j202_soc_core_j22_cpu_ml_M_macop_MAC_[4]), .B(n13322), .Y(n13328) );
  sky130_fd_sc_hd__o211ai_1 U20357 ( .A1(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[3]), .A2(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .B1(n24284), .C1(n13328), 
        .Y(n24283) );
  sky130_fd_sc_hd__nand2_1 U20358 ( .A(n23625), .B(n24283), .Y(n24672) );
  sky130_fd_sc_hd__nand2_1 U20360 ( .A(n13323), .B(n17355), .Y(n17351) );
  sky130_fd_sc_hd__inv_2 U20361 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), 
        .Y(n28435) );
  sky130_fd_sc_hd__nand2_2 U20362 ( .A(n28435), .B(n24677), .Y(n24674) );
  sky130_fd_sc_hd__nand2_1 U20363 ( .A(n17351), .B(n24674), .Y(n13333) );
  sky130_fd_sc_hd__inv_2 U20364 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]), 
        .Y(n18680) );
  sky130_fd_sc_hd__nor2_2 U20365 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[4]), .B(n18680), .Y(n24675) );
  sky130_fd_sc_hd__nand2_1 U20366 ( .A(n13333), .B(n24675), .Y(n13327) );
  sky130_fd_sc_hd__nand2_1 U20367 ( .A(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .Y(n17350) );
  sky130_fd_sc_hd__nand2_1 U20368 ( .A(n24675), .B(n13324), .Y(n28047) );
  sky130_fd_sc_hd__nand2_1 U20369 ( .A(j202_soc_core_j22_cpu_macop_MAC_[3]), 
        .B(j202_soc_core_j22_cpu_macop_MAC_[0]), .Y(n24286) );
  sky130_fd_sc_hd__nand2_1 U20370 ( .A(n24286), .B(n28053), .Y(n24288) );
  sky130_fd_sc_hd__nand2_1 U20371 ( .A(n24288), .B(
        j202_soc_core_j22_cpu_macop_MAC_[2]), .Y(n24428) );
  sky130_fd_sc_hd__nor2_1 U20372 ( .A(j202_soc_core_j22_cpu_macop_MAC_[4]), 
        .B(n24428), .Y(n24670) );
  sky130_fd_sc_hd__o21ai_1 U20373 ( .A1(n28053), .A2(n24286), .B1(n24670), .Y(
        n13326) );
  sky130_fd_sc_hd__nand3_1 U20374 ( .A(n24289), .B(
        j202_soc_core_j22_cpu_macop_MAC_[4]), .C(n28053), .Y(n24665) );
  sky130_fd_sc_hd__nand2_1 U20375 ( .A(n13326), .B(n24665), .Y(n27756) );
  sky130_fd_sc_hd__o2bb2ai_1 U20376 ( .B1(n24672), .B2(n13325), .A1_N(n13327), 
        .A2_N(n27756), .Y(n13329) );
  sky130_fd_sc_hd__nand2_1 U20377 ( .A(n13329), .B(n28538), .Y(n13334) );
  sky130_fd_sc_hd__nor2_1 U20378 ( .A(j202_soc_core_j22_cpu_macop_MAC_[4]), 
        .B(n28053), .Y(n13331) );
  sky130_fd_sc_hd__nand2_1 U20379 ( .A(n28435), .B(n11478), .Y(n13330) );
  sky130_fd_sc_hd__nand4_1 U20380 ( .A(n17965), .B(n24289), .C(n13331), .D(
        n13330), .Y(n13332) );
  sky130_fd_sc_hd__a2bb2oi_1 U20381 ( .B1(n13335), .B2(n13334), .A1_N(n13333), 
        .A2_N(n13332), .Y(n27757) );
  sky130_fd_sc_hd__inv_2 U20382 ( .A(j202_soc_core_j22_cpu_regop_other__1_), 
        .Y(n18859) );
  sky130_fd_sc_hd__inv_2 U20383 ( .A(n16487), .Y(n16533) );
  sky130_fd_sc_hd__nor2_1 U20384 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__2_), 
        .B(n13336), .Y(n23887) );
  sky130_fd_sc_hd__nand2_1 U20385 ( .A(n16533), .B(n23887), .Y(n16921) );
  sky130_fd_sc_hd__nand2_1 U20388 ( .A(n16491), .B(n22983), .Y(n13340) );
  sky130_fd_sc_hd__nand2_1 U20389 ( .A(n18859), .B(
        j202_soc_core_j22_cpu_regop_other__2_), .Y(n13425) );
  sky130_fd_sc_hd__nor2_1 U20390 ( .A(n18869), .B(n13425), .Y(n13338) );
  sky130_fd_sc_hd__nand2_1 U20391 ( .A(n13338), .B(n13431), .Y(n14373) );
  sky130_fd_sc_hd__nand2_1 U20392 ( .A(n13338), .B(n11094), .Y(n22894) );
  sky130_fd_sc_hd__nand2_1 U20393 ( .A(n14373), .B(n22894), .Y(n13339) );
  sky130_fd_sc_hd__mux2_2 U20394 ( .A0(n13340), .A1(n13339), .S(
        j202_soc_core_j22_cpu_regop_M_Wm__2_), .X(n13342) );
  sky130_fd_sc_hd__nor2_1 U20395 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__3_), 
        .B(n13341), .Y(n23840) );
  sky130_fd_sc_hd__nand3_1 U20396 ( .A(n13342), .B(
        j202_soc_core_j22_cpu_regop_M_Wm__1_), .C(n23840), .Y(n13343) );
  sky130_fd_sc_hd__nand3_1 U20397 ( .A(n27757), .B(n16921), .C(n13343), .Y(
        n13349) );
  sky130_fd_sc_hd__nor2_1 U20398 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .B(n21709), .Y(n26205) );
  sky130_fd_sc_hd__nand3_1 U20399 ( .A(n26205), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[5]), .C(n26270), .Y(n26373) );
  sky130_fd_sc_hd__nor2_1 U20400 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[0]), 
        .B(n26373), .Y(n26186) );
  sky130_fd_sc_hd__nand3_1 U20401 ( .A(n26205), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[0]), .C(n26142), .Y(n13345) );
  sky130_fd_sc_hd__nor2_1 U20402 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[2]), 
        .B(n18809), .Y(n26139) );
  sky130_fd_sc_hd__nand2_1 U20403 ( .A(n26295), .B(n26139), .Y(n13344) );
  sky130_fd_sc_hd__mux2i_1 U20404 ( .A0(n13345), .A1(n13344), .S(n26208), .Y(
        n13346) );
  sky130_fd_sc_hd__nor2_1 U20405 ( .A(n26186), .B(n13346), .Y(n13348) );
  sky130_fd_sc_hd__nor2_1 U20406 ( .A(n13348), .B(n13362), .Y(n24708) );
  sky130_fd_sc_hd__nor2_1 U20407 ( .A(n13349), .B(n24708), .Y(n13359) );
  sky130_fd_sc_hd__nor2_1 U20409 ( .A(n12030), .B(n12036), .Y(n13455) );
  sky130_fd_sc_hd__nand2_1 U20410 ( .A(n13483), .B(n13455), .Y(n13474) );
  sky130_fd_sc_hd__nor2_1 U20411 ( .A(n13474), .B(n13351), .Y(n23499) );
  sky130_fd_sc_hd__a22oi_1 U20412 ( .A1(n13352), .A2(
        j202_soc_core_j22_cpu_regop_Ra__0_), .B1(n24673), .B2(n23499), .Y(
        n13355) );
  sky130_fd_sc_hd__nor2_1 U20413 ( .A(j202_soc_core_j22_cpu_regop_Rm__0_), .B(
        j202_soc_core_j22_cpu_regop_Rm__1_), .Y(n13390) );
  sky130_fd_sc_hd__buf_2 U20414 ( .A(n11091), .X(n23500) );
  sky130_fd_sc_hd__nand2_1 U20415 ( .A(n13353), .B(n23500), .Y(n13354) );
  sky130_fd_sc_hd__nand3_1 U20416 ( .A(n13356), .B(n13355), .C(n13354), .Y(
        n13357) );
  sky130_fd_sc_hd__nor2_1 U20417 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__1_), 
        .B(j202_soc_core_j22_cpu_regop_M_Wm__0_), .Y(n23641) );
  sky130_fd_sc_hd__and3_1 U20418 ( .A(n23641), .B(
        j202_soc_core_j22_cpu_regop_M_Wm__2_), .C(n23831), .X(n23832) );
  sky130_fd_sc_hd__nand2_1 U20419 ( .A(n13357), .B(n23832), .Y(n13358) );
  sky130_fd_sc_hd__nand2_1 U20420 ( .A(n15656), .B(n15654), .Y(n24305) );
  sky130_fd_sc_hd__nand2_1 U20421 ( .A(n23643), .B(n24302), .Y(n13363) );
  sky130_fd_sc_hd__nor2_1 U20422 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[2]), 
        .B(n26374), .Y(n18825) );
  sky130_fd_sc_hd__nand2_1 U20423 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[2]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[4]), .Y(n18827) );
  sky130_fd_sc_hd__nand2_1 U20424 ( .A(n26148), .B(
        j202_soc_core_j22_cpu_rfuo_sr__t_), .Y(n13366) );
  sky130_fd_sc_hd__o21ai_1 U20425 ( .A1(j202_soc_core_j22_cpu_rfuo_sr__t_), 
        .A2(n25818), .B1(n13366), .Y(n13368) );
  sky130_fd_sc_hd__nand2_1 U20426 ( .A(n18825), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[4]), .Y(n13367) );
  sky130_fd_sc_hd__nand2_1 U20427 ( .A(n26148), .B(n26208), .Y(n26210) );
  sky130_fd_sc_hd__o22a_1 U20428 ( .A1(n13367), .A2(n26145), .B1(
        j202_soc_core_j22_cpu_exuop_EXU_[1]), .B2(n26210), .X(n28102) );
  sky130_fd_sc_hd__nor2_1 U20429 ( .A(n28104), .B(n13378), .Y(n24036) );
  sky130_fd_sc_hd__nand2b_4 U20430 ( .A_N(n14588), .B(n24036), .Y(n22705) );
  sky130_fd_sc_hd__nand2_1 U20431 ( .A(j202_soc_core_j22_cpu_pc[7]), .B(
        j202_soc_core_j22_cpu_pc[8]), .Y(n13369) );
  sky130_fd_sc_hd__nand2_1 U20432 ( .A(j202_soc_core_j22_cpu_pc[5]), .B(
        j202_soc_core_j22_cpu_pc[6]), .Y(n19099) );
  sky130_fd_sc_hd__nor2_1 U20433 ( .A(n13369), .B(n19099), .Y(n13371) );
  sky130_fd_sc_hd__nand2_1 U20434 ( .A(j202_soc_core_j22_cpu_pc[3]), .B(
        j202_soc_core_j22_cpu_pc[4]), .Y(n13370) );
  sky130_fd_sc_hd__nand2_1 U20435 ( .A(j202_soc_core_j22_cpu_pc[1]), .B(
        j202_soc_core_j22_cpu_pc[2]), .Y(n20445) );
  sky130_fd_sc_hd__nor2_1 U20436 ( .A(n13370), .B(n20445), .Y(n19098) );
  sky130_fd_sc_hd__nand2_1 U20437 ( .A(n13371), .B(n19098), .Y(n20929) );
  sky130_fd_sc_hd__nand2_1 U20438 ( .A(j202_soc_core_j22_cpu_pc[11]), .B(
        j202_soc_core_j22_cpu_pc[12]), .Y(n13372) );
  sky130_fd_sc_hd__nand2_1 U20439 ( .A(j202_soc_core_j22_cpu_pc[9]), .B(
        j202_soc_core_j22_cpu_pc[10]), .Y(n20930) );
  sky130_fd_sc_hd__nor2_1 U20440 ( .A(n13372), .B(n20930), .Y(n20960) );
  sky130_fd_sc_hd__nand2_1 U20441 ( .A(j202_soc_core_j22_cpu_pc[15]), .B(
        j202_soc_core_j22_cpu_pc[16]), .Y(n13373) );
  sky130_fd_sc_hd__nand2_1 U20442 ( .A(j202_soc_core_j22_cpu_pc[13]), .B(
        j202_soc_core_j22_cpu_pc[14]), .Y(n20976) );
  sky130_fd_sc_hd__nor2_1 U20443 ( .A(n13373), .B(n20976), .Y(n13374) );
  sky130_fd_sc_hd__nand2_1 U20444 ( .A(n20960), .B(n13374), .Y(n13375) );
  sky130_fd_sc_hd__nor2_1 U20445 ( .A(n20929), .B(n13375), .Y(n16095) );
  sky130_fd_sc_hd__nor2_1 U20446 ( .A(n22849), .B(n21026), .Y(n13376) );
  sky130_fd_sc_hd__xnor2_1 U20447 ( .A(n13377), .B(n13376), .Y(n25896) );
  sky130_fd_sc_hd__nand2_1 U20448 ( .A(n22747), .B(n25896), .Y(n17084) );
  sky130_fd_sc_hd__nor2_1 U20449 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[0]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[3]), .Y(n18837) );
  sky130_fd_sc_hd__nand2_1 U20450 ( .A(n18837), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[4]), .Y(n21201) );
  sky130_fd_sc_hd__nor2_1 U20451 ( .A(n21201), .B(n13378), .Y(n24033) );
  sky130_fd_sc_hd__nand2_4 U20452 ( .A(n22745), .B(n22743), .Y(n21924) );
  sky130_fd_sc_hd__nand2_1 U20453 ( .A(n13381), .B(
        j202_soc_core_j22_cpu_regop_Rm__0_), .Y(n13393) );
  sky130_fd_sc_hd__nand2_1 U20454 ( .A(n13380), .B(
        j202_soc_core_j22_cpu_regop_Rm__3_), .Y(n13394) );
  sky130_fd_sc_hd__nor2_1 U20455 ( .A(n13393), .B(n13394), .Y(n13838) );
  sky130_fd_sc_hd__inv_2 U20456 ( .A(n13631), .Y(n23781) );
  sky130_fd_sc_hd__nand2_1 U20457 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[306]), .Y(n13389) );
  sky130_fd_sc_hd__nand2_1 U20458 ( .A(j202_soc_core_j22_cpu_regop_Rm__3_), 
        .B(j202_soc_core_j22_cpu_regop_Rm__0_), .Y(n13382) );
  sky130_fd_sc_hd__nand2_1 U20459 ( .A(n13381), .B(
        j202_soc_core_j22_cpu_regop_Rm__2_), .Y(n13414) );
  sky130_fd_sc_hd__nor2_1 U20460 ( .A(n13382), .B(n13414), .Y(n13383) );
  sky130_fd_sc_hd__inv_2 U20461 ( .A(n13839), .Y(n23823) );
  sky130_fd_sc_hd__nand2_1 U20462 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[433]), .Y(n13388) );
  sky130_fd_sc_hd__nand2_1 U20463 ( .A(n13413), .B(
        j202_soc_core_j22_cpu_regop_Rm__0_), .Y(n13384) );
  sky130_fd_sc_hd__nor2_1 U20464 ( .A(n13384), .B(n13414), .Y(n13840) );
  sky130_fd_sc_hd__inv_2 U20465 ( .A(n13707), .Y(n23802) );
  sky130_fd_sc_hd__nand2_1 U20466 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[178]), .Y(n13387) );
  sky130_fd_sc_hd__nand2_1 U20469 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[114]), .Y(n13386) );
  sky130_fd_sc_hd__nand4_1 U20470 ( .A(n13389), .B(n13388), .C(n13387), .D(
        n13386), .Y(n13400) );
  sky130_fd_sc_hd__nor2_1 U20471 ( .A(n13391), .B(n13394), .Y(n13835) );
  sky130_fd_sc_hd__nand2_1 U20472 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[274]), .Y(n13398) );
  sky130_fd_sc_hd__nand2_1 U20474 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[50]), .Y(n13397) );
  sky130_fd_sc_hd__nor2_1 U20475 ( .A(n13403), .B(n13394), .Y(n13836) );
  sky130_fd_sc_hd__nand2_1 U20476 ( .A(n23776), .B(
        j202_soc_core_j22_cpu_rf_gpr[369]), .Y(n13396) );
  sky130_fd_sc_hd__inv_2 U20477 ( .A(j202_soc_core_j22_cpu_regop_Rm__0_), .Y(
        n13412) );
  sky130_fd_sc_hd__nor2_1 U20479 ( .A(n13409), .B(n13394), .Y(n13837) );
  sky130_fd_sc_hd__nand2_1 U20480 ( .A(n16064), .B(
        j202_soc_core_j22_cpu_rf_gpr[337]), .Y(n13395) );
  sky130_fd_sc_hd__nand4_1 U20481 ( .A(n13398), .B(n13397), .C(n13396), .D(
        n13395), .Y(n13399) );
  sky130_fd_sc_hd__nor2_1 U20482 ( .A(n13400), .B(n13399), .Y(n13424) );
  sky130_fd_sc_hd__nor2_1 U20483 ( .A(n13402), .B(n13409), .Y(n13818) );
  sky130_fd_sc_hd__nand2_1 U20484 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[210]), .Y(n13407) );
  sky130_fd_sc_hd__nand2_1 U20485 ( .A(j202_soc_core_j22_cpu_regop_Rm__2_), 
        .B(j202_soc_core_j22_cpu_regop_Rm__3_), .Y(n13401) );
  sky130_fd_sc_hd__nor2_1 U20486 ( .A(n13401), .B(n13409), .Y(n13819) );
  sky130_fd_sc_hd__nand2_1 U20487 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[465]), .Y(n13406) );
  sky130_fd_sc_hd__nand2_1 U20489 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[497]), .Y(n13405) );
  sky130_fd_sc_hd__nand2_1 U20490 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[242]), .Y(n13404) );
  sky130_fd_sc_hd__nand4_1 U20491 ( .A(n13407), .B(n13406), .C(n13405), .D(
        n13404), .Y(n13422) );
  sky130_fd_sc_hd__nand2_1 U20492 ( .A(n16506), .B(
        j202_soc_core_j22_cpu_rf_gpr[18]), .Y(n13420) );
  sky130_fd_sc_hd__nor2_1 U20493 ( .A(n13409), .B(n13408), .Y(n13826) );
  sky130_fd_sc_hd__nand2_1 U20494 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[82]), .Y(n13419) );
  sky130_fd_sc_hd__nand2_1 U20495 ( .A(n13412), .B(
        j202_soc_core_j22_cpu_regop_Rm__3_), .Y(n13410) );
  sky130_fd_sc_hd__nor2_1 U20496 ( .A(n13410), .B(n13414), .Y(n13411) );
  sky130_fd_sc_hd__nand2_1 U20497 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[401]), .Y(n13418) );
  sky130_fd_sc_hd__nand2_1 U20498 ( .A(n13413), .B(n13412), .Y(n13415) );
  sky130_fd_sc_hd__nand2_1 U20500 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[146]), .Y(n13417) );
  sky130_fd_sc_hd__nand4_1 U20501 ( .A(n13420), .B(n13419), .C(n13418), .D(
        n13417), .Y(n13421) );
  sky130_fd_sc_hd__nor2_1 U20502 ( .A(n13422), .B(n13421), .Y(n13423) );
  sky130_fd_sc_hd__nand2_1 U20503 ( .A(n13424), .B(n13423), .Y(n22375) );
  sky130_fd_sc_hd__nand2_1 U20504 ( .A(n22375), .B(n16523), .Y(n13442) );
  sky130_fd_sc_hd__nand3_1 U20505 ( .A(n18870), .B(n18869), .C(n13431), .Y(
        n14482) );
  sky130_fd_sc_hd__o21ai_0 U20506 ( .A1(n13427), .A2(n16525), .B1(n16524), .Y(
        n13435) );
  sky130_fd_sc_hd__nor2_1 U20507 ( .A(n18860), .B(n13428), .Y(n18865) );
  sky130_fd_sc_hd__nand2_1 U20508 ( .A(n18865), .B(n13431), .Y(n15886) );
  sky130_fd_sc_hd__nor2_1 U20509 ( .A(n18860), .B(n13430), .Y(n18868) );
  sky130_fd_sc_hd__o22ai_1 U20510 ( .A1(n13433), .A2(n16077), .B1(n13432), 
        .B2(n14477), .Y(n13434) );
  sky130_fd_sc_hd__nor2_1 U20511 ( .A(n13435), .B(n13434), .Y(n13441) );
  sky130_fd_sc_hd__inv_2 U20512 ( .A(n16488), .Y(n16531) );
  sky130_fd_sc_hd__nand2_1 U20513 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[18]), .Y(n13440) );
  sky130_fd_sc_hd__nand2_1 U20514 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[18]), .Y(n13439) );
  sky130_fd_sc_hd__nand2_1 U20515 ( .A(n16533), .B(
        j202_soc_core_j22_cpu_pc[18]), .Y(n13438) );
  sky130_fd_sc_hd__inv_2 U20516 ( .A(n16490), .Y(n16534) );
  sky130_fd_sc_hd__nand2_1 U20517 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[18]), .Y(n13437) );
  sky130_fd_sc_hd__nand2_1 U20518 ( .A(n21924), .B(n28519), .Y(n17083) );
  sky130_fd_sc_hd__nand3_1 U20519 ( .A(n13365), .B(
        j202_soc_core_j22_cpu_memop_Ma__0_), .C(n13443), .Y(n13444) );
  sky130_fd_sc_hd__nand2_1 U20521 ( .A(n13481), .B(n13455), .Y(n23809) );
  sky130_fd_sc_hd__nor2_1 U20522 ( .A(n13294), .B(n23809), .Y(n13445) );
  sky130_fd_sc_hd__inv_2 U20523 ( .A(n13445), .Y(n14033) );
  sky130_fd_sc_hd__nand2_1 U20524 ( .A(n16425), .B(
        j202_soc_core_j22_cpu_rf_gpr[146]), .Y(n13454) );
  sky130_fd_sc_hd__nor2_1 U20525 ( .A(n12036), .B(n12031), .Y(n13468) );
  sky130_fd_sc_hd__nand2_1 U20526 ( .A(n13468), .B(n13483), .Y(n23766) );
  sky130_fd_sc_hd__nor2_1 U20527 ( .A(n13294), .B(n23766), .Y(n13446) );
  sky130_fd_sc_hd__nand2_1 U20529 ( .A(n15796), .B(
        j202_soc_core_j22_cpu_rf_gpr[82]), .Y(n13453) );
  sky130_fd_sc_hd__nand2_1 U20530 ( .A(n13447), .B(n13455), .Y(n23819) );
  sky130_fd_sc_hd__nor2_1 U20531 ( .A(n13294), .B(n23819), .Y(n13448) );
  sky130_fd_sc_hd__nand2_1 U20532 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[401]), .Y(n13452) );
  sky130_fd_sc_hd__nor2_1 U20533 ( .A(n12032), .B(n12035), .Y(n13465) );
  sky130_fd_sc_hd__nand2_1 U20534 ( .A(n13465), .B(n13449), .Y(n23777) );
  sky130_fd_sc_hd__nor2_1 U20535 ( .A(n13294), .B(n23777), .Y(n13450) );
  sky130_fd_sc_hd__nand2_1 U20536 ( .A(n11196), .B(
        j202_soc_core_j22_cpu_rf_gpr[369]), .Y(n13451) );
  sky130_fd_sc_hd__nand4_1 U20537 ( .A(n13454), .B(n13453), .C(n13452), .D(
        n13451), .Y(n13463) );
  sky130_fd_sc_hd__nand2_1 U20538 ( .A(n13465), .B(n13455), .Y(n23814) );
  sky130_fd_sc_hd__nor2_1 U20539 ( .A(n13294), .B(n23814), .Y(n13456) );
  sky130_fd_sc_hd__nand2_1 U20540 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[274]), .Y(n13461) );
  sky130_fd_sc_hd__nor2_1 U20541 ( .A(n12030), .B(n12037), .Y(n13484) );
  sky130_fd_sc_hd__nand2_1 U20542 ( .A(n13465), .B(n13484), .Y(n23782) );
  sky130_fd_sc_hd__nor2_1 U20543 ( .A(n13294), .B(n23782), .Y(n13457) );
  sky130_fd_sc_hd__nand2_1 U20544 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[306]), .Y(n13460) );
  sky130_fd_sc_hd__nand2_1 U20545 ( .A(n13468), .B(n13447), .Y(n23788) );
  sky130_fd_sc_hd__nand2_1 U20546 ( .A(n15788), .B(
        j202_soc_core_j22_cpu_rf_gpr[465]), .Y(n13459) );
  sky130_fd_sc_hd__nand2_1 U20547 ( .A(n13484), .B(n13447), .Y(n23824) );
  sky130_fd_sc_hd__nor2_1 U20548 ( .A(n13294), .B(n23824), .Y(n13526) );
  sky130_fd_sc_hd__nand2_1 U20549 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[433]), .Y(n13458) );
  sky130_fd_sc_hd__nand4_1 U20550 ( .A(n13461), .B(n13460), .C(n13459), .D(
        n13458), .Y(n13462) );
  sky130_fd_sc_hd__nor2_1 U20551 ( .A(n13463), .B(n13462), .Y(n13493) );
  sky130_fd_sc_hd__nand2_1 U20552 ( .A(n13468), .B(n13465), .Y(n23797) );
  sky130_fd_sc_hd__nor2_1 U20553 ( .A(n13294), .B(n23797), .Y(n13466) );
  sky130_fd_sc_hd__inv_2 U20554 ( .A(n13466), .Y(n14082) );
  sky130_fd_sc_hd__nand2_1 U20555 ( .A(n16432), .B(
        j202_soc_core_j22_cpu_rf_gpr[337]), .Y(n13473) );
  sky130_fd_sc_hd__nand2_1 U20556 ( .A(n13481), .B(n13484), .Y(n23803) );
  sky130_fd_sc_hd__nor2_1 U20557 ( .A(n13294), .B(n23803), .Y(n13538) );
  sky130_fd_sc_hd__nand2_1 U20558 ( .A(n16410), .B(
        j202_soc_core_j22_cpu_rf_gpr[178]), .Y(n13472) );
  sky130_fd_sc_hd__nand2_1 U20559 ( .A(n13449), .B(n13483), .Y(n23761) );
  sky130_fd_sc_hd__nor2_1 U20560 ( .A(n13294), .B(n23761), .Y(n13467) );
  sky130_fd_sc_hd__nand2_1 U20561 ( .A(n14993), .B(
        j202_soc_core_j22_cpu_rf_gpr[114]), .Y(n13471) );
  sky130_fd_sc_hd__nand2_1 U20562 ( .A(n13481), .B(n13468), .Y(n23793) );
  sky130_fd_sc_hd__nor2_1 U20563 ( .A(n13294), .B(n23793), .Y(n13469) );
  sky130_fd_sc_hd__inv_2 U20564 ( .A(n13469), .Y(n13951) );
  sky130_fd_sc_hd__nand2_1 U20565 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[210]), .Y(n13470) );
  sky130_fd_sc_hd__nand2_1 U20566 ( .A(n13474), .B(n13477), .Y(n13475) );
  sky130_fd_sc_hd__nand2_1 U20567 ( .A(n13475), .B(
        j202_soc_core_j22_cpu_regop_Ra__0_), .Y(n13537) );
  sky130_fd_sc_hd__nor2_1 U20568 ( .A(n13476), .B(n14798), .Y(n13491) );
  sky130_fd_sc_hd__a21oi_1 U20569 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[18]), .B1(n14743), .Y(n13489) );
  sky130_fd_sc_hd__nand2_1 U20570 ( .A(n13481), .B(n13449), .Y(n23756) );
  sky130_fd_sc_hd__nor2_1 U20571 ( .A(n13294), .B(n23756), .Y(n13482) );
  sky130_fd_sc_hd__nand2_1 U20572 ( .A(n16043), .B(
        j202_soc_core_j22_cpu_rf_gpr[242]), .Y(n13488) );
  sky130_fd_sc_hd__nand2_1 U20573 ( .A(n13447), .B(n13449), .Y(n23843) );
  sky130_fd_sc_hd__nor2_1 U20574 ( .A(n13294), .B(n23843), .Y(n13546) );
  sky130_fd_sc_hd__nand2_1 U20575 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[497]), .Y(n13487) );
  sky130_fd_sc_hd__nand2_1 U20576 ( .A(n13484), .B(n13483), .Y(n23771) );
  sky130_fd_sc_hd__nor2_1 U20577 ( .A(n13294), .B(n23771), .Y(n13485) );
  sky130_fd_sc_hd__inv_2 U20578 ( .A(n13485), .Y(n13952) );
  sky130_fd_sc_hd__nand2_1 U20579 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[50]), .Y(n13486) );
  sky130_fd_sc_hd__nand4_1 U20580 ( .A(n13489), .B(n13488), .C(n13487), .D(
        n13486), .Y(n13490) );
  sky130_fd_sc_hd__nor2_1 U20581 ( .A(n13491), .B(n13490), .Y(n13492) );
  sky130_fd_sc_hd__nand2_1 U20582 ( .A(n21925), .B(n27115), .Y(n17082) );
  sky130_fd_sc_hd__and3_1 U20583 ( .A(n17084), .B(n17083), .C(n17082), .X(
        n14590) );
  sky130_fd_sc_hd__nor2_1 U20584 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[0]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[4]), .Y(n18826) );
  sky130_fd_sc_hd__o22ai_1 U20585 ( .A1(n21709), .A2(n26374), .B1(n26270), 
        .B2(n18826), .Y(n13495) );
  sky130_fd_sc_hd__nand2_1 U20586 ( .A(n26142), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[3]), .Y(n26266) );
  sky130_fd_sc_hd__nand2_1 U20587 ( .A(n26205), .B(n26295), .Y(n13494) );
  sky130_fd_sc_hd__nand3b_1 U20588 ( .A_N(n26149), .B(n26142), .C(n13494), .Y(
        n13790) );
  sky130_fd_sc_hd__nor2_1 U20589 ( .A(n13495), .B(n13790), .Y(n13555) );
  sky130_fd_sc_hd__and3_1 U20590 ( .A(n26142), .B(n18809), .C(
        j202_soc_core_j22_cpu_exuop_EXU_[0]), .X(n13498) );
  sky130_fd_sc_hd__nand3_1 U20591 ( .A(n26374), .B(n28104), .C(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n13497) );
  sky130_fd_sc_hd__nand2_1 U20592 ( .A(n26270), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[4]), .Y(n13496) );
  sky130_fd_sc_hd__nand3_1 U20593 ( .A(n13497), .B(n18827), .C(n13496), .Y(
        n13789) );
  sky130_fd_sc_hd__a21oi_1 U20594 ( .A1(n18825), .A2(n13498), .B1(n13789), .Y(
        n13787) );
  sky130_fd_sc_hd__nand2_1 U20595 ( .A(n18809), .B(n21709), .Y(n26341) );
  sky130_fd_sc_hd__nand2_1 U20596 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[1]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[0]), .Y(n25802) );
  sky130_fd_sc_hd__nand2_1 U20597 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[1]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[3]), .Y(n13499) );
  sky130_fd_sc_hd__nand3_1 U20598 ( .A(n24910), .B(n25802), .C(n13499), .Y(
        n13585) );
  sky130_fd_sc_hd__nand3_1 U20599 ( .A(n13555), .B(n13787), .C(n13585), .Y(
        n16424) );
  sky130_fd_sc_hd__inv_2 U20600 ( .A(n16424), .Y(n16501) );
  sky130_fd_sc_hd__nand2_1 U20601 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[198]), .Y(n13503) );
  sky130_fd_sc_hd__nand2_1 U20602 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[262]), .Y(n13502) );
  sky130_fd_sc_hd__nand2_1 U20603 ( .A(n14993), .B(
        j202_soc_core_j22_cpu_rf_gpr[102]), .Y(n13501) );
  sky130_fd_sc_hd__nand2_1 U20604 ( .A(n14985), .B(
        j202_soc_core_j22_cpu_rf_gpr[485]), .Y(n13500) );
  sky130_fd_sc_hd__nand4_1 U20605 ( .A(n13503), .B(n13502), .C(n13501), .D(
        n13500), .Y(n13509) );
  sky130_fd_sc_hd__nand2_1 U20606 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[134]), .Y(n13507) );
  sky130_fd_sc_hd__nand2_1 U20607 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[70]), .Y(n13506) );
  sky130_fd_sc_hd__nand2_1 U20608 ( .A(n11196), .B(
        j202_soc_core_j22_cpu_rf_gpr[357]), .Y(n13505) );
  sky130_fd_sc_hd__nand2_1 U20609 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[421]), .Y(n13504) );
  sky130_fd_sc_hd__nand4_1 U20610 ( .A(n13507), .B(n13506), .C(n13505), .D(
        n13504), .Y(n13508) );
  sky130_fd_sc_hd__nor2_1 U20611 ( .A(n13509), .B(n13508), .Y(n13525) );
  sky130_fd_sc_hd__nand2_1 U20612 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[294]), .Y(n13511) );
  sky130_fd_sc_hd__nand2_1 U20613 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[166]), .Y(n13510) );
  sky130_fd_sc_hd__nand2_1 U20614 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[325]), .Y(n13517) );
  sky130_fd_sc_hd__nand3_1 U20615 ( .A(n13477), .B(n13513), .C(
        j202_soc_core_intr_req_), .Y(n14196) );
  sky130_fd_sc_hd__o22ai_1 U20616 ( .A1(n14196), .A2(n29068), .B1(n13514), 
        .B2(n14312), .Y(n13515) );
  sky130_fd_sc_hd__a21oi_1 U20617 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[6]), .B1(n13515), .Y(n13516) );
  sky130_fd_sc_hd__nand2_1 U20618 ( .A(n13517), .B(n13516), .Y(n13523) );
  sky130_fd_sc_hd__nand2_1 U20619 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[230]), .Y(n13521) );
  sky130_fd_sc_hd__nand2_1 U20620 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[38]), .Y(n13520) );
  sky130_fd_sc_hd__nand2_1 U20621 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[389]), .Y(n13519) );
  sky130_fd_sc_hd__nand2_1 U20622 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[453]), .Y(n13518) );
  sky130_fd_sc_hd__nand4_1 U20623 ( .A(n13521), .B(n13520), .C(n13519), .D(
        n13518), .Y(n13522) );
  sky130_fd_sc_hd__nor2_1 U20624 ( .A(n13523), .B(n13522), .Y(n13524) );
  sky130_fd_sc_hd__nand2_1 U20625 ( .A(n16432), .B(
        j202_soc_core_j22_cpu_rf_gpr[324]), .Y(n13530) );
  sky130_fd_sc_hd__nand2_1 U20626 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[37]), .Y(n13529) );
  sky130_fd_sc_hd__nand2_1 U20627 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[388]), .Y(n13528) );
  sky130_fd_sc_hd__nand2_1 U20628 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[420]), .Y(n13527) );
  sky130_fd_sc_hd__nand4_1 U20629 ( .A(n13530), .B(n13529), .C(n13528), .D(
        n13527), .Y(n13536) );
  sky130_fd_sc_hd__nand2_1 U20630 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[356]), .Y(n13534) );
  sky130_fd_sc_hd__nand2_1 U20631 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[261]), .Y(n13533) );
  sky130_fd_sc_hd__nand2_1 U20632 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[229]), .Y(n13532) );
  sky130_fd_sc_hd__nand2_1 U20633 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[452]), .Y(n13531) );
  sky130_fd_sc_hd__nand4_1 U20634 ( .A(n13534), .B(n13533), .C(n13532), .D(
        n13531), .Y(n13535) );
  sky130_fd_sc_hd__nor2_1 U20635 ( .A(n13536), .B(n13535), .Y(n13554) );
  sky130_fd_sc_hd__nand2_1 U20636 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[165]), .Y(n13540) );
  sky130_fd_sc_hd__nand2_1 U20637 ( .A(n14993), .B(
        j202_soc_core_j22_cpu_rf_gpr[101]), .Y(n13539) );
  sky130_fd_sc_hd__nand2_1 U20638 ( .A(n16433), .B(
        j202_soc_core_j22_cpu_rf_gpr[197]), .Y(n13545) );
  sky130_fd_sc_hd__o22ai_1 U20639 ( .A1(n14196), .A2(n29071), .B1(n13542), 
        .B2(n14312), .Y(n13543) );
  sky130_fd_sc_hd__a21oi_1 U20640 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[5]), .B1(n13543), .Y(n13544) );
  sky130_fd_sc_hd__nand2_1 U20641 ( .A(n13545), .B(n13544), .Y(n13552) );
  sky130_fd_sc_hd__nand2_1 U20642 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[293]), .Y(n13550) );
  sky130_fd_sc_hd__nand2_1 U20643 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[69]), .Y(n13549) );
  sky130_fd_sc_hd__nand2_1 U20644 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[484]), .Y(n13548) );
  sky130_fd_sc_hd__nand2_1 U20645 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[133]), .Y(n13547) );
  sky130_fd_sc_hd__nand4_1 U20646 ( .A(n13550), .B(n13549), .C(n13548), .D(
        n13547), .Y(n13551) );
  sky130_fd_sc_hd__nor2_1 U20647 ( .A(n13552), .B(n13551), .Y(n13553) );
  sky130_fd_sc_hd__nor2_1 U20648 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .B(n26270), .Y(n16457) );
  sky130_fd_sc_hd__o22ai_1 U20649 ( .A1(n16501), .A2(n11191), .B1(n11189), 
        .B2(n16500), .Y(n13933) );
  sky130_fd_sc_hd__xnor2_1 U20650 ( .A(j202_soc_core_j22_cpu_rfuo_sr__q_), .B(
        j202_soc_core_j22_cpu_rfuo_sr__m_), .Y(n13586) );
  sky130_fd_sc_hd__nand2_1 U20651 ( .A(n13586), .B(n16457), .Y(n13792) );
  sky130_fd_sc_hd__nand2_1 U20652 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[198]), .Y(n13559) );
  sky130_fd_sc_hd__nand2_1 U20653 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[453]), .Y(n13558) );
  sky130_fd_sc_hd__nand2_1 U20654 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[485]), .Y(n13557) );
  sky130_fd_sc_hd__inv_2 U20655 ( .A(n13616), .Y(n16461) );
  sky130_fd_sc_hd__nand2_1 U20656 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[230]), .Y(n13556) );
  sky130_fd_sc_hd__nand4_1 U20657 ( .A(n13559), .B(n13558), .C(n13557), .D(
        n13556), .Y(n13565) );
  sky130_fd_sc_hd__nand2_1 U20658 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[6]), .Y(n13563) );
  sky130_fd_sc_hd__nand2_1 U20659 ( .A(n15984), .B(
        j202_soc_core_j22_cpu_rf_gpr[70]), .Y(n13562) );
  sky130_fd_sc_hd__nand2_1 U20660 ( .A(n16466), .B(
        j202_soc_core_j22_cpu_rf_gpr[389]), .Y(n13561) );
  sky130_fd_sc_hd__nand2_1 U20661 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[134]), .Y(n13560) );
  sky130_fd_sc_hd__nand4_1 U20662 ( .A(n13563), .B(n13562), .C(n13561), .D(
        n13560), .Y(n13564) );
  sky130_fd_sc_hd__nor2_1 U20663 ( .A(n13565), .B(n13564), .Y(n13574) );
  sky130_fd_sc_hd__a22oi_1 U20664 ( .A1(n23776), .A2(
        j202_soc_core_j22_cpu_rf_gpr[357]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[262]), .Y(n13573) );
  sky130_fd_sc_hd__a22oi_1 U20666 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[38]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_rf_gpr[325]), .Y(n13572) );
  sky130_fd_sc_hd__nand2_1 U20667 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[294]), .Y(n13570) );
  sky130_fd_sc_hd__nand2_1 U20668 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[421]), .Y(n13569) );
  sky130_fd_sc_hd__nand2_1 U20669 ( .A(n11199), .B(
        j202_soc_core_j22_cpu_rf_gpr[166]), .Y(n13568) );
  sky130_fd_sc_hd__nand4_1 U20672 ( .A(n13574), .B(n13573), .C(n13572), .D(
        n13571), .Y(n22161) );
  sky130_fd_sc_hd__o22ai_1 U20673 ( .A1(n22155), .A2(n15886), .B1(n22154), 
        .B2(n14373), .Y(n13578) );
  sky130_fd_sc_hd__o22ai_1 U20674 ( .A1(n13576), .A2(n16487), .B1(n14342), 
        .B2(n13575), .Y(n13577) );
  sky130_fd_sc_hd__nor2_1 U20675 ( .A(n13578), .B(n13577), .Y(n13583) );
  sky130_fd_sc_hd__nand2_1 U20676 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[6]), .Y(n13582) );
  sky130_fd_sc_hd__nand2_1 U20677 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[6]), .Y(n13581) );
  sky130_fd_sc_hd__a2bb2oi_1 U20678 ( .B1(n14378), .B2(
        j202_soc_core_j22_cpu_regop_imm__6_), .A1_N(n22151), .A2_N(n16525), 
        .Y(n13580) );
  sky130_fd_sc_hd__nand2_1 U20679 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[6]), .Y(n13579) );
  sky130_fd_sc_hd__o21a_1 U20680 ( .A1(n13587), .A2(n13586), .B1(n13585), .X(
        n13860) );
  sky130_fd_sc_hd__nand2_1 U20681 ( .A(n28495), .B(n16541), .Y(n13588) );
  sky130_fd_sc_hd__nor2_1 U20683 ( .A(n13933), .B(n13934), .Y(n21325) );
  sky130_fd_sc_hd__nand2_1 U20684 ( .A(n16410), .B(
        j202_soc_core_j22_cpu_rf_gpr[164]), .Y(n13592) );
  sky130_fd_sc_hd__nand2_1 U20685 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[419]), .Y(n13591) );
  sky130_fd_sc_hd__nand2_1 U20686 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[387]), .Y(n13590) );
  sky130_fd_sc_hd__nand2_1 U20687 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[483]), .Y(n13589) );
  sky130_fd_sc_hd__nand4_1 U20688 ( .A(n13592), .B(n13591), .C(n13590), .D(
        n13589), .Y(n13598) );
  sky130_fd_sc_hd__nand2_1 U20689 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[292]), .Y(n13596) );
  sky130_fd_sc_hd__nand2_1 U20690 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[323]), .Y(n13595) );
  sky130_fd_sc_hd__nand2_1 U20691 ( .A(n15796), .B(
        j202_soc_core_j22_cpu_rf_gpr[68]), .Y(n13594) );
  sky130_fd_sc_hd__nand2_1 U20692 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[260]), .Y(n13593) );
  sky130_fd_sc_hd__nand4_1 U20693 ( .A(n13596), .B(n13595), .C(n13594), .D(
        n13593), .Y(n13597) );
  sky130_fd_sc_hd__nor2_1 U20694 ( .A(n13598), .B(n13597), .Y(n13615) );
  sky130_fd_sc_hd__nand2_1 U20695 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[196]), .Y(n13602) );
  sky130_fd_sc_hd__o22ai_1 U20696 ( .A1(n14196), .A2(n24787), .B1(n13599), 
        .B2(n14312), .Y(n13600) );
  sky130_fd_sc_hd__a21oi_1 U20697 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[4]), .B1(n13600), .Y(n13601) );
  sky130_fd_sc_hd__nand2_1 U20698 ( .A(n13602), .B(n13601), .Y(n13608) );
  sky130_fd_sc_hd__nand2_1 U20699 ( .A(n16043), .B(
        j202_soc_core_j22_cpu_rf_gpr[228]), .Y(n13606) );
  sky130_fd_sc_hd__nand2_1 U20700 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[36]), .Y(n13605) );
  sky130_fd_sc_hd__nand2_1 U20701 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[132]), .Y(n13604) );
  sky130_fd_sc_hd__nand2_1 U20702 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[355]), .Y(n13603) );
  sky130_fd_sc_hd__nand4_1 U20703 ( .A(n13606), .B(n13605), .C(n13604), .D(
        n13603), .Y(n13607) );
  sky130_fd_sc_hd__nor2_1 U20704 ( .A(n13608), .B(n13607), .Y(n13614) );
  sky130_fd_sc_hd__nand2b_1 U20705 ( .A_N(n16444), .B(
        j202_soc_core_j22_cpu_rf_gpr[4]), .Y(n13611) );
  sky130_fd_sc_hd__nand2_1 U20706 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[451]), .Y(n13610) );
  sky130_fd_sc_hd__nand2_1 U20707 ( .A(n15783), .B(
        j202_soc_core_j22_cpu_rf_gpr[100]), .Y(n13609) );
  sky130_fd_sc_hd__nand3_1 U20708 ( .A(n13611), .B(n13610), .C(n13609), .Y(
        n13612) );
  sky130_fd_sc_hd__nand3_1 U20709 ( .A(n13615), .B(n13614), .C(n13613), .Y(
        n22136) );
  sky130_fd_sc_hd__inv_2 U20710 ( .A(n22136), .Y(n27365) );
  sky130_fd_sc_hd__o22ai_1 U20711 ( .A1(n16500), .A2(n27365), .B1(n11189), 
        .B2(n16501), .Y(n13931) );
  sky130_fd_sc_hd__nand2_1 U20712 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[197]), .Y(n13620) );
  sky130_fd_sc_hd__nand2_1 U20713 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[452]), .Y(n13619) );
  sky130_fd_sc_hd__nand2_1 U20714 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[484]), .Y(n13618) );
  sky130_fd_sc_hd__nand2_1 U20715 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[229]), .Y(n13617) );
  sky130_fd_sc_hd__nand4_1 U20716 ( .A(n13620), .B(n13619), .C(n13618), .D(
        n13617), .Y(n13626) );
  sky130_fd_sc_hd__nand2_1 U20717 ( .A(n16506), .B(
        j202_soc_core_j22_cpu_rf_gpr[5]), .Y(n13624) );
  sky130_fd_sc_hd__nand2_1 U20718 ( .A(n15984), .B(
        j202_soc_core_j22_cpu_rf_gpr[69]), .Y(n13623) );
  sky130_fd_sc_hd__nand2_1 U20719 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[388]), .Y(n13622) );
  sky130_fd_sc_hd__nand2_1 U20720 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[133]), .Y(n13621) );
  sky130_fd_sc_hd__nand4_1 U20721 ( .A(n13624), .B(n13623), .C(n13622), .D(
        n13621), .Y(n13625) );
  sky130_fd_sc_hd__nor2_1 U20722 ( .A(n13626), .B(n13625), .Y(n13638) );
  sky130_fd_sc_hd__nand2_1 U20723 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[261]), .Y(n13630) );
  sky130_fd_sc_hd__nand2_1 U20724 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[37]), .Y(n13629) );
  sky130_fd_sc_hd__nand2_1 U20725 ( .A(n15991), .B(
        j202_soc_core_j22_cpu_rf_gpr[356]), .Y(n13628) );
  sky130_fd_sc_hd__nand2_1 U20726 ( .A(n15017), .B(
        j202_soc_core_j22_cpu_rf_gpr[324]), .Y(n13627) );
  sky130_fd_sc_hd__and4_1 U20727 ( .A(n13630), .B(n13629), .C(n13628), .D(
        n13627), .X(n13637) );
  sky130_fd_sc_hd__nand2_1 U20728 ( .A(n15958), .B(
        j202_soc_core_j22_cpu_rf_gpr[293]), .Y(n13635) );
  sky130_fd_sc_hd__nand2_1 U20729 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[420]), .Y(n13634) );
  sky130_fd_sc_hd__nand2_1 U20730 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[165]), .Y(n13633) );
  sky130_fd_sc_hd__nand2_1 U20731 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[101]), .Y(n13632) );
  sky130_fd_sc_hd__and4_1 U20732 ( .A(n13635), .B(n13634), .C(n13633), .D(
        n13632), .X(n13636) );
  sky130_fd_sc_hd__o2bb2ai_1 U20733 ( .B1(n22283), .B2(n16525), .A1_N(n14378), 
        .A2_N(j202_soc_core_j22_cpu_regop_imm__5_), .Y(n13639) );
  sky130_fd_sc_hd__a21oi_1 U20734 ( .A1(n16534), .A2(
        j202_soc_core_j22_cpu_rf_gbr[5]), .B1(n13639), .Y(n13645) );
  sky130_fd_sc_hd__o22a_1 U20735 ( .A1(n22286), .A2(n14342), .B1(n22287), .B2(
        n14373), .X(n13644) );
  sky130_fd_sc_hd__o22a_1 U20736 ( .A1(n22288), .A2(n11202), .B1(n16487), .B2(
        n13640), .X(n13643) );
  sky130_fd_sc_hd__o22a_1 U20737 ( .A1(n13641), .A2(n16488), .B1(n22284), .B2(
        n16491), .X(n13642) );
  sky130_fd_sc_hd__nand4_1 U20738 ( .A(n13645), .B(n13644), .C(n13643), .D(
        n13642), .Y(n13646) );
  sky130_fd_sc_hd__a21oi_4 U20739 ( .A1(n22282), .A2(n16523), .B1(n13646), .Y(
        n26421) );
  sky130_fd_sc_hd__nand2_1 U20740 ( .A(n26421), .B(n16543), .Y(n13647) );
  sky130_fd_sc_hd__o21a_1 U20741 ( .A1(n26421), .A2(n16541), .B1(n13647), .X(
        n13932) );
  sky130_fd_sc_hd__nor2_1 U20742 ( .A(n21325), .B(n21663), .Y(n13936) );
  sky130_fd_sc_hd__nand2_1 U20743 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[35]), .Y(n13651) );
  sky130_fd_sc_hd__nand2_1 U20744 ( .A(n16425), .B(
        j202_soc_core_j22_cpu_rf_gpr[131]), .Y(n13650) );
  sky130_fd_sc_hd__nand2_1 U20745 ( .A(n11195), .B(
        j202_soc_core_j22_cpu_rf_gpr[386]), .Y(n13649) );
  sky130_fd_sc_hd__nand2_1 U20746 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[67]), .Y(n13648) );
  sky130_fd_sc_hd__nand4_1 U20747 ( .A(n13651), .B(n13650), .C(n13649), .D(
        n13648), .Y(n13657) );
  sky130_fd_sc_hd__nand2_1 U20748 ( .A(n16432), .B(
        j202_soc_core_j22_cpu_rf_gpr[322]), .Y(n13655) );
  sky130_fd_sc_hd__nand2_1 U20749 ( .A(n16410), .B(
        j202_soc_core_j22_cpu_rf_gpr[163]), .Y(n13654) );
  sky130_fd_sc_hd__nand2_1 U20750 ( .A(n15783), .B(
        j202_soc_core_j22_cpu_rf_gpr[99]), .Y(n13653) );
  sky130_fd_sc_hd__nand2_1 U20751 ( .A(n16433), .B(
        j202_soc_core_j22_cpu_rf_gpr[195]), .Y(n13652) );
  sky130_fd_sc_hd__nand4_1 U20752 ( .A(n13655), .B(n13654), .C(n13653), .D(
        n13652), .Y(n13656) );
  sky130_fd_sc_hd__nor2_1 U20753 ( .A(n13657), .B(n13656), .Y(n13672) );
  sky130_fd_sc_hd__nand2_1 U20754 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[291]), .Y(n13659) );
  sky130_fd_sc_hd__nand2_1 U20755 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[418]), .Y(n13658) );
  sky130_fd_sc_hd__nand2_1 U20756 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[450]), .Y(n13664) );
  sky130_fd_sc_hd__o22ai_1 U20757 ( .A1(n28366), .A2(n14196), .B1(n30017), 
        .B2(n14312), .Y(n13662) );
  sky130_fd_sc_hd__a21oi_1 U20758 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[3]), .B1(n13662), .Y(n13663) );
  sky130_fd_sc_hd__nand2_1 U20759 ( .A(n13664), .B(n13663), .Y(n13670) );
  sky130_fd_sc_hd__nand2_1 U20760 ( .A(n16043), .B(
        j202_soc_core_j22_cpu_rf_gpr[227]), .Y(n13668) );
  sky130_fd_sc_hd__nand2_1 U20761 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[259]), .Y(n13667) );
  sky130_fd_sc_hd__nand2_1 U20762 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[482]), .Y(n13666) );
  sky130_fd_sc_hd__nand2_1 U20763 ( .A(n11196), .B(
        j202_soc_core_j22_cpu_rf_gpr[354]), .Y(n13665) );
  sky130_fd_sc_hd__nand4_1 U20764 ( .A(n13668), .B(n13667), .C(n13666), .D(
        n13665), .Y(n13669) );
  sky130_fd_sc_hd__nor2_1 U20765 ( .A(n13670), .B(n13669), .Y(n13671) );
  sky130_fd_sc_hd__nand3_1 U20766 ( .A(n13672), .B(n13061), .C(n13671), .Y(
        n26334) );
  sky130_fd_sc_hd__nand2_1 U20767 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[290]), .Y(n13676) );
  sky130_fd_sc_hd__nand2_1 U20768 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[66]), .Y(n13675) );
  sky130_fd_sc_hd__nand2_1 U20769 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[385]), .Y(n13674) );
  sky130_fd_sc_hd__nand2_1 U20770 ( .A(n11196), .B(
        j202_soc_core_j22_cpu_rf_gpr[353]), .Y(n13673) );
  sky130_fd_sc_hd__nand4_1 U20771 ( .A(n13676), .B(n13675), .C(n13674), .D(
        n13673), .Y(n13682) );
  sky130_fd_sc_hd__nand2_1 U20772 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[258]), .Y(n13680) );
  sky130_fd_sc_hd__nand2_1 U20773 ( .A(n16432), .B(
        j202_soc_core_j22_cpu_rf_gpr[321]), .Y(n13679) );
  sky130_fd_sc_hd__nand2_1 U20774 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[449]), .Y(n13678) );
  sky130_fd_sc_hd__nand2_1 U20775 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[417]), .Y(n13677) );
  sky130_fd_sc_hd__nand4_1 U20776 ( .A(n13680), .B(n13679), .C(n13678), .D(
        n13677), .Y(n13681) );
  sky130_fd_sc_hd__nor2_1 U20777 ( .A(n13682), .B(n13681), .Y(n13696) );
  sky130_fd_sc_hd__nand2_1 U20778 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[162]), .Y(n13684) );
  sky130_fd_sc_hd__nand2_1 U20779 ( .A(n15783), .B(
        j202_soc_core_j22_cpu_rf_gpr[98]), .Y(n13683) );
  sky130_fd_sc_hd__nand2_1 U20780 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[194]), .Y(n13688) );
  sky130_fd_sc_hd__o22ai_1 U20781 ( .A1(n14196), .A2(n27348), .B1(n30018), 
        .B2(n14312), .Y(n13686) );
  sky130_fd_sc_hd__a21oi_1 U20782 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[2]), .B1(n13686), .Y(n13687) );
  sky130_fd_sc_hd__nand2_1 U20783 ( .A(n13688), .B(n13687), .Y(n13694) );
  sky130_fd_sc_hd__nand2_1 U20784 ( .A(n16425), .B(
        j202_soc_core_j22_cpu_rf_gpr[130]), .Y(n13692) );
  sky130_fd_sc_hd__nand2_1 U20785 ( .A(n16043), .B(
        j202_soc_core_j22_cpu_rf_gpr[226]), .Y(n13691) );
  sky130_fd_sc_hd__nand2_1 U20786 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[481]), .Y(n13690) );
  sky130_fd_sc_hd__nand2_1 U20787 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[34]), .Y(n13689) );
  sky130_fd_sc_hd__nand4_1 U20788 ( .A(n13692), .B(n13691), .C(n13690), .D(
        n13689), .Y(n13693) );
  sky130_fd_sc_hd__nor2_1 U20789 ( .A(n13694), .B(n13693), .Y(n13695) );
  sky130_fd_sc_hd__inv_2 U20790 ( .A(n26929), .Y(n27147) );
  sky130_fd_sc_hd__o22ai_1 U20791 ( .A1(n16501), .A2(n11190), .B1(n27147), 
        .B2(n16500), .Y(n13927) );
  sky130_fd_sc_hd__nand2_1 U20792 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[195]), .Y(n13700) );
  sky130_fd_sc_hd__nand2_1 U20793 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[450]), .Y(n13699) );
  sky130_fd_sc_hd__nand2_1 U20794 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[482]), .Y(n13698) );
  sky130_fd_sc_hd__nand2_1 U20795 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[227]), .Y(n13697) );
  sky130_fd_sc_hd__nand4_1 U20796 ( .A(n13700), .B(n13699), .C(n13698), .D(
        n13697), .Y(n13706) );
  sky130_fd_sc_hd__nand2_1 U20797 ( .A(n16506), .B(
        j202_soc_core_j22_cpu_rf_gpr[3]), .Y(n13704) );
  sky130_fd_sc_hd__nand2_1 U20798 ( .A(n15984), .B(
        j202_soc_core_j22_cpu_rf_gpr[67]), .Y(n13703) );
  sky130_fd_sc_hd__nand2_1 U20799 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[386]), .Y(n13702) );
  sky130_fd_sc_hd__inv_2 U20800 ( .A(n30190), .Y(n23808) );
  sky130_fd_sc_hd__nand2_1 U20801 ( .A(n23808), .B(
        j202_soc_core_j22_cpu_rf_gpr[131]), .Y(n13701) );
  sky130_fd_sc_hd__nand4_1 U20802 ( .A(n13704), .B(n13703), .C(n13702), .D(
        n13701), .Y(n13705) );
  sky130_fd_sc_hd__nor2_1 U20803 ( .A(n13706), .B(n13705), .Y(n13715) );
  sky130_fd_sc_hd__a22oi_1 U20804 ( .A1(n23776), .A2(
        j202_soc_core_j22_cpu_rf_gpr[354]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[259]), .Y(n13714) );
  sky130_fd_sc_hd__a22oi_1 U20805 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[35]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_rf_gpr[322]), .Y(n13713) );
  sky130_fd_sc_hd__nand2_1 U20806 ( .A(n15958), .B(
        j202_soc_core_j22_cpu_rf_gpr[291]), .Y(n13711) );
  sky130_fd_sc_hd__nand2_1 U20807 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[418]), .Y(n13710) );
  sky130_fd_sc_hd__nand2_1 U20808 ( .A(n11199), .B(
        j202_soc_core_j22_cpu_rf_gpr[163]), .Y(n13709) );
  sky130_fd_sc_hd__nand2_1 U20809 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[99]), .Y(n13708) );
  sky130_fd_sc_hd__and4_1 U20810 ( .A(n13711), .B(n13710), .C(n13709), .D(
        n13708), .X(n13712) );
  sky130_fd_sc_hd__nand4_1 U20811 ( .A(n13715), .B(n13714), .C(n13713), .D(
        n13712), .Y(n21242) );
  sky130_fd_sc_hd__o22ai_1 U20812 ( .A1(n21249), .A2(n16077), .B1(n21248), 
        .B2(n14342), .Y(n13716) );
  sky130_fd_sc_hd__nor2_1 U20813 ( .A(n13717), .B(n13716), .Y(n13722) );
  sky130_fd_sc_hd__nand2_1 U20814 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[3]), .Y(n13721) );
  sky130_fd_sc_hd__nand2_1 U20815 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[3]), .Y(n13720) );
  sky130_fd_sc_hd__nand2_1 U20816 ( .A(n16533), .B(j202_soc_core_j22_cpu_pc[3]), .Y(n13719) );
  sky130_fd_sc_hd__nand2_1 U20817 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[3]), .Y(n13718) );
  sky130_fd_sc_hd__nand2_1 U20818 ( .A(n28515), .B(n16541), .Y(n13724) );
  sky130_fd_sc_hd__o21ai_1 U20819 ( .A1(n16543), .A2(n28515), .B1(n13724), .Y(
        n13928) );
  sky130_fd_sc_hd__nor2_1 U20820 ( .A(n13927), .B(n13928), .Y(n20442) );
  sky130_fd_sc_hd__o22ai_1 U20821 ( .A1(n16501), .A2(n27365), .B1(n11190), 
        .B2(n16500), .Y(n13929) );
  sky130_fd_sc_hd__nand2_1 U20822 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[196]), .Y(n13731) );
  sky130_fd_sc_hd__nand2_1 U20823 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[451]), .Y(n13730) );
  sky130_fd_sc_hd__nand2_1 U20824 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[483]), .Y(n13729) );
  sky130_fd_sc_hd__nand2_1 U20825 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[228]), .Y(n13728) );
  sky130_fd_sc_hd__nand4_1 U20826 ( .A(n13731), .B(n13730), .C(n13729), .D(
        n13728), .Y(n13737) );
  sky130_fd_sc_hd__nand2_1 U20827 ( .A(n16506), .B(
        j202_soc_core_j22_cpu_rf_gpr[4]), .Y(n13735) );
  sky130_fd_sc_hd__nand2_1 U20828 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[68]), .Y(n13734) );
  sky130_fd_sc_hd__nand2_1 U20829 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[387]), .Y(n13733) );
  sky130_fd_sc_hd__nand2_1 U20830 ( .A(n23808), .B(
        j202_soc_core_j22_cpu_rf_gpr[132]), .Y(n13732) );
  sky130_fd_sc_hd__nand4_1 U20831 ( .A(n13735), .B(n13734), .C(n13733), .D(
        n13732), .Y(n13736) );
  sky130_fd_sc_hd__nor2_1 U20832 ( .A(n13737), .B(n13736), .Y(n13748) );
  sky130_fd_sc_hd__nand2_1 U20833 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[260]), .Y(n13741) );
  sky130_fd_sc_hd__nand2_1 U20834 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[36]), .Y(n13740) );
  sky130_fd_sc_hd__nand2_1 U20835 ( .A(n15991), .B(
        j202_soc_core_j22_cpu_rf_gpr[355]), .Y(n13739) );
  sky130_fd_sc_hd__nand2_1 U20836 ( .A(n15017), .B(
        j202_soc_core_j22_cpu_rf_gpr[323]), .Y(n13738) );
  sky130_fd_sc_hd__and4_1 U20837 ( .A(n13741), .B(n13740), .C(n13739), .D(
        n13738), .X(n13747) );
  sky130_fd_sc_hd__nand2_1 U20838 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[292]), .Y(n13745) );
  sky130_fd_sc_hd__nand2_1 U20839 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[419]), .Y(n13744) );
  sky130_fd_sc_hd__nand2_1 U20840 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[164]), .Y(n13743) );
  sky130_fd_sc_hd__nand2_1 U20841 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[100]), .Y(n13742) );
  sky130_fd_sc_hd__and4_1 U20842 ( .A(n13745), .B(n13744), .C(n13743), .D(
        n13742), .X(n13746) );
  sky130_fd_sc_hd__nand3_1 U20843 ( .A(n13748), .B(n13747), .C(n13746), .Y(
        n21797) );
  sky130_fd_sc_hd__o2bb2ai_1 U20844 ( .B1(n21798), .B2(n16525), .A1_N(n14378), 
        .A2_N(j202_soc_core_j22_cpu_regop_imm__4_), .Y(n13749) );
  sky130_fd_sc_hd__a21oi_1 U20845 ( .A1(n16534), .A2(
        j202_soc_core_j22_cpu_rf_gbr[4]), .B1(n13749), .Y(n13755) );
  sky130_fd_sc_hd__o22a_1 U20846 ( .A1(n21800), .A2(n14477), .B1(n21801), .B2(
        n14373), .X(n13754) );
  sky130_fd_sc_hd__o22a_1 U20847 ( .A1(n21802), .A2(n16077), .B1(n16487), .B2(
        n13750), .X(n13753) );
  sky130_fd_sc_hd__o22a_1 U20848 ( .A1(n13751), .A2(n16488), .B1(n21799), .B2(
        n16491), .X(n13752) );
  sky130_fd_sc_hd__nand4_1 U20849 ( .A(n13755), .B(n13754), .C(n13753), .D(
        n13752), .Y(n13756) );
  sky130_fd_sc_hd__mux2i_1 U20850 ( .A0(n16088), .A1(n16543), .S(n26240), .Y(
        n13930) );
  sky130_fd_sc_hd__nor2_1 U20851 ( .A(n13929), .B(n13930), .Y(n21789) );
  sky130_fd_sc_hd__nor2_1 U20852 ( .A(n20442), .B(n21789), .Y(n21329) );
  sky130_fd_sc_hd__nand2_1 U20853 ( .A(n13936), .B(n21329), .Y(n13938) );
  sky130_fd_sc_hd__nand2_1 U20854 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[193]), .Y(n13760) );
  sky130_fd_sc_hd__nand2_1 U20855 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[448]), .Y(n13759) );
  sky130_fd_sc_hd__nand2_1 U20856 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[480]), .Y(n13758) );
  sky130_fd_sc_hd__nand2_1 U20857 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[225]), .Y(n13757) );
  sky130_fd_sc_hd__nand4_1 U20858 ( .A(n13760), .B(n13759), .C(n13758), .D(
        n13757), .Y(n13767) );
  sky130_fd_sc_hd__nand2_1 U20859 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[1]), .Y(n13765) );
  sky130_fd_sc_hd__nand2_1 U20860 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[65]), .Y(n13764) );
  sky130_fd_sc_hd__nand2_1 U20861 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[384]), .Y(n13763) );
  sky130_fd_sc_hd__nand2_1 U20862 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[129]), .Y(n13762) );
  sky130_fd_sc_hd__nand4_1 U20863 ( .A(n13765), .B(n13764), .C(n13763), .D(
        n13762), .Y(n13766) );
  sky130_fd_sc_hd__nor2_1 U20864 ( .A(n13767), .B(n13766), .Y(n13776) );
  sky130_fd_sc_hd__a22oi_1 U20865 ( .A1(n23776), .A2(
        j202_soc_core_j22_cpu_rf_gpr[352]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[257]), .Y(n13775) );
  sky130_fd_sc_hd__a22oi_1 U20866 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[33]), .B1(n15017), .B2(
        j202_soc_core_j22_cpu_rf_gpr[320]), .Y(n13774) );
  sky130_fd_sc_hd__nand2_1 U20867 ( .A(n15958), .B(
        j202_soc_core_j22_cpu_rf_gpr[289]), .Y(n13771) );
  sky130_fd_sc_hd__nand2_1 U20868 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[416]), .Y(n13770) );
  sky130_fd_sc_hd__nand2_1 U20869 ( .A(n11199), .B(
        j202_soc_core_j22_cpu_rf_gpr[161]), .Y(n13769) );
  sky130_fd_sc_hd__nand2_1 U20870 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[97]), .Y(n13768) );
  sky130_fd_sc_hd__o22ai_1 U20872 ( .A1(n21987), .A2(n15886), .B1(n24668), 
        .B2(n14373), .Y(n13779) );
  sky130_fd_sc_hd__o22ai_1 U20873 ( .A1(n24792), .A2(n16487), .B1(n14342), 
        .B2(n13777), .Y(n13778) );
  sky130_fd_sc_hd__nor2_1 U20874 ( .A(n13779), .B(n13778), .Y(n13785) );
  sky130_fd_sc_hd__a2bb2oi_1 U20875 ( .B1(n14378), .B2(
        j202_soc_core_j22_cpu_regop_imm__1_), .A1_N(n21984), .A2_N(n16525), 
        .Y(n13780) );
  sky130_fd_sc_hd__o22ai_1 U20877 ( .A1(n13882), .A2(n16488), .B1(n16491), 
        .B2(n21985), .Y(n13782) );
  sky130_fd_sc_hd__nor2_1 U20878 ( .A(n13783), .B(n13782), .Y(n13784) );
  sky130_fd_sc_hd__o21ai_1 U20879 ( .A1(n13789), .A2(n28529), .B1(n13788), .Y(
        n13864) );
  sky130_fd_sc_hd__a21oi_1 U20880 ( .A1(n25802), .A2(
        j202_soc_core_j22_cpu_rfuo_sr__t_), .B1(n21709), .Y(n13791) );
  sky130_fd_sc_hd__a211oi_1 U20881 ( .A1(n26362), .A2(
        j202_soc_core_j22_cpu_rfuo_sr__t_), .B1(n13791), .C1(n13790), .Y(
        n13793) );
  sky130_fd_sc_hd__nand3_1 U20882 ( .A(n13864), .B(n13793), .C(n13792), .Y(
        n21702) );
  sky130_fd_sc_hd__nor2_1 U20883 ( .A(n13794), .B(n14798), .Y(n13802) );
  sky130_fd_sc_hd__nand2_1 U20884 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[128]), .Y(n13800) );
  sky130_fd_sc_hd__nand2_1 U20885 ( .A(n16043), .B(
        j202_soc_core_j22_cpu_rf_gpr[224]), .Y(n13799) );
  sky130_fd_sc_hd__a2bb2oi_1 U20886 ( .B1(j202_soc_core_j22_cpu_rf_tmp[0]), 
        .B2(n13053), .A1_N(n14312), .A2_N(n13795), .Y(n13798) );
  sky130_fd_sc_hd__nand2_1 U20887 ( .A(n14985), .B(
        j202_soc_core_j22_cpu_rf_gpr[479]), .Y(n13797) );
  sky130_fd_sc_hd__nand4_1 U20888 ( .A(n13800), .B(n13799), .C(n13798), .D(
        n13797), .Y(n13801) );
  sky130_fd_sc_hd__nand2_1 U20889 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[32]), .Y(n13806) );
  sky130_fd_sc_hd__nand2_1 U20890 ( .A(n15796), .B(
        j202_soc_core_j22_cpu_rf_gpr[64]), .Y(n13805) );
  sky130_fd_sc_hd__nand2_1 U20891 ( .A(n11195), .B(
        j202_soc_core_j22_cpu_rf_gpr[383]), .Y(n13804) );
  sky130_fd_sc_hd__nand2_1 U20892 ( .A(n11196), .B(
        j202_soc_core_j22_cpu_rf_gpr[351]), .Y(n13803) );
  sky130_fd_sc_hd__nand2_1 U20893 ( .A(n11194), .B(
        j202_soc_core_j22_cpu_rf_gpr[288]), .Y(n13810) );
  sky130_fd_sc_hd__nand2_1 U20894 ( .A(n16410), .B(
        j202_soc_core_j22_cpu_rf_gpr[160]), .Y(n13809) );
  sky130_fd_sc_hd__nand2_1 U20895 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[415]), .Y(n13808) );
  sky130_fd_sc_hd__nand2_1 U20896 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[256]), .Y(n13807) );
  sky130_fd_sc_hd__nand2_1 U20897 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[319]), .Y(n13814) );
  sky130_fd_sc_hd__nand2_1 U20898 ( .A(n16433), .B(
        j202_soc_core_j22_cpu_rf_gpr[192]), .Y(n13813) );
  sky130_fd_sc_hd__nand2_1 U20899 ( .A(n14993), .B(
        j202_soc_core_j22_cpu_rf_gpr[96]), .Y(n13812) );
  sky130_fd_sc_hd__nand2_1 U20900 ( .A(n15788), .B(
        j202_soc_core_j22_cpu_rf_gpr[447]), .Y(n13811) );
  sky130_fd_sc_hd__nand4_1 U20901 ( .A(n13814), .B(n13813), .C(n13812), .D(
        n13811), .Y(n13815) );
  sky130_fd_sc_hd__o22ai_1 U20902 ( .A1(n16500), .A2(n21717), .B1(n16501), 
        .B2(n11188), .Y(n13865) );
  sky130_fd_sc_hd__nand2_1 U20903 ( .A(n13818), .B(
        j202_soc_core_j22_cpu_rf_gpr[192]), .Y(n13825) );
  sky130_fd_sc_hd__nand2_1 U20904 ( .A(n13819), .B(
        j202_soc_core_j22_cpu_rf_gpr[447]), .Y(n13824) );
  sky130_fd_sc_hd__nand2_1 U20905 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[479]), .Y(n13823) );
  sky130_fd_sc_hd__nand2_1 U20906 ( .A(n13821), .B(
        j202_soc_core_j22_cpu_rf_gpr[224]), .Y(n13822) );
  sky130_fd_sc_hd__nand4_1 U20907 ( .A(n13825), .B(n13824), .C(n13823), .D(
        n13822), .Y(n13834) );
  sky130_fd_sc_hd__nand2_1 U20908 ( .A(n16506), .B(
        j202_soc_core_j22_cpu_rf_gpr[0]), .Y(n13832) );
  sky130_fd_sc_hd__nand2_1 U20909 ( .A(n13826), .B(
        j202_soc_core_j22_cpu_rf_gpr[64]), .Y(n13831) );
  sky130_fd_sc_hd__nand2_1 U20910 ( .A(n16466), .B(
        j202_soc_core_j22_cpu_rf_gpr[383]), .Y(n13830) );
  sky130_fd_sc_hd__nand2_1 U20911 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[128]), .Y(n13829) );
  sky130_fd_sc_hd__nand4_1 U20912 ( .A(n13832), .B(n13831), .C(n13830), .D(
        n13829), .Y(n13833) );
  sky130_fd_sc_hd__nor2_1 U20913 ( .A(n13834), .B(n13833), .Y(n13847) );
  sky130_fd_sc_hd__a22oi_1 U20914 ( .A1(n13836), .A2(
        j202_soc_core_j22_cpu_rf_gpr[351]), .B1(n13835), .B2(
        j202_soc_core_j22_cpu_rf_gpr[256]), .Y(n13846) );
  sky130_fd_sc_hd__a22oi_1 U20915 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[32]), .B1(n13837), .B2(
        j202_soc_core_j22_cpu_rf_gpr[319]), .Y(n13845) );
  sky130_fd_sc_hd__nand2_1 U20916 ( .A(n13838), .B(
        j202_soc_core_j22_cpu_rf_gpr[288]), .Y(n13844) );
  sky130_fd_sc_hd__nand2_1 U20917 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[415]), .Y(n13843) );
  sky130_fd_sc_hd__nand2_1 U20918 ( .A(n13840), .B(
        j202_soc_core_j22_cpu_rf_gpr[160]), .Y(n13842) );
  sky130_fd_sc_hd__nand2_1 U20919 ( .A(n14525), .B(
        j202_soc_core_j22_cpu_rf_gpr[96]), .Y(n13841) );
  sky130_fd_sc_hd__nand4_1 U20920 ( .A(n13847), .B(n13846), .C(n13845), .D(
        n13089), .Y(n21680) );
  sky130_fd_sc_hd__nand2_1 U20921 ( .A(n21680), .B(n16523), .Y(n13859) );
  sky130_fd_sc_hd__o22ai_1 U20922 ( .A1(n21674), .A2(n11202), .B1(n21717), 
        .B2(n14373), .Y(n13851) );
  sky130_fd_sc_hd__o22ai_1 U20923 ( .A1(n13849), .A2(n16487), .B1(n14342), 
        .B2(n13848), .Y(n13850) );
  sky130_fd_sc_hd__nor2_1 U20924 ( .A(n13851), .B(n13850), .Y(n13858) );
  sky130_fd_sc_hd__nand2_1 U20925 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[0]), .Y(n13855) );
  sky130_fd_sc_hd__nand2_1 U20926 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[0]), .Y(n13854) );
  sky130_fd_sc_hd__nand2_1 U20927 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[0]), .Y(n13852) );
  sky130_fd_sc_hd__nand4_1 U20928 ( .A(n13855), .B(n13854), .C(n13853), .D(
        n13852), .Y(n13856) );
  sky130_fd_sc_hd__nand3_2 U20929 ( .A(n13859), .B(n13858), .C(n13857), .Y(
        n28541) );
  sky130_fd_sc_hd__nand2_1 U20930 ( .A(n28541), .B(n13861), .Y(n13862) );
  sky130_fd_sc_hd__o21a_1 U20931 ( .A1(n16543), .A2(n28541), .B1(n13862), .X(
        n13863) );
  sky130_fd_sc_hd__nand2_1 U20932 ( .A(n13864), .B(n13863), .Y(n13866) );
  sky130_fd_sc_hd__nor2_1 U20933 ( .A(n13865), .B(n13866), .Y(n21698) );
  sky130_fd_sc_hd__nand2_1 U20934 ( .A(n13866), .B(n13865), .Y(n21699) );
  sky130_fd_sc_hd__o21ai_1 U20935 ( .A1(n13867), .A2(n21698), .B1(n21699), .Y(
        n17222) );
  sky130_fd_sc_hd__nand2_1 U20936 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[33]), .Y(n13871) );
  sky130_fd_sc_hd__nand2_1 U20937 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[65]), .Y(n13870) );
  sky130_fd_sc_hd__nand2_1 U20938 ( .A(n15783), .B(
        j202_soc_core_j22_cpu_rf_gpr[97]), .Y(n13869) );
  sky130_fd_sc_hd__nand2_1 U20939 ( .A(n11195), .B(
        j202_soc_core_j22_cpu_rf_gpr[384]), .Y(n13868) );
  sky130_fd_sc_hd__nand4_1 U20940 ( .A(n13871), .B(n13870), .C(n13869), .D(
        n13868), .Y(n13877) );
  sky130_fd_sc_hd__nand2_1 U20941 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[257]), .Y(n13875) );
  sky130_fd_sc_hd__nand2_1 U20942 ( .A(n11194), .B(
        j202_soc_core_j22_cpu_rf_gpr[289]), .Y(n13874) );
  sky130_fd_sc_hd__nand2_1 U20943 ( .A(n15788), .B(
        j202_soc_core_j22_cpu_rf_gpr[448]), .Y(n13873) );
  sky130_fd_sc_hd__nand2_1 U20944 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[129]), .Y(n13872) );
  sky130_fd_sc_hd__nand4_1 U20945 ( .A(n13875), .B(n13874), .C(n13873), .D(
        n13872), .Y(n13876) );
  sky130_fd_sc_hd__nor2_1 U20946 ( .A(n13877), .B(n13876), .Y(n13891) );
  sky130_fd_sc_hd__nand2_1 U20947 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[161]), .Y(n13881) );
  sky130_fd_sc_hd__nand2_1 U20948 ( .A(n16433), .B(
        j202_soc_core_j22_cpu_rf_gpr[193]), .Y(n13880) );
  sky130_fd_sc_hd__nand2_1 U20949 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[416]), .Y(n13879) );
  sky130_fd_sc_hd__nand2_1 U20950 ( .A(n16432), .B(
        j202_soc_core_j22_cpu_rf_gpr[320]), .Y(n13878) );
  sky130_fd_sc_hd__nor2_1 U20951 ( .A(n13882), .B(n14798), .Y(n13889) );
  sky130_fd_sc_hd__nand2_1 U20952 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[352]), .Y(n13887) );
  sky130_fd_sc_hd__nand2_1 U20953 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[225]), .Y(n13886) );
  sky130_fd_sc_hd__a2bb2oi_1 U20954 ( .B1(j202_soc_core_j22_cpu_rf_tmp[1]), 
        .B2(n13053), .A1_N(n14312), .A2_N(n13883), .Y(n13885) );
  sky130_fd_sc_hd__nand2_1 U20955 ( .A(n14985), .B(
        j202_soc_core_j22_cpu_rf_gpr[480]), .Y(n13884) );
  sky130_fd_sc_hd__nand4_1 U20956 ( .A(n13887), .B(n13886), .C(n13885), .D(
        n13884), .Y(n13888) );
  sky130_fd_sc_hd__nor2_1 U20957 ( .A(n13889), .B(n13888), .Y(n13890) );
  sky130_fd_sc_hd__nand3_1 U20958 ( .A(n13891), .B(n12120), .C(n13890), .Y(
        n26375) );
  sky130_fd_sc_hd__inv_2 U20959 ( .A(n26375), .Y(n26284) );
  sky130_fd_sc_hd__o22ai_1 U20960 ( .A1(n16501), .A2(n26284), .B1(n11188), 
        .B2(n16500), .Y(n13922) );
  sky130_fd_sc_hd__nor2_1 U20961 ( .A(n13922), .B(n11105), .Y(n20431) );
  sky130_fd_sc_hd__o22ai_1 U20962 ( .A1(n16500), .A2(n26284), .B1(n27147), 
        .B2(n16501), .Y(n13923) );
  sky130_fd_sc_hd__nand2_1 U20963 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[194]), .Y(n13895) );
  sky130_fd_sc_hd__nand2_1 U20964 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[449]), .Y(n13894) );
  sky130_fd_sc_hd__nand2_1 U20965 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[481]), .Y(n13893) );
  sky130_fd_sc_hd__nand2_1 U20966 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[226]), .Y(n13892) );
  sky130_fd_sc_hd__nand4_1 U20967 ( .A(n13895), .B(n13894), .C(n13893), .D(
        n13892), .Y(n13901) );
  sky130_fd_sc_hd__nand2_1 U20968 ( .A(n16506), .B(
        j202_soc_core_j22_cpu_rf_gpr[2]), .Y(n13899) );
  sky130_fd_sc_hd__nand2_1 U20969 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[66]), .Y(n13898) );
  sky130_fd_sc_hd__nand2_1 U20970 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[385]), .Y(n13897) );
  sky130_fd_sc_hd__nand2_1 U20971 ( .A(n23808), .B(
        j202_soc_core_j22_cpu_rf_gpr[130]), .Y(n13896) );
  sky130_fd_sc_hd__nand4_1 U20972 ( .A(n13899), .B(n13898), .C(n13897), .D(
        n13896), .Y(n13900) );
  sky130_fd_sc_hd__nor2_1 U20973 ( .A(n13901), .B(n13900), .Y(n13912) );
  sky130_fd_sc_hd__nand2_1 U20974 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[258]), .Y(n13905) );
  sky130_fd_sc_hd__nand2_1 U20975 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[34]), .Y(n13904) );
  sky130_fd_sc_hd__nand2_1 U20976 ( .A(n15991), .B(
        j202_soc_core_j22_cpu_rf_gpr[353]), .Y(n13903) );
  sky130_fd_sc_hd__nand2_1 U20977 ( .A(n16064), .B(
        j202_soc_core_j22_cpu_rf_gpr[321]), .Y(n13902) );
  sky130_fd_sc_hd__and4_1 U20978 ( .A(n13904), .B(n13905), .C(n13903), .D(
        n13902), .X(n13911) );
  sky130_fd_sc_hd__nand2_1 U20979 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[290]), .Y(n13909) );
  sky130_fd_sc_hd__nand2_1 U20980 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[417]), .Y(n13908) );
  sky130_fd_sc_hd__nand2_1 U20981 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[162]), .Y(n13907) );
  sky130_fd_sc_hd__nand2_1 U20982 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[98]), .Y(n13906) );
  sky130_fd_sc_hd__and4_1 U20983 ( .A(n13909), .B(n13908), .C(n13907), .D(
        n13906), .X(n13910) );
  sky130_fd_sc_hd__o22a_1 U20984 ( .A1(n19271), .A2(n11202), .B1(n19270), .B2(
        n14342), .X(n13919) );
  sky130_fd_sc_hd__o22a_1 U20985 ( .A1(n13914), .A2(n16488), .B1(n16487), .B2(
        n13913), .X(n13918) );
  sky130_fd_sc_hd__o22a_1 U20986 ( .A1(n19266), .A2(n16491), .B1(n16490), .B2(
        n13915), .X(n13917) );
  sky130_fd_sc_hd__nand4_1 U20987 ( .A(n13919), .B(n13918), .C(n13917), .D(
        n13916), .Y(n13920) );
  sky130_fd_sc_hd__nand2_1 U20988 ( .A(n26937), .B(n16086), .Y(n13921) );
  sky130_fd_sc_hd__nor2_1 U20991 ( .A(n20431), .B(n17219), .Y(n13926) );
  sky130_fd_sc_hd__nand2_1 U20992 ( .A(n11105), .B(n13922), .Y(n20432) );
  sky130_fd_sc_hd__nand2_1 U20993 ( .A(n13924), .B(n13923), .Y(n17220) );
  sky130_fd_sc_hd__o21ai_1 U20994 ( .A1(n20432), .A2(n17219), .B1(n17220), .Y(
        n13925) );
  sky130_fd_sc_hd__a21oi_1 U20995 ( .A1(n17222), .A2(n13926), .B1(n13925), .Y(
        n20443) );
  sky130_fd_sc_hd__nand2_1 U20996 ( .A(n13928), .B(n13927), .Y(n21785) );
  sky130_fd_sc_hd__nand2_1 U20997 ( .A(n13930), .B(n13929), .Y(n21790) );
  sky130_fd_sc_hd__o21ai_1 U20998 ( .A1(n21789), .A2(n21785), .B1(n21790), .Y(
        n21328) );
  sky130_fd_sc_hd__nand2_1 U20999 ( .A(n13932), .B(n13931), .Y(n21664) );
  sky130_fd_sc_hd__nand2_1 U21000 ( .A(n13934), .B(n13933), .Y(n21326) );
  sky130_fd_sc_hd__o21ai_1 U21001 ( .A1(n21664), .A2(n21325), .B1(n21326), .Y(
        n13935) );
  sky130_fd_sc_hd__a21oi_1 U21002 ( .A1(n13936), .A2(n21328), .B1(n13935), .Y(
        n13937) );
  sky130_fd_sc_hd__o21ai_1 U21003 ( .A1(n13938), .A2(n20443), .B1(n13937), .Y(
        n18815) );
  sky130_fd_sc_hd__nor2_1 U21004 ( .A(n14010), .B(n14798), .Y(n13945) );
  sky130_fd_sc_hd__nand2_1 U21005 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[235]), .Y(n13943) );
  sky130_fd_sc_hd__nand2_1 U21006 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[267]), .Y(n13942) );
  sky130_fd_sc_hd__a2bb2oi_1 U21007 ( .B1(j202_soc_core_j22_cpu_rf_tmp[11]), 
        .B2(n13053), .A1_N(n14312), .A2_N(n30012), .Y(n13941) );
  sky130_fd_sc_hd__nand2_1 U21008 ( .A(n11195), .B(
        j202_soc_core_j22_cpu_rf_gpr[394]), .Y(n13940) );
  sky130_fd_sc_hd__nand4_1 U21009 ( .A(n13943), .B(n13942), .C(n13941), .D(
        n13940), .Y(n13944) );
  sky130_fd_sc_hd__nor2_1 U21010 ( .A(n13945), .B(n13944), .Y(n13963) );
  sky130_fd_sc_hd__nand2_1 U21011 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[330]), .Y(n13950) );
  sky130_fd_sc_hd__nand2_1 U21012 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[171]), .Y(n13949) );
  sky130_fd_sc_hd__nand2_1 U21013 ( .A(n15783), .B(
        j202_soc_core_j22_cpu_rf_gpr[107]), .Y(n13948) );
  sky130_fd_sc_hd__nand2_1 U21014 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[490]), .Y(n13947) );
  sky130_fd_sc_hd__nand2_1 U21015 ( .A(n16433), .B(
        j202_soc_core_j22_cpu_rf_gpr[203]), .Y(n13956) );
  sky130_fd_sc_hd__nand2_1 U21016 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[43]), .Y(n13955) );
  sky130_fd_sc_hd__nand2_1 U21017 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[139]), .Y(n13954) );
  sky130_fd_sc_hd__nand2_1 U21018 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[75]), .Y(n13953) );
  sky130_fd_sc_hd__nand2_1 U21019 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[362]), .Y(n13962) );
  sky130_fd_sc_hd__nand2_1 U21020 ( .A(n11194), .B(
        j202_soc_core_j22_cpu_rf_gpr[299]), .Y(n13961) );
  sky130_fd_sc_hd__nand2_1 U21021 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[458]), .Y(n13960) );
  sky130_fd_sc_hd__nand2_1 U21022 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[426]), .Y(n13959) );
  sky130_fd_sc_hd__inv_2 U21023 ( .A(n26941), .Y(n27025) );
  sky130_fd_sc_hd__nand2_1 U21024 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[266]), .Y(n13967) );
  sky130_fd_sc_hd__nand2_1 U21025 ( .A(n15788), .B(
        j202_soc_core_j22_cpu_rf_gpr[457]), .Y(n13966) );
  sky130_fd_sc_hd__nand2_1 U21026 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[393]), .Y(n13965) );
  sky130_fd_sc_hd__nand2_1 U21027 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[138]), .Y(n13964) );
  sky130_fd_sc_hd__nand4_1 U21028 ( .A(n13967), .B(n13966), .C(n13965), .D(
        n13964), .Y(n13973) );
  sky130_fd_sc_hd__nand2_1 U21029 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[74]), .Y(n13971) );
  sky130_fd_sc_hd__nand2_1 U21030 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[361]), .Y(n13970) );
  sky130_fd_sc_hd__nand2_1 U21031 ( .A(n15783), .B(
        j202_soc_core_j22_cpu_rf_gpr[106]), .Y(n13969) );
  sky130_fd_sc_hd__nand2_1 U21032 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[425]), .Y(n13968) );
  sky130_fd_sc_hd__nand4_1 U21033 ( .A(n13971), .B(n13970), .C(n13969), .D(
        n13968), .Y(n13972) );
  sky130_fd_sc_hd__nor2_1 U21034 ( .A(n13973), .B(n13972), .Y(n13986) );
  sky130_fd_sc_hd__nand2_1 U21035 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[298]), .Y(n13977) );
  sky130_fd_sc_hd__nand2_1 U21036 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[170]), .Y(n13976) );
  sky130_fd_sc_hd__nand2_1 U21037 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[202]), .Y(n13975) );
  sky130_fd_sc_hd__nand2_1 U21038 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[329]), .Y(n13974) );
  sky130_fd_sc_hd__nor2_1 U21039 ( .A(n14346), .B(n14798), .Y(n13984) );
  sky130_fd_sc_hd__nand2_1 U21040 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[42]), .Y(n13982) );
  sky130_fd_sc_hd__nand2_1 U21041 ( .A(n16043), .B(
        j202_soc_core_j22_cpu_rf_gpr[234]), .Y(n13981) );
  sky130_fd_sc_hd__a2bb2oi_1 U21042 ( .B1(j202_soc_core_j22_cpu_rf_tmp[10]), 
        .B2(n13053), .A1_N(n14312), .A2_N(n13978), .Y(n13980) );
  sky130_fd_sc_hd__nand2_1 U21043 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[489]), .Y(n13979) );
  sky130_fd_sc_hd__nand4_1 U21044 ( .A(n13982), .B(n13981), .C(n13980), .D(
        n13979), .Y(n13983) );
  sky130_fd_sc_hd__nor2_1 U21045 ( .A(n13984), .B(n13983), .Y(n13985) );
  sky130_fd_sc_hd__nand3_1 U21046 ( .A(n13986), .B(n13038), .C(n13985), .Y(
        n26923) );
  sky130_fd_sc_hd__inv_2 U21047 ( .A(n26923), .Y(n27798) );
  sky130_fd_sc_hd__o22ai_1 U21048 ( .A1(n16501), .A2(n27025), .B1(n27798), 
        .B2(n16500), .Y(n14398) );
  sky130_fd_sc_hd__nand2_1 U21049 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[203]), .Y(n13990) );
  sky130_fd_sc_hd__nand2_1 U21050 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[458]), .Y(n13989) );
  sky130_fd_sc_hd__nand2_1 U21051 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[490]), .Y(n13988) );
  sky130_fd_sc_hd__nand2_1 U21052 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[235]), .Y(n13987) );
  sky130_fd_sc_hd__nand4_1 U21053 ( .A(n13990), .B(n13989), .C(n13988), .D(
        n13987), .Y(n13996) );
  sky130_fd_sc_hd__nand2_1 U21054 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[11]), .Y(n13994) );
  sky130_fd_sc_hd__nand2_1 U21055 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[75]), .Y(n13993) );
  sky130_fd_sc_hd__nand2_1 U21056 ( .A(n16466), .B(
        j202_soc_core_j22_cpu_rf_gpr[394]), .Y(n13992) );
  sky130_fd_sc_hd__nand2_1 U21057 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[139]), .Y(n13991) );
  sky130_fd_sc_hd__nand4_1 U21058 ( .A(n13994), .B(n13993), .C(n13992), .D(
        n13991), .Y(n13995) );
  sky130_fd_sc_hd__nor2_1 U21059 ( .A(n13996), .B(n13995), .Y(n14008) );
  sky130_fd_sc_hd__nand2_1 U21060 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[267]), .Y(n14000) );
  sky130_fd_sc_hd__nand2_1 U21061 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[43]), .Y(n13999) );
  sky130_fd_sc_hd__nand2_1 U21062 ( .A(n15991), .B(
        j202_soc_core_j22_cpu_rf_gpr[362]), .Y(n13998) );
  sky130_fd_sc_hd__nand2_1 U21063 ( .A(n15017), .B(
        j202_soc_core_j22_cpu_rf_gpr[330]), .Y(n13997) );
  sky130_fd_sc_hd__and4_1 U21064 ( .A(n14000), .B(n13999), .C(n13998), .D(
        n13997), .X(n14007) );
  sky130_fd_sc_hd__nand2_1 U21065 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[299]), .Y(n14005) );
  sky130_fd_sc_hd__nand2_1 U21066 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[426]), .Y(n14004) );
  sky130_fd_sc_hd__nand2_1 U21067 ( .A(n11199), .B(
        j202_soc_core_j22_cpu_rf_gpr[171]), .Y(n14003) );
  sky130_fd_sc_hd__nand2_1 U21068 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[107]), .Y(n14002) );
  sky130_fd_sc_hd__and4_1 U21069 ( .A(n14005), .B(n14004), .C(n14003), .D(
        n14002), .X(n14006) );
  sky130_fd_sc_hd__nand3_1 U21070 ( .A(n14008), .B(n14007), .C(n14006), .Y(
        n21291) );
  sky130_fd_sc_hd__o22a_1 U21071 ( .A1(n21298), .A2(n16077), .B1(n21297), .B2(
        n14342), .X(n14015) );
  sky130_fd_sc_hd__o22a_1 U21072 ( .A1(n14010), .A2(n16488), .B1(n16487), .B2(
        n14009), .X(n14014) );
  sky130_fd_sc_hd__o22a_1 U21073 ( .A1(n21293), .A2(n16491), .B1(n16490), .B2(
        n14011), .X(n14013) );
  sky130_fd_sc_hd__nand4_1 U21074 ( .A(n14015), .B(n14014), .C(n14013), .D(
        n14012), .Y(n14016) );
  sky130_fd_sc_hd__nand2_1 U21075 ( .A(n27023), .B(n16086), .Y(n14017) );
  sky130_fd_sc_hd__o21ai_1 U21076 ( .A1(n16088), .A2(n27023), .B1(n14017), .Y(
        n14399) );
  sky130_fd_sc_hd__nor2_1 U21077 ( .A(n14398), .B(n14399), .Y(n20938) );
  sky130_fd_sc_hd__nand2_1 U21078 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[44]), .Y(n14021) );
  sky130_fd_sc_hd__nand2_1 U21079 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[76]), .Y(n14020) );
  sky130_fd_sc_hd__nand2_1 U21080 ( .A(n11195), .B(
        j202_soc_core_j22_cpu_rf_gpr[395]), .Y(n14019) );
  sky130_fd_sc_hd__nand2_1 U21081 ( .A(n11196), .B(
        j202_soc_core_j22_cpu_rf_gpr[363]), .Y(n14018) );
  sky130_fd_sc_hd__nand4_1 U21082 ( .A(n14021), .B(n14020), .C(n14019), .D(
        n14018), .Y(n14027) );
  sky130_fd_sc_hd__nand2_1 U21083 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[300]), .Y(n14025) );
  sky130_fd_sc_hd__nand2_1 U21084 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[172]), .Y(n14024) );
  sky130_fd_sc_hd__nand2_1 U21085 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[427]), .Y(n14023) );
  sky130_fd_sc_hd__nand2_1 U21086 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[268]), .Y(n14022) );
  sky130_fd_sc_hd__nand4_1 U21087 ( .A(n14025), .B(n14024), .C(n14023), .D(
        n14022), .Y(n14026) );
  sky130_fd_sc_hd__nor2_1 U21088 ( .A(n14027), .B(n14026), .Y(n14041) );
  sky130_fd_sc_hd__nand2_1 U21089 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[331]), .Y(n14031) );
  sky130_fd_sc_hd__nand2_1 U21090 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[204]), .Y(n14030) );
  sky130_fd_sc_hd__nand2_1 U21091 ( .A(n15783), .B(
        j202_soc_core_j22_cpu_rf_gpr[108]), .Y(n14029) );
  sky130_fd_sc_hd__nand2_1 U21092 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[459]), .Y(n14028) );
  sky130_fd_sc_hd__nor2_1 U21093 ( .A(n14032), .B(n16444), .Y(n14039) );
  sky130_fd_sc_hd__a21oi_1 U21094 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[12]), .B1(n14743), .Y(n14037) );
  sky130_fd_sc_hd__nand2_1 U21095 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[491]), .Y(n14036) );
  sky130_fd_sc_hd__nand2_1 U21096 ( .A(n16425), .B(
        j202_soc_core_j22_cpu_rf_gpr[140]), .Y(n14035) );
  sky130_fd_sc_hd__nand2_1 U21097 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[236]), .Y(n14034) );
  sky130_fd_sc_hd__nand4_1 U21098 ( .A(n14037), .B(n14036), .C(n14035), .D(
        n14034), .Y(n14038) );
  sky130_fd_sc_hd__nor2_1 U21099 ( .A(n14039), .B(n14038), .Y(n14040) );
  sky130_fd_sc_hd__nand3_1 U21100 ( .A(n14041), .B(n13039), .C(n14040), .Y(
        n26946) );
  sky130_fd_sc_hd__inv_2 U21101 ( .A(n26946), .Y(n26318) );
  sky130_fd_sc_hd__o22ai_1 U21102 ( .A1(n16500), .A2(n27025), .B1(n26318), 
        .B2(n16501), .Y(n14400) );
  sky130_fd_sc_hd__nand2_1 U21103 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[204]), .Y(n14045) );
  sky130_fd_sc_hd__nand2_1 U21104 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[459]), .Y(n14044) );
  sky130_fd_sc_hd__nand2_1 U21105 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[491]), .Y(n14043) );
  sky130_fd_sc_hd__nand2_1 U21106 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[236]), .Y(n14042) );
  sky130_fd_sc_hd__nand4_1 U21107 ( .A(n14045), .B(n14044), .C(n14043), .D(
        n14042), .Y(n14051) );
  sky130_fd_sc_hd__nand2_1 U21108 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[12]), .Y(n14049) );
  sky130_fd_sc_hd__nand2_1 U21109 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[76]), .Y(n14048) );
  sky130_fd_sc_hd__nand2_1 U21110 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[395]), .Y(n14047) );
  sky130_fd_sc_hd__nand2_1 U21111 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[140]), .Y(n14046) );
  sky130_fd_sc_hd__nand4_1 U21112 ( .A(n14049), .B(n14048), .C(n14047), .D(
        n14046), .Y(n14050) );
  sky130_fd_sc_hd__nor2_1 U21113 ( .A(n14051), .B(n14050), .Y(n14061) );
  sky130_fd_sc_hd__a22oi_1 U21114 ( .A1(n23776), .A2(
        j202_soc_core_j22_cpu_rf_gpr[363]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[268]), .Y(n14060) );
  sky130_fd_sc_hd__a22oi_1 U21115 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[44]), .B1(n15017), .B2(
        j202_soc_core_j22_cpu_rf_gpr[331]), .Y(n14059) );
  sky130_fd_sc_hd__nand2_1 U21116 ( .A(n15958), .B(
        j202_soc_core_j22_cpu_rf_gpr[300]), .Y(n14057) );
  sky130_fd_sc_hd__nand2_1 U21117 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[427]), .Y(n14056) );
  sky130_fd_sc_hd__nand2_1 U21118 ( .A(n11199), .B(
        j202_soc_core_j22_cpu_rf_gpr[172]), .Y(n14055) );
  sky130_fd_sc_hd__nand2_1 U21119 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[108]), .Y(n14054) );
  sky130_fd_sc_hd__and4_1 U21120 ( .A(n14057), .B(n14056), .C(n14055), .D(
        n14054), .X(n14058) );
  sky130_fd_sc_hd__nand4_1 U21121 ( .A(n14061), .B(n14060), .C(n14059), .D(
        n14058), .Y(n21892) );
  sky130_fd_sc_hd__nand2_1 U21122 ( .A(n21892), .B(n16523), .Y(n14070) );
  sky130_fd_sc_hd__o21ai_0 U21123 ( .A1(n21884), .A2(n16525), .B1(n16524), .Y(
        n14064) );
  sky130_fd_sc_hd__o22ai_1 U21124 ( .A1(n14062), .A2(n16077), .B1(n11095), 
        .B2(n14477), .Y(n14063) );
  sky130_fd_sc_hd__nor2_1 U21125 ( .A(n14064), .B(n14063), .Y(n14069) );
  sky130_fd_sc_hd__nand2_1 U21126 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[12]), .Y(n14068) );
  sky130_fd_sc_hd__nand2_1 U21127 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[12]), .Y(n14067) );
  sky130_fd_sc_hd__nand2_1 U21128 ( .A(n16533), .B(
        j202_soc_core_j22_cpu_pc[12]), .Y(n14066) );
  sky130_fd_sc_hd__nand2_1 U21129 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[12]), .Y(n14065) );
  sky130_fd_sc_hd__nand2_1 U21130 ( .A(n28460), .B(n16541), .Y(n14071) );
  sky130_fd_sc_hd__nor2_1 U21132 ( .A(n14400), .B(n14401), .Y(n20940) );
  sky130_fd_sc_hd__nor2_1 U21133 ( .A(n20938), .B(n20940), .Y(n20964) );
  sky130_fd_sc_hd__nand2_1 U21134 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[302]), .Y(n14075) );
  sky130_fd_sc_hd__nand2_1 U21135 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[270]), .Y(n14074) );
  sky130_fd_sc_hd__nand2_1 U21136 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[397]), .Y(n14073) );
  sky130_fd_sc_hd__nand2_1 U21137 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[429]), .Y(n14072) );
  sky130_fd_sc_hd__nand4_1 U21138 ( .A(n14075), .B(n14074), .C(n14073), .D(
        n14072), .Y(n14081) );
  sky130_fd_sc_hd__nand2_1 U21139 ( .A(n16043), .B(
        j202_soc_core_j22_cpu_rf_gpr[238]), .Y(n14079) );
  sky130_fd_sc_hd__nand2_1 U21140 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[46]), .Y(n14078) );
  sky130_fd_sc_hd__nand2_1 U21141 ( .A(n14993), .B(
        j202_soc_core_j22_cpu_rf_gpr[110]), .Y(n14077) );
  sky130_fd_sc_hd__nand2_1 U21142 ( .A(n15796), .B(
        j202_soc_core_j22_cpu_rf_gpr[78]), .Y(n14076) );
  sky130_fd_sc_hd__nand4_1 U21143 ( .A(n14079), .B(n14078), .C(n14077), .D(
        n14076), .Y(n14080) );
  sky130_fd_sc_hd__nor2_1 U21144 ( .A(n14081), .B(n14080), .Y(n14094) );
  sky130_fd_sc_hd__nand2_1 U21145 ( .A(n16410), .B(
        j202_soc_core_j22_cpu_rf_gpr[174]), .Y(n14086) );
  sky130_fd_sc_hd__nand2_1 U21146 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[333]), .Y(n14085) );
  sky130_fd_sc_hd__nand2_1 U21147 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[461]), .Y(n14084) );
  sky130_fd_sc_hd__nand2_1 U21148 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[206]), .Y(n14083) );
  sky130_fd_sc_hd__nor2_1 U21149 ( .A(n14144), .B(n14798), .Y(n14092) );
  sky130_fd_sc_hd__a21oi_1 U21150 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[14]), .B1(n14743), .Y(n14090) );
  sky130_fd_sc_hd__nand2_1 U21151 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[142]), .Y(n14089) );
  sky130_fd_sc_hd__nand2_1 U21152 ( .A(n13546), .B(
        j202_soc_core_j22_cpu_rf_gpr[493]), .Y(n14088) );
  sky130_fd_sc_hd__nand2_1 U21153 ( .A(n11196), .B(
        j202_soc_core_j22_cpu_rf_gpr[365]), .Y(n14087) );
  sky130_fd_sc_hd__nand4_1 U21154 ( .A(n14090), .B(n14089), .C(n14088), .D(
        n14087), .Y(n14091) );
  sky130_fd_sc_hd__nor2_1 U21155 ( .A(n14092), .B(n14091), .Y(n14093) );
  sky130_fd_sc_hd__inv_2 U21156 ( .A(n26009), .Y(n26319) );
  sky130_fd_sc_hd__nand2_1 U21157 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[205]), .Y(n14099) );
  sky130_fd_sc_hd__nand2_1 U21158 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[141]), .Y(n14098) );
  sky130_fd_sc_hd__nand2_1 U21159 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[492]), .Y(n14097) );
  sky130_fd_sc_hd__nand2_1 U21160 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[237]), .Y(n14096) );
  sky130_fd_sc_hd__nand4_1 U21161 ( .A(n14099), .B(n14098), .C(n14097), .D(
        n14096), .Y(n14105) );
  sky130_fd_sc_hd__nand2_1 U21162 ( .A(n11194), .B(
        j202_soc_core_j22_cpu_rf_gpr[301]), .Y(n14103) );
  sky130_fd_sc_hd__nand2_1 U21163 ( .A(n16432), .B(
        j202_soc_core_j22_cpu_rf_gpr[332]), .Y(n14102) );
  sky130_fd_sc_hd__nand2_1 U21164 ( .A(n14993), .B(
        j202_soc_core_j22_cpu_rf_gpr[109]), .Y(n14101) );
  sky130_fd_sc_hd__nand2_1 U21165 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[173]), .Y(n14100) );
  sky130_fd_sc_hd__nand4_1 U21166 ( .A(n14103), .B(n14102), .C(n14101), .D(
        n14100), .Y(n14104) );
  sky130_fd_sc_hd__nor2_1 U21167 ( .A(n14105), .B(n14104), .Y(n14119) );
  sky130_fd_sc_hd__nand2_1 U21168 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[77]), .Y(n14111) );
  sky130_fd_sc_hd__nand2_1 U21169 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[269]), .Y(n14110) );
  sky130_fd_sc_hd__nand2_1 U21170 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[396]), .Y(n14109) );
  sky130_fd_sc_hd__nand2_1 U21171 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[460]), .Y(n14108) );
  sky130_fd_sc_hd__nor2_1 U21172 ( .A(n14176), .B(n14798), .Y(n14117) );
  sky130_fd_sc_hd__a21oi_1 U21173 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[13]), .B1(n14743), .Y(n14115) );
  sky130_fd_sc_hd__nand2_1 U21174 ( .A(n11196), .B(
        j202_soc_core_j22_cpu_rf_gpr[364]), .Y(n14114) );
  sky130_fd_sc_hd__nand2_1 U21175 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[45]), .Y(n14113) );
  sky130_fd_sc_hd__nand2_1 U21176 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[428]), .Y(n14112) );
  sky130_fd_sc_hd__nand4_1 U21177 ( .A(n14115), .B(n14114), .C(n14113), .D(
        n14112), .Y(n14116) );
  sky130_fd_sc_hd__nor2_1 U21178 ( .A(n14117), .B(n14116), .Y(n14118) );
  sky130_fd_sc_hd__nand3_1 U21179 ( .A(n14119), .B(n13093), .C(n14118), .Y(
        n26050) );
  sky130_fd_sc_hd__inv_2 U21180 ( .A(n26050), .Y(n26321) );
  sky130_fd_sc_hd__o22ai_1 U21181 ( .A1(n16501), .A2(n26319), .B1(n26321), 
        .B2(n16500), .Y(n14404) );
  sky130_fd_sc_hd__nand2_1 U21182 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[206]), .Y(n14123) );
  sky130_fd_sc_hd__nand2_1 U21183 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[461]), .Y(n14122) );
  sky130_fd_sc_hd__nand2_1 U21184 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[493]), .Y(n14121) );
  sky130_fd_sc_hd__nand2_1 U21185 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[238]), .Y(n14120) );
  sky130_fd_sc_hd__nand4_1 U21186 ( .A(n14123), .B(n14122), .C(n14121), .D(
        n14120), .Y(n14129) );
  sky130_fd_sc_hd__nand2_1 U21187 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[14]), .Y(n14127) );
  sky130_fd_sc_hd__nand2_1 U21188 ( .A(n15984), .B(
        j202_soc_core_j22_cpu_rf_gpr[78]), .Y(n14126) );
  sky130_fd_sc_hd__nand2_1 U21189 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[397]), .Y(n14125) );
  sky130_fd_sc_hd__nand2_1 U21190 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[142]), .Y(n14124) );
  sky130_fd_sc_hd__nand4_1 U21191 ( .A(n14127), .B(n14126), .C(n14125), .D(
        n14124), .Y(n14128) );
  sky130_fd_sc_hd__nor2_1 U21192 ( .A(n14129), .B(n14128), .Y(n14140) );
  sky130_fd_sc_hd__nand2_1 U21193 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[270]), .Y(n14133) );
  sky130_fd_sc_hd__nand2_1 U21194 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[46]), .Y(n14132) );
  sky130_fd_sc_hd__nand2_1 U21195 ( .A(n15991), .B(
        j202_soc_core_j22_cpu_rf_gpr[365]), .Y(n14131) );
  sky130_fd_sc_hd__nand2_1 U21196 ( .A(n15017), .B(
        j202_soc_core_j22_cpu_rf_gpr[333]), .Y(n14130) );
  sky130_fd_sc_hd__and4_1 U21197 ( .A(n14133), .B(n14132), .C(n14131), .D(
        n14130), .X(n14139) );
  sky130_fd_sc_hd__nand2_1 U21198 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[302]), .Y(n14137) );
  sky130_fd_sc_hd__nand2_1 U21199 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[429]), .Y(n14136) );
  sky130_fd_sc_hd__nand2_1 U21200 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[174]), .Y(n14135) );
  sky130_fd_sc_hd__nand2_1 U21201 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[110]), .Y(n14134) );
  sky130_fd_sc_hd__and4_1 U21202 ( .A(n14137), .B(n14136), .C(n14135), .D(
        n14134), .X(n14138) );
  sky130_fd_sc_hd__nand3_1 U21203 ( .A(n14140), .B(n14139), .C(n14138), .Y(
        n22580) );
  sky130_fd_sc_hd__o22a_1 U21204 ( .A1(n14142), .A2(n16077), .B1(n14141), .B2(
        n14342), .X(n14149) );
  sky130_fd_sc_hd__o22a_1 U21205 ( .A1(n14144), .A2(n16488), .B1(n16487), .B2(
        n14143), .X(n14148) );
  sky130_fd_sc_hd__o22a_1 U21206 ( .A1(n22573), .A2(n16491), .B1(n16490), .B2(
        n14145), .X(n14147) );
  sky130_fd_sc_hd__a21oi_1 U21207 ( .A1(n11201), .A2(
        j202_soc_core_j22_cpu_rf_gpr[493]), .B1(n16493), .Y(n14146) );
  sky130_fd_sc_hd__nand4_1 U21208 ( .A(n14149), .B(n14148), .C(n14147), .D(
        n14146), .Y(n14150) );
  sky130_fd_sc_hd__a21oi_1 U21209 ( .A1(n22580), .A2(n16523), .B1(n14150), .Y(
        n25973) );
  sky130_fd_sc_hd__nand2_1 U21210 ( .A(n25973), .B(n16086), .Y(n14151) );
  sky130_fd_sc_hd__o21ai_1 U21211 ( .A1(n16088), .A2(n25973), .B1(n14151), .Y(
        n14405) );
  sky130_fd_sc_hd__nor2_1 U21212 ( .A(n14404), .B(n14405), .Y(n21011) );
  sky130_fd_sc_hd__o22ai_1 U21213 ( .A1(n16501), .A2(n26321), .B1(n26318), 
        .B2(n16500), .Y(n14402) );
  sky130_fd_sc_hd__nand2_1 U21214 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[205]), .Y(n14155) );
  sky130_fd_sc_hd__nand2_1 U21215 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[460]), .Y(n14154) );
  sky130_fd_sc_hd__nand2_1 U21216 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[492]), .Y(n14153) );
  sky130_fd_sc_hd__nand2_1 U21217 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[237]), .Y(n14152) );
  sky130_fd_sc_hd__nand4_1 U21218 ( .A(n14155), .B(n14154), .C(n14153), .D(
        n14152), .Y(n14161) );
  sky130_fd_sc_hd__nand2_1 U21219 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[13]), .Y(n14159) );
  sky130_fd_sc_hd__nand2_1 U21220 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[77]), .Y(n14158) );
  sky130_fd_sc_hd__nand2_1 U21221 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[396]), .Y(n14157) );
  sky130_fd_sc_hd__nand2_1 U21222 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[141]), .Y(n14156) );
  sky130_fd_sc_hd__nand4_1 U21223 ( .A(n14159), .B(n14158), .C(n14157), .D(
        n14156), .Y(n14160) );
  sky130_fd_sc_hd__nor2_1 U21224 ( .A(n14161), .B(n14160), .Y(n14172) );
  sky130_fd_sc_hd__nand2_1 U21225 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[269]), .Y(n14165) );
  sky130_fd_sc_hd__nand2_1 U21226 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[45]), .Y(n14164) );
  sky130_fd_sc_hd__nand2_1 U21227 ( .A(n23776), .B(
        j202_soc_core_j22_cpu_rf_gpr[364]), .Y(n14163) );
  sky130_fd_sc_hd__nand2_1 U21228 ( .A(n15017), .B(
        j202_soc_core_j22_cpu_rf_gpr[332]), .Y(n14162) );
  sky130_fd_sc_hd__and4_1 U21229 ( .A(n14165), .B(n14164), .C(n14163), .D(
        n14162), .X(n14171) );
  sky130_fd_sc_hd__nand2_1 U21230 ( .A(n15958), .B(
        j202_soc_core_j22_cpu_rf_gpr[301]), .Y(n14169) );
  sky130_fd_sc_hd__nand2_1 U21231 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[428]), .Y(n14168) );
  sky130_fd_sc_hd__nand2_1 U21232 ( .A(n11199), .B(
        j202_soc_core_j22_cpu_rf_gpr[173]), .Y(n14167) );
  sky130_fd_sc_hd__nand2_1 U21233 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[109]), .Y(n14166) );
  sky130_fd_sc_hd__and4_1 U21234 ( .A(n14169), .B(n14168), .C(n14167), .D(
        n14166), .X(n14170) );
  sky130_fd_sc_hd__nand3_1 U21235 ( .A(n14172), .B(n14171), .C(n14170), .Y(
        n22997) );
  sky130_fd_sc_hd__o22a_1 U21236 ( .A1(n14176), .A2(n16488), .B1(n16487), .B2(
        n14175), .X(n14180) );
  sky130_fd_sc_hd__o22a_1 U21237 ( .A1(n22984), .A2(n16491), .B1(n16490), .B2(
        n14177), .X(n14179) );
  sky130_fd_sc_hd__a21oi_1 U21238 ( .A1(n11201), .A2(
        j202_soc_core_j22_cpu_rf_gpr[492]), .B1(n16493), .Y(n14178) );
  sky130_fd_sc_hd__nand4_1 U21239 ( .A(n14181), .B(n14180), .C(n14179), .D(
        n14178), .Y(n14182) );
  sky130_fd_sc_hd__nand2_1 U21240 ( .A(n25451), .B(n16086), .Y(n14183) );
  sky130_fd_sc_hd__o21ai_1 U21241 ( .A1(n16088), .A2(n25451), .B1(n14183), .Y(
        n14403) );
  sky130_fd_sc_hd__nor2_1 U21242 ( .A(n14402), .B(n14403), .Y(n20963) );
  sky130_fd_sc_hd__nor2_1 U21243 ( .A(n21011), .B(n20963), .Y(n14407) );
  sky130_fd_sc_hd__nand2_1 U21244 ( .A(n20964), .B(n14407), .Y(n14409) );
  sky130_fd_sc_hd__nand2_1 U21245 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[327]), .Y(n14187) );
  sky130_fd_sc_hd__nand2_1 U21246 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[455]), .Y(n14186) );
  sky130_fd_sc_hd__nand2_1 U21247 ( .A(n14993), .B(
        j202_soc_core_j22_cpu_rf_gpr[104]), .Y(n14185) );
  sky130_fd_sc_hd__nand2_1 U21248 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[423]), .Y(n14184) );
  sky130_fd_sc_hd__nand4_1 U21249 ( .A(n14187), .B(n14186), .C(n14185), .D(
        n14184), .Y(n14193) );
  sky130_fd_sc_hd__nand2_1 U21250 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[40]), .Y(n14191) );
  sky130_fd_sc_hd__nand2_1 U21251 ( .A(n11196), .B(
        j202_soc_core_j22_cpu_rf_gpr[359]), .Y(n14190) );
  sky130_fd_sc_hd__nand2_1 U21252 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[487]), .Y(n14189) );
  sky130_fd_sc_hd__nand2_1 U21253 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[264]), .Y(n14188) );
  sky130_fd_sc_hd__nand4_1 U21254 ( .A(n14191), .B(n14190), .C(n14189), .D(
        n14188), .Y(n14192) );
  sky130_fd_sc_hd__nor2_1 U21255 ( .A(n14193), .B(n14192), .Y(n14208) );
  sky130_fd_sc_hd__nand2_1 U21256 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[296]), .Y(n14195) );
  sky130_fd_sc_hd__nand2_1 U21257 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[168]), .Y(n14194) );
  sky130_fd_sc_hd__nand2_1 U21258 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[200]), .Y(n14199) );
  sky130_fd_sc_hd__o22ai_1 U21259 ( .A1(n14196), .A2(n29066), .B1(n14256), 
        .B2(n14312), .Y(n14197) );
  sky130_fd_sc_hd__a21oi_1 U21260 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[8]), .B1(n14197), .Y(n14198) );
  sky130_fd_sc_hd__nand2_1 U21261 ( .A(n14199), .B(n14198), .Y(n14206) );
  sky130_fd_sc_hd__nand2_1 U21262 ( .A(n16425), .B(
        j202_soc_core_j22_cpu_rf_gpr[136]), .Y(n14204) );
  sky130_fd_sc_hd__nand2_1 U21263 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[232]), .Y(n14203) );
  sky130_fd_sc_hd__nand2_1 U21264 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[391]), .Y(n14202) );
  sky130_fd_sc_hd__nand2_1 U21265 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[72]), .Y(n14201) );
  sky130_fd_sc_hd__nand4_1 U21266 ( .A(n14204), .B(n14203), .C(n14202), .D(
        n14201), .Y(n14205) );
  sky130_fd_sc_hd__nor2_1 U21267 ( .A(n14206), .B(n14205), .Y(n14207) );
  sky130_fd_sc_hd__inv_2 U21269 ( .A(n26945), .Y(n26317) );
  sky130_fd_sc_hd__nand2_1 U21270 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[39]), .Y(n14213) );
  sky130_fd_sc_hd__nand2_1 U21271 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[135]), .Y(n14212) );
  sky130_fd_sc_hd__nand2_1 U21272 ( .A(n16398), .B(
        j202_soc_core_j22_cpu_rf_gpr[103]), .Y(n14211) );
  sky130_fd_sc_hd__nand2_1 U21273 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[71]), .Y(n14210) );
  sky130_fd_sc_hd__nand4_1 U21274 ( .A(n14213), .B(n14212), .C(n14211), .D(
        n14210), .Y(n14219) );
  sky130_fd_sc_hd__nand2_1 U21275 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[295]), .Y(n14217) );
  sky130_fd_sc_hd__nand2_1 U21276 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[167]), .Y(n14216) );
  sky130_fd_sc_hd__nand2_1 U21277 ( .A(n11195), .B(
        j202_soc_core_j22_cpu_rf_gpr[390]), .Y(n14215) );
  sky130_fd_sc_hd__nand2_1 U21278 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[263]), .Y(n14214) );
  sky130_fd_sc_hd__nand4_1 U21279 ( .A(n14217), .B(n14216), .C(n14215), .D(
        n14214), .Y(n14218) );
  sky130_fd_sc_hd__nor2_1 U21280 ( .A(n14219), .B(n14218), .Y(n14233) );
  sky130_fd_sc_hd__nand2_1 U21281 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[199]), .Y(n14224) );
  sky130_fd_sc_hd__nand2_1 U21282 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[326]), .Y(n14223) );
  sky130_fd_sc_hd__nand2_1 U21283 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[422]), .Y(n14222) );
  sky130_fd_sc_hd__nand2_1 U21284 ( .A(n15788), .B(
        j202_soc_core_j22_cpu_rf_gpr[454]), .Y(n14221) );
  sky130_fd_sc_hd__nor2_1 U21285 ( .A(n18864), .B(n14798), .Y(n14231) );
  sky130_fd_sc_hd__nand2_1 U21286 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[231]), .Y(n14229) );
  sky130_fd_sc_hd__nand2_1 U21287 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[358]), .Y(n14228) );
  sky130_fd_sc_hd__a2bb2oi_1 U21288 ( .B1(j202_soc_core_j22_cpu_rf_tmp[7]), 
        .B2(n13053), .A1_N(n14312), .A2_N(n14225), .Y(n14227) );
  sky130_fd_sc_hd__nand2_1 U21289 ( .A(n14985), .B(
        j202_soc_core_j22_cpu_rf_gpr[486]), .Y(n14226) );
  sky130_fd_sc_hd__nand4_1 U21290 ( .A(n14229), .B(n14228), .C(n14227), .D(
        n14226), .Y(n14230) );
  sky130_fd_sc_hd__nor2_1 U21291 ( .A(n14231), .B(n14230), .Y(n14232) );
  sky130_fd_sc_hd__o22ai_1 U21292 ( .A1(n16501), .A2(n26317), .B1(n27616), 
        .B2(n16500), .Y(n14390) );
  sky130_fd_sc_hd__nand2_1 U21293 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[200]), .Y(n14237) );
  sky130_fd_sc_hd__nand2_1 U21294 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[455]), .Y(n14236) );
  sky130_fd_sc_hd__nand2_1 U21295 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[487]), .Y(n14235) );
  sky130_fd_sc_hd__nand2_1 U21296 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[232]), .Y(n14234) );
  sky130_fd_sc_hd__nand4_1 U21297 ( .A(n14237), .B(n14236), .C(n14235), .D(
        n14234), .Y(n14243) );
  sky130_fd_sc_hd__nand2_1 U21298 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[8]), .Y(n14241) );
  sky130_fd_sc_hd__nand2_1 U21299 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[72]), .Y(n14240) );
  sky130_fd_sc_hd__nand2_1 U21300 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[391]), .Y(n14239) );
  sky130_fd_sc_hd__nand2_1 U21301 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[136]), .Y(n14238) );
  sky130_fd_sc_hd__nand4_1 U21302 ( .A(n14241), .B(n14240), .C(n14239), .D(
        n14238), .Y(n14242) );
  sky130_fd_sc_hd__nor2_1 U21303 ( .A(n14243), .B(n14242), .Y(n14254) );
  sky130_fd_sc_hd__nand2_1 U21304 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[264]), .Y(n14247) );
  sky130_fd_sc_hd__nand2_1 U21305 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[40]), .Y(n14246) );
  sky130_fd_sc_hd__nand2_1 U21306 ( .A(n23776), .B(
        j202_soc_core_j22_cpu_rf_gpr[359]), .Y(n14245) );
  sky130_fd_sc_hd__nand2_1 U21307 ( .A(n16064), .B(
        j202_soc_core_j22_cpu_rf_gpr[327]), .Y(n14244) );
  sky130_fd_sc_hd__and4_1 U21308 ( .A(n14247), .B(n14246), .C(n14245), .D(
        n14244), .X(n14253) );
  sky130_fd_sc_hd__nand2_1 U21309 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[296]), .Y(n14251) );
  sky130_fd_sc_hd__nand2_1 U21310 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[423]), .Y(n14250) );
  sky130_fd_sc_hd__nand2_1 U21311 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[168]), .Y(n14249) );
  sky130_fd_sc_hd__nand2_1 U21312 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[104]), .Y(n14248) );
  sky130_fd_sc_hd__and4_1 U21313 ( .A(n14251), .B(n14250), .C(n14249), .D(
        n14248), .X(n14252) );
  sky130_fd_sc_hd__nand3_1 U21314 ( .A(n14254), .B(n14253), .C(n14252), .Y(
        n21744) );
  sky130_fd_sc_hd__o22ai_1 U21315 ( .A1(n14256), .A2(n14255), .B1(n14482), 
        .B2(n21734), .Y(n14257) );
  sky130_fd_sc_hd__a21oi_1 U21316 ( .A1(n16534), .A2(
        j202_soc_core_j22_cpu_rf_gbr[8]), .B1(n14257), .Y(n14263) );
  sky130_fd_sc_hd__o22a_1 U21317 ( .A1(n14258), .A2(n14342), .B1(n21737), .B2(
        n14373), .X(n14262) );
  sky130_fd_sc_hd__o22a_1 U21318 ( .A1(n14259), .A2(n16488), .B1(n21735), .B2(
        n16491), .X(n14260) );
  sky130_fd_sc_hd__nand4_1 U21319 ( .A(n14263), .B(n14262), .C(n14261), .D(
        n14260), .Y(n14264) );
  sky130_fd_sc_hd__mux2i_1 U21320 ( .A0(n16088), .A1(n16543), .S(n24931), .Y(
        n14391) );
  sky130_fd_sc_hd__nor2_1 U21321 ( .A(n14390), .B(n14391), .Y(n22748) );
  sky130_fd_sc_hd__o22ai_1 U21322 ( .A1(n16500), .A2(n11191), .B1(n27616), 
        .B2(n16501), .Y(n14388) );
  sky130_fd_sc_hd__nand2_1 U21323 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[199]), .Y(n14268) );
  sky130_fd_sc_hd__nand2_1 U21325 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[486]), .Y(n14266) );
  sky130_fd_sc_hd__nand2_1 U21326 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[231]), .Y(n14265) );
  sky130_fd_sc_hd__nand4_1 U21327 ( .A(n14268), .B(n14267), .C(n14266), .D(
        n14265), .Y(n14274) );
  sky130_fd_sc_hd__nand2_1 U21328 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[7]), .Y(n14272) );
  sky130_fd_sc_hd__nand2_1 U21329 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[71]), .Y(n14271) );
  sky130_fd_sc_hd__nand2_1 U21330 ( .A(n16466), .B(
        j202_soc_core_j22_cpu_rf_gpr[390]), .Y(n14270) );
  sky130_fd_sc_hd__nand2_1 U21331 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[135]), .Y(n14269) );
  sky130_fd_sc_hd__nand4_1 U21332 ( .A(n14272), .B(n14271), .C(n14270), .D(
        n14269), .Y(n14273) );
  sky130_fd_sc_hd__nor2_1 U21333 ( .A(n14274), .B(n14273), .Y(n14284) );
  sky130_fd_sc_hd__a22oi_1 U21334 ( .A1(n23776), .A2(
        j202_soc_core_j22_cpu_rf_gpr[358]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[263]), .Y(n14283) );
  sky130_fd_sc_hd__a22oi_1 U21335 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[39]), .B1(n15017), .B2(
        j202_soc_core_j22_cpu_rf_gpr[326]), .Y(n14282) );
  sky130_fd_sc_hd__nand2_1 U21336 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[295]), .Y(n14279) );
  sky130_fd_sc_hd__nand2_1 U21337 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[422]), .Y(n14278) );
  sky130_fd_sc_hd__nand2_1 U21338 ( .A(n11199), .B(
        j202_soc_core_j22_cpu_rf_gpr[167]), .Y(n14277) );
  sky130_fd_sc_hd__nand2_1 U21339 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[103]), .Y(n14276) );
  sky130_fd_sc_hd__nand4_1 U21341 ( .A(n14284), .B(n14283), .C(n14282), .D(
        n30024), .Y(n18858) );
  sky130_fd_sc_hd__o22ai_1 U21342 ( .A1(n18867), .A2(n11202), .B1(n16487), 
        .B2(n14285), .Y(n14287) );
  sky130_fd_sc_hd__o22ai_1 U21343 ( .A1(n18874), .A2(n14477), .B1(n14373), 
        .B2(n18866), .Y(n14286) );
  sky130_fd_sc_hd__nor2_1 U21344 ( .A(n14287), .B(n14286), .Y(n14294) );
  sky130_fd_sc_hd__o21ai_0 U21345 ( .A1(n14289), .A2(n16490), .B1(n14288), .Y(
        n14292) );
  sky130_fd_sc_hd__o22ai_1 U21346 ( .A1(n18864), .A2(n16488), .B1(n16491), 
        .B2(n14290), .Y(n14291) );
  sky130_fd_sc_hd__nor2_1 U21347 ( .A(n14292), .B(n14291), .Y(n14293) );
  sky130_fd_sc_hd__mux2i_1 U21348 ( .A0(n16543), .A1(n16088), .S(n28489), .Y(
        n14389) );
  sky130_fd_sc_hd__nor2_1 U21349 ( .A(n14388), .B(n14389), .Y(n22753) );
  sky130_fd_sc_hd__nor2_1 U21350 ( .A(n22748), .B(n22753), .Y(n21341) );
  sky130_fd_sc_hd__nand2_1 U21351 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[424]), .Y(n14299) );
  sky130_fd_sc_hd__nand2_1 U21352 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[265]), .Y(n14298) );
  sky130_fd_sc_hd__nand2_1 U21353 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[392]), .Y(n14297) );
  sky130_fd_sc_hd__nand2_1 U21354 ( .A(n16398), .B(
        j202_soc_core_j22_cpu_rf_gpr[105]), .Y(n14296) );
  sky130_fd_sc_hd__nand4_1 U21355 ( .A(n14299), .B(n14298), .C(n14297), .D(
        n14296), .Y(n14305) );
  sky130_fd_sc_hd__nand2_1 U21356 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[201]), .Y(n14303) );
  sky130_fd_sc_hd__nand2_1 U21357 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[233]), .Y(n14302) );
  sky130_fd_sc_hd__nand2_1 U21358 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[488]), .Y(n14301) );
  sky130_fd_sc_hd__nand2_1 U21359 ( .A(n15796), .B(
        j202_soc_core_j22_cpu_rf_gpr[73]), .Y(n14300) );
  sky130_fd_sc_hd__nand4_1 U21360 ( .A(n14303), .B(n14302), .C(n14301), .D(
        n14300), .Y(n14304) );
  sky130_fd_sc_hd__nor2_1 U21361 ( .A(n14305), .B(n14304), .Y(n14320) );
  sky130_fd_sc_hd__nand2_1 U21362 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[328]), .Y(n14309) );
  sky130_fd_sc_hd__nand2_1 U21363 ( .A(n16410), .B(
        j202_soc_core_j22_cpu_rf_gpr[169]), .Y(n14308) );
  sky130_fd_sc_hd__nand2_1 U21364 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[360]), .Y(n14307) );
  sky130_fd_sc_hd__nand2_1 U21365 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[456]), .Y(n14306) );
  sky130_fd_sc_hd__nor2_1 U21366 ( .A(n14310), .B(n16444), .Y(n14318) );
  sky130_fd_sc_hd__nand2_1 U21367 ( .A(n11194), .B(
        j202_soc_core_j22_cpu_rf_gpr[297]), .Y(n14316) );
  sky130_fd_sc_hd__nand2_1 U21368 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[41]), .Y(n14315) );
  sky130_fd_sc_hd__a2bb2oi_1 U21369 ( .B1(j202_soc_core_j22_cpu_rf_tmp[9]), 
        .B2(n13053), .A1_N(n14312), .A2_N(n30027), .Y(n14314) );
  sky130_fd_sc_hd__nand2_1 U21370 ( .A(n16425), .B(
        j202_soc_core_j22_cpu_rf_gpr[137]), .Y(n14313) );
  sky130_fd_sc_hd__nand4_1 U21371 ( .A(n14316), .B(n14315), .C(n14314), .D(
        n14313), .Y(n14317) );
  sky130_fd_sc_hd__nor2_1 U21372 ( .A(n14318), .B(n14317), .Y(n14319) );
  sky130_fd_sc_hd__nand3_1 U21373 ( .A(n14320), .B(n13064), .C(n14319), .Y(
        n25916) );
  sky130_fd_sc_hd__inv_2 U21374 ( .A(n25916), .Y(n26944) );
  sky130_fd_sc_hd__o22ai_1 U21375 ( .A1(n16500), .A2(n26944), .B1(n27798), 
        .B2(n16501), .Y(n14394) );
  sky130_fd_sc_hd__nand2_1 U21376 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[202]), .Y(n14324) );
  sky130_fd_sc_hd__nand2_1 U21377 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[457]), .Y(n14323) );
  sky130_fd_sc_hd__nand2_1 U21378 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[489]), .Y(n14322) );
  sky130_fd_sc_hd__nand2_1 U21379 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[234]), .Y(n14321) );
  sky130_fd_sc_hd__nand4_1 U21380 ( .A(n14324), .B(n14323), .C(n14322), .D(
        n14321), .Y(n14330) );
  sky130_fd_sc_hd__nand2_1 U21381 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[10]), .Y(n14328) );
  sky130_fd_sc_hd__nand2_1 U21382 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[74]), .Y(n14327) );
  sky130_fd_sc_hd__nand2_1 U21383 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[393]), .Y(n14326) );
  sky130_fd_sc_hd__nand2_1 U21384 ( .A(n23808), .B(
        j202_soc_core_j22_cpu_rf_gpr[138]), .Y(n14325) );
  sky130_fd_sc_hd__nand4_1 U21385 ( .A(n14328), .B(n14327), .C(n14326), .D(
        n14325), .Y(n14329) );
  sky130_fd_sc_hd__nor2_1 U21386 ( .A(n14330), .B(n14329), .Y(n14341) );
  sky130_fd_sc_hd__nand2_1 U21387 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[266]), .Y(n14334) );
  sky130_fd_sc_hd__nand2_1 U21388 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[42]), .Y(n14333) );
  sky130_fd_sc_hd__nand2_1 U21389 ( .A(n23776), .B(
        j202_soc_core_j22_cpu_rf_gpr[361]), .Y(n14332) );
  sky130_fd_sc_hd__nand2_1 U21390 ( .A(n16064), .B(
        j202_soc_core_j22_cpu_rf_gpr[329]), .Y(n14331) );
  sky130_fd_sc_hd__and4_1 U21391 ( .A(n14334), .B(n14333), .C(n14332), .D(
        n14331), .X(n14340) );
  sky130_fd_sc_hd__nand2_1 U21392 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[298]), .Y(n14338) );
  sky130_fd_sc_hd__nand2_1 U21393 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[425]), .Y(n14337) );
  sky130_fd_sc_hd__nand2_1 U21394 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[170]), .Y(n14336) );
  sky130_fd_sc_hd__nand2_1 U21395 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[106]), .Y(n14335) );
  sky130_fd_sc_hd__and4_1 U21396 ( .A(n14338), .B(n14337), .C(n14336), .D(
        n14335), .X(n14339) );
  sky130_fd_sc_hd__nand3_1 U21397 ( .A(n14341), .B(n14340), .C(n14339), .Y(
        n19290) );
  sky130_fd_sc_hd__o22a_1 U21398 ( .A1(n14346), .A2(n16488), .B1(n16487), .B2(
        n14345), .X(n14350) );
  sky130_fd_sc_hd__o22a_1 U21399 ( .A1(n19283), .A2(n16491), .B1(n16490), .B2(
        n14347), .X(n14349) );
  sky130_fd_sc_hd__nand4_1 U21400 ( .A(n14351), .B(n14350), .C(n14349), .D(
        n14348), .Y(n14352) );
  sky130_fd_sc_hd__a21oi_1 U21401 ( .A1(n19290), .A2(n16523), .B1(n14352), .Y(
        n27816) );
  sky130_fd_sc_hd__nand2_1 U21402 ( .A(n27816), .B(n16086), .Y(n14353) );
  sky130_fd_sc_hd__nor2_1 U21404 ( .A(n14394), .B(n14395), .Y(n22693) );
  sky130_fd_sc_hd__o22ai_1 U21405 ( .A1(n16501), .A2(n26944), .B1(n26317), 
        .B2(n16500), .Y(n14392) );
  sky130_fd_sc_hd__nand2_1 U21406 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[201]), .Y(n14357) );
  sky130_fd_sc_hd__nand2_1 U21407 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[456]), .Y(n14356) );
  sky130_fd_sc_hd__nand2_1 U21408 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[488]), .Y(n14355) );
  sky130_fd_sc_hd__nand2_1 U21409 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[233]), .Y(n14354) );
  sky130_fd_sc_hd__nand4_1 U21410 ( .A(n14357), .B(n14356), .C(n14355), .D(
        n14354), .Y(n14363) );
  sky130_fd_sc_hd__nand2_1 U21411 ( .A(n16506), .B(
        j202_soc_core_j22_cpu_rf_gpr[9]), .Y(n14361) );
  sky130_fd_sc_hd__nand2_1 U21412 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[73]), .Y(n14360) );
  sky130_fd_sc_hd__nand2_1 U21413 ( .A(n16466), .B(
        j202_soc_core_j22_cpu_rf_gpr[392]), .Y(n14359) );
  sky130_fd_sc_hd__nand2_1 U21414 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[137]), .Y(n14358) );
  sky130_fd_sc_hd__nand4_1 U21415 ( .A(n14361), .B(n14360), .C(n14359), .D(
        n14358), .Y(n14362) );
  sky130_fd_sc_hd__nor2_1 U21416 ( .A(n14363), .B(n14362), .Y(n14372) );
  sky130_fd_sc_hd__a22oi_1 U21417 ( .A1(n23776), .A2(
        j202_soc_core_j22_cpu_rf_gpr[360]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[265]), .Y(n14371) );
  sky130_fd_sc_hd__a22oi_1 U21418 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[41]), .B1(n15017), .B2(
        j202_soc_core_j22_cpu_rf_gpr[328]), .Y(n14370) );
  sky130_fd_sc_hd__nand2_1 U21419 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[297]), .Y(n14368) );
  sky130_fd_sc_hd__nand2_1 U21420 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[424]), .Y(n14367) );
  sky130_fd_sc_hd__nand2_1 U21421 ( .A(n11199), .B(
        j202_soc_core_j22_cpu_rf_gpr[169]), .Y(n14366) );
  sky130_fd_sc_hd__nand2_1 U21422 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[105]), .Y(n14365) );
  sky130_fd_sc_hd__and4_1 U21423 ( .A(n14368), .B(n14367), .C(n14366), .D(
        n14365), .X(n14369) );
  sky130_fd_sc_hd__nand4_1 U21424 ( .A(n14372), .B(n14371), .C(n14370), .D(
        n14369), .Y(n22903) );
  sky130_fd_sc_hd__nand2_1 U21425 ( .A(n22903), .B(n16523), .Y(n14386) );
  sky130_fd_sc_hd__o22ai_1 U21426 ( .A1(n22896), .A2(n11202), .B1(n22895), 
        .B2(n14373), .Y(n14377) );
  sky130_fd_sc_hd__o22ai_1 U21427 ( .A1(n14375), .A2(n16487), .B1(n14477), 
        .B2(n14374), .Y(n14376) );
  sky130_fd_sc_hd__nor2_1 U21428 ( .A(n14377), .B(n14376), .Y(n14385) );
  sky130_fd_sc_hd__nand2_1 U21429 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[9]), .Y(n14382) );
  sky130_fd_sc_hd__nand2_1 U21430 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[9]), .Y(n14381) );
  sky130_fd_sc_hd__nand2_1 U21431 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[9]), .Y(n14379) );
  sky130_fd_sc_hd__nand4_1 U21432 ( .A(n14382), .B(n14381), .C(n14380), .D(
        n14379), .Y(n14383) );
  sky130_fd_sc_hd__nand3_1 U21433 ( .A(n14386), .B(n14385), .C(n14384), .Y(
        n28478) );
  sky130_fd_sc_hd__nand2_1 U21434 ( .A(n28478), .B(n16541), .Y(n14387) );
  sky130_fd_sc_hd__o21ai_1 U21435 ( .A1(n16543), .A2(n28478), .B1(n14387), .Y(
        n14393) );
  sky130_fd_sc_hd__nor2_1 U21436 ( .A(n14392), .B(n14393), .Y(n21340) );
  sky130_fd_sc_hd__nor2_1 U21437 ( .A(n22693), .B(n21340), .Y(n14397) );
  sky130_fd_sc_hd__nand2_1 U21438 ( .A(n21341), .B(n14397), .Y(n20937) );
  sky130_fd_sc_hd__nor2_1 U21439 ( .A(n14409), .B(n20937), .Y(n14411) );
  sky130_fd_sc_hd__nand2_1 U21440 ( .A(n14389), .B(n14388), .Y(n22751) );
  sky130_fd_sc_hd__nand2_1 U21441 ( .A(n14391), .B(n14390), .Y(n22749) );
  sky130_fd_sc_hd__nand2_1 U21443 ( .A(n14393), .B(n14392), .Y(n22689) );
  sky130_fd_sc_hd__nand2_1 U21444 ( .A(n14395), .B(n14394), .Y(n22694) );
  sky130_fd_sc_hd__o21ai_1 U21445 ( .A1(n22689), .A2(n22693), .B1(n22694), .Y(
        n14396) );
  sky130_fd_sc_hd__a21oi_1 U21446 ( .A1(n14397), .A2(n21342), .B1(n14396), .Y(
        n20936) );
  sky130_fd_sc_hd__nand2_1 U21447 ( .A(n14399), .B(n14398), .Y(n21180) );
  sky130_fd_sc_hd__nand2_1 U21448 ( .A(n14401), .B(n14400), .Y(n20941) );
  sky130_fd_sc_hd__o21ai_1 U21449 ( .A1(n21180), .A2(n20940), .B1(n20941), .Y(
        n20966) );
  sky130_fd_sc_hd__nand2_1 U21450 ( .A(n14403), .B(n14402), .Y(n21007) );
  sky130_fd_sc_hd__nand2_1 U21451 ( .A(n14405), .B(n14404), .Y(n21012) );
  sky130_fd_sc_hd__a21oi_1 U21453 ( .A1(n14407), .A2(n20966), .B1(n14406), .Y(
        n14408) );
  sky130_fd_sc_hd__o21ai_1 U21454 ( .A1(n14409), .A2(n20936), .B1(n14408), .Y(
        n14410) );
  sky130_fd_sc_hd__nand2_1 U21455 ( .A(n16425), .B(
        j202_soc_core_j22_cpu_rf_gpr[145]), .Y(n14415) );
  sky130_fd_sc_hd__nand2_1 U21456 ( .A(n15796), .B(
        j202_soc_core_j22_cpu_rf_gpr[81]), .Y(n14414) );
  sky130_fd_sc_hd__nand2_1 U21457 ( .A(n11195), .B(
        j202_soc_core_j22_cpu_rf_gpr[400]), .Y(n14413) );
  sky130_fd_sc_hd__nand2_1 U21458 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[368]), .Y(n14412) );
  sky130_fd_sc_hd__nand4_1 U21459 ( .A(n14415), .B(n14414), .C(n14413), .D(
        n14412), .Y(n14421) );
  sky130_fd_sc_hd__nand2_1 U21460 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[273]), .Y(n14419) );
  sky130_fd_sc_hd__nand2_1 U21461 ( .A(n11194), .B(
        j202_soc_core_j22_cpu_rf_gpr[305]), .Y(n14418) );
  sky130_fd_sc_hd__nand2_1 U21462 ( .A(n15788), .B(
        j202_soc_core_j22_cpu_rf_gpr[464]), .Y(n14417) );
  sky130_fd_sc_hd__nand2_1 U21463 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[432]), .Y(n14416) );
  sky130_fd_sc_hd__nand4_1 U21464 ( .A(n14419), .B(n14418), .C(n14417), .D(
        n14416), .Y(n14420) );
  sky130_fd_sc_hd__nor2_1 U21465 ( .A(n14421), .B(n14420), .Y(n14433) );
  sky130_fd_sc_hd__nand2_1 U21466 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[336]), .Y(n14425) );
  sky130_fd_sc_hd__nand2_1 U21467 ( .A(n16410), .B(
        j202_soc_core_j22_cpu_rf_gpr[177]), .Y(n14424) );
  sky130_fd_sc_hd__nand2_1 U21468 ( .A(n16398), .B(
        j202_soc_core_j22_cpu_rf_gpr[113]), .Y(n14423) );
  sky130_fd_sc_hd__nand2_1 U21469 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[209]), .Y(n14422) );
  sky130_fd_sc_hd__nor2_1 U21470 ( .A(n14480), .B(n14798), .Y(n14431) );
  sky130_fd_sc_hd__a21oi_1 U21471 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[17]), .B1(n14743), .Y(n14429) );
  sky130_fd_sc_hd__nand2_1 U21472 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[241]), .Y(n14428) );
  sky130_fd_sc_hd__nand2_1 U21473 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[496]), .Y(n14427) );
  sky130_fd_sc_hd__nand2_1 U21474 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[49]), .Y(n14426) );
  sky130_fd_sc_hd__nand4_1 U21475 ( .A(n14429), .B(n14428), .C(n14427), .D(
        n14426), .Y(n14430) );
  sky130_fd_sc_hd__nor2_1 U21476 ( .A(n14431), .B(n14430), .Y(n14432) );
  sky130_fd_sc_hd__inv_2 U21477 ( .A(n26051), .Y(n26320) );
  sky130_fd_sc_hd__nand2_1 U21478 ( .A(n16425), .B(
        j202_soc_core_j22_cpu_rf_gpr[144]), .Y(n14437) );
  sky130_fd_sc_hd__nand2_1 U21479 ( .A(n15796), .B(
        j202_soc_core_j22_cpu_rf_gpr[80]), .Y(n14436) );
  sky130_fd_sc_hd__nand2_1 U21480 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[399]), .Y(n14435) );
  sky130_fd_sc_hd__nand2_1 U21481 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[367]), .Y(n14434) );
  sky130_fd_sc_hd__nand4_1 U21482 ( .A(n14437), .B(n14436), .C(n14435), .D(
        n14434), .Y(n14443) );
  sky130_fd_sc_hd__nand2_1 U21483 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[272]), .Y(n14441) );
  sky130_fd_sc_hd__nand2_1 U21484 ( .A(n11194), .B(
        j202_soc_core_j22_cpu_rf_gpr[304]), .Y(n14440) );
  sky130_fd_sc_hd__nand2_1 U21485 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[463]), .Y(n14439) );
  sky130_fd_sc_hd__nand2_1 U21486 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[431]), .Y(n14438) );
  sky130_fd_sc_hd__nand4_1 U21487 ( .A(n14441), .B(n14440), .C(n14439), .D(
        n14438), .Y(n14442) );
  sky130_fd_sc_hd__nor2_1 U21488 ( .A(n14443), .B(n14442), .Y(n14455) );
  sky130_fd_sc_hd__nand2_1 U21489 ( .A(n16432), .B(
        j202_soc_core_j22_cpu_rf_gpr[335]), .Y(n14447) );
  sky130_fd_sc_hd__nand2_1 U21490 ( .A(n16410), .B(
        j202_soc_core_j22_cpu_rf_gpr[176]), .Y(n14446) );
  sky130_fd_sc_hd__nand2_1 U21491 ( .A(n14993), .B(
        j202_soc_core_j22_cpu_rf_gpr[112]), .Y(n14445) );
  sky130_fd_sc_hd__nand2_1 U21492 ( .A(n16433), .B(
        j202_soc_core_j22_cpu_rf_gpr[208]), .Y(n14444) );
  sky130_fd_sc_hd__nor2_1 U21493 ( .A(n14536), .B(n14798), .Y(n14453) );
  sky130_fd_sc_hd__a21oi_1 U21494 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[16]), .B1(n14743), .Y(n14451) );
  sky130_fd_sc_hd__nand2_1 U21495 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[240]), .Y(n14450) );
  sky130_fd_sc_hd__nand2_1 U21496 ( .A(n14985), .B(
        j202_soc_core_j22_cpu_rf_gpr[495]), .Y(n14449) );
  sky130_fd_sc_hd__nand2_1 U21497 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[48]), .Y(n14448) );
  sky130_fd_sc_hd__nand4_1 U21498 ( .A(n14451), .B(n14450), .C(n14449), .D(
        n14448), .Y(n14452) );
  sky130_fd_sc_hd__nor2_1 U21499 ( .A(n14453), .B(n14452), .Y(n14454) );
  sky130_fd_sc_hd__inv_2 U21500 ( .A(n27111), .Y(n26322) );
  sky130_fd_sc_hd__o22ai_1 U21501 ( .A1(n16501), .A2(n26320), .B1(n26322), 
        .B2(n16500), .Y(n14577) );
  sky130_fd_sc_hd__nand2_1 U21502 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[209]), .Y(n14459) );
  sky130_fd_sc_hd__nand2_1 U21503 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[464]), .Y(n14458) );
  sky130_fd_sc_hd__nand2_1 U21504 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[496]), .Y(n14457) );
  sky130_fd_sc_hd__nand2_1 U21505 ( .A(n13821), .B(
        j202_soc_core_j22_cpu_rf_gpr[241]), .Y(n14456) );
  sky130_fd_sc_hd__nand4_1 U21506 ( .A(n14459), .B(n14458), .C(n14457), .D(
        n14456), .Y(n14465) );
  sky130_fd_sc_hd__nand2_1 U21507 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[17]), .Y(n14463) );
  sky130_fd_sc_hd__nand2_1 U21508 ( .A(n15984), .B(
        j202_soc_core_j22_cpu_rf_gpr[81]), .Y(n14462) );
  sky130_fd_sc_hd__nand2_1 U21509 ( .A(n13411), .B(
        j202_soc_core_j22_cpu_rf_gpr[400]), .Y(n14461) );
  sky130_fd_sc_hd__nand2_1 U21510 ( .A(n23808), .B(
        j202_soc_core_j22_cpu_rf_gpr[145]), .Y(n14460) );
  sky130_fd_sc_hd__nand4_1 U21511 ( .A(n14463), .B(n14462), .C(n14461), .D(
        n14460), .Y(n14464) );
  sky130_fd_sc_hd__nor2_1 U21512 ( .A(n14465), .B(n14464), .Y(n14476) );
  sky130_fd_sc_hd__nand2_1 U21513 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[273]), .Y(n14469) );
  sky130_fd_sc_hd__nand2_1 U21514 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[49]), .Y(n14468) );
  sky130_fd_sc_hd__nand2_1 U21515 ( .A(n23776), .B(
        j202_soc_core_j22_cpu_rf_gpr[368]), .Y(n14467) );
  sky130_fd_sc_hd__nand2_1 U21516 ( .A(n16064), .B(
        j202_soc_core_j22_cpu_rf_gpr[336]), .Y(n14466) );
  sky130_fd_sc_hd__and4_1 U21517 ( .A(n14469), .B(n14468), .C(n14467), .D(
        n14466), .X(n14475) );
  sky130_fd_sc_hd__nand2_1 U21518 ( .A(n15958), .B(
        j202_soc_core_j22_cpu_rf_gpr[305]), .Y(n14473) );
  sky130_fd_sc_hd__nand2_1 U21519 ( .A(n13383), .B(
        j202_soc_core_j22_cpu_rf_gpr[432]), .Y(n14472) );
  sky130_fd_sc_hd__nand2_1 U21520 ( .A(n11199), .B(
        j202_soc_core_j22_cpu_rf_gpr[177]), .Y(n14471) );
  sky130_fd_sc_hd__nand2_1 U21521 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[113]), .Y(n14470) );
  sky130_fd_sc_hd__and4_1 U21522 ( .A(n14473), .B(n14472), .C(n14471), .D(
        n14470), .X(n14474) );
  sky130_fd_sc_hd__nand3_1 U21523 ( .A(n14476), .B(n14475), .C(n14474), .Y(
        n22855) );
  sky130_fd_sc_hd__o22a_1 U21524 ( .A1(n14480), .A2(n16488), .B1(n16487), .B2(
        n22849), .X(n14485) );
  sky130_fd_sc_hd__o22a_1 U21525 ( .A1(n14481), .A2(n16491), .B1(n16490), .B2(
        n22856), .X(n14484) );
  sky130_fd_sc_hd__a21oi_1 U21526 ( .A1(n11201), .A2(
        j202_soc_core_j22_cpu_rf_gpr[496]), .B1(n16493), .Y(n14483) );
  sky130_fd_sc_hd__nand4_1 U21527 ( .A(n14486), .B(n14485), .C(n14484), .D(
        n14483), .Y(n14487) );
  sky130_fd_sc_hd__nand2_1 U21528 ( .A(n26285), .B(n16086), .Y(n14488) );
  sky130_fd_sc_hd__nor2_1 U21530 ( .A(n14577), .B(n14578), .Y(n21032) );
  sky130_fd_sc_hd__nand2_1 U21531 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[47]), .Y(n14492) );
  sky130_fd_sc_hd__nand2_1 U21532 ( .A(n16410), .B(
        j202_soc_core_j22_cpu_rf_gpr[175]), .Y(n14491) );
  sky130_fd_sc_hd__nand2_1 U21533 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[462]), .Y(n14490) );
  sky130_fd_sc_hd__nand2_1 U21534 ( .A(n11196), .B(
        j202_soc_core_j22_cpu_rf_gpr[366]), .Y(n14489) );
  sky130_fd_sc_hd__nand4_1 U21535 ( .A(n14492), .B(n14491), .C(n14490), .D(
        n14489), .Y(n14498) );
  sky130_fd_sc_hd__nand2_1 U21536 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[334]), .Y(n14496) );
  sky130_fd_sc_hd__nand2_1 U21537 ( .A(n11194), .B(
        j202_soc_core_j22_cpu_rf_gpr[303]), .Y(n14495) );
  sky130_fd_sc_hd__nand2_1 U21538 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[239]), .Y(n14494) );
  sky130_fd_sc_hd__nand2_1 U21539 ( .A(n15796), .B(
        j202_soc_core_j22_cpu_rf_gpr[79]), .Y(n14493) );
  sky130_fd_sc_hd__nand4_1 U21540 ( .A(n14496), .B(n14495), .C(n14494), .D(
        n14493), .Y(n14497) );
  sky130_fd_sc_hd__nor2_1 U21541 ( .A(n14498), .B(n14497), .Y(n14510) );
  sky130_fd_sc_hd__nand2_1 U21542 ( .A(n16433), .B(
        j202_soc_core_j22_cpu_rf_gpr[207]), .Y(n14502) );
  sky130_fd_sc_hd__nand2_1 U21543 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[430]), .Y(n14501) );
  sky130_fd_sc_hd__nand2_1 U21544 ( .A(n16398), .B(
        j202_soc_core_j22_cpu_rf_gpr[111]), .Y(n14500) );
  sky130_fd_sc_hd__nand2_1 U21545 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[271]), .Y(n14499) );
  sky130_fd_sc_hd__nor2_1 U21546 ( .A(n14564), .B(n14798), .Y(n14508) );
  sky130_fd_sc_hd__a21oi_1 U21547 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[15]), .B1(n14743), .Y(n14506) );
  sky130_fd_sc_hd__nand2_1 U21548 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[143]), .Y(n14505) );
  sky130_fd_sc_hd__nand2_1 U21549 ( .A(n14985), .B(
        j202_soc_core_j22_cpu_rf_gpr[494]), .Y(n14504) );
  sky130_fd_sc_hd__nand2_1 U21550 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[398]), .Y(n14503) );
  sky130_fd_sc_hd__nand4_1 U21551 ( .A(n14506), .B(n14505), .C(n14504), .D(
        n14503), .Y(n14507) );
  sky130_fd_sc_hd__nor2_1 U21552 ( .A(n14508), .B(n14507), .Y(n14509) );
  sky130_fd_sc_hd__inv_2 U21553 ( .A(n26064), .Y(n26430) );
  sky130_fd_sc_hd__nand2_1 U21555 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[208]), .Y(n14514) );
  sky130_fd_sc_hd__nand2_1 U21556 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[463]), .Y(n14513) );
  sky130_fd_sc_hd__nand2_1 U21557 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[495]), .Y(n14512) );
  sky130_fd_sc_hd__nand2_1 U21558 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[240]), .Y(n14511) );
  sky130_fd_sc_hd__nand4_1 U21559 ( .A(n14514), .B(n14513), .C(n14512), .D(
        n14511), .Y(n14520) );
  sky130_fd_sc_hd__nand2_1 U21560 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[16]), .Y(n14518) );
  sky130_fd_sc_hd__nand2_1 U21561 ( .A(n15984), .B(
        j202_soc_core_j22_cpu_rf_gpr[80]), .Y(n14517) );
  sky130_fd_sc_hd__nand2_1 U21562 ( .A(n16466), .B(
        j202_soc_core_j22_cpu_rf_gpr[399]), .Y(n14516) );
  sky130_fd_sc_hd__nand2_1 U21563 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[144]), .Y(n14515) );
  sky130_fd_sc_hd__nand4_1 U21564 ( .A(n14518), .B(n14517), .C(n14516), .D(
        n14515), .Y(n14519) );
  sky130_fd_sc_hd__nor2_1 U21565 ( .A(n14520), .B(n14519), .Y(n14532) );
  sky130_fd_sc_hd__nand2_1 U21566 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[272]), .Y(n14524) );
  sky130_fd_sc_hd__nand2_1 U21567 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[48]), .Y(n14523) );
  sky130_fd_sc_hd__nand2_1 U21568 ( .A(n15991), .B(
        j202_soc_core_j22_cpu_rf_gpr[367]), .Y(n14522) );
  sky130_fd_sc_hd__nand2_1 U21569 ( .A(n16064), .B(
        j202_soc_core_j22_cpu_rf_gpr[335]), .Y(n14521) );
  sky130_fd_sc_hd__and4_1 U21570 ( .A(n14524), .B(n14523), .C(n14522), .D(
        n14521), .X(n14531) );
  sky130_fd_sc_hd__nand2_1 U21571 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[304]), .Y(n14529) );
  sky130_fd_sc_hd__nand2_1 U21572 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[431]), .Y(n14528) );
  sky130_fd_sc_hd__nand2_1 U21573 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[176]), .Y(n14527) );
  sky130_fd_sc_hd__nand2_1 U21574 ( .A(n14525), .B(
        j202_soc_core_j22_cpu_rf_gpr[112]), .Y(n14526) );
  sky130_fd_sc_hd__and4_1 U21575 ( .A(n14529), .B(n14528), .C(n14527), .D(
        n14526), .X(n14530) );
  sky130_fd_sc_hd__nand3_1 U21576 ( .A(n14532), .B(n14531), .C(n14530), .Y(
        n22777) );
  sky130_fd_sc_hd__o22a_1 U21577 ( .A1(n14534), .A2(n16077), .B1(n14533), .B2(
        n14477), .X(n14540) );
  sky130_fd_sc_hd__o22a_1 U21578 ( .A1(n14535), .A2(n16491), .B1(n16487), .B2(
        n22769), .X(n14539) );
  sky130_fd_sc_hd__o22a_1 U21579 ( .A1(n14536), .A2(n16488), .B1(n16490), .B2(
        n22771), .X(n14538) );
  sky130_fd_sc_hd__a21oi_1 U21580 ( .A1(n11201), .A2(
        j202_soc_core_j22_cpu_rf_gpr[495]), .B1(n16493), .Y(n14537) );
  sky130_fd_sc_hd__nand4_1 U21581 ( .A(n14540), .B(n14539), .C(n14538), .D(
        n14537), .Y(n14541) );
  sky130_fd_sc_hd__mux2i_1 U21582 ( .A0(n16088), .A1(n16543), .S(n28532), .Y(
        n14576) );
  sky130_fd_sc_hd__o22ai_1 U21583 ( .A1(n16500), .A2(n26319), .B1(n26430), 
        .B2(n16501), .Y(n14573) );
  sky130_fd_sc_hd__nand2_1 U21584 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[207]), .Y(n14545) );
  sky130_fd_sc_hd__nand2_1 U21585 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[462]), .Y(n14544) );
  sky130_fd_sc_hd__nand2_1 U21586 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[494]), .Y(n14543) );
  sky130_fd_sc_hd__nand2_1 U21587 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[239]), .Y(n14542) );
  sky130_fd_sc_hd__nand4_1 U21588 ( .A(n14545), .B(n14544), .C(n14543), .D(
        n14542), .Y(n14551) );
  sky130_fd_sc_hd__nand2_1 U21589 ( .A(n16506), .B(
        j202_soc_core_j22_cpu_rf_gpr[15]), .Y(n14549) );
  sky130_fd_sc_hd__nand2_1 U21590 ( .A(n15984), .B(
        j202_soc_core_j22_cpu_rf_gpr[79]), .Y(n14548) );
  sky130_fd_sc_hd__nand2_1 U21591 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[398]), .Y(n14547) );
  sky130_fd_sc_hd__nand2_1 U21592 ( .A(n23808), .B(
        j202_soc_core_j22_cpu_rf_gpr[143]), .Y(n14546) );
  sky130_fd_sc_hd__nand4_1 U21593 ( .A(n14549), .B(n14548), .C(n14547), .D(
        n14546), .Y(n14550) );
  sky130_fd_sc_hd__nor2_1 U21594 ( .A(n14551), .B(n14550), .Y(n14562) );
  sky130_fd_sc_hd__nand2_1 U21595 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[271]), .Y(n14555) );
  sky130_fd_sc_hd__nand2_1 U21596 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[47]), .Y(n14554) );
  sky130_fd_sc_hd__nand2_1 U21597 ( .A(n15991), .B(
        j202_soc_core_j22_cpu_rf_gpr[366]), .Y(n14553) );
  sky130_fd_sc_hd__nand2_1 U21598 ( .A(n15017), .B(
        j202_soc_core_j22_cpu_rf_gpr[334]), .Y(n14552) );
  sky130_fd_sc_hd__and4_1 U21599 ( .A(n14555), .B(n14554), .C(n14553), .D(
        n14552), .X(n14561) );
  sky130_fd_sc_hd__nand2_1 U21600 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[303]), .Y(n14559) );
  sky130_fd_sc_hd__nand2_1 U21601 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[430]), .Y(n14558) );
  sky130_fd_sc_hd__nand2_1 U21602 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[175]), .Y(n14557) );
  sky130_fd_sc_hd__nand2_1 U21603 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[111]), .Y(n14556) );
  sky130_fd_sc_hd__and4_1 U21604 ( .A(n14559), .B(n14558), .C(n14557), .D(
        n14556), .X(n14560) );
  sky130_fd_sc_hd__nand3_1 U21605 ( .A(n14562), .B(n14561), .C(n14560), .Y(
        n18889) );
  sky130_fd_sc_hd__o22a_1 U21606 ( .A1(n18896), .A2(n15886), .B1(n18895), .B2(
        n14477), .X(n14569) );
  sky130_fd_sc_hd__o22a_1 U21607 ( .A1(n14564), .A2(n16488), .B1(n16487), .B2(
        n14563), .X(n14568) );
  sky130_fd_sc_hd__o22a_1 U21608 ( .A1(n18891), .A2(n16491), .B1(n16490), .B2(
        n14565), .X(n14567) );
  sky130_fd_sc_hd__a21oi_1 U21609 ( .A1(n11201), .A2(
        j202_soc_core_j22_cpu_rf_gpr[494]), .B1(n16493), .Y(n14566) );
  sky130_fd_sc_hd__nand4_1 U21610 ( .A(n14569), .B(n14568), .C(n14567), .D(
        n14566), .Y(n14570) );
  sky130_fd_sc_hd__nand2_1 U21611 ( .A(n26311), .B(n16086), .Y(n14571) );
  sky130_fd_sc_hd__o21ai_1 U21612 ( .A1(n16088), .A2(n26311), .B1(n14571), .Y(
        n14574) );
  sky130_fd_sc_hd__nor2_1 U21613 ( .A(n14573), .B(n14574), .Y(n20982) );
  sky130_fd_sc_hd__nor2_1 U21614 ( .A(n21032), .B(n14572), .Y(n14581) );
  sky130_fd_sc_hd__nand2_1 U21615 ( .A(n14574), .B(n14573), .Y(n20995) );
  sky130_fd_sc_hd__nand2_1 U21616 ( .A(n14576), .B(n14575), .Y(n20985) );
  sky130_fd_sc_hd__o21ai_2 U21617 ( .A1(n20995), .A2(n20984), .B1(n20985), .Y(
        n21029) );
  sky130_fd_sc_hd__nand2_1 U21618 ( .A(n14578), .B(n14577), .Y(n21033) );
  sky130_fd_sc_hd__o21ai_1 U21619 ( .A1(n21032), .A2(n14579), .B1(n21033), .Y(
        n14580) );
  sky130_fd_sc_hd__a21oi_1 U21620 ( .A1(n17040), .A2(n14581), .B1(n14580), .Y(
        n14587) );
  sky130_fd_sc_hd__o22ai_1 U21621 ( .A1(n16501), .A2(n27800), .B1(n26320), 
        .B2(n16500), .Y(n14583) );
  sky130_fd_sc_hd__nand2_1 U21622 ( .A(n28519), .B(n16541), .Y(n14582) );
  sky130_fd_sc_hd__nor2_1 U21624 ( .A(n14583), .B(n14584), .Y(n15069) );
  sky130_fd_sc_hd__nand2_1 U21625 ( .A(n14584), .B(n14583), .Y(n15068) );
  sky130_fd_sc_hd__nand2_1 U21626 ( .A(n14585), .B(n15068), .Y(n14586) );
  sky130_fd_sc_hd__xor2_1 U21627 ( .A(n14587), .B(n14586), .X(n25899) );
  sky130_fd_sc_hd__nor2_1 U21628 ( .A(n24034), .B(n14588), .Y(n14589) );
  sky130_fd_sc_hd__nand2_1 U21629 ( .A(n25899), .B(n17225), .Y(n17085) );
  sky130_fd_sc_hd__nand2_1 U21630 ( .A(n18764), .B(n19140), .Y(n14591) );
  sky130_fd_sc_hd__nand2_1 U21631 ( .A(n21101), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n17239) );
  sky130_fd_sc_hd__nand2_1 U21632 ( .A(n21104), .B(n20485), .Y(n14636) );
  sky130_fd_sc_hd__nor2_1 U21633 ( .A(n14591), .B(n14636), .Y(n14596) );
  sky130_fd_sc_hd__nand2_1 U21634 ( .A(n14596), .B(n21088), .Y(n16749) );
  sky130_fd_sc_hd__nor2_1 U21635 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n21145), .Y(n17242) );
  sky130_fd_sc_hd__nor2_1 U21636 ( .A(n20485), .B(n18697), .Y(n16757) );
  sky130_fd_sc_hd__nand2_1 U21637 ( .A(n16757), .B(n14592), .Y(n16274) );
  sky130_fd_sc_hd__nand2_1 U21638 ( .A(n16126), .B(n19130), .Y(n16742) );
  sky130_fd_sc_hd__nand3_1 U21639 ( .A(n13179), .B(n21145), .C(n13199), .Y(
        n14635) );
  sky130_fd_sc_hd__nand3_1 U21640 ( .A(n14621), .B(n18764), .C(n18744), .Y(
        n16266) );
  sky130_fd_sc_hd__nand3_1 U21641 ( .A(n16749), .B(n16742), .C(n16266), .Y(
        n14594) );
  sky130_fd_sc_hd__nand2_1 U21642 ( .A(n18764), .B(n21088), .Y(n21595) );
  sky130_fd_sc_hd__nor2_1 U21643 ( .A(n20485), .B(n21595), .Y(n19132) );
  sky130_fd_sc_hd__nand2_1 U21644 ( .A(n19132), .B(n21104), .Y(n16745) );
  sky130_fd_sc_hd__nor2_1 U21645 ( .A(n21088), .B(n18712), .Y(n21074) );
  sky130_fd_sc_hd__nand2_1 U21646 ( .A(n21074), .B(n18744), .Y(n14612) );
  sky130_fd_sc_hd__nand2_1 U21647 ( .A(n16764), .B(n14621), .Y(n16845) );
  sky130_fd_sc_hd__o21a_1 U21648 ( .A1(n19140), .A2(n16745), .B1(n16845), .X(
        n16259) );
  sky130_fd_sc_hd__nand3_1 U21650 ( .A(n20485), .B(n21145), .C(n21359), .Y(
        n14646) );
  sky130_fd_sc_hd__nand2_1 U21651 ( .A(n16764), .B(n16850), .Y(n16857) );
  sky130_fd_sc_hd__nand2_1 U21652 ( .A(n14596), .B(n19130), .Y(n14609) );
  sky130_fd_sc_hd__nand4_1 U21653 ( .A(n16259), .B(n16274), .C(n16857), .D(
        n14609), .Y(n14593) );
  sky130_fd_sc_hd__a22oi_1 U21654 ( .A1(n14594), .A2(n20368), .B1(n14593), 
        .B2(n20393), .Y(n14607) );
  sky130_fd_sc_hd__nand2_1 U21655 ( .A(n13199), .B(n21359), .Y(n14602) );
  sky130_fd_sc_hd__nand2b_1 U21656 ( .A_N(n14612), .B(n14595), .Y(n16740) );
  sky130_fd_sc_hd__nand2_1 U21657 ( .A(n16757), .B(n16764), .Y(n16746) );
  sky130_fd_sc_hd__nand3_1 U21658 ( .A(n16740), .B(n14706), .C(n16746), .Y(
        n14599) );
  sky130_fd_sc_hd__nor2_1 U21659 ( .A(n13199), .B(n21595), .Y(n20809) );
  sky130_fd_sc_hd__nand2_1 U21660 ( .A(n20809), .B(n17242), .Y(n16267) );
  sky130_fd_sc_hd__nor2_1 U21661 ( .A(n18744), .B(n21595), .Y(n14600) );
  sky130_fd_sc_hd__nand2_1 U21662 ( .A(n14600), .B(n16850), .Y(n16865) );
  sky130_fd_sc_hd__nand2_1 U21663 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .B(n19148), .Y(n16139) );
  sky130_fd_sc_hd__nand2_1 U21664 ( .A(n16207), .B(n16139), .Y(n19394) );
  sky130_fd_sc_hd__a21oi_1 U21665 ( .A1(n16267), .A2(n16865), .B1(n19394), .Y(
        n14598) );
  sky130_fd_sc_hd__a21oi_1 U21666 ( .A1(n14599), .A2(n20385), .B1(n14598), .Y(
        n14606) );
  sky130_fd_sc_hd__nor2_1 U21667 ( .A(n19140), .B(n21595), .Y(n16851) );
  sky130_fd_sc_hd__nand2_1 U21668 ( .A(n19132), .B(n15577), .Y(n16117) );
  sky130_fd_sc_hd__nand2b_1 U21669 ( .A_N(n16117), .B(n13179), .Y(n16846) );
  sky130_fd_sc_hd__nor2_1 U21670 ( .A(n18744), .B(n21132), .Y(n16747) );
  sky130_fd_sc_hd__nand3_1 U21671 ( .A(n20485), .B(n13179), .C(n21145), .Y(
        n14619) );
  sky130_fd_sc_hd__nand2_1 U21672 ( .A(n14600), .B(n14698), .Y(n16741) );
  sky130_fd_sc_hd__o21a_1 U21673 ( .A1(n14646), .A2(n16271), .B1(n16741), .X(
        n14703) );
  sky130_fd_sc_hd__o211ai_1 U21674 ( .A1(n14601), .A2(n14646), .B1(n16846), 
        .C1(n14703), .Y(n16113) );
  sky130_fd_sc_hd__nand2_1 U21675 ( .A(n16113), .B(n20374), .Y(n14605) );
  sky130_fd_sc_hd__nor2_1 U21676 ( .A(n20485), .B(n17239), .Y(n16763) );
  sky130_fd_sc_hd__nand2_1 U21677 ( .A(n16763), .B(n16747), .Y(n14694) );
  sky130_fd_sc_hd__nor2_1 U21678 ( .A(n21101), .B(n14602), .Y(n16161) );
  sky130_fd_sc_hd__nand2_1 U21679 ( .A(n16764), .B(n16161), .Y(n16858) );
  sky130_fd_sc_hd__nand2_1 U21680 ( .A(n14694), .B(n16858), .Y(n16125) );
  sky130_fd_sc_hd__nand2b_1 U21681 ( .A_N(n16117), .B(n21359), .Y(n16258) );
  sky130_fd_sc_hd__nand2_1 U21682 ( .A(n16747), .B(n14698), .Y(n16864) );
  sky130_fd_sc_hd__nand4b_1 U21683 ( .A_N(n16125), .B(n16258), .C(n16864), .D(
        n16746), .Y(n14603) );
  sky130_fd_sc_hd__nand2_1 U21684 ( .A(n14603), .B(n19394), .Y(n14604) );
  sky130_fd_sc_hd__nand4_1 U21685 ( .A(n14607), .B(n14606), .C(n14605), .D(
        n14604), .Y(n14618) );
  sky130_fd_sc_hd__nand2_1 U21686 ( .A(n16851), .B(n16161), .Y(n16275) );
  sky130_fd_sc_hd__nand2_1 U21687 ( .A(n21074), .B(n13199), .Y(n19145) );
  sky130_fd_sc_hd__nor2_1 U21688 ( .A(n15106), .B(n19145), .Y(n14610) );
  sky130_fd_sc_hd__nand2_1 U21689 ( .A(n14610), .B(n13179), .Y(n16859) );
  sky130_fd_sc_hd__nand2_1 U21690 ( .A(n20485), .B(n18744), .Y(n17007) );
  sky130_fd_sc_hd__nor2_1 U21691 ( .A(n18712), .B(n17007), .Y(n17156) );
  sky130_fd_sc_hd__nand2_1 U21692 ( .A(n17156), .B(n17242), .Y(n16268) );
  sky130_fd_sc_hd__nand2_1 U21693 ( .A(n16859), .B(n16268), .Y(n16761) );
  sky130_fd_sc_hd__nor2_1 U21694 ( .A(n14608), .B(n16761), .Y(n16260) );
  sky130_fd_sc_hd__nor2_1 U21695 ( .A(n13199), .B(n18744), .Y(n16994) );
  sky130_fd_sc_hd__nand3_1 U21696 ( .A(n16994), .B(n18764), .C(n17242), .Y(
        n16755) );
  sky130_fd_sc_hd__nor2_1 U21697 ( .A(n13199), .B(n18697), .Y(n14658) );
  sky130_fd_sc_hd__nand2_1 U21698 ( .A(n14658), .B(n16764), .Y(n16759) );
  sky130_fd_sc_hd__nand3_1 U21699 ( .A(n14609), .B(n16755), .C(n16759), .Y(
        n16277) );
  sky130_fd_sc_hd__a31oi_1 U21700 ( .A1(n16759), .A2(n16755), .A3(n16262), 
        .B1(n16207), .Y(n14611) );
  sky130_fd_sc_hd__a21oi_1 U21701 ( .A1(n16277), .A2(n20374), .B1(n14611), .Y(
        n14617) );
  sky130_fd_sc_hd__nand2_1 U21702 ( .A(n16851), .B(n14621), .Y(n16754) );
  sky130_fd_sc_hd__nand4b_1 U21703 ( .A_N(n16125), .B(n16859), .C(n16754), .D(
        n16746), .Y(n14615) );
  sky130_fd_sc_hd__nor2_1 U21704 ( .A(n14636), .B(n14612), .Y(n16782) );
  sky130_fd_sc_hd__nand2_1 U21705 ( .A(n14657), .B(n16851), .Y(n16842) );
  sky130_fd_sc_hd__nand3b_1 U21706 ( .A_N(n16782), .B(n16842), .C(n16268), .Y(
        n14613) );
  sky130_fd_sc_hd__nand2_1 U21707 ( .A(n20809), .B(n16205), .Y(n16756) );
  sky130_fd_sc_hd__nand2b_1 U21708 ( .A_N(n16756), .B(n13179), .Y(n16204) );
  sky130_fd_sc_hd__nand2_1 U21709 ( .A(n16749), .B(n16204), .Y(n14702) );
  sky130_fd_sc_hd__nor2_1 U21710 ( .A(n14613), .B(n14702), .Y(n16264) );
  sky130_fd_sc_hd__nand2b_1 U21711 ( .A_N(n16745), .B(n19140), .Y(n14614) );
  sky130_fd_sc_hd__nand2_1 U21712 ( .A(n16264), .B(n14614), .Y(n16743) );
  sky130_fd_sc_hd__o211ai_1 U21714 ( .A1(n16260), .A2(n16206), .B1(n14617), 
        .C1(n14616), .Y(n16129) );
  sky130_fd_sc_hd__nor2_1 U21715 ( .A(n11150), .B(
        j202_soc_core_bootrom_00_address_w[8]), .Y(n16770) );
  sky130_fd_sc_hd__nand2_1 U21717 ( .A(n18712), .B(n21088), .Y(n19125) );
  sky130_fd_sc_hd__nor2_1 U21718 ( .A(n19140), .B(n19125), .Y(n14665) );
  sky130_fd_sc_hd__nand2_1 U21719 ( .A(n14665), .B(n16161), .Y(n16785) );
  sky130_fd_sc_hd__nor2_1 U21720 ( .A(n18744), .B(n19125), .Y(n14677) );
  sky130_fd_sc_hd__nand2_1 U21721 ( .A(n14677), .B(n14698), .Y(n16809) );
  sky130_fd_sc_hd__nand2_1 U21722 ( .A(n16785), .B(n16809), .Y(n16831) );
  sky130_fd_sc_hd__nor2_4 U21723 ( .A(n21088), .B(n18764), .Y(n17251) );
  sky130_fd_sc_hd__nand2_1 U21724 ( .A(n17251), .B(n19140), .Y(n16135) );
  sky130_fd_sc_hd__nor2_1 U21725 ( .A(n14619), .B(n16135), .Y(n16149) );
  sky130_fd_sc_hd__nand2_1 U21726 ( .A(n14677), .B(n16850), .Y(n16246) );
  sky130_fd_sc_hd__nor2_1 U21727 ( .A(n16149), .B(n14620), .Y(n14622) );
  sky130_fd_sc_hd__nand3_1 U21728 ( .A(n20303), .B(n19140), .C(n17242), .Y(
        n16827) );
  sky130_fd_sc_hd__nand2_1 U21729 ( .A(n14677), .B(n14621), .Y(n16823) );
  sky130_fd_sc_hd__nand4_1 U21730 ( .A(n14641), .B(n14622), .C(n16827), .D(
        n16823), .Y(n14627) );
  sky130_fd_sc_hd__nand2_1 U21731 ( .A(n14677), .B(n14657), .Y(n14642) );
  sky130_fd_sc_hd__nand2_1 U21732 ( .A(n14698), .B(n16160), .Y(n16776) );
  sky130_fd_sc_hd__nor2_1 U21733 ( .A(n19130), .B(n16776), .Y(n14647) );
  sky130_fd_sc_hd__nor2_1 U21734 ( .A(n14623), .B(n14647), .Y(n16227) );
  sky130_fd_sc_hd__nor2_1 U21735 ( .A(n14635), .B(n14632), .Y(n16226) );
  sky130_fd_sc_hd__nand2_1 U21736 ( .A(n14665), .B(n16763), .Y(n16154) );
  sky130_fd_sc_hd__nand3_1 U21737 ( .A(n16227), .B(n16775), .C(n16154), .Y(
        n16223) );
  sky130_fd_sc_hd__nand2_1 U21738 ( .A(n14677), .B(n16161), .Y(n14678) );
  sky130_fd_sc_hd__nand2_1 U21739 ( .A(n14658), .B(n14677), .Y(n16816) );
  sky130_fd_sc_hd__nand2_1 U21740 ( .A(n16161), .B(n17251), .Y(n14624) );
  sky130_fd_sc_hd__nand2_1 U21741 ( .A(n16816), .B(n14624), .Y(n16240) );
  sky130_fd_sc_hd__nand2b_1 U21742 ( .A_N(n14636), .B(n14665), .Y(n14656) );
  sky130_fd_sc_hd__nand2_1 U21743 ( .A(n16757), .B(n14665), .Y(n16242) );
  sky130_fd_sc_hd__nand2_1 U21744 ( .A(n14656), .B(n16242), .Y(n14650) );
  sky130_fd_sc_hd__nor3_1 U21745 ( .A(n16803), .B(n16240), .C(n14650), .Y(
        n14625) );
  sky130_fd_sc_hd__nand2_1 U21746 ( .A(n14626), .B(n14625), .Y(n16133) );
  sky130_fd_sc_hd__o21ai_1 U21747 ( .A1(n14627), .A2(n16133), .B1(n20393), .Y(
        n14663) );
  sky130_fd_sc_hd__nand2_1 U21748 ( .A(n17251), .B(n18744), .Y(n16820) );
  sky130_fd_sc_hd__nor2_1 U21749 ( .A(n14628), .B(n16820), .Y(n14667) );
  sky130_fd_sc_hd__nand2_1 U21750 ( .A(n14629), .B(n14642), .Y(n14630) );
  sky130_fd_sc_hd__nand2_1 U21751 ( .A(n16226), .B(n21088), .Y(n16243) );
  sky130_fd_sc_hd__nand4b_1 U21752 ( .A_N(n14630), .B(n16842), .C(n16154), .D(
        n16243), .Y(n14634) );
  sky130_fd_sc_hd__nor2_1 U21753 ( .A(n16149), .B(n14631), .Y(n16229) );
  sky130_fd_sc_hd__nor2_1 U21754 ( .A(n14646), .B(n14632), .Y(n14686) );
  sky130_fd_sc_hd__nand2_1 U21755 ( .A(n14686), .B(n21088), .Y(n14633) );
  sky130_fd_sc_hd__nand2_1 U21756 ( .A(n16229), .B(n14633), .Y(n16238) );
  sky130_fd_sc_hd__nor2_1 U21757 ( .A(n14634), .B(n16238), .Y(n16774) );
  sky130_fd_sc_hd__nor2_1 U21758 ( .A(n14635), .B(n16135), .Y(n16780) );
  sky130_fd_sc_hd__nor2_1 U21759 ( .A(n16780), .B(n16803), .Y(n14664) );
  sky130_fd_sc_hd__nand2_1 U21760 ( .A(n14656), .B(n14664), .Y(n14637) );
  sky130_fd_sc_hd__nand2b_1 U21761 ( .A_N(n14636), .B(n17251), .Y(n16221) );
  sky130_fd_sc_hd__nand2_1 U21762 ( .A(n16221), .B(n16816), .Y(n16158) );
  sky130_fd_sc_hd__nor3_1 U21763 ( .A(n16782), .B(n14637), .C(n16158), .Y(
        n14638) );
  sky130_fd_sc_hd__nand2_1 U21764 ( .A(n16774), .B(n14638), .Y(n14639) );
  sky130_fd_sc_hd__nand2_1 U21765 ( .A(n14639), .B(n20385), .Y(n14662) );
  sky130_fd_sc_hd__nor2_1 U21766 ( .A(n16149), .B(n16782), .Y(n14640) );
  sky130_fd_sc_hd__nand4_1 U21767 ( .A(n14641), .B(n14640), .C(n16827), .D(
        n14642), .Y(n14653) );
  sky130_fd_sc_hd__nand2b_1 U21768 ( .A_N(n16135), .B(n16763), .Y(n14654) );
  sky130_fd_sc_hd__nand2_1 U21769 ( .A(n16140), .B(n19130), .Y(n14668) );
  sky130_fd_sc_hd__nor2_1 U21770 ( .A(n20485), .B(n16820), .Y(n17101) );
  sky130_fd_sc_hd__nand2_1 U21771 ( .A(n17101), .B(n21101), .Y(n16828) );
  sky130_fd_sc_hd__nand3_1 U21772 ( .A(n14668), .B(n16828), .C(n14642), .Y(
        n16814) );
  sky130_fd_sc_hd__nor2_1 U21773 ( .A(n14644), .B(n14643), .Y(n16808) );
  sky130_fd_sc_hd__nand2_1 U21774 ( .A(n14682), .B(n14657), .Y(n16150) );
  sky130_fd_sc_hd__nand2_1 U21775 ( .A(n14682), .B(n17242), .Y(n14645) );
  sky130_fd_sc_hd__nand2_1 U21776 ( .A(n16150), .B(n14645), .Y(n16788) );
  sky130_fd_sc_hd__nor2_1 U21777 ( .A(n16808), .B(n16788), .Y(n16834) );
  sky130_fd_sc_hd__nor2_1 U21778 ( .A(n14646), .B(n16135), .Y(n16167) );
  sky130_fd_sc_hd__nor2_1 U21779 ( .A(n16167), .B(n14647), .Y(n14648) );
  sky130_fd_sc_hd__nand3_1 U21780 ( .A(n14649), .B(n16834), .C(n14648), .Y(
        n16220) );
  sky130_fd_sc_hd__nor4_1 U21781 ( .A(n16149), .B(n14686), .C(n14650), .D(
        n16220), .Y(n14651) );
  sky130_fd_sc_hd__a21oi_1 U21782 ( .A1(n14654), .A2(n14651), .B1(n16139), .Y(
        n14652) );
  sky130_fd_sc_hd__a21oi_1 U21783 ( .A1(n14653), .A2(n20368), .B1(n14652), .Y(
        n16144) );
  sky130_fd_sc_hd__nand2_1 U21784 ( .A(n16757), .B(n14677), .Y(n14684) );
  sky130_fd_sc_hd__nand2_1 U21785 ( .A(n14654), .B(n14684), .Y(n16216) );
  sky130_fd_sc_hd__nand2_1 U21786 ( .A(n14655), .B(n16154), .Y(n16162) );
  sky130_fd_sc_hd__nand2_1 U21787 ( .A(n14676), .B(n14657), .Y(n16826) );
  sky130_fd_sc_hd__nand2_1 U21788 ( .A(n14658), .B(n16160), .Y(n16789) );
  sky130_fd_sc_hd__nand4b_1 U21789 ( .A_N(n16780), .B(n16784), .C(n16826), .D(
        n16789), .Y(n16239) );
  sky130_fd_sc_hd__nor2_1 U21790 ( .A(n16162), .B(n16239), .Y(n14660) );
  sky130_fd_sc_hd__nor2_1 U21791 ( .A(n18697), .B(n16820), .Y(n16166) );
  sky130_fd_sc_hd__nand2_1 U21792 ( .A(n16166), .B(n20485), .Y(n16818) );
  sky130_fd_sc_hd__nand2_1 U21793 ( .A(n16818), .B(n16246), .Y(n16241) );
  sky130_fd_sc_hd__nor2_1 U21794 ( .A(n16247), .B(n16241), .Y(n14659) );
  sky130_fd_sc_hd__o22a_1 U21795 ( .A1(n16207), .A2(n14660), .B1(n16139), .B2(
        n14659), .X(n14661) );
  sky130_fd_sc_hd__nand4_1 U21796 ( .A(n14663), .B(n14662), .C(n16144), .D(
        n14661), .Y(n14693) );
  sky130_fd_sc_hd__nor2_1 U21797 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .B(n13182), .Y(n16801) );
  sky130_fd_sc_hd__nand2b_1 U21798 ( .A_N(n16149), .B(n14664), .Y(n16786) );
  sky130_fd_sc_hd__nor2_1 U21799 ( .A(n16831), .B(n16786), .Y(n14670) );
  sky130_fd_sc_hd__nand2_1 U21800 ( .A(n14686), .B(n19130), .Y(n16792) );
  sky130_fd_sc_hd__o21a_1 U21801 ( .A1(n18697), .A2(n14666), .B1(n16792), .X(
        n16147) );
  sky130_fd_sc_hd__nor2_1 U21802 ( .A(n16167), .B(n14667), .Y(n14669) );
  sky130_fd_sc_hd__nand4_1 U21803 ( .A(n14670), .B(n16147), .C(n14669), .D(
        n14668), .Y(n14671) );
  sky130_fd_sc_hd__nor2_1 U21805 ( .A(n16808), .B(n14672), .Y(n14675) );
  sky130_fd_sc_hd__nor2_1 U21806 ( .A(n13199), .B(n19125), .Y(n19143) );
  sky130_fd_sc_hd__nand2_1 U21807 ( .A(n19143), .B(n15516), .Y(n16778) );
  sky130_fd_sc_hd__nand2_1 U21808 ( .A(n14673), .B(n16778), .Y(n16832) );
  sky130_fd_sc_hd__nand4_1 U21809 ( .A(n14675), .B(n14674), .C(n16826), .D(
        n16823), .Y(n14681) );
  sky130_fd_sc_hd__a31oi_1 U21811 ( .A1(n14679), .A2(n16809), .A3(n14678), 
        .B1(n17102), .Y(n14680) );
  sky130_fd_sc_hd__a21oi_1 U21812 ( .A1(n14681), .A2(n20385), .B1(n14680), .Y(
        n14690) );
  sky130_fd_sc_hd__nand2_1 U21813 ( .A(n14682), .B(n16757), .Y(n16214) );
  sky130_fd_sc_hd__nand3_1 U21814 ( .A(n16243), .B(n16816), .C(n16214), .Y(
        n14683) );
  sky130_fd_sc_hd__nor2_1 U21815 ( .A(n14683), .B(n16239), .Y(n16153) );
  sky130_fd_sc_hd__nor2_1 U21816 ( .A(n16167), .B(n14685), .Y(n16249) );
  sky130_fd_sc_hd__nand2_1 U21817 ( .A(n16763), .B(n17251), .Y(n16131) );
  sky130_fd_sc_hd__nor2b_1 U21818 ( .B_N(n16131), .A(n14686), .Y(n14687) );
  sky130_fd_sc_hd__nand4_1 U21819 ( .A(n16153), .B(n16249), .C(n14687), .D(
        n16785), .Y(n14688) );
  sky130_fd_sc_hd__nand2_1 U21820 ( .A(n14688), .B(n20374), .Y(n14689) );
  sky130_fd_sc_hd__nand2_1 U21821 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .B(n11150), .Y(n16255) );
  sky130_fd_sc_hd__a31oi_1 U21822 ( .A1(n14691), .A2(n14690), .A3(n14689), 
        .B1(n16255), .Y(n14692) );
  sky130_fd_sc_hd__a21oi_1 U21823 ( .A1(n14693), .A2(n16801), .B1(n14692), .Y(
        n14719) );
  sky130_fd_sc_hd__nand2_1 U21824 ( .A(n16756), .B(n16741), .Y(n16273) );
  sky130_fd_sc_hd__nand3_1 U21825 ( .A(n16745), .B(n16754), .C(n16755), .Y(
        n14695) );
  sky130_fd_sc_hd__nand2_1 U21826 ( .A(n16742), .B(n14694), .Y(n16124) );
  sky130_fd_sc_hd__nor2_1 U21827 ( .A(n14695), .B(n16124), .Y(n16866) );
  sky130_fd_sc_hd__nand2_1 U21828 ( .A(n16866), .B(n16746), .Y(n16112) );
  sky130_fd_sc_hd__o31a_1 U21829 ( .A1(n16116), .A2(n16273), .A3(n16112), .B1(
        n20368), .X(n14717) );
  sky130_fd_sc_hd__nor2_1 U21830 ( .A(n19140), .B(n16267), .Y(n14697) );
  sky130_fd_sc_hd__nor2_1 U21831 ( .A(n14697), .B(n14696), .Y(n16211) );
  sky130_fd_sc_hd__nand2_1 U21832 ( .A(n16764), .B(n14698), .Y(n16263) );
  sky130_fd_sc_hd__nand2_1 U21833 ( .A(n16263), .B(n16865), .Y(n14699) );
  sky130_fd_sc_hd__nor2_1 U21834 ( .A(n14700), .B(n14699), .Y(n14701) );
  sky130_fd_sc_hd__nand3b_1 U21835 ( .A_N(n14702), .B(n16211), .C(n14701), .Y(
        n14712) );
  sky130_fd_sc_hd__nand3_1 U21836 ( .A(n16749), .B(n14703), .C(n16275), .Y(
        n14704) );
  sky130_fd_sc_hd__nand2_1 U21837 ( .A(n14704), .B(n20385), .Y(n14710) );
  sky130_fd_sc_hd__nand2_1 U21838 ( .A(n14705), .B(n19130), .Y(n14707) );
  sky130_fd_sc_hd__nand4_1 U21839 ( .A(n14707), .B(n14706), .C(n16263), .D(
        n16858), .Y(n14708) );
  sky130_fd_sc_hd__nand2_1 U21840 ( .A(n14708), .B(n20393), .Y(n14709) );
  sky130_fd_sc_hd__nand2_1 U21841 ( .A(n14710), .B(n14709), .Y(n14711) );
  sky130_fd_sc_hd__a21oi_1 U21842 ( .A1(n14712), .A2(n20374), .B1(n14711), .Y(
        n16870) );
  sky130_fd_sc_hd__nand2_1 U21843 ( .A(n16267), .B(n16745), .Y(n14713) );
  sky130_fd_sc_hd__nand2_1 U21844 ( .A(n14713), .B(n18744), .Y(n16856) );
  sky130_fd_sc_hd__nand3_1 U21845 ( .A(n16856), .B(n16842), .C(n16741), .Y(
        n14715) );
  sky130_fd_sc_hd__a21oi_1 U21846 ( .A1(n16267), .A2(n16117), .B1(n16206), .Y(
        n14714) );
  sky130_fd_sc_hd__a21oi_1 U21847 ( .A1(n14715), .A2(n20393), .B1(n14714), .Y(
        n14716) );
  sky130_fd_sc_hd__nand2_1 U21848 ( .A(n16870), .B(n14716), .Y(n16122) );
  sky130_fd_sc_hd__nor2_1 U21849 ( .A(n11150), .B(n17264), .Y(n16871) );
  sky130_fd_sc_hd__o21ai_1 U21850 ( .A1(n14717), .A2(n16122), .B1(n16871), .Y(
        n14718) );
  sky130_fd_sc_hd__nand3_1 U21851 ( .A(n14720), .B(n14719), .C(n14718), .Y(
        n14721) );
  sky130_fd_sc_hd__nand2_1 U21852 ( .A(n14721), .B(n21629), .Y(n14724) );
  sky130_fd_sc_hd__a22oi_1 U21853 ( .A1(n21516), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[24]), .B1(n20759), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[88]), .Y(n14723) );
  sky130_fd_sc_hd__a22oi_1 U21854 ( .A1(n20540), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[56]), .B1(n21513), .B2(
        j202_soc_core_uart_div0[0]), .Y(n14722) );
  sky130_fd_sc_hd__nand3_1 U21855 ( .A(n14724), .B(n14723), .C(n14722), .Y(
        n14725) );
  sky130_fd_sc_hd__a21oi_1 U21856 ( .A1(j202_soc_core_memory0_ram_dout0[504]), 
        .A2(n11207), .B1(n14725), .Y(n14727) );
  sky130_fd_sc_hd__nand2_1 U21857 ( .A(j202_soc_core_memory0_ram_dout0[88]), 
        .B(n20458), .Y(n14726) );
  sky130_fd_sc_hd__nand2_1 U21858 ( .A(n21020), .B(n21768), .Y(n16294) );
  sky130_fd_sc_hd__nand2_1 U21859 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[56]), .Y(n14731) );
  sky130_fd_sc_hd__nand2_1 U21860 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[248]), .Y(n14730) );
  sky130_fd_sc_hd__nand2_1 U21861 ( .A(n11195), .B(
        j202_soc_core_j22_cpu_rf_gpr[407]), .Y(n14729) );
  sky130_fd_sc_hd__nand2_1 U21862 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[375]), .Y(n14728) );
  sky130_fd_sc_hd__nand4_1 U21863 ( .A(n14731), .B(n14730), .C(n14729), .D(
        n14728), .Y(n14737) );
  sky130_fd_sc_hd__nand2_1 U21864 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[343]), .Y(n14735) );
  sky130_fd_sc_hd__nand2_1 U21865 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[184]), .Y(n14734) );
  sky130_fd_sc_hd__nand2_1 U21866 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[439]), .Y(n14733) );
  sky130_fd_sc_hd__nand2_1 U21867 ( .A(n15788), .B(
        j202_soc_core_j22_cpu_rf_gpr[471]), .Y(n14732) );
  sky130_fd_sc_hd__nand4_1 U21868 ( .A(n14735), .B(n14734), .C(n14733), .D(
        n14732), .Y(n14736) );
  sky130_fd_sc_hd__nor2_1 U21869 ( .A(n14737), .B(n14736), .Y(n14752) );
  sky130_fd_sc_hd__nand2_1 U21870 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[312]), .Y(n14741) );
  sky130_fd_sc_hd__nand2_1 U21871 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[216]), .Y(n14740) );
  sky130_fd_sc_hd__nand2_1 U21872 ( .A(n16398), .B(
        j202_soc_core_j22_cpu_rf_gpr[120]), .Y(n14739) );
  sky130_fd_sc_hd__nand2_1 U21873 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[280]), .Y(n14738) );
  sky130_fd_sc_hd__and4_1 U21874 ( .A(n14741), .B(n14740), .C(n14739), .D(
        n14738), .X(n14751) );
  sky130_fd_sc_hd__nor2_1 U21875 ( .A(n14742), .B(n14798), .Y(n14749) );
  sky130_fd_sc_hd__a21oi_1 U21876 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[24]), .B1(n14743), .Y(n14747) );
  sky130_fd_sc_hd__nand2_1 U21877 ( .A(n16425), .B(
        j202_soc_core_j22_cpu_rf_gpr[152]), .Y(n14746) );
  sky130_fd_sc_hd__nand2_1 U21878 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[503]), .Y(n14745) );
  sky130_fd_sc_hd__nand2_1 U21879 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[88]), .Y(n14744) );
  sky130_fd_sc_hd__nand4_1 U21880 ( .A(n14747), .B(n14746), .C(n14745), .D(
        n14744), .Y(n14748) );
  sky130_fd_sc_hd__nor2_1 U21881 ( .A(n14749), .B(n14748), .Y(n14750) );
  sky130_fd_sc_hd__nand2_1 U21882 ( .A(j202_soc_core_j22_cpu_pc[19]), .B(
        j202_soc_core_j22_cpu_pc[20]), .Y(n14753) );
  sky130_fd_sc_hd__nand2_1 U21883 ( .A(j202_soc_core_j22_cpu_pc[17]), .B(
        j202_soc_core_j22_cpu_pc[18]), .Y(n15376) );
  sky130_fd_sc_hd__nor2_1 U21884 ( .A(n14753), .B(n15376), .Y(n15175) );
  sky130_fd_sc_hd__nand2_1 U21885 ( .A(j202_soc_core_j22_cpu_pc[21]), .B(
        j202_soc_core_j22_cpu_pc[22]), .Y(n15258) );
  sky130_fd_sc_hd__nor2_1 U21886 ( .A(n15260), .B(n15258), .Y(n14754) );
  sky130_fd_sc_hd__nand2_1 U21887 ( .A(n15175), .B(n14754), .Y(n16094) );
  sky130_fd_sc_hd__nor2_1 U21888 ( .A(n16094), .B(n21026), .Y(n14755) );
  sky130_fd_sc_hd__xnor2_1 U21889 ( .A(n22725), .B(n14755), .Y(n26455) );
  sky130_fd_sc_hd__nand2_1 U21890 ( .A(n22747), .B(n26455), .Y(n14787) );
  sky130_fd_sc_hd__nand2_1 U21891 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[216]), .Y(n14759) );
  sky130_fd_sc_hd__nand2_1 U21892 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[471]), .Y(n14758) );
  sky130_fd_sc_hd__nand2_1 U21893 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[503]), .Y(n14757) );
  sky130_fd_sc_hd__nand2_1 U21894 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[248]), .Y(n14756) );
  sky130_fd_sc_hd__nand4_1 U21895 ( .A(n14759), .B(n14758), .C(n14757), .D(
        n14756), .Y(n14765) );
  sky130_fd_sc_hd__nand2_1 U21896 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[24]), .Y(n14763) );
  sky130_fd_sc_hd__nand2_1 U21897 ( .A(n15984), .B(
        j202_soc_core_j22_cpu_rf_gpr[88]), .Y(n14762) );
  sky130_fd_sc_hd__nand2_1 U21898 ( .A(n16466), .B(
        j202_soc_core_j22_cpu_rf_gpr[407]), .Y(n14761) );
  sky130_fd_sc_hd__nand2_1 U21899 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[152]), .Y(n14760) );
  sky130_fd_sc_hd__nand4_1 U21900 ( .A(n14763), .B(n14762), .C(n14761), .D(
        n14760), .Y(n14764) );
  sky130_fd_sc_hd__nor2_1 U21901 ( .A(n14765), .B(n14764), .Y(n14773) );
  sky130_fd_sc_hd__a22oi_1 U21902 ( .A1(n23776), .A2(
        j202_soc_core_j22_cpu_rf_gpr[375]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[280]), .Y(n14772) );
  sky130_fd_sc_hd__a22oi_1 U21903 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[56]), .B1(n15017), .B2(
        j202_soc_core_j22_cpu_rf_gpr[343]), .Y(n14771) );
  sky130_fd_sc_hd__nand2_1 U21904 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[312]), .Y(n14769) );
  sky130_fd_sc_hd__nand2_1 U21905 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[439]), .Y(n14768) );
  sky130_fd_sc_hd__nand2_1 U21906 ( .A(n11199), .B(
        j202_soc_core_j22_cpu_rf_gpr[184]), .Y(n14767) );
  sky130_fd_sc_hd__nand2_1 U21907 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[120]), .Y(n14766) );
  sky130_fd_sc_hd__and4_1 U21908 ( .A(n14769), .B(n14768), .C(n14767), .D(
        n14766), .X(n14770) );
  sky130_fd_sc_hd__nand4_1 U21909 ( .A(n14773), .B(n14772), .C(n14771), .D(
        n14770), .Y(n22730) );
  sky130_fd_sc_hd__nand2_1 U21910 ( .A(n22730), .B(n16523), .Y(n14785) );
  sky130_fd_sc_hd__o21ai_0 U21911 ( .A1(n14774), .A2(n16525), .B1(n16524), .Y(
        n14779) );
  sky130_fd_sc_hd__o22ai_1 U21912 ( .A1(n14777), .A2(n11202), .B1(n14776), 
        .B2(n14477), .Y(n14778) );
  sky130_fd_sc_hd__nor2_1 U21913 ( .A(n14779), .B(n14778), .Y(n14784) );
  sky130_fd_sc_hd__nand2_1 U21914 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[24]), .Y(n14783) );
  sky130_fd_sc_hd__nand2_1 U21915 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[24]), .Y(n14782) );
  sky130_fd_sc_hd__nand2_1 U21916 ( .A(n16533), .B(
        j202_soc_core_j22_cpu_pc[24]), .Y(n14781) );
  sky130_fd_sc_hd__nand2_1 U21917 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[24]), .Y(n14780) );
  sky130_fd_sc_hd__nand2_1 U21918 ( .A(n21924), .B(n24929), .Y(n14786) );
  sky130_fd_sc_hd__nand2_1 U21920 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[438]), .Y(n14791) );
  sky130_fd_sc_hd__nand2_1 U21921 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[279]), .Y(n14790) );
  sky130_fd_sc_hd__nand2_1 U21922 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[406]), .Y(n14789) );
  sky130_fd_sc_hd__nand2_1 U21923 ( .A(n16398), .B(
        j202_soc_core_j22_cpu_rf_gpr[119]), .Y(n14788) );
  sky130_fd_sc_hd__nand4_1 U21924 ( .A(n14791), .B(n14790), .C(n14789), .D(
        n14788), .Y(n14797) );
  sky130_fd_sc_hd__nand2_1 U21925 ( .A(n16433), .B(
        j202_soc_core_j22_cpu_rf_gpr[215]), .Y(n14795) );
  sky130_fd_sc_hd__nand2_1 U21926 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[151]), .Y(n14794) );
  sky130_fd_sc_hd__nand2_1 U21927 ( .A(n14985), .B(
        j202_soc_core_j22_cpu_rf_gpr[502]), .Y(n14793) );
  sky130_fd_sc_hd__nand2_1 U21928 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[247]), .Y(n14792) );
  sky130_fd_sc_hd__nand4_1 U21929 ( .A(n14795), .B(n14794), .C(n14793), .D(
        n14792), .Y(n14796) );
  sky130_fd_sc_hd__nor2_1 U21930 ( .A(n14797), .B(n14796), .Y(n14812) );
  sky130_fd_sc_hd__nor2_1 U21931 ( .A(n14799), .B(n14798), .Y(n14805) );
  sky130_fd_sc_hd__a21oi_1 U21932 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[23]), .B1(n14743), .Y(n14803) );
  sky130_fd_sc_hd__nand2_1 U21933 ( .A(n11194), .B(
        j202_soc_core_j22_cpu_rf_gpr[311]), .Y(n14802) );
  sky130_fd_sc_hd__nand2_1 U21934 ( .A(n15796), .B(
        j202_soc_core_j22_cpu_rf_gpr[87]), .Y(n14801) );
  sky130_fd_sc_hd__nand2_1 U21935 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[55]), .Y(n14800) );
  sky130_fd_sc_hd__nand4_1 U21936 ( .A(n14803), .B(n14802), .C(n14801), .D(
        n14800), .Y(n14804) );
  sky130_fd_sc_hd__nor2_1 U21937 ( .A(n14805), .B(n14804), .Y(n14811) );
  sky130_fd_sc_hd__nand2_1 U21938 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[183]), .Y(n14809) );
  sky130_fd_sc_hd__nand2_1 U21939 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[342]), .Y(n14808) );
  sky130_fd_sc_hd__nand2_1 U21940 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[374]), .Y(n14807) );
  sky130_fd_sc_hd__nand2_1 U21941 ( .A(n15788), .B(
        j202_soc_core_j22_cpu_rf_gpr[470]), .Y(n14806) );
  sky130_fd_sc_hd__and4_1 U21942 ( .A(n14809), .B(n14808), .C(n14807), .D(
        n14806), .X(n14810) );
  sky130_fd_sc_hd__o22ai_1 U21943 ( .A1(n16500), .A2(n26431), .B1(n26323), 
        .B2(n16501), .Y(n14814) );
  sky130_fd_sc_hd__nand2_1 U21944 ( .A(n24929), .B(n16541), .Y(n14813) );
  sky130_fd_sc_hd__o21ai_1 U21945 ( .A1(n16543), .A2(n24929), .B1(n14813), .Y(
        n14815) );
  sky130_fd_sc_hd__nor2_1 U21946 ( .A(n14814), .B(n14815), .Y(n16013) );
  sky130_fd_sc_hd__nand2_1 U21947 ( .A(n14815), .B(n14814), .Y(n16012) );
  sky130_fd_sc_hd__nand2_1 U21948 ( .A(n14816), .B(n16012), .Y(n15089) );
  sky130_fd_sc_hd__nand2_1 U21949 ( .A(n16425), .B(
        j202_soc_core_j22_cpu_rf_gpr[150]), .Y(n14820) );
  sky130_fd_sc_hd__nand2_1 U21950 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[86]), .Y(n14819) );
  sky130_fd_sc_hd__nand2_1 U21951 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[405]), .Y(n14818) );
  sky130_fd_sc_hd__nand2_1 U21952 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[373]), .Y(n14817) );
  sky130_fd_sc_hd__nand4_1 U21953 ( .A(n14820), .B(n14819), .C(n14818), .D(
        n14817), .Y(n14827) );
  sky130_fd_sc_hd__nand2_1 U21954 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[278]), .Y(n14825) );
  sky130_fd_sc_hd__nand2_1 U21955 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[310]), .Y(n14824) );
  sky130_fd_sc_hd__nand2_1 U21956 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[469]), .Y(n14823) );
  sky130_fd_sc_hd__nand2_1 U21957 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[437]), .Y(n14822) );
  sky130_fd_sc_hd__nand4_1 U21958 ( .A(n14825), .B(n14824), .C(n14823), .D(
        n14822), .Y(n14826) );
  sky130_fd_sc_hd__nor2_1 U21959 ( .A(n14827), .B(n14826), .Y(n14842) );
  sky130_fd_sc_hd__nand2_1 U21960 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[341]), .Y(n14832) );
  sky130_fd_sc_hd__nand2_1 U21961 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[182]), .Y(n14831) );
  sky130_fd_sc_hd__nand2_1 U21962 ( .A(n16398), .B(
        j202_soc_core_j22_cpu_rf_gpr[118]), .Y(n14830) );
  sky130_fd_sc_hd__nand2_1 U21963 ( .A(n16433), .B(
        j202_soc_core_j22_cpu_rf_gpr[214]), .Y(n14829) );
  sky130_fd_sc_hd__nor2_1 U21964 ( .A(n14834), .B(n16444), .Y(n14840) );
  sky130_fd_sc_hd__a21oi_1 U21965 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[22]), .B1(n14743), .Y(n14838) );
  sky130_fd_sc_hd__nand2_1 U21966 ( .A(n16043), .B(
        j202_soc_core_j22_cpu_rf_gpr[246]), .Y(n14837) );
  sky130_fd_sc_hd__nand2_1 U21967 ( .A(n14985), .B(
        j202_soc_core_j22_cpu_rf_gpr[501]), .Y(n14836) );
  sky130_fd_sc_hd__nand2_1 U21968 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[54]), .Y(n14835) );
  sky130_fd_sc_hd__nand4_1 U21969 ( .A(n14838), .B(n14837), .C(n14836), .D(
        n14835), .Y(n14839) );
  sky130_fd_sc_hd__nor2_1 U21970 ( .A(n14840), .B(n14839), .Y(n14841) );
  sky130_fd_sc_hd__nand3_1 U21971 ( .A(n14842), .B(n14833), .C(n14841), .Y(
        n25642) );
  sky130_fd_sc_hd__inv_2 U21972 ( .A(n25642), .Y(n26324) );
  sky130_fd_sc_hd__o22ai_1 U21973 ( .A1(n16501), .A2(n26431), .B1(n26324), 
        .B2(n16500), .Y(n15084) );
  sky130_fd_sc_hd__nand2_1 U21974 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[215]), .Y(n14846) );
  sky130_fd_sc_hd__nand2_1 U21975 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[470]), .Y(n14845) );
  sky130_fd_sc_hd__nand2_1 U21976 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[502]), .Y(n14844) );
  sky130_fd_sc_hd__nand2_1 U21977 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[247]), .Y(n14843) );
  sky130_fd_sc_hd__nand4_1 U21978 ( .A(n14846), .B(n14845), .C(n14844), .D(
        n14843), .Y(n14852) );
  sky130_fd_sc_hd__nand2_1 U21979 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[23]), .Y(n14850) );
  sky130_fd_sc_hd__nand2_1 U21980 ( .A(n15984), .B(
        j202_soc_core_j22_cpu_rf_gpr[87]), .Y(n14849) );
  sky130_fd_sc_hd__nand2_1 U21981 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[406]), .Y(n14848) );
  sky130_fd_sc_hd__nand2_1 U21982 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[151]), .Y(n14847) );
  sky130_fd_sc_hd__nand4_1 U21983 ( .A(n14850), .B(n14849), .C(n14848), .D(
        n14847), .Y(n14851) );
  sky130_fd_sc_hd__nor2_1 U21984 ( .A(n14852), .B(n14851), .Y(n14860) );
  sky130_fd_sc_hd__a22oi_1 U21985 ( .A1(n23776), .A2(
        j202_soc_core_j22_cpu_rf_gpr[374]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[279]), .Y(n14859) );
  sky130_fd_sc_hd__a22oi_1 U21986 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[55]), .B1(n15017), .B2(
        j202_soc_core_j22_cpu_rf_gpr[342]), .Y(n14858) );
  sky130_fd_sc_hd__nand2_1 U21987 ( .A(n15958), .B(
        j202_soc_core_j22_cpu_rf_gpr[311]), .Y(n14856) );
  sky130_fd_sc_hd__nand2_1 U21988 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[438]), .Y(n14855) );
  sky130_fd_sc_hd__nand2_1 U21989 ( .A(n11199), .B(
        j202_soc_core_j22_cpu_rf_gpr[183]), .Y(n14854) );
  sky130_fd_sc_hd__nand2_1 U21990 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[119]), .Y(n14853) );
  sky130_fd_sc_hd__and4_1 U21991 ( .A(n14856), .B(n14855), .C(n14854), .D(
        n14853), .X(n14857) );
  sky130_fd_sc_hd__nand4_1 U21992 ( .A(n14860), .B(n14859), .C(n14858), .D(
        n14857), .Y(n22095) );
  sky130_fd_sc_hd__nand2_1 U21993 ( .A(n22095), .B(n16523), .Y(n14872) );
  sky130_fd_sc_hd__o21ai_0 U21994 ( .A1(n14861), .A2(n16525), .B1(n16524), .Y(
        n14866) );
  sky130_fd_sc_hd__o22ai_1 U21995 ( .A1(n14864), .A2(n15886), .B1(n14862), 
        .B2(n14342), .Y(n14865) );
  sky130_fd_sc_hd__nor2_1 U21996 ( .A(n14866), .B(n14865), .Y(n14871) );
  sky130_fd_sc_hd__nand2_1 U21997 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[23]), .Y(n14870) );
  sky130_fd_sc_hd__nand2_1 U21998 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[23]), .Y(n14869) );
  sky130_fd_sc_hd__nand2_1 U21999 ( .A(n16533), .B(
        j202_soc_core_j22_cpu_pc[23]), .Y(n14868) );
  sky130_fd_sc_hd__nand2_1 U22000 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[23]), .Y(n14867) );
  sky130_fd_sc_hd__nand3_1 U22001 ( .A(n14872), .B(n14871), .C(n13060), .Y(
        n25230) );
  sky130_fd_sc_hd__nand2_1 U22002 ( .A(n25230), .B(n16541), .Y(n14873) );
  sky130_fd_sc_hd__nor2_1 U22004 ( .A(n15084), .B(n15085), .Y(n15896) );
  sky130_fd_sc_hd__nand2_1 U22005 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[338]), .Y(n14877) );
  sky130_fd_sc_hd__nand2_1 U22006 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[179]), .Y(n14876) );
  sky130_fd_sc_hd__nand2_1 U22007 ( .A(n14993), .B(
        j202_soc_core_j22_cpu_rf_gpr[115]), .Y(n14875) );
  sky130_fd_sc_hd__nand2_1 U22008 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[434]), .Y(n14874) );
  sky130_fd_sc_hd__nand4_1 U22009 ( .A(n14877), .B(n14876), .C(n14875), .D(
        n14874), .Y(n14883) );
  sky130_fd_sc_hd__nand2_1 U22010 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[51]), .Y(n14881) );
  sky130_fd_sc_hd__nand2_1 U22011 ( .A(n16433), .B(
        j202_soc_core_j22_cpu_rf_gpr[211]), .Y(n14880) );
  sky130_fd_sc_hd__nand2_1 U22012 ( .A(n15796), .B(
        j202_soc_core_j22_cpu_rf_gpr[83]), .Y(n14879) );
  sky130_fd_sc_hd__nand2_1 U22013 ( .A(n11196), .B(
        j202_soc_core_j22_cpu_rf_gpr[370]), .Y(n14878) );
  sky130_fd_sc_hd__nand4_1 U22014 ( .A(n14881), .B(n14880), .C(n14879), .D(
        n14878), .Y(n14882) );
  sky130_fd_sc_hd__nor2_1 U22015 ( .A(n14883), .B(n14882), .Y(n14898) );
  sky130_fd_sc_hd__nand2_1 U22016 ( .A(n16043), .B(
        j202_soc_core_j22_cpu_rf_gpr[243]), .Y(n14887) );
  sky130_fd_sc_hd__nand2_1 U22017 ( .A(n16425), .B(
        j202_soc_core_j22_cpu_rf_gpr[147]), .Y(n14886) );
  sky130_fd_sc_hd__nand2_1 U22018 ( .A(n11195), .B(
        j202_soc_core_j22_cpu_rf_gpr[402]), .Y(n14885) );
  sky130_fd_sc_hd__nand2_1 U22019 ( .A(n14985), .B(
        j202_soc_core_j22_cpu_rf_gpr[498]), .Y(n14884) );
  sky130_fd_sc_hd__nand4_1 U22020 ( .A(n14887), .B(n14886), .C(n14885), .D(
        n14884), .Y(n14888) );
  sky130_fd_sc_hd__nor2_1 U22021 ( .A(n14889), .B(n16444), .Y(n14895) );
  sky130_fd_sc_hd__a21oi_1 U22022 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[19]), .B1(n14743), .Y(n14893) );
  sky130_fd_sc_hd__nand2_1 U22023 ( .A(n11194), .B(
        j202_soc_core_j22_cpu_rf_gpr[307]), .Y(n14892) );
  sky130_fd_sc_hd__nand2_1 U22024 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[275]), .Y(n14891) );
  sky130_fd_sc_hd__nand2_1 U22025 ( .A(n15788), .B(
        j202_soc_core_j22_cpu_rf_gpr[466]), .Y(n14890) );
  sky130_fd_sc_hd__nand4_1 U22026 ( .A(n14893), .B(n14892), .C(n14891), .D(
        n14890), .Y(n14894) );
  sky130_fd_sc_hd__nor2_1 U22027 ( .A(n14895), .B(n14894), .Y(n14896) );
  sky130_fd_sc_hd__nand3_1 U22028 ( .A(n14898), .B(n14897), .C(n14896), .Y(
        n25697) );
  sky130_fd_sc_hd__inv_2 U22029 ( .A(n25697), .Y(n27027) );
  sky130_fd_sc_hd__o22ai_1 U22030 ( .A1(n16500), .A2(n27800), .B1(n27027), 
        .B2(n16501), .Y(n15072) );
  sky130_fd_sc_hd__nand2_1 U22031 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[211]), .Y(n14902) );
  sky130_fd_sc_hd__nand2_1 U22032 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[466]), .Y(n14901) );
  sky130_fd_sc_hd__nand2_1 U22033 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[498]), .Y(n14900) );
  sky130_fd_sc_hd__nand2_1 U22034 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[243]), .Y(n14899) );
  sky130_fd_sc_hd__nand4_1 U22035 ( .A(n14902), .B(n14901), .C(n14900), .D(
        n14899), .Y(n14908) );
  sky130_fd_sc_hd__nand2_1 U22036 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[19]), .Y(n14906) );
  sky130_fd_sc_hd__nand2_1 U22037 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[83]), .Y(n14905) );
  sky130_fd_sc_hd__nand2_1 U22038 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[402]), .Y(n14904) );
  sky130_fd_sc_hd__nand2_1 U22039 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[147]), .Y(n14903) );
  sky130_fd_sc_hd__nand4_1 U22040 ( .A(n14906), .B(n14905), .C(n14904), .D(
        n14903), .Y(n14907) );
  sky130_fd_sc_hd__nor2_1 U22041 ( .A(n14908), .B(n14907), .Y(n14916) );
  sky130_fd_sc_hd__a22oi_1 U22042 ( .A1(n15991), .A2(
        j202_soc_core_j22_cpu_rf_gpr[370]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[275]), .Y(n14915) );
  sky130_fd_sc_hd__a22oi_1 U22043 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[51]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_rf_gpr[338]), .Y(n14914) );
  sky130_fd_sc_hd__nand2_1 U22044 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[307]), .Y(n14912) );
  sky130_fd_sc_hd__nand2_1 U22045 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[434]), .Y(n14911) );
  sky130_fd_sc_hd__nand2_1 U22046 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[179]), .Y(n14910) );
  sky130_fd_sc_hd__nand2_1 U22047 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[115]), .Y(n14909) );
  sky130_fd_sc_hd__nand4_1 U22048 ( .A(n14916), .B(n14915), .C(n14914), .D(
        n14913), .Y(n22824) );
  sky130_fd_sc_hd__nand2_1 U22049 ( .A(n22824), .B(n16523), .Y(n14927) );
  sky130_fd_sc_hd__o21ai_0 U22050 ( .A1(n14917), .A2(n16525), .B1(n16524), .Y(
        n14921) );
  sky130_fd_sc_hd__o22ai_1 U22051 ( .A1(n14919), .A2(n16077), .B1(n14918), 
        .B2(n14342), .Y(n14920) );
  sky130_fd_sc_hd__nor2_1 U22052 ( .A(n14921), .B(n14920), .Y(n14926) );
  sky130_fd_sc_hd__nand2_1 U22053 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[19]), .Y(n14925) );
  sky130_fd_sc_hd__nand2_1 U22054 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[19]), .Y(n14924) );
  sky130_fd_sc_hd__nand2_1 U22055 ( .A(n16533), .B(
        j202_soc_core_j22_cpu_pc[19]), .Y(n14923) );
  sky130_fd_sc_hd__nand2_1 U22056 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[19]), .Y(n14922) );
  sky130_fd_sc_hd__nand2_1 U22057 ( .A(n25692), .B(n16541), .Y(n14928) );
  sky130_fd_sc_hd__nor2_1 U22059 ( .A(n15072), .B(n15073), .Y(n15489) );
  sky130_fd_sc_hd__nand2_1 U22060 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[148]), .Y(n14932) );
  sky130_fd_sc_hd__nand2_1 U22061 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[84]), .Y(n14931) );
  sky130_fd_sc_hd__nand2_1 U22062 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[403]), .Y(n14930) );
  sky130_fd_sc_hd__nand2_1 U22063 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[371]), .Y(n14929) );
  sky130_fd_sc_hd__nand4_1 U22064 ( .A(n14932), .B(n14931), .C(n14930), .D(
        n14929), .Y(n14938) );
  sky130_fd_sc_hd__nand2_1 U22065 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[276]), .Y(n14936) );
  sky130_fd_sc_hd__nand2_1 U22066 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[308]), .Y(n14935) );
  sky130_fd_sc_hd__nand2_1 U22067 ( .A(n15788), .B(
        j202_soc_core_j22_cpu_rf_gpr[467]), .Y(n14934) );
  sky130_fd_sc_hd__nand2_1 U22068 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[435]), .Y(n14933) );
  sky130_fd_sc_hd__nand4_1 U22069 ( .A(n14936), .B(n14935), .C(n14934), .D(
        n14933), .Y(n14937) );
  sky130_fd_sc_hd__nor2_1 U22070 ( .A(n14938), .B(n14937), .Y(n14950) );
  sky130_fd_sc_hd__nand2_1 U22071 ( .A(n16432), .B(
        j202_soc_core_j22_cpu_rf_gpr[339]), .Y(n14942) );
  sky130_fd_sc_hd__nand2_1 U22072 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[180]), .Y(n14941) );
  sky130_fd_sc_hd__nand2_1 U22073 ( .A(n15783), .B(
        j202_soc_core_j22_cpu_rf_gpr[116]), .Y(n14940) );
  sky130_fd_sc_hd__nand2_1 U22074 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[212]), .Y(n14939) );
  sky130_fd_sc_hd__nor2_1 U22075 ( .A(n14975), .B(n14798), .Y(n14948) );
  sky130_fd_sc_hd__a21oi_1 U22076 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[20]), .B1(n14743), .Y(n14946) );
  sky130_fd_sc_hd__nand2_1 U22077 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[244]), .Y(n14945) );
  sky130_fd_sc_hd__nand2_1 U22078 ( .A(n14985), .B(
        j202_soc_core_j22_cpu_rf_gpr[499]), .Y(n14944) );
  sky130_fd_sc_hd__nand2_1 U22079 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[52]), .Y(n14943) );
  sky130_fd_sc_hd__nand4_1 U22080 ( .A(n14946), .B(n14945), .C(n14944), .D(
        n14943), .Y(n14947) );
  sky130_fd_sc_hd__nor2_1 U22081 ( .A(n14948), .B(n14947), .Y(n14949) );
  sky130_fd_sc_hd__inv_2 U22082 ( .A(n26331), .Y(n27383) );
  sky130_fd_sc_hd__o22ai_1 U22083 ( .A1(n16501), .A2(n27383), .B1(n27027), 
        .B2(n16500), .Y(n15074) );
  sky130_fd_sc_hd__nand2_1 U22084 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[212]), .Y(n14954) );
  sky130_fd_sc_hd__nand2_1 U22085 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[467]), .Y(n14953) );
  sky130_fd_sc_hd__nand2_1 U22086 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[499]), .Y(n14952) );
  sky130_fd_sc_hd__nand2_1 U22087 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[244]), .Y(n14951) );
  sky130_fd_sc_hd__nand4_1 U22088 ( .A(n14954), .B(n14953), .C(n14952), .D(
        n14951), .Y(n14960) );
  sky130_fd_sc_hd__nand2_1 U22089 ( .A(n16506), .B(
        j202_soc_core_j22_cpu_rf_gpr[20]), .Y(n14958) );
  sky130_fd_sc_hd__nand2_1 U22090 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[84]), .Y(n14957) );
  sky130_fd_sc_hd__nand2_1 U22091 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[403]), .Y(n14956) );
  sky130_fd_sc_hd__nand2_1 U22092 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[148]), .Y(n14955) );
  sky130_fd_sc_hd__nand4_1 U22093 ( .A(n14958), .B(n14957), .C(n14956), .D(
        n14955), .Y(n14959) );
  sky130_fd_sc_hd__nor2_1 U22094 ( .A(n14960), .B(n14959), .Y(n14971) );
  sky130_fd_sc_hd__nand2_1 U22095 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[276]), .Y(n14964) );
  sky130_fd_sc_hd__nand2_1 U22096 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[52]), .Y(n14963) );
  sky130_fd_sc_hd__nand2_1 U22097 ( .A(n23776), .B(
        j202_soc_core_j22_cpu_rf_gpr[371]), .Y(n14962) );
  sky130_fd_sc_hd__nand2_1 U22098 ( .A(n16064), .B(
        j202_soc_core_j22_cpu_rf_gpr[339]), .Y(n14961) );
  sky130_fd_sc_hd__and4_1 U22099 ( .A(n14964), .B(n14963), .C(n14962), .D(
        n14961), .X(n14970) );
  sky130_fd_sc_hd__nand2_1 U22100 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[308]), .Y(n14968) );
  sky130_fd_sc_hd__nand2_1 U22101 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[435]), .Y(n14967) );
  sky130_fd_sc_hd__nand2_1 U22102 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[180]), .Y(n14966) );
  sky130_fd_sc_hd__nand2_1 U22103 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[116]), .Y(n14965) );
  sky130_fd_sc_hd__and4_1 U22104 ( .A(n14968), .B(n14967), .C(n14966), .D(
        n14965), .X(n14969) );
  sky130_fd_sc_hd__nand3_1 U22105 ( .A(n14971), .B(n14970), .C(n14969), .Y(
        n22326) );
  sky130_fd_sc_hd__o22a_1 U22106 ( .A1(n14974), .A2(n16491), .B1(n16487), .B2(
        n22322), .X(n14978) );
  sky130_fd_sc_hd__o22a_1 U22107 ( .A1(n14975), .A2(n16488), .B1(n16490), .B2(
        n22321), .X(n14977) );
  sky130_fd_sc_hd__a21oi_1 U22108 ( .A1(n11201), .A2(
        j202_soc_core_j22_cpu_rf_gpr[499]), .B1(n16493), .Y(n14976) );
  sky130_fd_sc_hd__nand4_1 U22109 ( .A(n14979), .B(n14978), .C(n14977), .D(
        n14976), .Y(n14980) );
  sky130_fd_sc_hd__a21oi_2 U22110 ( .A1(n22326), .A2(n16523), .B1(n14980), .Y(
        n28506) );
  sky130_fd_sc_hd__mux2i_1 U22111 ( .A0(n16088), .A1(n16543), .S(n28506), .Y(
        n15075) );
  sky130_fd_sc_hd__nor2_1 U22112 ( .A(n15074), .B(n15075), .Y(n15384) );
  sky130_fd_sc_hd__nand2_1 U22113 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[181]), .Y(n14984) );
  sky130_fd_sc_hd__nand2_1 U22114 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[436]), .Y(n14983) );
  sky130_fd_sc_hd__nand2_1 U22115 ( .A(n11195), .B(
        j202_soc_core_j22_cpu_rf_gpr[404]), .Y(n14982) );
  sky130_fd_sc_hd__nand2_1 U22116 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[277]), .Y(n14981) );
  sky130_fd_sc_hd__nand4_1 U22117 ( .A(n14984), .B(n14983), .C(n14982), .D(
        n14981), .Y(n14992) );
  sky130_fd_sc_hd__nand2_1 U22118 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[213]), .Y(n14990) );
  sky130_fd_sc_hd__nand2_1 U22119 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[53]), .Y(n14989) );
  sky130_fd_sc_hd__nand2_1 U22120 ( .A(n14985), .B(
        j202_soc_core_j22_cpu_rf_gpr[500]), .Y(n14988) );
  sky130_fd_sc_hd__nand2_1 U22121 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[149]), .Y(n14987) );
  sky130_fd_sc_hd__nand4_1 U22122 ( .A(n14990), .B(n14989), .C(n14988), .D(
        n14987), .Y(n14991) );
  sky130_fd_sc_hd__nor2_1 U22123 ( .A(n14992), .B(n14991), .Y(n15006) );
  sky130_fd_sc_hd__nand2_1 U22124 ( .A(n16432), .B(
        j202_soc_core_j22_cpu_rf_gpr[340]), .Y(n14997) );
  sky130_fd_sc_hd__nand2_1 U22125 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[372]), .Y(n14996) );
  sky130_fd_sc_hd__nand2_1 U22126 ( .A(n14993), .B(
        j202_soc_core_j22_cpu_rf_gpr[117]), .Y(n14995) );
  sky130_fd_sc_hd__nand2_1 U22127 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[468]), .Y(n14994) );
  sky130_fd_sc_hd__nor2_1 U22128 ( .A(n14998), .B(n14798), .Y(n15004) );
  sky130_fd_sc_hd__a21oi_1 U22129 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[21]), .B1(n14743), .Y(n15002) );
  sky130_fd_sc_hd__nand2_1 U22130 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[309]), .Y(n15001) );
  sky130_fd_sc_hd__nand2_1 U22131 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[85]), .Y(n15000) );
  sky130_fd_sc_hd__nand2_1 U22132 ( .A(n16043), .B(
        j202_soc_core_j22_cpu_rf_gpr[245]), .Y(n14999) );
  sky130_fd_sc_hd__nand4_1 U22133 ( .A(n15002), .B(n15001), .C(n15000), .D(
        n14999), .Y(n15003) );
  sky130_fd_sc_hd__nor2_1 U22134 ( .A(n15004), .B(n15003), .Y(n15005) );
  sky130_fd_sc_hd__o22ai_1 U22135 ( .A1(n16501), .A2(n26324), .B1(n26280), 
        .B2(n16500), .Y(n15078) );
  sky130_fd_sc_hd__nand2_1 U22136 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[214]), .Y(n15010) );
  sky130_fd_sc_hd__nand2_1 U22137 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[469]), .Y(n15009) );
  sky130_fd_sc_hd__nand2_1 U22138 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[501]), .Y(n15008) );
  sky130_fd_sc_hd__nand2_1 U22139 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[246]), .Y(n15007) );
  sky130_fd_sc_hd__nand4_1 U22140 ( .A(n15010), .B(n15009), .C(n15008), .D(
        n15007), .Y(n15016) );
  sky130_fd_sc_hd__nand2_1 U22141 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[22]), .Y(n15014) );
  sky130_fd_sc_hd__nand2_1 U22142 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[86]), .Y(n15013) );
  sky130_fd_sc_hd__nand2_1 U22143 ( .A(n16466), .B(
        j202_soc_core_j22_cpu_rf_gpr[405]), .Y(n15012) );
  sky130_fd_sc_hd__nand2_1 U22144 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[150]), .Y(n15011) );
  sky130_fd_sc_hd__nand4_1 U22145 ( .A(n15014), .B(n15013), .C(n15012), .D(
        n15011), .Y(n15015) );
  sky130_fd_sc_hd__nor2_1 U22146 ( .A(n15016), .B(n15015), .Y(n15025) );
  sky130_fd_sc_hd__a22oi_1 U22147 ( .A1(n15991), .A2(
        j202_soc_core_j22_cpu_rf_gpr[373]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[278]), .Y(n15024) );
  sky130_fd_sc_hd__a22oi_1 U22148 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[54]), .B1(n15017), .B2(
        j202_soc_core_j22_cpu_rf_gpr[341]), .Y(n15023) );
  sky130_fd_sc_hd__nand2_1 U22149 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[310]), .Y(n15021) );
  sky130_fd_sc_hd__nand2_1 U22150 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[437]), .Y(n15020) );
  sky130_fd_sc_hd__nand2_1 U22151 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[182]), .Y(n15019) );
  sky130_fd_sc_hd__nand2_1 U22152 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[118]), .Y(n15018) );
  sky130_fd_sc_hd__nand4_1 U22153 ( .A(n15025), .B(n15024), .C(n15023), .D(
        n15022), .Y(n22169) );
  sky130_fd_sc_hd__nand2_1 U22154 ( .A(n22169), .B(n16523), .Y(n15036) );
  sky130_fd_sc_hd__o21ai_0 U22155 ( .A1(n15026), .A2(n16525), .B1(n16524), .Y(
        n15030) );
  sky130_fd_sc_hd__o22ai_1 U22156 ( .A1(n15028), .A2(n16077), .B1(n15027), 
        .B2(n14477), .Y(n15029) );
  sky130_fd_sc_hd__nor2_1 U22157 ( .A(n15030), .B(n15029), .Y(n15035) );
  sky130_fd_sc_hd__nand2_1 U22158 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[22]), .Y(n15034) );
  sky130_fd_sc_hd__nand2_1 U22159 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[22]), .Y(n15033) );
  sky130_fd_sc_hd__nand2_1 U22160 ( .A(n16533), .B(
        j202_soc_core_j22_cpu_pc[22]), .Y(n15032) );
  sky130_fd_sc_hd__nand2_1 U22161 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[22]), .Y(n15031) );
  sky130_fd_sc_hd__nand3_1 U22162 ( .A(n15036), .B(n15035), .C(n13084), .Y(
        n28493) );
  sky130_fd_sc_hd__nand2_1 U22163 ( .A(n28493), .B(n16541), .Y(n15037) );
  sky130_fd_sc_hd__nor2_1 U22165 ( .A(n15078), .B(n15079), .Y(n15184) );
  sky130_fd_sc_hd__o22ai_1 U22166 ( .A1(n16501), .A2(n26280), .B1(n27383), 
        .B2(n16500), .Y(n15076) );
  sky130_fd_sc_hd__nand2_1 U22167 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[213]), .Y(n15041) );
  sky130_fd_sc_hd__nand2_1 U22168 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[468]), .Y(n15040) );
  sky130_fd_sc_hd__nand2_1 U22169 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[500]), .Y(n15039) );
  sky130_fd_sc_hd__nand2_1 U22170 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[245]), .Y(n15038) );
  sky130_fd_sc_hd__nand4_1 U22171 ( .A(n15041), .B(n15040), .C(n15039), .D(
        n15038), .Y(n15047) );
  sky130_fd_sc_hd__nand2_1 U22172 ( .A(n16506), .B(
        j202_soc_core_j22_cpu_rf_gpr[21]), .Y(n15045) );
  sky130_fd_sc_hd__nand2_1 U22173 ( .A(n15984), .B(
        j202_soc_core_j22_cpu_rf_gpr[85]), .Y(n15044) );
  sky130_fd_sc_hd__nand2_1 U22174 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[404]), .Y(n15043) );
  sky130_fd_sc_hd__nand2_1 U22175 ( .A(n23808), .B(
        j202_soc_core_j22_cpu_rf_gpr[149]), .Y(n15042) );
  sky130_fd_sc_hd__nand4_1 U22176 ( .A(n15045), .B(n15044), .C(n15043), .D(
        n15042), .Y(n15046) );
  sky130_fd_sc_hd__nor2_1 U22177 ( .A(n15047), .B(n15046), .Y(n15055) );
  sky130_fd_sc_hd__a22oi_1 U22178 ( .A1(n23776), .A2(
        j202_soc_core_j22_cpu_rf_gpr[372]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[277]), .Y(n15054) );
  sky130_fd_sc_hd__a22oi_1 U22179 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[53]), .B1(n15017), .B2(
        j202_soc_core_j22_cpu_rf_gpr[340]), .Y(n15053) );
  sky130_fd_sc_hd__nand2_1 U22180 ( .A(n15958), .B(
        j202_soc_core_j22_cpu_rf_gpr[309]), .Y(n15051) );
  sky130_fd_sc_hd__nand2_1 U22181 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[436]), .Y(n15050) );
  sky130_fd_sc_hd__nand2_1 U22182 ( .A(n11199), .B(
        j202_soc_core_j22_cpu_rf_gpr[181]), .Y(n15049) );
  sky130_fd_sc_hd__nand2_1 U22183 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[117]), .Y(n15048) );
  sky130_fd_sc_hd__nand4_1 U22184 ( .A(n15055), .B(n15054), .C(n15053), .D(
        n15052), .Y(n22306) );
  sky130_fd_sc_hd__nand2_1 U22185 ( .A(n22306), .B(n16523), .Y(n15066) );
  sky130_fd_sc_hd__o21ai_0 U22186 ( .A1(n15056), .A2(n16525), .B1(n16524), .Y(
        n15060) );
  sky130_fd_sc_hd__o22ai_1 U22187 ( .A1(n15058), .A2(n16077), .B1(n15057), 
        .B2(n14477), .Y(n15059) );
  sky130_fd_sc_hd__nor2_1 U22188 ( .A(n15060), .B(n15059), .Y(n15065) );
  sky130_fd_sc_hd__nand2_1 U22189 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[21]), .Y(n15064) );
  sky130_fd_sc_hd__nand2_1 U22190 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[21]), .Y(n15063) );
  sky130_fd_sc_hd__nand2_1 U22191 ( .A(n16533), .B(
        j202_soc_core_j22_cpu_pc[21]), .Y(n15062) );
  sky130_fd_sc_hd__nand2_1 U22192 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[21]), .Y(n15061) );
  sky130_fd_sc_hd__nand2_1 U22193 ( .A(n28499), .B(n16541), .Y(n15067) );
  sky130_fd_sc_hd__nor2_1 U22195 ( .A(n15076), .B(n15077), .Y(n15639) );
  sky130_fd_sc_hd__nor2_1 U22196 ( .A(n15184), .B(n15639), .Y(n15081) );
  sky130_fd_sc_hd__nand2_1 U22197 ( .A(n15181), .B(n15081), .Y(n15083) );
  sky130_fd_sc_hd__nor2_1 U22198 ( .A(n15069), .B(n21032), .Y(n15071) );
  sky130_fd_sc_hd__nand2_1 U22199 ( .A(n21030), .B(n15071), .Y(n15380) );
  sky130_fd_sc_hd__inv_2 U22200 ( .A(n16545), .Y(n17030) );
  sky130_fd_sc_hd__nor2_1 U22201 ( .A(n15896), .B(n17030), .Y(n15087) );
  sky130_fd_sc_hd__o21ai_1 U22202 ( .A1(n21033), .A2(n15069), .B1(n15068), .Y(
        n15070) );
  sky130_fd_sc_hd__nand2_1 U22204 ( .A(n15073), .B(n15072), .Y(n15490) );
  sky130_fd_sc_hd__nand2_1 U22205 ( .A(n15075), .B(n15074), .Y(n15385) );
  sky130_fd_sc_hd__nand2_1 U22207 ( .A(n15077), .B(n15076), .Y(n15640) );
  sky130_fd_sc_hd__nand2_1 U22208 ( .A(n15079), .B(n15078), .Y(n15185) );
  sky130_fd_sc_hd__a21oi_1 U22210 ( .A1(n15081), .A2(n15180), .B1(n15080), .Y(
        n15082) );
  sky130_fd_sc_hd__o21ai_2 U22211 ( .A1(n15083), .A2(n15381), .B1(n15082), .Y(
        n16555) );
  sky130_fd_sc_hd__inv_2 U22212 ( .A(n16555), .Y(n17036) );
  sky130_fd_sc_hd__nand2_1 U22213 ( .A(n15085), .B(n15084), .Y(n16014) );
  sky130_fd_sc_hd__o21ai_1 U22214 ( .A1(n15896), .A2(n17036), .B1(n16014), .Y(
        n15086) );
  sky130_fd_sc_hd__a21oi_1 U22215 ( .A1(n17040), .A2(n15087), .B1(n15086), .Y(
        n15088) );
  sky130_fd_sc_hd__xor2_1 U22216 ( .A(n15089), .B(n15088), .X(n26461) );
  sky130_fd_sc_hd__nand2_1 U22217 ( .A(n26461), .B(n17225), .Y(n15090) );
  sky130_fd_sc_hd__nand2_1 U22218 ( .A(j202_soc_core_memory0_ram_dout0[86]), 
        .B(n20458), .Y(n15092) );
  sky130_fd_sc_hd__and2_0 U22219 ( .A(n15093), .B(n20454), .X(n15094) );
  sky130_fd_sc_hd__nand2_1 U22220 ( .A(n15684), .B(n20485), .Y(n15119) );
  sky130_fd_sc_hd__nand2_1 U22221 ( .A(n17241), .B(
        j202_soc_core_bootrom_00_address_w[8]), .Y(n15096) );
  sky130_fd_sc_hd__nor2_1 U22222 ( .A(n15119), .B(n15096), .Y(n15340) );
  sky130_fd_sc_hd__nor2_1 U22223 ( .A(n15678), .B(n15111), .Y(n15597) );
  sky130_fd_sc_hd__nor2_1 U22224 ( .A(n15685), .B(n15149), .Y(n15148) );
  sky130_fd_sc_hd__nand2_1 U22225 ( .A(n15303), .B(n20196), .Y(n15585) );
  sky130_fd_sc_hd__nand2_1 U22226 ( .A(n15597), .B(n15684), .Y(n15098) );
  sky130_fd_sc_hd__nand2_1 U22227 ( .A(n15585), .B(n15098), .Y(n15518) );
  sky130_fd_sc_hd__nor2_1 U22228 ( .A(n15148), .B(n15518), .Y(n15540) );
  sky130_fd_sc_hd__nand2_1 U22229 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .B(n13199), .Y(n21580) );
  sky130_fd_sc_hd__nand2_1 U22230 ( .A(n15685), .B(n21580), .Y(n15133) );
  sky130_fd_sc_hd__nand3_1 U22231 ( .A(n15133), .B(n17250), .C(
        j202_soc_core_bootrom_00_address_w[8]), .Y(n15095) );
  sky130_fd_sc_hd__nand2_1 U22232 ( .A(n15540), .B(n15095), .Y(n15604) );
  sky130_fd_sc_hd__o21ai_1 U22233 ( .A1(n15340), .A2(n15604), .B1(n19816), .Y(
        n15103) );
  sky130_fd_sc_hd__nand2_1 U22234 ( .A(n19124), .B(n20485), .Y(n20603) );
  sky130_fd_sc_hd__nand2b_1 U22235 ( .A_N(n20603), .B(
        j202_soc_core_bootrom_00_address_w[8]), .Y(n15307) );
  sky130_fd_sc_hd__nand2_1 U22236 ( .A(n19504), .B(n16871), .Y(n15509) );
  sky130_fd_sc_hd__nand2b_1 U22237 ( .A_N(n15509), .B(n13199), .Y(n15328) );
  sky130_fd_sc_hd__nand2_1 U22238 ( .A(n19129), .B(n20485), .Y(n15120) );
  sky130_fd_sc_hd__nand2_1 U22239 ( .A(n15097), .B(n15153), .Y(n15495) );
  sky130_fd_sc_hd__nand3_1 U22240 ( .A(n15307), .B(n15328), .C(n15495), .Y(
        n15602) );
  sky130_fd_sc_hd__nand2_1 U22241 ( .A(n15602), .B(n21103), .Y(n15102) );
  sky130_fd_sc_hd__nand2_1 U22242 ( .A(n15303), .B(n20235), .Y(n15566) );
  sky130_fd_sc_hd__nand2_1 U22243 ( .A(n15566), .B(n15098), .Y(n15329) );
  sky130_fd_sc_hd__nand2b_1 U22244 ( .A_N(n15509), .B(n20485), .Y(n15584) );
  sky130_fd_sc_hd__nand2_1 U22245 ( .A(n15585), .B(n15584), .Y(n15275) );
  sky130_fd_sc_hd__nand2b_1 U22246 ( .A_N(n20603), .B(n17264), .Y(n15559) );
  sky130_fd_sc_hd__nand2b_1 U22247 ( .A_N(n19120), .B(n20194), .Y(n15277) );
  sky130_fd_sc_hd__nand2_1 U22248 ( .A(n17250), .B(n19119), .Y(n15677) );
  sky130_fd_sc_hd__nand2b_1 U22249 ( .A_N(n15677), .B(n20126), .Y(n15327) );
  sky130_fd_sc_hd__and3_1 U22250 ( .A(n15277), .B(n15327), .C(n15495), .X(
        n15099) );
  sky130_fd_sc_hd__nand3_1 U22251 ( .A(n15100), .B(n15559), .C(n15099), .Y(
        n15354) );
  sky130_fd_sc_hd__o21ai_1 U22252 ( .A1(n15329), .A2(n15354), .B1(n17237), .Y(
        n15101) );
  sky130_fd_sc_hd__nand3_1 U22253 ( .A(n15103), .B(n15102), .C(n15101), .Y(
        n15108) );
  sky130_fd_sc_hd__nand2_1 U22254 ( .A(n19124), .B(n20235), .Y(n15589) );
  sky130_fd_sc_hd__nand2_1 U22255 ( .A(n17250), .B(n20235), .Y(n15109) );
  sky130_fd_sc_hd__nand2b_1 U22256 ( .A_N(n15109), .B(n19129), .Y(n15568) );
  sky130_fd_sc_hd__nand2_1 U22257 ( .A(n15589), .B(n15568), .Y(n15280) );
  sky130_fd_sc_hd__nand2_1 U22258 ( .A(n19124), .B(n20196), .Y(n15283) );
  sky130_fd_sc_hd__nand2b_1 U22259 ( .A_N(n15280), .B(n15283), .Y(n15564) );
  sky130_fd_sc_hd__nand2b_1 U22260 ( .A_N(n15120), .B(n17250), .Y(n15555) );
  sky130_fd_sc_hd__nor2_1 U22261 ( .A(n17264), .B(n15555), .Y(n15294) );
  sky130_fd_sc_hd__nand2b_1 U22262 ( .A_N(n15677), .B(n20196), .Y(n15547) );
  sky130_fd_sc_hd__nand2_1 U22263 ( .A(n15584), .B(n15547), .Y(n15211) );
  sky130_fd_sc_hd__o21ai_1 U22265 ( .A1(n15568), .A2(n19726), .B1(n15104), .Y(
        n15105) );
  sky130_fd_sc_hd__a21oi_1 U22266 ( .A1(n15564), .A2(n19804), .B1(n15105), .Y(
        n15107) );
  sky130_fd_sc_hd__a2bb2oi_1 U22267 ( .B1(n15610), .B2(n15108), .A1_N(n15107), 
        .A2_N(n15106), .Y(n15240) );
  sky130_fd_sc_hd__nand2b_1 U22268 ( .A_N(n15109), .B(n20531), .Y(n15304) );
  sky130_fd_sc_hd__nand2_1 U22269 ( .A(n15568), .B(n15304), .Y(n15352) );
  sky130_fd_sc_hd__nor2_1 U22270 ( .A(n15138), .B(n15352), .Y(n15587) );
  sky130_fd_sc_hd__nand2_1 U22271 ( .A(n15303), .B(n20126), .Y(n15295) );
  sky130_fd_sc_hd__nand3_1 U22272 ( .A(n15587), .B(n15589), .C(n15295), .Y(
        n15110) );
  sky130_fd_sc_hd__nand2_1 U22273 ( .A(n15110), .B(n21103), .Y(n15116) );
  sky130_fd_sc_hd__nand2_1 U22274 ( .A(n15303), .B(n15111), .Y(n15112) );
  sky130_fd_sc_hd__nand3_1 U22275 ( .A(n15310), .B(n15495), .C(n15112), .Y(
        n15219) );
  sky130_fd_sc_hd__nand2b_1 U22276 ( .A_N(n15219), .B(n15277), .Y(n15350) );
  sky130_fd_sc_hd__nand2_1 U22277 ( .A(n15350), .B(n19804), .Y(n15115) );
  sky130_fd_sc_hd__nor2_1 U22278 ( .A(n19816), .B(n17237), .Y(n19468) );
  sky130_fd_sc_hd__nand3_1 U22279 ( .A(n17250), .B(n20531), .C(n20126), .Y(
        n15546) );
  sky130_fd_sc_hd__o22ai_1 U22280 ( .A1(n19468), .A2(n15546), .B1(n19726), 
        .B2(n15327), .Y(n15113) );
  sky130_fd_sc_hd__a21oi_1 U22281 ( .A1(n17237), .A2(n15148), .B1(n15113), .Y(
        n15114) );
  sky130_fd_sc_hd__nand3_1 U22282 ( .A(n15116), .B(n15115), .C(n15114), .Y(
        n15129) );
  sky130_fd_sc_hd__nand2_1 U22283 ( .A(n19119), .B(n13199), .Y(n21150) );
  sky130_fd_sc_hd__nor2_1 U22284 ( .A(n21150), .B(n17100), .Y(n19131) );
  sky130_fd_sc_hd__nand2_1 U22285 ( .A(n19131), .B(
        j202_soc_core_bootrom_00_address_w[8]), .Y(n15599) );
  sky130_fd_sc_hd__nand2_1 U22286 ( .A(n15559), .B(n15599), .Y(n15284) );
  sky130_fd_sc_hd__o21ai_0 U22287 ( .A1(n15117), .A2(n15284), .B1(n17237), .Y(
        n15127) );
  sky130_fd_sc_hd__nand2_1 U22288 ( .A(n20531), .B(n13199), .Y(n15118) );
  sky130_fd_sc_hd__nand2_1 U22289 ( .A(n15153), .B(n15118), .Y(n15139) );
  sky130_fd_sc_hd__nand2b_1 U22290 ( .A_N(n15139), .B(n15119), .Y(n15567) );
  sky130_fd_sc_hd__nand3_1 U22291 ( .A(n15559), .B(n15310), .C(n15567), .Y(
        n15122) );
  sky130_fd_sc_hd__nand2_1 U22292 ( .A(n15153), .B(n15120), .Y(n15554) );
  sky130_fd_sc_hd__a31oi_1 U22293 ( .A1(n20603), .A2(n15547), .A3(n15554), 
        .B1(n19726), .Y(n15121) );
  sky130_fd_sc_hd__a21oi_1 U22294 ( .A1(n15122), .A2(n19804), .B1(n15121), .Y(
        n15126) );
  sky130_fd_sc_hd__nand2_1 U22295 ( .A(n19712), .B(n20194), .Y(n15504) );
  sky130_fd_sc_hd__nand2_1 U22296 ( .A(n15277), .B(n15504), .Y(n15593) );
  sky130_fd_sc_hd__nor2_1 U22297 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n15327), .Y(n15130) );
  sky130_fd_sc_hd__nor2_1 U22298 ( .A(n15593), .B(n15130), .Y(n15503) );
  sky130_fd_sc_hd__nand2_1 U22299 ( .A(n15304), .B(n15495), .Y(n15123) );
  sky130_fd_sc_hd__nand3_1 U22300 ( .A(n15153), .B(n19129), .C(n13199), .Y(
        n15508) );
  sky130_fd_sc_hd__nand2_1 U22301 ( .A(n15535), .B(n15508), .Y(n15526) );
  sky130_fd_sc_hd__nor2_1 U22302 ( .A(n15123), .B(n15526), .Y(n15317) );
  sky130_fd_sc_hd__nor2_1 U22303 ( .A(n19839), .B(n19120), .Y(n15595) );
  sky130_fd_sc_hd__and3_1 U22304 ( .A(n15562), .B(n15590), .C(n15546), .X(
        n15278) );
  sky130_fd_sc_hd__nand3_1 U22305 ( .A(n15503), .B(n15317), .C(n15278), .Y(
        n15124) );
  sky130_fd_sc_hd__nand2_1 U22306 ( .A(n15124), .B(n21103), .Y(n15125) );
  sky130_fd_sc_hd__nand3_1 U22307 ( .A(n15127), .B(n15126), .C(n15125), .Y(
        n15128) );
  sky130_fd_sc_hd__a22oi_1 U22308 ( .A1(n15610), .A2(n15129), .B1(n15128), 
        .B2(n15577), .Y(n15167) );
  sky130_fd_sc_hd__nand2_1 U22309 ( .A(n15599), .B(n15310), .Y(n15549) );
  sky130_fd_sc_hd__nand2_1 U22310 ( .A(n20485), .B(
        j202_soc_core_bootrom_00_address_w[4]), .Y(n21395) );
  sky130_fd_sc_hd__nand2b_1 U22311 ( .A_N(n17100), .B(n21603), .Y(n20520) );
  sky130_fd_sc_hd__nand3_1 U22312 ( .A(n15344), .B(n15504), .C(n20520), .Y(
        n15537) );
  sky130_fd_sc_hd__nand2_1 U22313 ( .A(n19131), .B(n17264), .Y(n15557) );
  sky130_fd_sc_hd__nand2b_1 U22314 ( .A_N(n19120), .B(n20126), .Y(n15583) );
  sky130_fd_sc_hd__nand2_1 U22315 ( .A(n15557), .B(n15583), .Y(n15321) );
  sky130_fd_sc_hd__nor2_1 U22316 ( .A(n15537), .B(n15321), .Y(n15131) );
  sky130_fd_sc_hd__nor2_1 U22317 ( .A(n15596), .B(n15605), .Y(n15342) );
  sky130_fd_sc_hd__nand4_1 U22318 ( .A(n15131), .B(n15342), .C(n15585), .D(
        n15328), .Y(n15132) );
  sky130_fd_sc_hd__nor3_1 U22319 ( .A(n15280), .B(n15549), .C(n15132), .Y(
        n15146) );
  sky130_fd_sc_hd__nand2_1 U22320 ( .A(n15153), .B(n15133), .Y(n15134) );
  sky130_fd_sc_hd__nand2_1 U22321 ( .A(n15134), .B(n15546), .Y(n15135) );
  sky130_fd_sc_hd__nand2_1 U22322 ( .A(n17241), .B(n20235), .Y(n15225) );
  sky130_fd_sc_hd__nand2b_1 U22323 ( .A_N(n15225), .B(n19129), .Y(n15532) );
  sky130_fd_sc_hd__nor2_1 U22324 ( .A(n15135), .B(n15347), .Y(n15136) );
  sky130_fd_sc_hd__nand4_1 U22325 ( .A(n15152), .B(n15307), .C(n15136), .D(
        n15599), .Y(n15143) );
  sky130_fd_sc_hd__nand2_1 U22326 ( .A(n19712), .B(n20235), .Y(n15598) );
  sky130_fd_sc_hd__nor2_1 U22327 ( .A(n15138), .B(n15137), .Y(n15140) );
  sky130_fd_sc_hd__nand2_1 U22328 ( .A(n19119), .B(n20485), .Y(n21412) );
  sky130_fd_sc_hd__nand2b_1 U22329 ( .A_N(n15139), .B(n21412), .Y(n15325) );
  sky130_fd_sc_hd__nand4_1 U22330 ( .A(n15140), .B(n15589), .C(n15557), .D(
        n15325), .Y(n15141) );
  sky130_fd_sc_hd__o2bb2ai_1 U22331 ( .B1(n19468), .B2(n15295), .A1_N(n19816), 
        .A2_N(n15141), .Y(n15142) );
  sky130_fd_sc_hd__a21oi_1 U22332 ( .A1(n15143), .A2(n21103), .B1(n15142), .Y(
        n15145) );
  sky130_fd_sc_hd__nand2_1 U22333 ( .A(n15559), .B(n15504), .Y(n15299) );
  sky130_fd_sc_hd__nand4_1 U22334 ( .A(n15540), .B(n15342), .C(n15344), .D(
        n15599), .Y(n15291) );
  sky130_fd_sc_hd__o211ai_1 U22336 ( .A1(n12089), .A2(n15146), .B1(n15145), 
        .C1(n15144), .Y(n15147) );
  sky130_fd_sc_hd__nand2_1 U22337 ( .A(n15147), .B(n16205), .Y(n15166) );
  sky130_fd_sc_hd__nand3_1 U22338 ( .A(n15559), .B(n15590), .C(n15570), .Y(
        n15501) );
  sky130_fd_sc_hd__nor2_1 U22339 ( .A(n15150), .B(n15149), .Y(n15339) );
  sky130_fd_sc_hd__nand2_1 U22340 ( .A(n15295), .B(n15569), .Y(n15221) );
  sky130_fd_sc_hd__nor2_1 U22341 ( .A(n15594), .B(n15593), .Y(n15151) );
  sky130_fd_sc_hd__nand3_1 U22342 ( .A(n15152), .B(n15499), .C(n15151), .Y(
        n15311) );
  sky130_fd_sc_hd__nor3_1 U22343 ( .A(n15595), .B(n15501), .C(n15311), .Y(
        n15163) );
  sky130_fd_sc_hd__nand2_1 U22344 ( .A(n15344), .B(n15598), .Y(n15232) );
  sky130_fd_sc_hd__nand3_1 U22345 ( .A(n15153), .B(n20531), .C(n20485), .Y(
        n15341) );
  sky130_fd_sc_hd__nand3_1 U22346 ( .A(n20603), .B(n15341), .C(n15304), .Y(
        n15154) );
  sky130_fd_sc_hd__o31a_1 U22347 ( .A1(n15232), .A2(n15321), .A3(n15154), .B1(
        n17237), .X(n15158) );
  sky130_fd_sc_hd__nor2_1 U22348 ( .A(n19816), .B(n21103), .Y(n15274) );
  sky130_fd_sc_hd__nand2_1 U22349 ( .A(n16801), .B(n20485), .Y(n15270) );
  sky130_fd_sc_hd__nor2_1 U22350 ( .A(n15155), .B(n15270), .Y(n15510) );
  sky130_fd_sc_hd__nor3_1 U22351 ( .A(n15339), .B(n15510), .C(n15280), .Y(
        n15156) );
  sky130_fd_sc_hd__o22ai_1 U22352 ( .A1(n16986), .A2(n15503), .B1(n15274), 
        .B2(n15156), .Y(n15157) );
  sky130_fd_sc_hd__nor2_1 U22353 ( .A(n15158), .B(n15157), .Y(n15162) );
  sky130_fd_sc_hd__nor2_1 U22355 ( .A(n15160), .B(n15284), .Y(n15272) );
  sky130_fd_sc_hd__nand2b_1 U22356 ( .A_N(n17100), .B(n20126), .Y(n15563) );
  sky130_fd_sc_hd__nand4_1 U22357 ( .A(n15272), .B(n15590), .C(n15563), .D(
        n15508), .Y(n15200) );
  sky130_fd_sc_hd__nand2_1 U22358 ( .A(n15200), .B(n19816), .Y(n15161) );
  sky130_fd_sc_hd__o211ai_1 U22359 ( .A1(n12089), .A2(n15163), .B1(n15162), 
        .C1(n15161), .Y(n15164) );
  sky130_fd_sc_hd__nand2_1 U22360 ( .A(n15164), .B(n15516), .Y(n15165) );
  sky130_fd_sc_hd__nand4_1 U22361 ( .A(n15240), .B(n15167), .C(n15166), .D(
        n15165), .Y(n15168) );
  sky130_fd_sc_hd__nand2_1 U22362 ( .A(n15168), .B(n21629), .Y(n15172) );
  sky130_fd_sc_hd__a22oi_1 U22363 ( .A1(n21516), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[22]), .B1(n20759), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[86]), .Y(n15171) );
  sky130_fd_sc_hd__a22oi_1 U22364 ( .A1(n20540), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[54]), .B1(n21513), .B2(
        j202_soc_core_uart_div1[6]), .Y(n15170) );
  sky130_fd_sc_hd__nand2_1 U22365 ( .A(n20786), .B(
        j202_soc_core_bldc_core_00_pwm_duty[10]), .Y(n15169) );
  sky130_fd_sc_hd__nand4_1 U22366 ( .A(n15172), .B(n15171), .C(n15170), .D(
        n15169), .Y(n15173) );
  sky130_fd_sc_hd__a21oi_1 U22367 ( .A1(j202_soc_core_memory0_ram_dout0[502]), 
        .A2(n11207), .B1(n15173), .Y(n15174) );
  sky130_fd_sc_hd__nor2_1 U22368 ( .A(n15176), .B(n21026), .Y(n15257) );
  sky130_fd_sc_hd__nand2_1 U22369 ( .A(n15257), .B(
        j202_soc_core_j22_cpu_pc[21]), .Y(n15177) );
  sky130_fd_sc_hd__xor2_1 U22370 ( .A(n15177), .B(n22164), .X(n25595) );
  sky130_fd_sc_hd__nand2_1 U22371 ( .A(n22747), .B(n25595), .Y(n15179) );
  sky130_fd_sc_hd__nand2_1 U22372 ( .A(n21924), .B(n28493), .Y(n15178) );
  sky130_fd_sc_hd__o211a_2 U22373 ( .A1(n26324), .A2(n11186), .B1(n15179), 
        .C1(n15178), .X(n15190) );
  sky130_fd_sc_hd__nand2_1 U22374 ( .A(n15488), .B(n15181), .Y(n15635) );
  sky130_fd_sc_hd__nor2_1 U22375 ( .A(n15639), .B(n15635), .Y(n15183) );
  sky130_fd_sc_hd__inv_1 U22376 ( .A(n15381), .Y(n15487) );
  sky130_fd_sc_hd__a21oi_1 U22377 ( .A1(n15487), .A2(n15181), .B1(n15180), .Y(
        n15636) );
  sky130_fd_sc_hd__a21oi_1 U22379 ( .A1(n17040), .A2(n15183), .B1(n15182), .Y(
        n15188) );
  sky130_fd_sc_hd__nand2_1 U22380 ( .A(n15186), .B(n15185), .Y(n15187) );
  sky130_fd_sc_hd__xor2_1 U22381 ( .A(n15188), .B(n15187), .X(n25601) );
  sky130_fd_sc_hd__nand2_1 U22382 ( .A(n25601), .B(n17225), .Y(n15189) );
  sky130_fd_sc_hd__nand2_1 U22383 ( .A(n15584), .B(n15341), .Y(n15201) );
  sky130_fd_sc_hd__o21ai_1 U22384 ( .A1(n15201), .A2(n15200), .B1(n19816), .Y(
        n15208) );
  sky130_fd_sc_hd__nand3_1 U22385 ( .A(n15230), .B(n15555), .C(n15495), .Y(
        n15203) );
  sky130_fd_sc_hd__nand3_1 U22386 ( .A(n15344), .B(n15504), .C(n15341), .Y(
        n15533) );
  sky130_fd_sc_hd__nand2_1 U22387 ( .A(n15307), .B(n15583), .Y(n15505) );
  sky130_fd_sc_hd__o31a_1 U22388 ( .A1(n19131), .A2(n15533), .A3(n15505), .B1(
        n17237), .X(n15202) );
  sky130_fd_sc_hd__a21oi_1 U22389 ( .A1(n21103), .A2(n15203), .B1(n15202), .Y(
        n15207) );
  sky130_fd_sc_hd__and3_1 U22390 ( .A(n15277), .B(n15583), .C(n15598), .X(
        n15204) );
  sky130_fd_sc_hd__nand4_1 U22391 ( .A(n15588), .B(n15204), .C(n15283), .D(
        n15566), .Y(n15205) );
  sky130_fd_sc_hd__nand3_1 U22393 ( .A(n15208), .B(n15207), .C(n15206), .Y(
        n15209) );
  sky130_fd_sc_hd__nand2_1 U22394 ( .A(n15209), .B(n15516), .Y(n15241) );
  sky130_fd_sc_hd__nand2_1 U22395 ( .A(n15307), .B(n15295), .Y(n15226) );
  sky130_fd_sc_hd__nand2_1 U22396 ( .A(n15226), .B(n17237), .Y(n15215) );
  sky130_fd_sc_hd__a21oi_1 U22397 ( .A1(n15277), .A2(n15225), .B1(n19726), .Y(
        n15210) );
  sky130_fd_sc_hd__a21oi_1 U22398 ( .A1(n15211), .A2(n19804), .B1(n15210), .Y(
        n15214) );
  sky130_fd_sc_hd__nand4b_1 U22399 ( .A_N(n15232), .B(n15502), .C(n15557), .D(
        n15328), .Y(n15212) );
  sky130_fd_sc_hd__nand2_1 U22400 ( .A(n15212), .B(n21103), .Y(n15213) );
  sky130_fd_sc_hd__nand3_1 U22401 ( .A(n15215), .B(n15214), .C(n15213), .Y(
        n15217) );
  sky130_fd_sc_hd__nand2_1 U22402 ( .A(n21103), .B(n20196), .Y(n15216) );
  sky130_fd_sc_hd__nand3_1 U22404 ( .A(n15599), .B(n15295), .C(n15277), .Y(
        n15218) );
  sky130_fd_sc_hd__nor2_1 U22405 ( .A(n15219), .B(n15218), .Y(n15582) );
  sky130_fd_sc_hd__nand2_1 U22406 ( .A(n15582), .B(n15570), .Y(n15220) );
  sky130_fd_sc_hd__nand2_1 U22407 ( .A(n15220), .B(n19804), .Y(n15224) );
  sky130_fd_sc_hd__a2bb2oi_1 U22408 ( .B1(n19816), .B2(n15339), .A1_N(n15410), 
        .A2_N(n15508), .Y(n15223) );
  sky130_fd_sc_hd__o21ai_1 U22409 ( .A1(n15595), .A2(n15221), .B1(n21103), .Y(
        n15222) );
  sky130_fd_sc_hd__nand3_1 U22410 ( .A(n15224), .B(n15223), .C(n15222), .Y(
        n15237) );
  sky130_fd_sc_hd__nand2b_1 U22411 ( .A_N(n15225), .B(n19119), .Y(n15536) );
  sky130_fd_sc_hd__nand4b_1 U22412 ( .A_N(n15294), .B(n15283), .C(n15509), .D(
        n15536), .Y(n15227) );
  sky130_fd_sc_hd__nand3_1 U22414 ( .A(n15589), .B(n15532), .C(n15504), .Y(
        n15293) );
  sky130_fd_sc_hd__nand3_1 U22415 ( .A(n15498), .B(n15228), .C(n15283), .Y(
        n15229) );
  sky130_fd_sc_hd__nand2_1 U22416 ( .A(n15229), .B(n21103), .Y(n15234) );
  sky130_fd_sc_hd__nand4_1 U22417 ( .A(n15230), .B(n15570), .C(n15557), .D(
        n20520), .Y(n15231) );
  sky130_fd_sc_hd__nand2_1 U22418 ( .A(n15231), .B(n19816), .Y(n15521) );
  sky130_fd_sc_hd__nand4_1 U22420 ( .A(n15235), .B(n15234), .C(n15521), .D(
        n15233), .Y(n15236) );
  sky130_fd_sc_hd__a22oi_1 U22421 ( .A1(n15237), .A2(n15610), .B1(n15236), 
        .B2(n16205), .Y(n15238) );
  sky130_fd_sc_hd__nand4_1 U22422 ( .A(n15241), .B(n15240), .C(n15239), .D(
        n15238), .Y(n15242) );
  sky130_fd_sc_hd__nand2_1 U22423 ( .A(n15242), .B(n21629), .Y(n15253) );
  sky130_fd_sc_hd__nand2_1 U22424 ( .A(n20759), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[87]), .Y(n15249) );
  sky130_fd_sc_hd__nand2_1 U22425 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[23]), .Y(n15248) );
  sky130_fd_sc_hd__nand3_1 U22426 ( .A(n15249), .B(n21768), .C(n15248), .Y(
        n15245) );
  sky130_fd_sc_hd__nand2_1 U22427 ( .A(n20540), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[55]), .Y(n15244) );
  sky130_fd_sc_hd__nand2_1 U22428 ( .A(n21513), .B(j202_soc_core_uart_div1[7]), 
        .Y(n15243) );
  sky130_fd_sc_hd__nand2_1 U22429 ( .A(n15244), .B(n15243), .Y(n15250) );
  sky130_fd_sc_hd__nor2_1 U22430 ( .A(n15245), .B(n15250), .Y(n15246) );
  sky130_fd_sc_hd__nand2_1 U22431 ( .A(n20786), .B(
        j202_soc_core_bldc_core_00_pwm_duty[11]), .Y(n15252) );
  sky130_fd_sc_hd__nand2_1 U22433 ( .A(j202_soc_core_memory0_ram_dout0[503]), 
        .B(n21650), .Y(n15255) );
  sky130_fd_sc_hd__nand3_1 U22434 ( .A(n15249), .B(n21653), .C(n15248), .Y(
        n15251) );
  sky130_fd_sc_hd__nor2_1 U22435 ( .A(n15251), .B(n15250), .Y(n15254) );
  sky130_fd_sc_hd__nand4_1 U22436 ( .A(n15255), .B(n15254), .C(n15253), .D(
        n15252), .Y(n15256) );
  sky130_fd_sc_hd__nor2_1 U22437 ( .A(n15258), .B(n15631), .Y(n15259) );
  sky130_fd_sc_hd__xnor2_1 U22438 ( .A(n15260), .B(n15259), .Y(n25247) );
  sky130_fd_sc_hd__nand2_1 U22439 ( .A(n22747), .B(n25247), .Y(n15262) );
  sky130_fd_sc_hd__nand2_1 U22440 ( .A(n21924), .B(n25230), .Y(n15261) );
  sky130_fd_sc_hd__o211a_2 U22441 ( .A1(n26431), .A2(n11186), .B1(n15262), 
        .C1(n15261), .X(n15267) );
  sky130_fd_sc_hd__a21oi_1 U22442 ( .A1(n17040), .A2(n16545), .B1(n16555), .Y(
        n15265) );
  sky130_fd_sc_hd__nand2_1 U22443 ( .A(n15263), .B(n16014), .Y(n15264) );
  sky130_fd_sc_hd__xor2_1 U22444 ( .A(n15265), .B(n15264), .X(n25252) );
  sky130_fd_sc_hd__nand2_1 U22445 ( .A(n25252), .B(n17225), .Y(n15266) );
  sky130_fd_sc_hd__o21a_1 U22446 ( .A1(n15270), .A2(n15269), .B1(n15563), .X(
        n15271) );
  sky130_fd_sc_hd__nand3_1 U22447 ( .A(n15272), .B(n15271), .C(n15585), .Y(
        n15511) );
  sky130_fd_sc_hd__o21ai_1 U22448 ( .A1(n15273), .A2(n15511), .B1(n19816), .Y(
        n15289) );
  sky130_fd_sc_hd__o31a_1 U22449 ( .A1(n15605), .A2(n15537), .A3(n15275), .B1(
        n21103), .X(n15276) );
  sky130_fd_sc_hd__a21oi_1 U22450 ( .A1(n15564), .A2(n15525), .B1(n15276), .Y(
        n15288) );
  sky130_fd_sc_hd__nand3_1 U22451 ( .A(n15278), .B(n20603), .C(n15277), .Y(
        n15279) );
  sky130_fd_sc_hd__nor2_1 U22452 ( .A(n15280), .B(n15279), .Y(n15281) );
  sky130_fd_sc_hd__nand2_1 U22453 ( .A(n15540), .B(n15281), .Y(n15282) );
  sky130_fd_sc_hd__nand2_1 U22454 ( .A(n15282), .B(n19804), .Y(n15287) );
  sky130_fd_sc_hd__nand3_1 U22455 ( .A(n15570), .B(n15283), .C(n15304), .Y(
        n15285) );
  sky130_fd_sc_hd__nand4_1 U22457 ( .A(n15289), .B(n15288), .C(n15287), .D(
        n15286), .Y(n15290) );
  sky130_fd_sc_hd__nand2_1 U22458 ( .A(n15290), .B(n15516), .Y(n15363) );
  sky130_fd_sc_hd__nand2_1 U22459 ( .A(n15499), .B(n15589), .Y(n15292) );
  sky130_fd_sc_hd__o21ai_1 U22460 ( .A1(n15292), .A2(n15291), .B1(n17237), .Y(
        n15316) );
  sky130_fd_sc_hd__nand2_1 U22462 ( .A(n15295), .B(n15328), .Y(n15296) );
  sky130_fd_sc_hd__nand2_1 U22463 ( .A(n15296), .B(n19804), .Y(n15297) );
  sky130_fd_sc_hd__nand2_1 U22464 ( .A(n15298), .B(n15297), .Y(n15522) );
  sky130_fd_sc_hd__o31a_1 U22465 ( .A1(n15301), .A2(n15300), .A3(n15299), .B1(
        n19804), .X(n15302) );
  sky130_fd_sc_hd__nor2_1 U22466 ( .A(n15522), .B(n15302), .Y(n15315) );
  sky130_fd_sc_hd__nand2_1 U22467 ( .A(n15303), .B(n17237), .Y(n16655) );
  sky130_fd_sc_hd__nor2_1 U22468 ( .A(n15595), .B(n15305), .Y(n15306) );
  sky130_fd_sc_hd__nand4_1 U22469 ( .A(n15307), .B(n15559), .C(n15306), .D(
        n15535), .Y(n15308) );
  sky130_fd_sc_hd__a22oi_1 U22470 ( .A1(n20235), .A2(n15309), .B1(n15308), 
        .B2(n21103), .Y(n15314) );
  sky130_fd_sc_hd__nand3_1 U22471 ( .A(n15310), .B(n15557), .C(n15341), .Y(
        n15312) );
  sky130_fd_sc_hd__o21ai_1 U22472 ( .A1(n15312), .A2(n15311), .B1(n19816), .Y(
        n15313) );
  sky130_fd_sc_hd__nand4_1 U22473 ( .A(n15316), .B(n15315), .C(n15314), .D(
        n15313), .Y(n15338) );
  sky130_fd_sc_hd__nand3_1 U22474 ( .A(n15317), .B(n15547), .C(n15341), .Y(
        n15318) );
  sky130_fd_sc_hd__o21ai_1 U22475 ( .A1(n15318), .A2(n15564), .B1(n19804), .Y(
        n15334) );
  sky130_fd_sc_hd__nand3_1 U22476 ( .A(n15319), .B(n15555), .C(n15547), .Y(
        n15320) );
  sky130_fd_sc_hd__nor2_1 U22477 ( .A(n15321), .B(n15320), .Y(n15322) );
  sky130_fd_sc_hd__nand4_1 U22478 ( .A(n15540), .B(n15322), .C(n15499), .D(
        n15559), .Y(n15323) );
  sky130_fd_sc_hd__nand2_1 U22479 ( .A(n15323), .B(n17237), .Y(n15333) );
  sky130_fd_sc_hd__nand2b_1 U22480 ( .A_N(n19120), .B(n21103), .Y(n16654) );
  sky130_fd_sc_hd__nor2_1 U22481 ( .A(n15596), .B(n15597), .Y(n15324) );
  sky130_fd_sc_hd__nand4_1 U22482 ( .A(n15590), .B(n15325), .C(n15324), .D(
        n15568), .Y(n15326) );
  sky130_fd_sc_hd__a22oi_1 U22483 ( .A1(n13199), .A2(n15666), .B1(n15326), 
        .B2(n19816), .Y(n15332) );
  sky130_fd_sc_hd__nand2_1 U22484 ( .A(n15597), .B(n13179), .Y(n15556) );
  sky130_fd_sc_hd__nand4_1 U22485 ( .A(n15328), .B(n15556), .C(n15327), .D(
        n15508), .Y(n15330) );
  sky130_fd_sc_hd__nand4_1 U22487 ( .A(n15334), .B(n15333), .C(n15332), .D(
        n15331), .Y(n15335) );
  sky130_fd_sc_hd__nand2_1 U22488 ( .A(n15335), .B(n15577), .Y(n15336) );
  sky130_fd_sc_hd__o31ai_1 U22489 ( .A1(n20485), .A2(n16986), .A3(n19728), 
        .B1(n15336), .Y(n15337) );
  sky130_fd_sc_hd__a21oi_1 U22490 ( .A1(n15338), .A2(n16205), .B1(n15337), .Y(
        n15362) );
  sky130_fd_sc_hd__nor2_1 U22491 ( .A(n15340), .B(n15339), .Y(n15343) );
  sky130_fd_sc_hd__nand4_1 U22492 ( .A(n15343), .B(n15342), .C(n15557), .D(
        n15341), .Y(n15345) );
  sky130_fd_sc_hd__nand3_1 U22493 ( .A(n15344), .B(n15589), .C(n15599), .Y(
        n15351) );
  sky130_fd_sc_hd__or3_1 U22494 ( .A(n15345), .B(n15604), .C(n15351), .X(
        n15346) );
  sky130_fd_sc_hd__nand2_1 U22495 ( .A(n15346), .B(n19816), .Y(n15359) );
  sky130_fd_sc_hd__nor2_1 U22496 ( .A(n15526), .B(n15602), .Y(n15552) );
  sky130_fd_sc_hd__nor2_1 U22497 ( .A(n15595), .B(n15347), .Y(n15348) );
  sky130_fd_sc_hd__nand4_1 U22498 ( .A(n15552), .B(n15348), .C(n15559), .D(
        n15583), .Y(n15349) );
  sky130_fd_sc_hd__nand2_1 U22499 ( .A(n15349), .B(n21103), .Y(n15358) );
  sky130_fd_sc_hd__o21ai_1 U22500 ( .A1(n15351), .A2(n15350), .B1(n19804), .Y(
        n15357) );
  sky130_fd_sc_hd__nor2_1 U22501 ( .A(n15526), .B(n15352), .Y(n15353) );
  sky130_fd_sc_hd__nand4_1 U22502 ( .A(n15353), .B(n15570), .C(n15504), .D(
        n15562), .Y(n15355) );
  sky130_fd_sc_hd__nand4_1 U22504 ( .A(n15359), .B(n15358), .C(n15357), .D(
        n15356), .Y(n15360) );
  sky130_fd_sc_hd__nand2_1 U22505 ( .A(n15360), .B(n15610), .Y(n15361) );
  sky130_fd_sc_hd__nand3_1 U22506 ( .A(n15363), .B(n15362), .C(n15361), .Y(
        n15364) );
  sky130_fd_sc_hd__nand2_1 U22507 ( .A(n15364), .B(n21629), .Y(n15368) );
  sky130_fd_sc_hd__a22oi_1 U22508 ( .A1(n21516), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[20]), .B1(n20540), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[52]), .Y(n15367) );
  sky130_fd_sc_hd__a22oi_1 U22509 ( .A1(n20759), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[84]), .B1(n21513), .B2(
        j202_soc_core_uart_div1[4]), .Y(n15366) );
  sky130_fd_sc_hd__nand2_1 U22510 ( .A(n20786), .B(
        j202_soc_core_bldc_core_00_pwm_duty[8]), .Y(n15365) );
  sky130_fd_sc_hd__nand4_1 U22511 ( .A(n15368), .B(n15367), .C(n15366), .D(
        n15365), .Y(n15369) );
  sky130_fd_sc_hd__a21oi_1 U22512 ( .A1(j202_soc_core_memory0_ram_dout0[500]), 
        .A2(n11207), .B1(n15369), .Y(n15375) );
  sky130_fd_sc_hd__a22oi_1 U22513 ( .A1(j202_soc_core_memory0_ram_dout0[244]), 
        .A2(j202_soc_core_memory0_ram_dout0_sel[7]), .B1(n20455), .B2(
        j202_soc_core_memory0_ram_dout0[212]), .Y(n15373) );
  sky130_fd_sc_hd__nand2_1 U22514 ( .A(j202_soc_core_memory0_ram_dout0[84]), 
        .B(n20458), .Y(n15371) );
  sky130_fd_sc_hd__nand4_1 U22515 ( .A(n15373), .B(n15372), .C(n15370), .D(
        n15371), .Y(n15374) );
  sky130_fd_sc_hd__nor2_1 U22516 ( .A(n15376), .B(n21026), .Y(n15483) );
  sky130_fd_sc_hd__nand2_1 U22517 ( .A(n15483), .B(
        j202_soc_core_j22_cpu_pc[19]), .Y(n15377) );
  sky130_fd_sc_hd__xor2_1 U22518 ( .A(n15377), .B(n22322), .X(n25666) );
  sky130_fd_sc_hd__o22a_1 U22519 ( .A1(n28506), .A2(n22743), .B1(n27383), .B2(
        n11186), .X(n15378) );
  sky130_fd_sc_hd__a21oi_1 U22521 ( .A1(n25666), .A2(n22747), .B1(n15379), .Y(
        n15390) );
  sky130_fd_sc_hd__nor2_1 U22522 ( .A(n15489), .B(n15380), .Y(n15383) );
  sky130_fd_sc_hd__o21ai_1 U22523 ( .A1(n15489), .A2(n15381), .B1(n15490), .Y(
        n15382) );
  sky130_fd_sc_hd__a21oi_1 U22524 ( .A1(n17040), .A2(n15383), .B1(n15382), .Y(
        n15388) );
  sky130_fd_sc_hd__nand2_1 U22525 ( .A(n15386), .B(n15385), .Y(n15387) );
  sky130_fd_sc_hd__xor2_1 U22526 ( .A(n15388), .B(n15387), .X(n25674) );
  sky130_fd_sc_hd__nand2_1 U22527 ( .A(n25674), .B(n17225), .Y(n15389) );
  sky130_fd_sc_hd__nand4_1 U22528 ( .A(n19440), .B(n19783), .C(n19814), .D(
        n19729), .Y(n15392) );
  sky130_fd_sc_hd__nor2_1 U22529 ( .A(n15392), .B(n15391), .Y(n15406) );
  sky130_fd_sc_hd__o2bb2ai_1 U22530 ( .B1(n15394), .B2(n19504), .A1_N(n18699), 
        .A2_N(n19810), .Y(n19778) );
  sky130_fd_sc_hd__nand4_1 U22531 ( .A(n15395), .B(n19695), .C(n19801), .D(
        n19778), .Y(n15401) );
  sky130_fd_sc_hd__nand2_1 U22532 ( .A(n19810), .B(n15396), .Y(n15397) );
  sky130_fd_sc_hd__nor2_1 U22533 ( .A(n15397), .B(n15409), .Y(n15398) );
  sky130_fd_sc_hd__nand4_1 U22534 ( .A(n15398), .B(n19813), .C(n19432), .D(
        n19770), .Y(n15399) );
  sky130_fd_sc_hd__nor2_1 U22535 ( .A(n19698), .B(n15399), .Y(n19830) );
  sky130_fd_sc_hd__nand3_1 U22536 ( .A(n19830), .B(n19518), .C(n19812), .Y(
        n15400) );
  sky130_fd_sc_hd__a22oi_1 U22537 ( .A1(n15401), .A2(n19816), .B1(n15400), 
        .B2(n21103), .Y(n15405) );
  sky130_fd_sc_hd__nand2_1 U22538 ( .A(n18695), .B(n18764), .Y(n18694) );
  sky130_fd_sc_hd__nor2_1 U22539 ( .A(n21145), .B(n18694), .Y(n18751) );
  sky130_fd_sc_hd__nand2_1 U22540 ( .A(n18751), .B(n15684), .Y(n19734) );
  sky130_fd_sc_hd__nand2_1 U22541 ( .A(n19771), .B(n19734), .Y(n15402) );
  sky130_fd_sc_hd__nor2_1 U22542 ( .A(n15402), .B(n19821), .Y(n19768) );
  sky130_fd_sc_hd__nand3_1 U22543 ( .A(n19715), .B(n19753), .C(n19809), .Y(
        n19699) );
  sky130_fd_sc_hd__nand3_1 U22544 ( .A(n19768), .B(n19719), .C(n19744), .Y(
        n15447) );
  sky130_fd_sc_hd__o21ai_1 U22545 ( .A1(n15403), .A2(n15447), .B1(n17237), .Y(
        n15404) );
  sky130_fd_sc_hd__o211ai_1 U22546 ( .A1(n12089), .A2(n15406), .B1(n15405), 
        .C1(n15404), .Y(n15407) );
  sky130_fd_sc_hd__nand2_1 U22547 ( .A(n15407), .B(n20126), .Y(n15465) );
  sky130_fd_sc_hd__nand4_1 U22548 ( .A(n19738), .B(n19707), .C(n19811), .D(
        n19777), .Y(n15408) );
  sky130_fd_sc_hd__nand2_1 U22549 ( .A(n19801), .B(n19714), .Y(n15450) );
  sky130_fd_sc_hd__nand2b_1 U22550 ( .A_N(n15450), .B(n19467), .Y(n19817) );
  sky130_fd_sc_hd__o21ai_1 U22551 ( .A1(n15408), .A2(n19817), .B1(n19816), .Y(
        n15418) );
  sky130_fd_sc_hd__nor2_1 U22552 ( .A(n19507), .B(n15409), .Y(n15436) );
  sky130_fd_sc_hd__nand2_1 U22553 ( .A(n19825), .B(n19814), .Y(n19761) );
  sky130_fd_sc_hd__nand2b_1 U22554 ( .A_N(n19733), .B(n19765), .Y(n19482) );
  sky130_fd_sc_hd__nor4b_1 U22555 ( .D_N(n15436), .A(n19716), .B(n19761), .C(
        n19482), .Y(n15411) );
  sky130_fd_sc_hd__a2bb2oi_1 U22556 ( .B1(n19486), .B2(n15412), .A1_N(n15411), 
        .A2_N(n15410), .Y(n15417) );
  sky130_fd_sc_hd__nor2_1 U22557 ( .A(n19507), .B(n15413), .Y(n15429) );
  sky130_fd_sc_hd__nand4_1 U22558 ( .A(n19441), .B(n19512), .C(n15429), .D(
        n19770), .Y(n15414) );
  sky130_fd_sc_hd__nand2_1 U22559 ( .A(n15414), .B(n21103), .Y(n15416) );
  sky130_fd_sc_hd__nand4_1 U22560 ( .A(n19765), .B(n19754), .C(n19782), .D(
        n19728), .Y(n19732) );
  sky130_fd_sc_hd__o21ai_0 U22561 ( .A1(n19797), .A2(n19732), .B1(n19804), .Y(
        n15415) );
  sky130_fd_sc_hd__nand4_1 U22562 ( .A(n15418), .B(n15417), .C(n15416), .D(
        n15415), .Y(n15419) );
  sky130_fd_sc_hd__nand2_1 U22563 ( .A(n15419), .B(n20196), .Y(n15464) );
  sky130_fd_sc_hd__nor2_1 U22564 ( .A(n15420), .B(n19521), .Y(n15421) );
  sky130_fd_sc_hd__nand4b_1 U22565 ( .A_N(n15422), .B(n15421), .C(n19754), .D(
        n19812), .Y(n15423) );
  sky130_fd_sc_hd__and3_1 U22566 ( .A(n19777), .B(n19734), .C(n19782), .X(
        n15456) );
  sky130_fd_sc_hd__nand3_1 U22567 ( .A(n19759), .B(n15456), .C(n19770), .Y(
        n19696) );
  sky130_fd_sc_hd__o21ai_1 U22568 ( .A1(n15423), .A2(n19696), .B1(n19816), .Y(
        n15445) );
  sky130_fd_sc_hd__o211ai_1 U22569 ( .A1(n20810), .A2(n18694), .B1(n19774), 
        .C1(n15425), .Y(n15427) );
  sky130_fd_sc_hd__o21ai_1 U22570 ( .A1(n15427), .A2(n15426), .B1(n19804), .Y(
        n15444) );
  sky130_fd_sc_hd__nor2_1 U22571 ( .A(n19699), .B(n15428), .Y(n19496) );
  sky130_fd_sc_hd__nand4_1 U22572 ( .A(n19706), .B(n15430), .C(n15429), .D(
        n19782), .Y(n15432) );
  sky130_fd_sc_hd__nand2_1 U22573 ( .A(n19764), .B(n15431), .Y(n19819) );
  sky130_fd_sc_hd__nor2_1 U22574 ( .A(n15432), .B(n19819), .Y(n15433) );
  sky130_fd_sc_hd__nand2_1 U22575 ( .A(n19496), .B(n15433), .Y(n15434) );
  sky130_fd_sc_hd__nand2_1 U22576 ( .A(n15434), .B(n17237), .Y(n15443) );
  sky130_fd_sc_hd__nor2_1 U22577 ( .A(n19521), .B(n15435), .Y(n15437) );
  sky130_fd_sc_hd__nand3_1 U22578 ( .A(n19715), .B(n15437), .C(n15436), .Y(
        n15439) );
  sky130_fd_sc_hd__nor2_1 U22579 ( .A(n15439), .B(n15438), .Y(n15440) );
  sky130_fd_sc_hd__nand2_1 U22580 ( .A(n19481), .B(n15440), .Y(n15441) );
  sky130_fd_sc_hd__nand2_1 U22581 ( .A(n15441), .B(n21103), .Y(n15442) );
  sky130_fd_sc_hd__nand4_1 U22582 ( .A(n15445), .B(n15444), .C(n15443), .D(
        n15442), .Y(n15446) );
  sky130_fd_sc_hd__nand2_1 U22583 ( .A(n15446), .B(n20235), .Y(n15463) );
  sky130_fd_sc_hd__nand3_1 U22584 ( .A(n19801), .B(n19490), .C(n19781), .Y(
        n15448) );
  sky130_fd_sc_hd__nor2_1 U22586 ( .A(n19708), .B(n19516), .Y(n15449) );
  sky130_fd_sc_hd__nand4b_1 U22587 ( .A_N(n15450), .B(n15449), .C(n19767), .D(
        n15456), .Y(n15454) );
  sky130_fd_sc_hd__nand2_1 U22588 ( .A(n19712), .B(n21145), .Y(n15451) );
  sky130_fd_sc_hd__nand3_1 U22589 ( .A(n19810), .B(n19782), .C(n15451), .Y(
        n15452) );
  sky130_fd_sc_hd__nand3_1 U22590 ( .A(n19715), .B(n19432), .C(n19753), .Y(
        n19742) );
  sky130_fd_sc_hd__nand2_1 U22591 ( .A(n19693), .B(n19734), .Y(n19700) );
  sky130_fd_sc_hd__nor3_1 U22592 ( .A(n15452), .B(n19742), .C(n19700), .Y(
        n15453) );
  sky130_fd_sc_hd__a2bb2oi_1 U22593 ( .B1(n21103), .B2(n15454), .A1_N(n12089), 
        .A2_N(n15453), .Y(n15459) );
  sky130_fd_sc_hd__nor2_1 U22594 ( .A(n19797), .B(n19779), .Y(n19721) );
  sky130_fd_sc_hd__nor2_1 U22595 ( .A(n15455), .B(n19795), .Y(n19450) );
  sky130_fd_sc_hd__nand3_1 U22596 ( .A(n19721), .B(n15456), .C(n19450), .Y(
        n15457) );
  sky130_fd_sc_hd__nand2_1 U22597 ( .A(n15457), .B(n19816), .Y(n15458) );
  sky130_fd_sc_hd__nand3_1 U22598 ( .A(n15460), .B(n15459), .C(n15458), .Y(
        n15461) );
  sky130_fd_sc_hd__nand2_1 U22599 ( .A(n15461), .B(n20194), .Y(n15462) );
  sky130_fd_sc_hd__nand4_1 U22600 ( .A(n15465), .B(n15464), .C(n15463), .D(
        n15462), .Y(n15466) );
  sky130_fd_sc_hd__nand2_1 U22601 ( .A(n15466), .B(n21629), .Y(n15479) );
  sky130_fd_sc_hd__nand2_1 U22602 ( .A(n20759), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[83]), .Y(n15474) );
  sky130_fd_sc_hd__nand2_1 U22603 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[19]), .Y(n15473) );
  sky130_fd_sc_hd__nand3_1 U22604 ( .A(n15474), .B(n21768), .C(n15473), .Y(
        n15469) );
  sky130_fd_sc_hd__nand2_1 U22605 ( .A(n20540), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[51]), .Y(n15468) );
  sky130_fd_sc_hd__nand2_1 U22606 ( .A(n21513), .B(j202_soc_core_uart_div1[3]), 
        .Y(n15467) );
  sky130_fd_sc_hd__nand2_1 U22607 ( .A(n15468), .B(n15467), .Y(n15472) );
  sky130_fd_sc_hd__nor2_1 U22608 ( .A(n15469), .B(n15472), .Y(n15470) );
  sky130_fd_sc_hd__nand2_1 U22609 ( .A(n20786), .B(
        j202_soc_core_bldc_core_00_pwm_duty[7]), .Y(n15476) );
  sky130_fd_sc_hd__nand2_1 U22610 ( .A(j202_soc_core_memory0_ram_dout0[499]), 
        .B(n21650), .Y(n15481) );
  sky130_fd_sc_hd__nand4_1 U22611 ( .A(n15475), .B(n21653), .C(n15474), .D(
        n15473), .Y(n15478) );
  sky130_fd_sc_hd__nor2_1 U22612 ( .A(n15478), .B(n15477), .Y(n15480) );
  sky130_fd_sc_hd__nand3_1 U22613 ( .A(n15481), .B(n15480), .C(n15479), .Y(
        n15482) );
  sky130_fd_sc_hd__xnor2_1 U22614 ( .A(n15484), .B(n15483), .Y(n25710) );
  sky130_fd_sc_hd__nand2_1 U22615 ( .A(n22747), .B(n25710), .Y(n15486) );
  sky130_fd_sc_hd__nand2_1 U22616 ( .A(n21924), .B(n25692), .Y(n15485) );
  sky130_fd_sc_hd__nand2_1 U22618 ( .A(n15491), .B(n15490), .Y(n15492) );
  sky130_fd_sc_hd__xor2_1 U22619 ( .A(n15493), .B(n15492), .X(n25715) );
  sky130_fd_sc_hd__nand2_1 U22620 ( .A(n25715), .B(n17225), .Y(n15494) );
  sky130_fd_sc_hd__nand2_1 U22621 ( .A(n15495), .B(n15508), .Y(n15496) );
  sky130_fd_sc_hd__nor2_1 U22622 ( .A(n21359), .B(n15547), .Y(n15580) );
  sky130_fd_sc_hd__nor2_1 U22623 ( .A(n15496), .B(n15580), .Y(n15497) );
  sky130_fd_sc_hd__nand3_1 U22624 ( .A(n15499), .B(n15498), .C(n15497), .Y(
        n15500) );
  sky130_fd_sc_hd__nor3_1 U22625 ( .A(n15501), .B(n15505), .C(n15500), .Y(
        n15515) );
  sky130_fd_sc_hd__nand4_1 U22626 ( .A(n15503), .B(n15502), .C(n15563), .D(
        n15590), .Y(n15507) );
  sky130_fd_sc_hd__nand3b_1 U22627 ( .A_N(n15505), .B(n15584), .C(n15504), .Y(
        n15506) );
  sky130_fd_sc_hd__a22oi_1 U22628 ( .A1(n15507), .A2(n21103), .B1(n15506), 
        .B2(n17237), .Y(n15514) );
  sky130_fd_sc_hd__nand3b_1 U22629 ( .A_N(n15510), .B(n15509), .C(n15508), .Y(
        n15512) );
  sky130_fd_sc_hd__o211ai_1 U22631 ( .A1(n15515), .A2(n12089), .B1(n15514), 
        .C1(n15513), .Y(n15517) );
  sky130_fd_sc_hd__nand2_1 U22632 ( .A(n15517), .B(n15516), .Y(n15614) );
  sky130_fd_sc_hd__o21ai_1 U22633 ( .A1(n15519), .A2(n15518), .B1(n21103), .Y(
        n15520) );
  sky130_fd_sc_hd__nand2_1 U22634 ( .A(n15521), .B(n15520), .Y(n15523) );
  sky130_fd_sc_hd__nor2_1 U22635 ( .A(n15523), .B(n15522), .Y(n15545) );
  sky130_fd_sc_hd__nand2_1 U22636 ( .A(n15584), .B(n15598), .Y(n15524) );
  sky130_fd_sc_hd__nand2_1 U22637 ( .A(n15524), .B(n19816), .Y(n15530) );
  sky130_fd_sc_hd__nand2_1 U22638 ( .A(n15526), .B(n15525), .Y(n15529) );
  sky130_fd_sc_hd__nor2_1 U22639 ( .A(n15527), .B(n16654), .Y(n15560) );
  sky130_fd_sc_hd__nand3_1 U22640 ( .A(n15530), .B(n15529), .C(n15528), .Y(
        n15531) );
  sky130_fd_sc_hd__a21oi_1 U22641 ( .A1(n15549), .A2(n19486), .B1(n15531), .Y(
        n15544) );
  sky130_fd_sc_hd__nand2_1 U22642 ( .A(n15585), .B(n15532), .Y(n15548) );
  sky130_fd_sc_hd__nand2b_1 U22643 ( .A_N(n15548), .B(n15570), .Y(n15534) );
  sky130_fd_sc_hd__o21ai_1 U22644 ( .A1(n15534), .A2(n15533), .B1(n19804), .Y(
        n15543) );
  sky130_fd_sc_hd__nand2_1 U22645 ( .A(n15536), .B(n15535), .Y(n15538) );
  sky130_fd_sc_hd__nor2_1 U22646 ( .A(n15538), .B(n15537), .Y(n15539) );
  sky130_fd_sc_hd__nand3_1 U22647 ( .A(n15540), .B(n15539), .C(n15559), .Y(
        n15541) );
  sky130_fd_sc_hd__nand2_1 U22648 ( .A(n15541), .B(n17237), .Y(n15542) );
  sky130_fd_sc_hd__nand4_1 U22649 ( .A(n15545), .B(n15544), .C(n15543), .D(
        n15542), .Y(n15579) );
  sky130_fd_sc_hd__nand3_1 U22650 ( .A(n15590), .B(n15547), .C(n15546), .Y(
        n15550) );
  sky130_fd_sc_hd__nor3_1 U22651 ( .A(n15550), .B(n15549), .C(n15548), .Y(
        n15551) );
  sky130_fd_sc_hd__nand2_1 U22652 ( .A(n15552), .B(n15551), .Y(n15553) );
  sky130_fd_sc_hd__nand2_1 U22653 ( .A(n15553), .B(n17237), .Y(n15576) );
  sky130_fd_sc_hd__and4_1 U22654 ( .A(n15556), .B(n15555), .C(n15598), .D(
        n15554), .X(n15558) );
  sky130_fd_sc_hd__nand3_1 U22655 ( .A(n15559), .B(n15558), .C(n15557), .Y(
        n15561) );
  sky130_fd_sc_hd__a21oi_1 U22656 ( .A1(n15561), .A2(n21103), .B1(n15560), .Y(
        n15575) );
  sky130_fd_sc_hd__nand3_1 U22657 ( .A(n15567), .B(n15563), .C(n15562), .Y(
        n15565) );
  sky130_fd_sc_hd__o21ai_1 U22658 ( .A1(n15565), .A2(n15564), .B1(n19804), .Y(
        n15574) );
  sky130_fd_sc_hd__nand2_1 U22659 ( .A(n15567), .B(n15566), .Y(n15572) );
  sky130_fd_sc_hd__nand4_1 U22660 ( .A(n15570), .B(n15569), .C(n15568), .D(
        n15585), .Y(n15571) );
  sky130_fd_sc_hd__o21ai_1 U22661 ( .A1(n15572), .A2(n15571), .B1(n19816), .Y(
        n15573) );
  sky130_fd_sc_hd__nand4_1 U22662 ( .A(n15576), .B(n15575), .C(n15574), .D(
        n15573), .Y(n15578) );
  sky130_fd_sc_hd__a22oi_1 U22663 ( .A1(n15579), .A2(n16205), .B1(n15578), 
        .B2(n15577), .Y(n15613) );
  sky130_fd_sc_hd__a31oi_1 U22664 ( .A1(n15582), .A2(n15598), .A3(n15581), 
        .B1(n12089), .Y(n15609) );
  sky130_fd_sc_hd__and3_1 U22665 ( .A(n15585), .B(n15584), .C(n15583), .X(
        n15586) );
  sky130_fd_sc_hd__nand3_1 U22666 ( .A(n15588), .B(n15587), .C(n15586), .Y(
        n15592) );
  sky130_fd_sc_hd__a21oi_1 U22667 ( .A1(n15590), .A2(n15589), .B1(n19468), .Y(
        n15591) );
  sky130_fd_sc_hd__a21oi_1 U22668 ( .A1(n15592), .A2(n17237), .B1(n15591), .Y(
        n15608) );
  sky130_fd_sc_hd__nor3_1 U22669 ( .A(n15595), .B(n15594), .C(n15593), .Y(
        n15601) );
  sky130_fd_sc_hd__a21oi_1 U22670 ( .A1(n15597), .A2(n19119), .B1(n15596), .Y(
        n15600) );
  sky130_fd_sc_hd__nand4_1 U22671 ( .A(n15601), .B(n15600), .C(n15599), .D(
        n15598), .Y(n15603) );
  sky130_fd_sc_hd__o21ai_1 U22672 ( .A1(n15603), .A2(n15602), .B1(n21103), .Y(
        n15607) );
  sky130_fd_sc_hd__nand4b_1 U22674 ( .A_N(n15609), .B(n15608), .C(n15607), .D(
        n15606), .Y(n15611) );
  sky130_fd_sc_hd__nand2_1 U22675 ( .A(n15611), .B(n15610), .Y(n15612) );
  sky130_fd_sc_hd__nand3_1 U22676 ( .A(n15614), .B(n15613), .C(n15612), .Y(
        n15615) );
  sky130_fd_sc_hd__nand2_1 U22677 ( .A(n15615), .B(n21629), .Y(n15626) );
  sky130_fd_sc_hd__nand2_1 U22678 ( .A(n20759), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[85]), .Y(n15622) );
  sky130_fd_sc_hd__nand2_1 U22679 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[21]), .Y(n15621) );
  sky130_fd_sc_hd__nand3_1 U22680 ( .A(n15622), .B(n21768), .C(n15621), .Y(
        n15618) );
  sky130_fd_sc_hd__nand2_1 U22681 ( .A(n20540), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[53]), .Y(n15617) );
  sky130_fd_sc_hd__nand2_1 U22682 ( .A(n21513), .B(j202_soc_core_uart_div1[5]), 
        .Y(n15616) );
  sky130_fd_sc_hd__nand2_1 U22683 ( .A(n15617), .B(n15616), .Y(n15623) );
  sky130_fd_sc_hd__nor2_1 U22684 ( .A(n15618), .B(n15623), .Y(n15619) );
  sky130_fd_sc_hd__nand2_1 U22685 ( .A(n20786), .B(
        j202_soc_core_bldc_core_00_pwm_duty[9]), .Y(n15625) );
  sky130_fd_sc_hd__nand3_1 U22686 ( .A(n15626), .B(n15619), .C(n15625), .Y(
        n15620) );
  sky130_fd_sc_hd__nand2_1 U22687 ( .A(j202_soc_core_memory0_ram_dout0[501]), 
        .B(n21650), .Y(n15628) );
  sky130_fd_sc_hd__nand3_1 U22688 ( .A(n15622), .B(n21653), .C(n15621), .Y(
        n15624) );
  sky130_fd_sc_hd__nor2_1 U22689 ( .A(n15624), .B(n15623), .Y(n15627) );
  sky130_fd_sc_hd__nand4_1 U22690 ( .A(n15628), .B(n15627), .C(n15626), .D(
        n15625), .Y(n15629) );
  sky130_fd_sc_hd__nand2_1 U22692 ( .A(n22226), .B(n22739), .Y(n15645) );
  sky130_fd_sc_hd__o22ai_1 U22693 ( .A1(n13047), .A2(n13365), .B1(n26280), 
        .B2(n11186), .Y(n15632) );
  sky130_fd_sc_hd__a21oi_1 U22694 ( .A1(n22701), .A2(n28499), .B1(n15632), .Y(
        n15634) );
  sky130_fd_sc_hd__nand2_1 U22695 ( .A(n22702), .B(n28499), .Y(n15633) );
  sky130_fd_sc_hd__a21oi_1 U22696 ( .A1(n17040), .A2(n15638), .B1(n15637), .Y(
        n15643) );
  sky130_fd_sc_hd__nand2_1 U22697 ( .A(n15641), .B(n15640), .Y(n15642) );
  sky130_fd_sc_hd__xor2_1 U22698 ( .A(n15643), .B(n15642), .X(n25385) );
  sky130_fd_sc_hd__nand2_1 U22699 ( .A(n25385), .B(n17225), .Y(n15644) );
  sky130_fd_sc_hd__a21oi_1 U22700 ( .A1(n29746), .A2(
        j202_soc_core_j22_cpu_ifetchl), .B1(j202_soc_core_j22_cpu_id_op2_v_), 
        .Y(n15653) );
  sky130_fd_sc_hd__nand2_1 U22701 ( .A(n15647), .B(n15646), .Y(n23885) );
  sky130_fd_sc_hd__nand2_1 U22702 ( .A(j202_soc_core_j22_cpu_opst[3]), .B(
        j202_soc_core_j22_cpu_opst[2]), .Y(n15649) );
  sky130_fd_sc_hd__nand2_1 U22703 ( .A(n23413), .B(n28355), .Y(n15648) );
  sky130_fd_sc_hd__nor2_1 U22704 ( .A(n15649), .B(n15648), .Y(n28401) );
  sky130_fd_sc_hd__nand2_1 U22705 ( .A(n28401), .B(n28373), .Y(n28071) );
  sky130_fd_sc_hd__nand3_1 U22706 ( .A(n15650), .B(
        j202_soc_core_j22_cpu_opst[0]), .C(n23413), .Y(n24394) );
  sky130_fd_sc_hd__nand2_1 U22707 ( .A(n28071), .B(n24394), .Y(n28340) );
  sky130_fd_sc_hd__nor2_1 U22708 ( .A(j202_soc_core_j22_cpu_opst[3]), .B(
        n23413), .Y(n22011) );
  sky130_fd_sc_hd__nor2_1 U22709 ( .A(j202_soc_core_j22_cpu_opst[0]), .B(
        j202_soc_core_j22_cpu_opst[2]), .Y(n28085) );
  sky130_fd_sc_hd__nand2_1 U22710 ( .A(n22011), .B(n28085), .Y(n24703) );
  sky130_fd_sc_hd__nand2_1 U22711 ( .A(n24703), .B(n15651), .Y(n24418) );
  sky130_fd_sc_hd__nand2_1 U22712 ( .A(n24418), .B(
        j202_soc_core_j22_cpu_opst[1]), .Y(n24540) );
  sky130_fd_sc_hd__nand2_1 U22713 ( .A(n23413), .B(
        j202_soc_core_j22_cpu_opst[1]), .Y(n28072) );
  sky130_fd_sc_hd__nor2_1 U22714 ( .A(n20428), .B(n28072), .Y(n23417) );
  sky130_fd_sc_hd__nand2_1 U22715 ( .A(n23417), .B(n28402), .Y(n23998) );
  sky130_fd_sc_hd__nand4b_1 U22716 ( .A_N(n28340), .B(n28103), .C(n24540), .D(
        n23998), .Y(n15652) );
  sky130_fd_sc_hd__nand2_1 U22717 ( .A(n28109), .B(
        j202_soc_core_j22_cpu_pc_hold), .Y(n24704) );
  sky130_fd_sc_hd__o22ai_1 U22718 ( .A1(n15653), .A2(n23885), .B1(n15652), 
        .B2(n24704), .Y(n29484) );
  sky130_fd_sc_hd__nand3_1 U22719 ( .A(n24647), .B(
        j202_soc_core_j22_cpu_memop_MEM__0_), .C(n12040), .Y(n24303) );
  sky130_fd_sc_hd__nand2_1 U22720 ( .A(n15654), .B(n12040), .Y(n24300) );
  sky130_fd_sc_hd__nand3_1 U22721 ( .A(n24590), .B(n24587), .C(
        j202_soc_core_j22_cpu_memop_MEM__3_), .Y(n23963) );
  sky130_fd_sc_hd__o21a_1 U22722 ( .A1(n24590), .A2(n24300), .B1(n23963), .X(
        n18855) );
  sky130_fd_sc_hd__nand2_1 U22723 ( .A(j202_soc_core_j22_cpu_memop_MEM__3_), 
        .B(j202_soc_core_j22_cpu_memop_MEM__1_), .Y(n23961) );
  sky130_fd_sc_hd__nand3_1 U22724 ( .A(n15655), .B(n12041), .C(n24587), .Y(
        n24304) );
  sky130_fd_sc_hd__nand2_1 U22725 ( .A(n15656), .B(
        j202_soc_core_j22_cpu_memop_MEM__3_), .Y(n22779) );
  sky130_fd_sc_hd__nand2_1 U22726 ( .A(n24304), .B(n22779), .Y(n22452) );
  sky130_fd_sc_hd__nand2_1 U22728 ( .A(j202_soc_core_memory0_ram_dout0[61]), 
        .B(n21633), .Y(n15658) );
  sky130_fd_sc_hd__nand2_1 U22729 ( .A(j202_soc_core_memory0_ram_dout0[93]), 
        .B(n21642), .Y(n15660) );
  sky130_fd_sc_hd__nand2_1 U22730 ( .A(j202_soc_core_memory0_ram_dout0[157]), 
        .B(n21489), .Y(n15659) );
  sky130_fd_sc_hd__nand2_1 U22731 ( .A(j202_soc_core_memory0_ram_dout0[253]), 
        .B(n21641), .Y(n15662) );
  sky130_fd_sc_hd__nand2_1 U22732 ( .A(j202_soc_core_memory0_ram_dout0[317]), 
        .B(n21503), .Y(n15661) );
  sky130_fd_sc_hd__nand2_1 U22733 ( .A(j202_soc_core_memory0_ram_dout0[29]), 
        .B(n21639), .Y(n15663) );
  sky130_fd_sc_hd__a2bb2oi_1 U22734 ( .B1(j202_soc_core_uart_div0[5]), .B2(
        n21513), .A1_N(n21512), .A2_N(n15664), .Y(n15774) );
  sky130_fd_sc_hd__nand2b_1 U22735 ( .A_N(n21515), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[61]), .Y(n15773) );
  sky130_fd_sc_hd__nand2_1 U22736 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[29]), .Y(n15772) );
  sky130_fd_sc_hd__nand4_1 U22737 ( .A(n15774), .B(n21768), .C(n15773), .D(
        n15772), .Y(n15695) );
  sky130_fd_sc_hd__nor2_1 U22738 ( .A(n15678), .B(n18730), .Y(n16638) );
  sky130_fd_sc_hd__nor2_1 U22739 ( .A(n19119), .B(n15665), .Y(n15696) );
  sky130_fd_sc_hd__nor2_1 U22740 ( .A(n15666), .B(n15696), .Y(n15705) );
  sky130_fd_sc_hd__nor2_1 U22741 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n14597), .Y(n21075) );
  sky130_fd_sc_hd__nand3_1 U22742 ( .A(n17241), .B(n21075), .C(n19119), .Y(
        n16349) );
  sky130_fd_sc_hd__nand2_1 U22743 ( .A(n15727), .B(n19130), .Y(n16686) );
  sky130_fd_sc_hd__nand3_1 U22744 ( .A(n15705), .B(n16655), .C(n16686), .Y(
        n15670) );
  sky130_fd_sc_hd__nand2_1 U22745 ( .A(n19124), .B(n21088), .Y(n20467) );
  sky130_fd_sc_hd__nand2b_1 U22746 ( .A_N(n20467), .B(n19148), .Y(n16663) );
  sky130_fd_sc_hd__nand2_1 U22747 ( .A(n11150), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n17108) );
  sky130_fd_sc_hd__nand2_1 U22748 ( .A(n20304), .B(n19148), .Y(n17269) );
  sky130_fd_sc_hd__nor2_1 U22749 ( .A(n17108), .B(n17269), .Y(n15733) );
  sky130_fd_sc_hd__nand2_1 U22750 ( .A(n15733), .B(n19119), .Y(n16989) );
  sky130_fd_sc_hd__nand2_1 U22751 ( .A(n16663), .B(n16989), .Y(n16981) );
  sky130_fd_sc_hd__nand2_1 U22752 ( .A(n19124), .B(n19804), .Y(n16963) );
  sky130_fd_sc_hd__nand2_1 U22753 ( .A(n19816), .B(n19119), .Y(n15667) );
  sky130_fd_sc_hd__nor2_1 U22754 ( .A(n15678), .B(n15667), .Y(n15718) );
  sky130_fd_sc_hd__nand2_1 U22755 ( .A(n15718), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n15699) );
  sky130_fd_sc_hd__nand2_1 U22756 ( .A(n16963), .B(n15699), .Y(n16575) );
  sky130_fd_sc_hd__nand2_1 U22757 ( .A(n21109), .B(n20464), .Y(n16960) );
  sky130_fd_sc_hd__nor2_1 U22758 ( .A(n20464), .B(n19130), .Y(n20210) );
  sky130_fd_sc_hd__nand2_1 U22759 ( .A(n16638), .B(n20210), .Y(n16577) );
  sky130_fd_sc_hd__nand2_1 U22760 ( .A(n16960), .B(n16577), .Y(n15730) );
  sky130_fd_sc_hd__nand3_1 U22761 ( .A(n15668), .B(n20374), .C(n19130), .Y(
        n16576) );
  sky130_fd_sc_hd__nor2_1 U22762 ( .A(n20464), .B(n11150), .Y(n19146) );
  sky130_fd_sc_hd__nand3_1 U22763 ( .A(n21075), .B(n18764), .C(n19146), .Y(
        n16372) );
  sky130_fd_sc_hd__nand2b_1 U22764 ( .A_N(n16372), .B(n19130), .Y(n16334) );
  sky130_fd_sc_hd__nand2_1 U22765 ( .A(n16576), .B(n16334), .Y(n15712) );
  sky130_fd_sc_hd__nor2_1 U22766 ( .A(n15730), .B(n15712), .Y(n15669) );
  sky130_fd_sc_hd__nand3_1 U22767 ( .A(n16623), .B(n16311), .C(n15669), .Y(
        n16608) );
  sky130_fd_sc_hd__nand2_1 U22768 ( .A(n19140), .B(n13199), .Y(n16950) );
  sky130_fd_sc_hd__o21a_1 U22769 ( .A1(n15670), .A2(n16608), .B1(n16980), .X(
        n15694) );
  sky130_fd_sc_hd__nand3_1 U22770 ( .A(n17241), .B(
        j202_soc_core_bootrom_00_address_w[4]), .C(n21075), .Y(n16573) );
  sky130_fd_sc_hd__nand2_1 U22771 ( .A(n15671), .B(n21088), .Y(n16617) );
  sky130_fd_sc_hd__nand2b_1 U22772 ( .A_N(n16985), .B(n15672), .Y(n16610) );
  sky130_fd_sc_hd__nand3_1 U22773 ( .A(n16617), .B(n16610), .C(n16577), .Y(
        n15673) );
  sky130_fd_sc_hd__nor2_1 U22774 ( .A(n21088), .B(n16346), .Y(n16679) );
  sky130_fd_sc_hd__nor2_1 U22775 ( .A(n15673), .B(n16679), .Y(n16657) );
  sky130_fd_sc_hd__nand2_1 U22776 ( .A(n21103), .B(n21359), .Y(n15674) );
  sky130_fd_sc_hd__nor2_1 U22777 ( .A(n15674), .B(n16985), .Y(n15697) );
  sky130_fd_sc_hd__nand2_1 U22778 ( .A(n15718), .B(n13179), .Y(n16694) );
  sky130_fd_sc_hd__nor2_1 U22779 ( .A(n15697), .B(n16642), .Y(n16990) );
  sky130_fd_sc_hd__nand2b_1 U22780 ( .A_N(n16356), .B(n15684), .Y(n15715) );
  sky130_fd_sc_hd__nand3_1 U22781 ( .A(n16657), .B(n16990), .C(n15715), .Y(
        n15680) );
  sky130_fd_sc_hd__nand2_1 U22782 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .B(j202_soc_core_bootrom_00_address_w[2]), .Y(n18731) );
  sky130_fd_sc_hd__nor2_1 U22783 ( .A(n18731), .B(n15677), .Y(n16637) );
  sky130_fd_sc_hd__nand2_1 U22784 ( .A(n16637), .B(n19130), .Y(n16678) );
  sky130_fd_sc_hd__nand2_1 U22785 ( .A(n16678), .B(n16654), .Y(n16945) );
  sky130_fd_sc_hd__nor2_1 U22786 ( .A(n16641), .B(n16945), .Y(n16965) );
  sky130_fd_sc_hd__nor2_1 U22787 ( .A(n19130), .B(n16372), .Y(n16376) );
  sky130_fd_sc_hd__nand2_1 U22788 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .B(n21088), .Y(n20200) );
  sky130_fd_sc_hd__nand2b_1 U22789 ( .A_N(n17100), .B(n20179), .Y(n19203) );
  sky130_fd_sc_hd__nor2_1 U22790 ( .A(n21088), .B(n15678), .Y(n20532) );
  sky130_fd_sc_hd__nand2_1 U22791 ( .A(n20532), .B(n20374), .Y(n16698) );
  sky130_fd_sc_hd__nand2_1 U22792 ( .A(n16689), .B(n16698), .Y(n15737) );
  sky130_fd_sc_hd__nor2_1 U22793 ( .A(n16376), .B(n15737), .Y(n15679) );
  sky130_fd_sc_hd__nand3_1 U22794 ( .A(n16623), .B(n16965), .C(n15679), .Y(
        n15749) );
  sky130_fd_sc_hd__o21a_1 U22795 ( .A1(n15680), .A2(n15749), .B1(n16994), .X(
        n15693) );
  sky130_fd_sc_hd__nand2_1 U22796 ( .A(n20532), .B(n21075), .Y(n17288) );
  sky130_fd_sc_hd__nor2_1 U22797 ( .A(n16637), .B(n16611), .Y(n15681) );
  sky130_fd_sc_hd__nand2_1 U22798 ( .A(n21102), .B(n19129), .Y(n16938) );
  sky130_fd_sc_hd__nand4_1 U22799 ( .A(n16314), .B(n15681), .C(n16372), .D(
        n16938), .Y(n15688) );
  sky130_fd_sc_hd__nor2_1 U22800 ( .A(n12089), .B(n16985), .Y(n15710) );
  sky130_fd_sc_hd__nor2_1 U22801 ( .A(n15710), .B(n15755), .Y(n15682) );
  sky130_fd_sc_hd__nor2_1 U22802 ( .A(n16206), .B(n17100), .Y(n15751) );
  sky130_fd_sc_hd__nand2_1 U22803 ( .A(n15751), .B(n21088), .Y(n17003) );
  sky130_fd_sc_hd__nand4_1 U22804 ( .A(n15682), .B(n15699), .C(n16959), .D(
        n17003), .Y(n16661) );
  sky130_fd_sc_hd__nor2_1 U22805 ( .A(n15747), .B(n15683), .Y(n16345) );
  sky130_fd_sc_hd__nand2_1 U22806 ( .A(n15684), .B(n11150), .Y(n19185) );
  sky130_fd_sc_hd__o22ai_1 U22807 ( .A1(n18700), .A2(n19185), .B1(n15685), 
        .B2(n16356), .Y(n15686) );
  sky130_fd_sc_hd__nor2_1 U22808 ( .A(n16345), .B(n15686), .Y(n15687) );
  sky130_fd_sc_hd__nand4_1 U22809 ( .A(n15687), .B(n16617), .C(n16694), .D(
        n16689), .Y(n16674) );
  sky130_fd_sc_hd__nor3_1 U22810 ( .A(n15688), .B(n16661), .C(n16674), .Y(
        n15691) );
  sky130_fd_sc_hd__nand4_1 U22811 ( .A(n17003), .B(n16694), .C(n16654), .D(
        n16577), .Y(n16336) );
  sky130_fd_sc_hd__nand4_1 U22812 ( .A(n16617), .B(n16576), .C(n15715), .D(
        n17288), .Y(n15689) );
  sky130_fd_sc_hd__nor3_1 U22813 ( .A(n16336), .B(n15689), .C(n16981), .Y(
        n15690) );
  sky130_fd_sc_hd__nand2_1 U22814 ( .A(n18744), .B(n13199), .Y(n17009) );
  sky130_fd_sc_hd__o22ai_1 U22815 ( .A1(n17007), .A2(n15691), .B1(n15690), 
        .B2(n17009), .Y(n15692) );
  sky130_fd_sc_hd__o31a_1 U22816 ( .A1(n15694), .A2(n15693), .A3(n15692), .B1(
        n20784), .X(n15771) );
  sky130_fd_sc_hd__nor2_1 U22817 ( .A(n15695), .B(n15771), .Y(n15770) );
  sky130_fd_sc_hd__nand2_1 U22818 ( .A(n15696), .B(n21088), .Y(n16987) );
  sky130_fd_sc_hd__nand2_1 U22819 ( .A(n19712), .B(n19130), .Y(n20814) );
  sky130_fd_sc_hd__nand2_1 U22820 ( .A(n16987), .B(n16321), .Y(n16310) );
  sky130_fd_sc_hd__nand2b_1 U22821 ( .A_N(n19120), .B(n19130), .Y(n16619) );
  sky130_fd_sc_hd__nand3_1 U22822 ( .A(n16619), .B(n16578), .C(n16372), .Y(
        n16341) );
  sky130_fd_sc_hd__nand2b_1 U22823 ( .A_N(n16356), .B(n20531), .Y(n17002) );
  sky130_fd_sc_hd__nand2_1 U22824 ( .A(n16637), .B(n21088), .Y(n16350) );
  sky130_fd_sc_hd__nand4_1 U22825 ( .A(n15719), .B(n17002), .C(n16689), .D(
        n16350), .Y(n15698) );
  sky130_fd_sc_hd__nor3_1 U22826 ( .A(n16310), .B(n16341), .C(n15698), .Y(
        n15704) );
  sky130_fd_sc_hd__nand3_1 U22827 ( .A(n15700), .B(n19148), .C(n17251), .Y(
        n16977) );
  sky130_fd_sc_hd__nand3_1 U22828 ( .A(n16655), .B(n16617), .C(n16977), .Y(
        n16609) );
  sky130_fd_sc_hd__nor2_1 U22829 ( .A(n16335), .B(n16609), .Y(n16326) );
  sky130_fd_sc_hd__nand4_1 U22830 ( .A(n16648), .B(n16960), .C(n16610), .D(
        n16989), .Y(n15701) );
  sky130_fd_sc_hd__nand4_1 U22831 ( .A(n17003), .B(n16694), .C(n16349), .D(
        n16654), .Y(n16597) );
  sky130_fd_sc_hd__nor2_1 U22832 ( .A(n15701), .B(n16597), .Y(n15702) );
  sky130_fd_sc_hd__nand2_1 U22833 ( .A(n16326), .B(n15702), .Y(n15703) );
  sky130_fd_sc_hd__nand2_1 U22834 ( .A(n15703), .B(n16980), .Y(n17010) );
  sky130_fd_sc_hd__o21a_1 U22835 ( .A1(n16950), .A2(n15704), .B1(n17010), .X(
        n15724) );
  sky130_fd_sc_hd__nor2_1 U22836 ( .A(n18731), .B(n16985), .Y(n15756) );
  sky130_fd_sc_hd__nor2_1 U22837 ( .A(n16631), .B(n15756), .Y(n16673) );
  sky130_fd_sc_hd__nand4_1 U22838 ( .A(n15705), .B(n16655), .C(n17003), .D(
        n16673), .Y(n15716) );
  sky130_fd_sc_hd__nand2b_1 U22839 ( .A_N(n16356), .B(n20464), .Y(n16632) );
  sky130_fd_sc_hd__nand3_1 U22840 ( .A(n16694), .B(n16632), .C(n16349), .Y(
        n15706) );
  sky130_fd_sc_hd__nor3_1 U22841 ( .A(n16341), .B(n15706), .C(n15737), .Y(
        n15707) );
  sky130_fd_sc_hd__nand3_1 U22842 ( .A(n16623), .B(n15708), .C(n15707), .Y(
        n15709) );
  sky130_fd_sc_hd__nand2_1 U22843 ( .A(n15709), .B(n16994), .Y(n15723) );
  sky130_fd_sc_hd__nand3_1 U22844 ( .A(n15715), .B(n15711), .C(n16577), .Y(
        n16983) );
  sky130_fd_sc_hd__nor3_1 U22845 ( .A(n15751), .B(n16983), .C(n16609), .Y(
        n16692) );
  sky130_fd_sc_hd__nand2_1 U22846 ( .A(n16367), .B(n16610), .Y(n16696) );
  sky130_fd_sc_hd__nand3_1 U22847 ( .A(n16689), .B(n16694), .C(n16346), .Y(
        n16976) );
  sky130_fd_sc_hd__nor2_1 U22848 ( .A(n16696), .B(n16976), .Y(n16582) );
  sky130_fd_sc_hd__nand3_1 U22849 ( .A(n16692), .B(n16582), .C(n15713), .Y(
        n15714) );
  sky130_fd_sc_hd__nand2_1 U22850 ( .A(n15714), .B(n16992), .Y(n15722) );
  sky130_fd_sc_hd__nand4_1 U22851 ( .A(n16576), .B(n16610), .C(n16573), .D(
        n15715), .Y(n15717) );
  sky130_fd_sc_hd__nor2_1 U22852 ( .A(n15717), .B(n15716), .Y(n16594) );
  sky130_fd_sc_hd__nand4_1 U22853 ( .A(n16594), .B(n15719), .C(n15736), .D(
        n17002), .Y(n15720) );
  sky130_fd_sc_hd__nand2_1 U22854 ( .A(n15720), .B(n17099), .Y(n15721) );
  sky130_fd_sc_hd__nand4_1 U22855 ( .A(n15724), .B(n15723), .C(n15722), .D(
        n15721), .Y(n15725) );
  sky130_fd_sc_hd__nand2_1 U22856 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .B(n21145), .Y(n20823) );
  sky130_fd_sc_hd__nand2_1 U22857 ( .A(n15725), .B(n20508), .Y(n15745) );
  sky130_fd_sc_hd__nand2_1 U22858 ( .A(n15756), .B(n21088), .Y(n16618) );
  sky130_fd_sc_hd__nand2_1 U22859 ( .A(n16618), .B(n16577), .Y(n15726) );
  sky130_fd_sc_hd__nor2_1 U22860 ( .A(n15726), .B(n16945), .Y(n16368) );
  sky130_fd_sc_hd__nand2_1 U22861 ( .A(n15727), .B(n21088), .Y(n16672) );
  sky130_fd_sc_hd__nand2_1 U22862 ( .A(n15759), .B(n16672), .Y(n15728) );
  sky130_fd_sc_hd__nand2_1 U22863 ( .A(n16350), .B(n16334), .Y(n16660) );
  sky130_fd_sc_hd__nor2_1 U22864 ( .A(n15728), .B(n16660), .Y(n16691) );
  sky130_fd_sc_hd__nand4_1 U22865 ( .A(n16368), .B(n16691), .C(n16644), .D(
        n16694), .Y(n15729) );
  sky130_fd_sc_hd__nand2_1 U22866 ( .A(n15729), .B(n16994), .Y(n15742) );
  sky130_fd_sc_hd__nor2_1 U22867 ( .A(n16700), .B(n15730), .Y(n15731) );
  sky130_fd_sc_hd__nand4_1 U22868 ( .A(n16965), .B(n16326), .C(n16644), .D(
        n15731), .Y(n15732) );
  sky130_fd_sc_hd__nand2_1 U22869 ( .A(n15732), .B(n17099), .Y(n15741) );
  sky130_fd_sc_hd__nor2_1 U22870 ( .A(n15737), .B(n16597), .Y(n15734) );
  sky130_fd_sc_hd__nand4_1 U22871 ( .A(n15734), .B(n16311), .C(n16657), .D(
        n16639), .Y(n15735) );
  sky130_fd_sc_hd__nand2_1 U22872 ( .A(n15735), .B(n16992), .Y(n15740) );
  sky130_fd_sc_hd__nand4_1 U22873 ( .A(n16672), .B(n16977), .C(n15736), .D(
        n16632), .Y(n15738) );
  sky130_fd_sc_hd__nand3_1 U22874 ( .A(n16617), .B(n16686), .C(n16578), .Y(
        n15754) );
  sky130_fd_sc_hd__o31ai_1 U22875 ( .A1(n15738), .A2(n15754), .A3(n15737), 
        .B1(n16980), .Y(n15739) );
  sky130_fd_sc_hd__nand4_1 U22876 ( .A(n15742), .B(n15741), .C(n15740), .D(
        n15739), .Y(n15743) );
  sky130_fd_sc_hd__nand2_1 U22877 ( .A(n21101), .B(
        j202_soc_core_bootrom_00_address_w[8]), .Y(n20858) );
  sky130_fd_sc_hd__nand2_1 U22878 ( .A(n15743), .B(n20505), .Y(n15744) );
  sky130_fd_sc_hd__nand2_1 U22879 ( .A(n15745), .B(n15744), .Y(n15746) );
  sky130_fd_sc_hd__nand2_1 U22880 ( .A(n15746), .B(n21629), .Y(n15780) );
  sky130_fd_sc_hd__nand3_1 U22881 ( .A(n16648), .B(n16672), .C(n16963), .Y(
        n16701) );
  sky130_fd_sc_hd__nor2_1 U22882 ( .A(n11150), .B(n15747), .Y(n19144) );
  sky130_fd_sc_hd__nand2_1 U22883 ( .A(n19144), .B(n21358), .Y(n20656) );
  sky130_fd_sc_hd__nand3_1 U22884 ( .A(n16326), .B(n15748), .C(n20656), .Y(
        n15750) );
  sky130_fd_sc_hd__o21ai_1 U22885 ( .A1(n15750), .A2(n15749), .B1(n16980), .Y(
        n15768) );
  sky130_fd_sc_hd__nand2_1 U22886 ( .A(n16694), .B(n16334), .Y(n15752) );
  sky130_fd_sc_hd__nand2_1 U22887 ( .A(n16374), .B(n19203), .Y(n16944) );
  sky130_fd_sc_hd__nor3_1 U22888 ( .A(n16631), .B(n15752), .C(n16944), .Y(
        n15753) );
  sky130_fd_sc_hd__nand4_1 U22889 ( .A(n15753), .B(n16663), .C(n16678), .D(
        n16618), .Y(n15757) );
  sky130_fd_sc_hd__nor2_1 U22890 ( .A(n15755), .B(n15754), .Y(n16636) );
  sky130_fd_sc_hd__nand2_1 U22891 ( .A(n15756), .B(n19130), .Y(n16988) );
  sky130_fd_sc_hd__nand3_1 U22892 ( .A(n16636), .B(n16672), .C(n16988), .Y(
        n16995) );
  sky130_fd_sc_hd__nand2_1 U22894 ( .A(n16655), .B(n16959), .Y(n16357) );
  sky130_fd_sc_hd__nor2_1 U22895 ( .A(n15758), .B(n16357), .Y(n16347) );
  sky130_fd_sc_hd__nand3_1 U22896 ( .A(n16618), .B(n15759), .C(n16334), .Y(
        n16943) );
  sky130_fd_sc_hd__nor2_1 U22897 ( .A(n16968), .B(n16983), .Y(n15760) );
  sky130_fd_sc_hd__nand4_1 U22898 ( .A(n16347), .B(n16636), .C(n16605), .D(
        n15760), .Y(n15761) );
  sky130_fd_sc_hd__nand2_1 U22899 ( .A(n15761), .B(n16992), .Y(n15766) );
  sky130_fd_sc_hd__nand3_1 U22900 ( .A(n16672), .B(n16632), .C(n17288), .Y(
        n15762) );
  sky130_fd_sc_hd__nor2_1 U22901 ( .A(n15762), .B(n16661), .Y(n16622) );
  sky130_fd_sc_hd__nand2_1 U22902 ( .A(n16960), .B(n20656), .Y(n16697) );
  sky130_fd_sc_hd__nor2_1 U22903 ( .A(n16697), .B(n16309), .Y(n15763) );
  sky130_fd_sc_hd__nand4_1 U22904 ( .A(n16622), .B(n16308), .C(n15763), .D(
        n19120), .Y(n15764) );
  sky130_fd_sc_hd__nand2_1 U22905 ( .A(n15764), .B(n16994), .Y(n15765) );
  sky130_fd_sc_hd__nand4_1 U22906 ( .A(n15768), .B(n15767), .C(n15766), .D(
        n15765), .Y(n15769) );
  sky130_fd_sc_hd__nor2_1 U22907 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .B(n21101), .Y(n16996) );
  sky130_fd_sc_hd__nand2_1 U22908 ( .A(n15769), .B(n20757), .Y(n15778) );
  sky130_fd_sc_hd__nand2_1 U22909 ( .A(j202_soc_core_memory0_ram_dout0[509]), 
        .B(n21650), .Y(n15782) );
  sky130_fd_sc_hd__nand3_1 U22910 ( .A(n15773), .B(n21653), .C(n15772), .Y(
        n15776) );
  sky130_fd_sc_hd__nor2_1 U22911 ( .A(n15776), .B(n15775), .Y(n15777) );
  sky130_fd_sc_hd__and3_1 U22912 ( .A(n15779), .B(n15778), .C(n15777), .X(
        n15781) );
  sky130_fd_sc_hd__nand3_1 U22913 ( .A(n15782), .B(n15781), .C(n15780), .Y(
        n19855) );
  sky130_fd_sc_hd__nand2_1 U22914 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[58]), .Y(n15787) );
  sky130_fd_sc_hd__nand2_1 U22915 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[250]), .Y(n15786) );
  sky130_fd_sc_hd__nand2_1 U22916 ( .A(n15783), .B(
        j202_soc_core_j22_cpu_rf_gpr[122]), .Y(n15785) );
  sky130_fd_sc_hd__nand2_1 U22917 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[505]), .Y(n15784) );
  sky130_fd_sc_hd__nand4_1 U22918 ( .A(n15787), .B(n15786), .C(n15785), .D(
        n15784), .Y(n15794) );
  sky130_fd_sc_hd__nand2_1 U22919 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[345]), .Y(n15792) );
  sky130_fd_sc_hd__nand2_1 U22920 ( .A(n15788), .B(
        j202_soc_core_j22_cpu_rf_gpr[473]), .Y(n15791) );
  sky130_fd_sc_hd__nand2_1 U22921 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[409]), .Y(n15790) );
  sky130_fd_sc_hd__nand2_1 U22922 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[441]), .Y(n15789) );
  sky130_fd_sc_hd__nand4_1 U22923 ( .A(n15792), .B(n15791), .C(n15790), .D(
        n15789), .Y(n15793) );
  sky130_fd_sc_hd__nor2_1 U22924 ( .A(n15794), .B(n15793), .Y(n15809) );
  sky130_fd_sc_hd__nor2_1 U22925 ( .A(n15795), .B(n14798), .Y(n15802) );
  sky130_fd_sc_hd__a21oi_1 U22926 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[26]), .B1(n14743), .Y(n15800) );
  sky130_fd_sc_hd__nand2_1 U22927 ( .A(n15796), .B(
        j202_soc_core_j22_cpu_rf_gpr[90]), .Y(n15799) );
  sky130_fd_sc_hd__nand2_1 U22928 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[154]), .Y(n15798) );
  sky130_fd_sc_hd__nand2_1 U22929 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[282]), .Y(n15797) );
  sky130_fd_sc_hd__nand4_1 U22930 ( .A(n15800), .B(n15799), .C(n15798), .D(
        n15797), .Y(n15801) );
  sky130_fd_sc_hd__nor2_1 U22931 ( .A(n15802), .B(n15801), .Y(n15808) );
  sky130_fd_sc_hd__nand2_1 U22932 ( .A(n11194), .B(
        j202_soc_core_j22_cpu_rf_gpr[314]), .Y(n15806) );
  sky130_fd_sc_hd__nand2_1 U22933 ( .A(n16410), .B(
        j202_soc_core_j22_cpu_rf_gpr[186]), .Y(n15805) );
  sky130_fd_sc_hd__nand2_1 U22934 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[377]), .Y(n15804) );
  sky130_fd_sc_hd__nand2_1 U22935 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[218]), .Y(n15803) );
  sky130_fd_sc_hd__and4_1 U22936 ( .A(n15806), .B(n15805), .C(n15804), .D(
        n15803), .X(n15807) );
  sky130_fd_sc_hd__nand3_1 U22937 ( .A(n15809), .B(n15808), .C(n15807), .Y(
        n27788) );
  sky130_fd_sc_hd__inv_2 U22938 ( .A(n27788), .Y(n27825) );
  sky130_fd_sc_hd__nand2_1 U22939 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[313]), .Y(n15813) );
  sky130_fd_sc_hd__nand2_1 U22940 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[281]), .Y(n15812) );
  sky130_fd_sc_hd__nand2_1 U22941 ( .A(n11195), .B(
        j202_soc_core_j22_cpu_rf_gpr[408]), .Y(n15811) );
  sky130_fd_sc_hd__nand2_1 U22942 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[440]), .Y(n15810) );
  sky130_fd_sc_hd__nand4_1 U22943 ( .A(n15813), .B(n15812), .C(n15811), .D(
        n15810), .Y(n15819) );
  sky130_fd_sc_hd__nand2_1 U22944 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[472]), .Y(n15817) );
  sky130_fd_sc_hd__nand2_1 U22945 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[57]), .Y(n15816) );
  sky130_fd_sc_hd__nand2_1 U22946 ( .A(n14985), .B(
        j202_soc_core_j22_cpu_rf_gpr[504]), .Y(n15815) );
  sky130_fd_sc_hd__nand2_1 U22947 ( .A(n15796), .B(
        j202_soc_core_j22_cpu_rf_gpr[89]), .Y(n15814) );
  sky130_fd_sc_hd__nand4_1 U22948 ( .A(n15817), .B(n15816), .C(n15815), .D(
        n15814), .Y(n15818) );
  sky130_fd_sc_hd__nor2_1 U22949 ( .A(n15819), .B(n15818), .Y(n15832) );
  sky130_fd_sc_hd__nand2_1 U22950 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[344]), .Y(n15823) );
  sky130_fd_sc_hd__nand2_1 U22951 ( .A(n16410), .B(
        j202_soc_core_j22_cpu_rf_gpr[185]), .Y(n15822) );
  sky130_fd_sc_hd__nand2_1 U22952 ( .A(n15783), .B(
        j202_soc_core_j22_cpu_rf_gpr[121]), .Y(n15821) );
  sky130_fd_sc_hd__nand2_1 U22953 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[217]), .Y(n15820) );
  sky130_fd_sc_hd__and4_1 U22954 ( .A(n15823), .B(n15822), .C(n15821), .D(
        n15820), .X(n15831) );
  sky130_fd_sc_hd__nor2_1 U22955 ( .A(n15888), .B(n14798), .Y(n15829) );
  sky130_fd_sc_hd__a21oi_1 U22956 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[25]), .B1(n14743), .Y(n15827) );
  sky130_fd_sc_hd__nand2_1 U22957 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[153]), .Y(n15826) );
  sky130_fd_sc_hd__nand2_1 U22958 ( .A(n16043), .B(
        j202_soc_core_j22_cpu_rf_gpr[249]), .Y(n15825) );
  sky130_fd_sc_hd__nand2_1 U22959 ( .A(n11196), .B(
        j202_soc_core_j22_cpu_rf_gpr[376]), .Y(n15824) );
  sky130_fd_sc_hd__nand4_1 U22960 ( .A(n15827), .B(n15826), .C(n15825), .D(
        n15824), .Y(n15828) );
  sky130_fd_sc_hd__nor2_1 U22961 ( .A(n15829), .B(n15828), .Y(n15830) );
  sky130_fd_sc_hd__nand3_1 U22962 ( .A(n15832), .B(n15831), .C(n15830), .Y(
        n27032) );
  sky130_fd_sc_hd__inv_2 U22963 ( .A(n27032), .Y(n27796) );
  sky130_fd_sc_hd__o22ai_1 U22964 ( .A1(n16501), .A2(n27825), .B1(n27796), 
        .B2(n16500), .Y(n16017) );
  sky130_fd_sc_hd__nand2_1 U22965 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[218]), .Y(n15836) );
  sky130_fd_sc_hd__nand2_1 U22966 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[473]), .Y(n15835) );
  sky130_fd_sc_hd__nand2_1 U22967 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[505]), .Y(n15834) );
  sky130_fd_sc_hd__nand2_1 U22968 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[250]), .Y(n15833) );
  sky130_fd_sc_hd__nand4_1 U22969 ( .A(n15836), .B(n15835), .C(n15834), .D(
        n15833), .Y(n15842) );
  sky130_fd_sc_hd__nand2_1 U22970 ( .A(n16506), .B(
        j202_soc_core_j22_cpu_rf_gpr[26]), .Y(n15840) );
  sky130_fd_sc_hd__nand2_1 U22971 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[90]), .Y(n15839) );
  sky130_fd_sc_hd__nand2_1 U22972 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[409]), .Y(n15838) );
  sky130_fd_sc_hd__nand2_1 U22973 ( .A(n23808), .B(
        j202_soc_core_j22_cpu_rf_gpr[154]), .Y(n15837) );
  sky130_fd_sc_hd__nand4_1 U22974 ( .A(n15840), .B(n15839), .C(n15838), .D(
        n15837), .Y(n15841) );
  sky130_fd_sc_hd__nor2_1 U22975 ( .A(n15842), .B(n15841), .Y(n15851) );
  sky130_fd_sc_hd__a22oi_1 U22976 ( .A1(n23776), .A2(
        j202_soc_core_j22_cpu_rf_gpr[377]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[282]), .Y(n15850) );
  sky130_fd_sc_hd__a22oi_1 U22977 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[58]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_rf_gpr[345]), .Y(n15849) );
  sky130_fd_sc_hd__nand2_1 U22978 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[314]), .Y(n15847) );
  sky130_fd_sc_hd__nand2_1 U22979 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[441]), .Y(n15846) );
  sky130_fd_sc_hd__nand2_1 U22980 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[186]), .Y(n15845) );
  sky130_fd_sc_hd__nand2_1 U22981 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[122]), .Y(n15844) );
  sky130_fd_sc_hd__and4_1 U22982 ( .A(n15847), .B(n15846), .C(n15845), .D(
        n15844), .X(n15848) );
  sky130_fd_sc_hd__nand4_1 U22983 ( .A(n15851), .B(n15850), .C(n15849), .D(
        n15848), .Y(n22662) );
  sky130_fd_sc_hd__nand2_1 U22984 ( .A(n22662), .B(n16523), .Y(n15862) );
  sky130_fd_sc_hd__o21ai_0 U22985 ( .A1(n15852), .A2(n16525), .B1(n16524), .Y(
        n15856) );
  sky130_fd_sc_hd__o22ai_1 U22986 ( .A1(n15854), .A2(n16077), .B1(n15853), 
        .B2(n14342), .Y(n15855) );
  sky130_fd_sc_hd__nor2_1 U22987 ( .A(n15856), .B(n15855), .Y(n15861) );
  sky130_fd_sc_hd__nand2_1 U22988 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[26]), .Y(n15860) );
  sky130_fd_sc_hd__nand2_1 U22989 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[26]), .Y(n15859) );
  sky130_fd_sc_hd__nand2_1 U22990 ( .A(n16533), .B(
        j202_soc_core_j22_cpu_pc[26]), .Y(n15858) );
  sky130_fd_sc_hd__nand2_1 U22991 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[26]), .Y(n15857) );
  sky130_fd_sc_hd__nand3_1 U22992 ( .A(n15862), .B(n15861), .C(n13107), .Y(
        n28471) );
  sky130_fd_sc_hd__nand2_1 U22993 ( .A(n28471), .B(n16541), .Y(n15863) );
  sky130_fd_sc_hd__o21ai_1 U22994 ( .A1(n16543), .A2(n28471), .B1(n15863), .Y(
        n16018) );
  sky130_fd_sc_hd__nor2_1 U22995 ( .A(n16017), .B(n16018), .Y(n16901) );
  sky130_fd_sc_hd__o22ai_1 U22996 ( .A1(n16501), .A2(n27796), .B1(n26323), 
        .B2(n16500), .Y(n16015) );
  sky130_fd_sc_hd__nand2_1 U22997 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[217]), .Y(n15867) );
  sky130_fd_sc_hd__nand2_1 U22998 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[472]), .Y(n15866) );
  sky130_fd_sc_hd__nand2_1 U22999 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[504]), .Y(n15865) );
  sky130_fd_sc_hd__nand2_1 U23000 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[249]), .Y(n15864) );
  sky130_fd_sc_hd__nand4_1 U23001 ( .A(n15867), .B(n15866), .C(n15865), .D(
        n15864), .Y(n15873) );
  sky130_fd_sc_hd__nand2_1 U23002 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[25]), .Y(n15871) );
  sky130_fd_sc_hd__nand2_1 U23003 ( .A(n15984), .B(
        j202_soc_core_j22_cpu_rf_gpr[89]), .Y(n15870) );
  sky130_fd_sc_hd__nand2_1 U23004 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[408]), .Y(n15869) );
  sky130_fd_sc_hd__nand2_1 U23005 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[153]), .Y(n15868) );
  sky130_fd_sc_hd__nand4_1 U23006 ( .A(n15871), .B(n15870), .C(n15869), .D(
        n15868), .Y(n15872) );
  sky130_fd_sc_hd__nor2_1 U23007 ( .A(n15873), .B(n15872), .Y(n15884) );
  sky130_fd_sc_hd__nand2_1 U23008 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[281]), .Y(n15877) );
  sky130_fd_sc_hd__nand2_1 U23009 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[57]), .Y(n15876) );
  sky130_fd_sc_hd__nand2_1 U23010 ( .A(n15991), .B(
        j202_soc_core_j22_cpu_rf_gpr[376]), .Y(n15875) );
  sky130_fd_sc_hd__nand2_1 U23011 ( .A(n16064), .B(
        j202_soc_core_j22_cpu_rf_gpr[344]), .Y(n15874) );
  sky130_fd_sc_hd__and4_1 U23012 ( .A(n15877), .B(n15876), .C(n15875), .D(
        n15874), .X(n15883) );
  sky130_fd_sc_hd__nand2_1 U23013 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[313]), .Y(n15881) );
  sky130_fd_sc_hd__nand2_1 U23014 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[440]), .Y(n15880) );
  sky130_fd_sc_hd__nand2_1 U23015 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[185]), .Y(n15879) );
  sky130_fd_sc_hd__nand2_1 U23016 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[121]), .Y(n15878) );
  sky130_fd_sc_hd__and4_1 U23017 ( .A(n15881), .B(n15880), .C(n15879), .D(
        n15878), .X(n15882) );
  sky130_fd_sc_hd__nand3_1 U23018 ( .A(n15884), .B(n15883), .C(n15882), .Y(
        n22908) );
  sky130_fd_sc_hd__o22a_1 U23019 ( .A1(n15888), .A2(n16488), .B1(n16487), .B2(
        n22905), .X(n15892) );
  sky130_fd_sc_hd__o22a_1 U23020 ( .A1(n15889), .A2(n16491), .B1(n16490), .B2(
        n22904), .X(n15891) );
  sky130_fd_sc_hd__a21oi_1 U23021 ( .A1(n11201), .A2(
        j202_soc_core_j22_cpu_rf_gpr[504]), .B1(n16493), .Y(n15890) );
  sky130_fd_sc_hd__nand4_1 U23022 ( .A(n15893), .B(n15892), .C(n15891), .D(
        n15890), .Y(n15894) );
  sky130_fd_sc_hd__nand2_1 U23023 ( .A(n26276), .B(n16086), .Y(n15895) );
  sky130_fd_sc_hd__nor2_1 U23025 ( .A(n16015), .B(n16016), .Y(n16299) );
  sky130_fd_sc_hd__nor2_1 U23026 ( .A(n16901), .B(n16299), .Y(n16020) );
  sky130_fd_sc_hd__nor2_1 U23027 ( .A(n16013), .B(n15896), .Y(n16892) );
  sky130_fd_sc_hd__nand2_1 U23028 ( .A(n16020), .B(n16892), .Y(n16544) );
  sky130_fd_sc_hd__nand2_1 U23029 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[156]), .Y(n15900) );
  sky130_fd_sc_hd__nand2_1 U23030 ( .A(n15796), .B(
        j202_soc_core_j22_cpu_rf_gpr[92]), .Y(n15899) );
  sky130_fd_sc_hd__nand2_1 U23031 ( .A(n11195), .B(
        j202_soc_core_j22_cpu_rf_gpr[411]), .Y(n15898) );
  sky130_fd_sc_hd__nand2_1 U23032 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[379]), .Y(n15897) );
  sky130_fd_sc_hd__nand4_1 U23033 ( .A(n15900), .B(n15899), .C(n15898), .D(
        n15897), .Y(n15906) );
  sky130_fd_sc_hd__nand2_1 U23034 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[284]), .Y(n15904) );
  sky130_fd_sc_hd__nand2_1 U23035 ( .A(n11194), .B(n12245), .Y(n15903) );
  sky130_fd_sc_hd__nand2_1 U23036 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[475]), .Y(n15902) );
  sky130_fd_sc_hd__nand2_1 U23037 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[443]), .Y(n15901) );
  sky130_fd_sc_hd__nand4_1 U23038 ( .A(n15904), .B(n15903), .C(n15902), .D(
        n15901), .Y(n15905) );
  sky130_fd_sc_hd__nor2_1 U23039 ( .A(n15906), .B(n15905), .Y(n15920) );
  sky130_fd_sc_hd__nand2_1 U23040 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[347]), .Y(n15911) );
  sky130_fd_sc_hd__nand2_1 U23041 ( .A(n16410), .B(
        j202_soc_core_j22_cpu_rf_gpr[188]), .Y(n15910) );
  sky130_fd_sc_hd__nand2_1 U23042 ( .A(n15783), .B(
        j202_soc_core_j22_cpu_rf_gpr[124]), .Y(n15909) );
  sky130_fd_sc_hd__nand2_1 U23043 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[220]), .Y(n15908) );
  sky130_fd_sc_hd__nor2_1 U23044 ( .A(n15912), .B(n14798), .Y(n15918) );
  sky130_fd_sc_hd__a21oi_1 U23045 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[28]), .B1(n14743), .Y(n15916) );
  sky130_fd_sc_hd__nand2_1 U23046 ( .A(n16043), .B(
        j202_soc_core_j22_cpu_rf_gpr[252]), .Y(n15915) );
  sky130_fd_sc_hd__nand2_1 U23047 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[507]), .Y(n15914) );
  sky130_fd_sc_hd__nand2_1 U23048 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[60]), .Y(n15913) );
  sky130_fd_sc_hd__nand4_1 U23049 ( .A(n15916), .B(n15915), .C(n15914), .D(
        n15913), .Y(n15917) );
  sky130_fd_sc_hd__nor2_1 U23050 ( .A(n15918), .B(n15917), .Y(n15919) );
  sky130_fd_sc_hd__nand2_1 U23051 ( .A(n16433), .B(
        j202_soc_core_j22_cpu_rf_gpr[219]), .Y(n15924) );
  sky130_fd_sc_hd__nand2_1 U23052 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[59]), .Y(n15923) );
  sky130_fd_sc_hd__nand2_1 U23053 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[506]), .Y(n15922) );
  sky130_fd_sc_hd__nand2_1 U23054 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[251]), .Y(n15921) );
  sky130_fd_sc_hd__nand4_1 U23055 ( .A(n15924), .B(n15923), .C(n15922), .D(
        n15921), .Y(n15931) );
  sky130_fd_sc_hd__nand2_1 U23056 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[187]), .Y(n15929) );
  sky130_fd_sc_hd__nand2_1 U23057 ( .A(n16432), .B(
        j202_soc_core_j22_cpu_rf_gpr[346]), .Y(n15928) );
  sky130_fd_sc_hd__nand2_1 U23058 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[378]), .Y(n15927) );
  sky130_fd_sc_hd__nand2_1 U23059 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[442]), .Y(n15926) );
  sky130_fd_sc_hd__nand4_1 U23060 ( .A(n15929), .B(n15928), .C(n15927), .D(
        n15926), .Y(n15930) );
  sky130_fd_sc_hd__nor2_1 U23061 ( .A(n15931), .B(n15930), .Y(n15945) );
  sky130_fd_sc_hd__nand2_1 U23062 ( .A(n15796), .B(
        j202_soc_core_j22_cpu_rf_gpr[91]), .Y(n15935) );
  sky130_fd_sc_hd__nand2_1 U23063 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[283]), .Y(n15934) );
  sky130_fd_sc_hd__nand2_1 U23064 ( .A(n16398), .B(
        j202_soc_core_j22_cpu_rf_gpr[123]), .Y(n15933) );
  sky130_fd_sc_hd__nand2_1 U23065 ( .A(n15788), .B(
        j202_soc_core_j22_cpu_rf_gpr[474]), .Y(n15932) );
  sky130_fd_sc_hd__nor2_1 U23066 ( .A(n15936), .B(n16444), .Y(n15943) );
  sky130_fd_sc_hd__a21oi_1 U23067 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[27]), .B1(n14743), .Y(n15941) );
  sky130_fd_sc_hd__nand2_1 U23068 ( .A(n11194), .B(
        j202_soc_core_j22_cpu_rf_gpr[315]), .Y(n15940) );
  sky130_fd_sc_hd__nand2_1 U23069 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[410]), .Y(n15939) );
  sky130_fd_sc_hd__nand2_1 U23070 ( .A(n16425), .B(
        j202_soc_core_j22_cpu_rf_gpr[155]), .Y(n15938) );
  sky130_fd_sc_hd__nand4_1 U23071 ( .A(n15941), .B(n15940), .C(n15939), .D(
        n15938), .Y(n15942) );
  sky130_fd_sc_hd__nor2_1 U23072 ( .A(n15943), .B(n15942), .Y(n15944) );
  sky130_fd_sc_hd__nand3_1 U23073 ( .A(n15945), .B(n13049), .C(n15944), .Y(
        n27042) );
  sky130_fd_sc_hd__nand2_1 U23075 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[220]), .Y(n15949) );
  sky130_fd_sc_hd__nand2_1 U23076 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[475]), .Y(n15948) );
  sky130_fd_sc_hd__nand2_1 U23077 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[507]), .Y(n15947) );
  sky130_fd_sc_hd__nand2_1 U23078 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[252]), .Y(n15946) );
  sky130_fd_sc_hd__nand4_1 U23079 ( .A(n15949), .B(n15948), .C(n15947), .D(
        n15946), .Y(n15957) );
  sky130_fd_sc_hd__nand2_1 U23080 ( .A(n16506), .B(
        j202_soc_core_j22_cpu_rf_gpr[28]), .Y(n15955) );
  sky130_fd_sc_hd__nand2_1 U23081 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[92]), .Y(n15954) );
  sky130_fd_sc_hd__nand2_1 U23082 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[411]), .Y(n15953) );
  sky130_fd_sc_hd__nand2_1 U23083 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[156]), .Y(n15952) );
  sky130_fd_sc_hd__nand4_1 U23084 ( .A(n15955), .B(n15954), .C(n15953), .D(
        n15952), .Y(n15956) );
  sky130_fd_sc_hd__nor2_1 U23085 ( .A(n15957), .B(n15956), .Y(n15965) );
  sky130_fd_sc_hd__a22oi_1 U23086 ( .A1(n23776), .A2(
        j202_soc_core_j22_cpu_rf_gpr[379]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[284]), .Y(n15964) );
  sky130_fd_sc_hd__a22oi_1 U23087 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[60]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_rf_gpr[347]), .Y(n15963) );
  sky130_fd_sc_hd__nand2_1 U23088 ( .A(n15958), .B(n12245), .Y(n15962) );
  sky130_fd_sc_hd__nand2_1 U23089 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[443]), .Y(n15961) );
  sky130_fd_sc_hd__nand2_1 U23090 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[188]), .Y(n15960) );
  sky130_fd_sc_hd__nand2_1 U23091 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[124]), .Y(n15959) );
  sky130_fd_sc_hd__nand4_1 U23092 ( .A(n15965), .B(n15964), .C(n15963), .D(
        n13067), .Y(n22644) );
  sky130_fd_sc_hd__nand2_1 U23093 ( .A(n22644), .B(n16523), .Y(n15976) );
  sky130_fd_sc_hd__o21ai_0 U23094 ( .A1(n15966), .A2(n16525), .B1(n16524), .Y(
        n15970) );
  sky130_fd_sc_hd__o22ai_1 U23095 ( .A1(n15968), .A2(n11202), .B1(n15967), 
        .B2(n14477), .Y(n15969) );
  sky130_fd_sc_hd__nor2_1 U23096 ( .A(n15970), .B(n15969), .Y(n15975) );
  sky130_fd_sc_hd__nand2_1 U23097 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[28]), .Y(n15974) );
  sky130_fd_sc_hd__nand2_1 U23098 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[28]), .Y(n15973) );
  sky130_fd_sc_hd__nand2_1 U23099 ( .A(n16533), .B(
        j202_soc_core_j22_cpu_pc[28]), .Y(n15972) );
  sky130_fd_sc_hd__nand2_1 U23100 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[28]), .Y(n15971) );
  sky130_fd_sc_hd__nand3_1 U23101 ( .A(n15976), .B(n15975), .C(n13091), .Y(
        n25825) );
  sky130_fd_sc_hd__nand2_1 U23102 ( .A(n25825), .B(n16541), .Y(n15977) );
  sky130_fd_sc_hd__nor2_1 U23104 ( .A(n16023), .B(n16024), .Y(n17041) );
  sky130_fd_sc_hd__o22ai_1 U23105 ( .A1(n16500), .A2(n27825), .B1(n27804), 
        .B2(n16501), .Y(n16021) );
  sky130_fd_sc_hd__nand2_1 U23106 ( .A(n13818), .B(
        j202_soc_core_j22_cpu_rf_gpr[219]), .Y(n15983) );
  sky130_fd_sc_hd__nand2_1 U23107 ( .A(n13819), .B(
        j202_soc_core_j22_cpu_rf_gpr[474]), .Y(n15982) );
  sky130_fd_sc_hd__nand2_1 U23108 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[506]), .Y(n15981) );
  sky130_fd_sc_hd__nand2_1 U23109 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[251]), .Y(n15980) );
  sky130_fd_sc_hd__nand4_1 U23110 ( .A(n15983), .B(n15982), .C(n15981), .D(
        n15980), .Y(n15990) );
  sky130_fd_sc_hd__nand2_1 U23111 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[27]), .Y(n15988) );
  sky130_fd_sc_hd__nand2_1 U23112 ( .A(n15984), .B(
        j202_soc_core_j22_cpu_rf_gpr[91]), .Y(n15987) );
  sky130_fd_sc_hd__nand2_1 U23113 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[410]), .Y(n15986) );
  sky130_fd_sc_hd__nand2_1 U23114 ( .A(n23808), .B(
        j202_soc_core_j22_cpu_rf_gpr[155]), .Y(n15985) );
  sky130_fd_sc_hd__nand4_1 U23115 ( .A(n15988), .B(n15987), .C(n15986), .D(
        n15985), .Y(n15989) );
  sky130_fd_sc_hd__nor2_1 U23116 ( .A(n15990), .B(n15989), .Y(n15999) );
  sky130_fd_sc_hd__a22oi_1 U23117 ( .A1(n15991), .A2(
        j202_soc_core_j22_cpu_rf_gpr[378]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[283]), .Y(n15998) );
  sky130_fd_sc_hd__a22oi_1 U23118 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[59]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_rf_gpr[346]), .Y(n15997) );
  sky130_fd_sc_hd__nand2_1 U23119 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[315]), .Y(n15996) );
  sky130_fd_sc_hd__nand2_1 U23120 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[442]), .Y(n15995) );
  sky130_fd_sc_hd__nand2_1 U23121 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[187]), .Y(n15994) );
  sky130_fd_sc_hd__nand2_1 U23122 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[123]), .Y(n15993) );
  sky130_fd_sc_hd__nand4_1 U23123 ( .A(n15999), .B(n15998), .C(n15997), .D(
        n13058), .Y(n22532) );
  sky130_fd_sc_hd__nand2_1 U23124 ( .A(n22532), .B(n16523), .Y(n16010) );
  sky130_fd_sc_hd__o21ai_0 U23125 ( .A1(n16000), .A2(n16525), .B1(n16524), .Y(
        n16004) );
  sky130_fd_sc_hd__o22ai_1 U23126 ( .A1(n16002), .A2(n11202), .B1(n30075), 
        .B2(n14477), .Y(n16003) );
  sky130_fd_sc_hd__nor2_1 U23127 ( .A(n16004), .B(n16003), .Y(n16009) );
  sky130_fd_sc_hd__nand2_1 U23128 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[27]), .Y(n16008) );
  sky130_fd_sc_hd__nand2_1 U23129 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[27]), .Y(n16007) );
  sky130_fd_sc_hd__nand2_1 U23130 ( .A(n16533), .B(
        j202_soc_core_j22_cpu_pc[27]), .Y(n16006) );
  sky130_fd_sc_hd__nand2_1 U23131 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[27]), .Y(n16005) );
  sky130_fd_sc_hd__nand3_1 U23132 ( .A(n16010), .B(n16009), .C(n13099), .Y(
        n28463) );
  sky130_fd_sc_hd__nand2_1 U23133 ( .A(n28463), .B(n16541), .Y(n16011) );
  sky130_fd_sc_hd__o21ai_1 U23134 ( .A1(n16543), .A2(n28463), .B1(n16011), .Y(
        n16022) );
  sky130_fd_sc_hd__nor2_1 U23135 ( .A(n16021), .B(n16022), .Y(n16194) );
  sky130_fd_sc_hd__nand2_1 U23136 ( .A(n17029), .B(n16718), .Y(n16026) );
  sky130_fd_sc_hd__nor2_1 U23137 ( .A(n16026), .B(n17030), .Y(n16028) );
  sky130_fd_sc_hd__nand2_1 U23138 ( .A(n16016), .B(n16015), .Y(n16893) );
  sky130_fd_sc_hd__nand2_1 U23139 ( .A(n16018), .B(n16017), .Y(n16902) );
  sky130_fd_sc_hd__a21oi_1 U23141 ( .A1(n16020), .A2(n16896), .B1(n16019), .Y(
        n16551) );
  sky130_fd_sc_hd__nand2_1 U23142 ( .A(n16022), .B(n16021), .Y(n17031) );
  sky130_fd_sc_hd__nand2_1 U23143 ( .A(n16024), .B(n16023), .Y(n17042) );
  sky130_fd_sc_hd__a21oi_1 U23145 ( .A1(n17034), .A2(n16718), .B1(n16720), .Y(
        n16025) );
  sky130_fd_sc_hd__o21ai_1 U23146 ( .A1(n16026), .A2(n17036), .B1(n16025), .Y(
        n16027) );
  sky130_fd_sc_hd__nand2_1 U23148 ( .A(n14986), .B(
        j202_soc_core_j22_cpu_rf_gpr[157]), .Y(n16032) );
  sky130_fd_sc_hd__nand2_1 U23149 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[93]), .Y(n16031) );
  sky130_fd_sc_hd__nand2_1 U23150 ( .A(n11195), .B(
        j202_soc_core_j22_cpu_rf_gpr[412]), .Y(n16030) );
  sky130_fd_sc_hd__nand2_1 U23151 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[380]), .Y(n16029) );
  sky130_fd_sc_hd__nand4_1 U23152 ( .A(n16032), .B(n16031), .C(n16030), .D(
        n16029), .Y(n16038) );
  sky130_fd_sc_hd__nand2_1 U23153 ( .A(n11197), .B(
        j202_soc_core_j22_cpu_rf_gpr[285]), .Y(n16036) );
  sky130_fd_sc_hd__nand2_1 U23154 ( .A(n11194), .B(
        j202_soc_core_j22_cpu_rf_gpr[316]), .Y(n16035) );
  sky130_fd_sc_hd__nand2_1 U23155 ( .A(n15788), .B(
        j202_soc_core_j22_cpu_rf_gpr[476]), .Y(n16034) );
  sky130_fd_sc_hd__nand2_1 U23156 ( .A(n15925), .B(
        j202_soc_core_j22_cpu_rf_gpr[444]), .Y(n16033) );
  sky130_fd_sc_hd__nand4_1 U23157 ( .A(n16036), .B(n16035), .C(n16034), .D(
        n16033), .Y(n16037) );
  sky130_fd_sc_hd__nor2_1 U23158 ( .A(n16038), .B(n16037), .Y(n16053) );
  sky130_fd_sc_hd__nand2_1 U23159 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[348]), .Y(n16042) );
  sky130_fd_sc_hd__nand2_1 U23160 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[189]), .Y(n16041) );
  sky130_fd_sc_hd__nand2_1 U23161 ( .A(n16398), .B(
        j202_soc_core_j22_cpu_rf_gpr[125]), .Y(n16040) );
  sky130_fd_sc_hd__nand2_1 U23162 ( .A(n16433), .B(
        j202_soc_core_j22_cpu_rf_gpr[221]), .Y(n16039) );
  sky130_fd_sc_hd__and4_1 U23163 ( .A(n16042), .B(n16041), .C(n16040), .D(
        n16039), .X(n16052) );
  sky130_fd_sc_hd__nor2_1 U23164 ( .A(n16080), .B(n16444), .Y(n16050) );
  sky130_fd_sc_hd__a21oi_1 U23165 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[29]), .B1(n14743), .Y(n16048) );
  sky130_fd_sc_hd__nand2_1 U23166 ( .A(n16043), .B(
        j202_soc_core_j22_cpu_rf_gpr[253]), .Y(n16047) );
  sky130_fd_sc_hd__nand2_1 U23167 ( .A(n13546), .B(
        j202_soc_core_j22_cpu_rf_gpr[508]), .Y(n16046) );
  sky130_fd_sc_hd__nand2_1 U23168 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[61]), .Y(n16045) );
  sky130_fd_sc_hd__nand4_1 U23169 ( .A(n16048), .B(n16047), .C(n16046), .D(
        n16045), .Y(n16049) );
  sky130_fd_sc_hd__nor2_1 U23170 ( .A(n16050), .B(n16049), .Y(n16051) );
  sky130_fd_sc_hd__nand3_1 U23171 ( .A(n16053), .B(n16052), .C(n16051), .Y(
        n27033) );
  sky130_fd_sc_hd__o22ai_1 U23172 ( .A1(n16501), .A2(n26296), .B1(n27026), 
        .B2(n16500), .Y(n16089) );
  sky130_fd_sc_hd__nand2_1 U23173 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[221]), .Y(n16057) );
  sky130_fd_sc_hd__nand2_1 U23174 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[476]), .Y(n16056) );
  sky130_fd_sc_hd__nand2_1 U23175 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[508]), .Y(n16055) );
  sky130_fd_sc_hd__nand2_1 U23176 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[253]), .Y(n16054) );
  sky130_fd_sc_hd__nand4_1 U23177 ( .A(n16057), .B(n16056), .C(n16055), .D(
        n16054), .Y(n16063) );
  sky130_fd_sc_hd__nand2_1 U23178 ( .A(n16506), .B(
        j202_soc_core_j22_cpu_rf_gpr[29]), .Y(n16061) );
  sky130_fd_sc_hd__nand2_1 U23179 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[93]), .Y(n16060) );
  sky130_fd_sc_hd__nand2_1 U23180 ( .A(n16466), .B(
        j202_soc_core_j22_cpu_rf_gpr[412]), .Y(n16059) );
  sky130_fd_sc_hd__nand2_1 U23181 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[157]), .Y(n16058) );
  sky130_fd_sc_hd__nand4_1 U23182 ( .A(n16061), .B(n16060), .C(n16059), .D(
        n16058), .Y(n16062) );
  sky130_fd_sc_hd__nor2_1 U23183 ( .A(n16063), .B(n16062), .Y(n16075) );
  sky130_fd_sc_hd__nand2_1 U23184 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[285]), .Y(n16068) );
  sky130_fd_sc_hd__nand2_1 U23185 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[61]), .Y(n16067) );
  sky130_fd_sc_hd__nand2_1 U23186 ( .A(n23776), .B(
        j202_soc_core_j22_cpu_rf_gpr[380]), .Y(n16066) );
  sky130_fd_sc_hd__nand2_1 U23187 ( .A(n16064), .B(
        j202_soc_core_j22_cpu_rf_gpr[348]), .Y(n16065) );
  sky130_fd_sc_hd__and4_1 U23188 ( .A(n16068), .B(n16067), .C(n16066), .D(
        n16065), .X(n16074) );
  sky130_fd_sc_hd__nand2_1 U23189 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[316]), .Y(n16072) );
  sky130_fd_sc_hd__nand2_1 U23190 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[444]), .Y(n16071) );
  sky130_fd_sc_hd__nand2_1 U23191 ( .A(n11199), .B(
        j202_soc_core_j22_cpu_rf_gpr[189]), .Y(n16070) );
  sky130_fd_sc_hd__nand2_1 U23192 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[125]), .Y(n16069) );
  sky130_fd_sc_hd__and4_1 U23193 ( .A(n16072), .B(n16071), .C(n16070), .D(
        n16069), .X(n16073) );
  sky130_fd_sc_hd__nand3_1 U23194 ( .A(n16075), .B(n16074), .C(n16073), .Y(
        n23011) );
  sky130_fd_sc_hd__o22a_1 U23195 ( .A1(n16078), .A2(n16077), .B1(n16076), .B2(
        n14342), .X(n16084) );
  sky130_fd_sc_hd__o22a_1 U23196 ( .A1(n16079), .A2(n16491), .B1(n16487), .B2(
        n23001), .X(n16083) );
  sky130_fd_sc_hd__o22a_1 U23197 ( .A1(n16080), .A2(n16488), .B1(n16490), .B2(
        n22999), .X(n16082) );
  sky130_fd_sc_hd__a21oi_1 U23198 ( .A1(n11201), .A2(
        j202_soc_core_j22_cpu_rf_gpr[508]), .B1(n16493), .Y(n16081) );
  sky130_fd_sc_hd__nand4_1 U23199 ( .A(n16084), .B(n16083), .C(n16082), .D(
        n16081), .Y(n16085) );
  sky130_fd_sc_hd__a21oi_1 U23200 ( .A1(n23011), .A2(n16523), .B1(n16085), .Y(
        n28451) );
  sky130_fd_sc_hd__nand2_1 U23201 ( .A(n28451), .B(n16086), .Y(n16087) );
  sky130_fd_sc_hd__nor2_1 U23203 ( .A(n16089), .B(n16090), .Y(n16723) );
  sky130_fd_sc_hd__nand2_1 U23204 ( .A(n16090), .B(n16089), .Y(n16721) );
  sky130_fd_sc_hd__nand2_1 U23205 ( .A(n16091), .B(n16721), .Y(n16092) );
  sky130_fd_sc_hd__o22a_1 U23207 ( .A1(n28451), .A2(n22743), .B1(n26296), .B2(
        n11186), .X(n16098) );
  sky130_fd_sc_hd__nor2_1 U23208 ( .A(n22725), .B(n16094), .Y(n16096) );
  sky130_fd_sc_hd__nand2_1 U23209 ( .A(n25465), .B(n22747), .Y(n16097) );
  sky130_fd_sc_hd__o211ai_1 U23210 ( .A1(n28451), .A2(n22745), .B1(n16098), 
        .C1(n16097), .Y(n16099) );
  sky130_fd_sc_hd__nand2_1 U23211 ( .A(j202_soc_core_memory0_ram_dout0[475]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n16104) );
  sky130_fd_sc_hd__nand2_1 U23212 ( .A(j202_soc_core_memory0_ram_dout0[251]), 
        .B(n21641), .Y(n16103) );
  sky130_fd_sc_hd__nand2_1 U23213 ( .A(j202_soc_core_memory0_ram_dout0[27]), 
        .B(n21639), .Y(n16102) );
  sky130_fd_sc_hd__nand2_1 U23214 ( .A(j202_soc_core_memory0_ram_dout0[315]), 
        .B(n21503), .Y(n16101) );
  sky130_fd_sc_hd__nand4_1 U23215 ( .A(n16104), .B(n16103), .C(n16102), .D(
        n16101), .Y(n16110) );
  sky130_fd_sc_hd__nand2_1 U23216 ( .A(j202_soc_core_memory0_ram_dout0[59]), 
        .B(n21633), .Y(n16108) );
  sky130_fd_sc_hd__nand2_1 U23217 ( .A(j202_soc_core_memory0_ram_dout0[347]), 
        .B(n21490), .Y(n16107) );
  sky130_fd_sc_hd__nand2_1 U23218 ( .A(j202_soc_core_memory0_ram_dout0[283]), 
        .B(n21634), .Y(n16106) );
  sky130_fd_sc_hd__nand2_1 U23219 ( .A(j202_soc_core_memory0_ram_dout0[411]), 
        .B(n21496), .Y(n16105) );
  sky130_fd_sc_hd__nand4_1 U23220 ( .A(n16108), .B(n16107), .C(n16106), .D(
        n16105), .Y(n16109) );
  sky130_fd_sc_hd__a2bb2oi_1 U23221 ( .B1(j202_soc_core_uart_div0[3]), .B2(
        n21513), .A1_N(n21512), .A2_N(n16111), .Y(n16183) );
  sky130_fd_sc_hd__nand2b_1 U23222 ( .A_N(n21515), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[59]), .Y(n16182) );
  sky130_fd_sc_hd__nand2_1 U23223 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[27]), .Y(n16181) );
  sky130_fd_sc_hd__nand4_1 U23224 ( .A(n16183), .B(n21768), .C(n16182), .D(
        n16181), .Y(n16179) );
  sky130_fd_sc_hd__o2bb2ai_1 U23225 ( .B1(n16206), .B2(n16842), .A1_N(n20368), 
        .A2_N(n16112), .Y(n16213) );
  sky130_fd_sc_hd__o21ai_1 U23226 ( .A1(n16114), .A2(n16113), .B1(n20368), .Y(
        n16121) );
  sky130_fd_sc_hd__o22ai_1 U23227 ( .A1(n16206), .A2(n16262), .B1(n16139), 
        .B2(n16858), .Y(n16115) );
  sky130_fd_sc_hd__a21oi_1 U23228 ( .A1(n16116), .A2(n19394), .B1(n16115), .Y(
        n16120) );
  sky130_fd_sc_hd__nand2_1 U23229 ( .A(n16117), .B(n16754), .Y(n16118) );
  sky130_fd_sc_hd__nand3_1 U23231 ( .A(n16121), .B(n16120), .C(n16119), .Y(
        n16123) );
  sky130_fd_sc_hd__o31a_1 U23232 ( .A1(n16213), .A2(n16123), .A3(n16122), .B1(
        n16871), .X(n16178) );
  sky130_fd_sc_hd__nand2_1 U23233 ( .A(n16124), .B(n20374), .Y(n16128) );
  sky130_fd_sc_hd__o21ai_1 U23234 ( .A1(n16126), .A2(n16125), .B1(n20368), .Y(
        n16127) );
  sky130_fd_sc_hd__nand2_1 U23235 ( .A(n16128), .B(n16127), .Y(n16130) );
  sky130_fd_sc_hd__nand4_1 U23237 ( .A(n16249), .B(n16150), .C(n16132), .D(
        n16131), .Y(n16134) );
  sky130_fd_sc_hd__nor2_1 U23239 ( .A(n16135), .B(n16819), .Y(n16804) );
  sky130_fd_sc_hd__nor2_1 U23240 ( .A(n16136), .B(n16804), .Y(n16137) );
  sky130_fd_sc_hd__nand4_1 U23241 ( .A(n16774), .B(n16137), .C(n16150), .D(
        n16823), .Y(n16138) );
  sky130_fd_sc_hd__nand2_1 U23242 ( .A(n16138), .B(n20385), .Y(n16145) );
  sky130_fd_sc_hd__a21oi_1 U23243 ( .A1(n16154), .A2(n16809), .B1(n16139), .Y(
        n16142) );
  sky130_fd_sc_hd__o21a_1 U23244 ( .A1(n16140), .A2(n16241), .B1(n20368), .X(
        n16141) );
  sky130_fd_sc_hd__nor2_1 U23245 ( .A(n16142), .B(n16141), .Y(n16143) );
  sky130_fd_sc_hd__nand4_1 U23246 ( .A(n16146), .B(n16145), .C(n16144), .D(
        n16143), .Y(n16174) );
  sky130_fd_sc_hd__a211o_1 U23247 ( .A1(n17242), .A2(n20303), .B1(n16803), 
        .C1(n16148), .X(n16772) );
  sky130_fd_sc_hd__nor3_1 U23248 ( .A(n16149), .B(n16247), .C(n16216), .Y(
        n16151) );
  sky130_fd_sc_hd__nand4_1 U23249 ( .A(n16151), .B(n16828), .C(n16150), .D(
        n16776), .Y(n16152) );
  sky130_fd_sc_hd__nand3_1 U23251 ( .A(n16229), .B(n16153), .C(n16242), .Y(
        n16156) );
  sky130_fd_sc_hd__o31a_1 U23252 ( .A1(n16804), .A2(n16156), .A3(n16155), .B1(
        n20374), .X(n16157) );
  sky130_fd_sc_hd__a21oi_1 U23253 ( .A1(n16159), .A2(n16158), .B1(n16157), .Y(
        n16171) );
  sky130_fd_sc_hd__nand2_1 U23254 ( .A(n16161), .B(n16160), .Y(n16777) );
  sky130_fd_sc_hd__nand3_1 U23255 ( .A(n16246), .B(n16777), .C(n16163), .Y(
        n16164) );
  sky130_fd_sc_hd__o31a_1 U23256 ( .A1(n16166), .A2(n16165), .A3(n16164), .B1(
        n20393), .X(n16169) );
  sky130_fd_sc_hd__o31a_1 U23257 ( .A1(n16808), .A2(n16167), .A3(n16832), .B1(
        n20385), .X(n16168) );
  sky130_fd_sc_hd__nor2_1 U23258 ( .A(n16169), .B(n16168), .Y(n16170) );
  sky130_fd_sc_hd__a31oi_1 U23259 ( .A1(n16172), .A2(n16171), .A3(n16170), 
        .B1(n16255), .Y(n16173) );
  sky130_fd_sc_hd__a21oi_1 U23260 ( .A1(n16174), .A2(n16801), .B1(n16173), .Y(
        n16175) );
  sky130_fd_sc_hd__nand2_1 U23261 ( .A(n16176), .B(n16175), .Y(n16177) );
  sky130_fd_sc_hd__o21a_1 U23262 ( .A1(n16178), .A2(n16177), .B1(n21629), .X(
        n16186) );
  sky130_fd_sc_hd__nor2_1 U23263 ( .A(n16179), .B(n16186), .Y(n16180) );
  sky130_fd_sc_hd__nand2_1 U23264 ( .A(j202_soc_core_memory0_ram_dout0[507]), 
        .B(n21650), .Y(n16189) );
  sky130_fd_sc_hd__nand3_1 U23265 ( .A(n16182), .B(n21653), .C(n16181), .Y(
        n16185) );
  sky130_fd_sc_hd__nor2_1 U23266 ( .A(n16185), .B(n16184), .Y(n16188) );
  sky130_fd_sc_hd__nand3_1 U23267 ( .A(n16189), .B(n16188), .C(n16187), .Y(
        n20719) );
  sky130_fd_sc_hd__ha_1 U23269 ( .A(n16190), .B(j202_soc_core_j22_cpu_pc[27]), 
        .COUT(n17046), .SUM(n16191) );
  sky130_fd_sc_hd__o22ai_1 U23270 ( .A1(n27064), .A2(n13365), .B1(n27804), 
        .B2(n11186), .Y(n17061) );
  sky130_fd_sc_hd__nor2_1 U23271 ( .A(n16544), .B(n17030), .Y(n16193) );
  sky130_fd_sc_hd__o21ai_1 U23272 ( .A1(n16544), .A2(n17036), .B1(n16551), .Y(
        n16192) );
  sky130_fd_sc_hd__nand2_1 U23273 ( .A(n17033), .B(n17031), .Y(n16195) );
  sky130_fd_sc_hd__o2bb2ai_1 U23275 ( .B1(n22705), .B2(n27064), .A1_N(n28463), 
        .A2_N(n21924), .Y(n16197) );
  sky130_fd_sc_hd__inv_1 U23276 ( .A(n16199), .Y(n16569) );
  sky130_fd_sc_hd__nand2_1 U23277 ( .A(j202_soc_core_memory0_ram_dout0[249]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[7]), .Y(n16200) );
  sky130_fd_sc_hd__nand2_1 U23278 ( .A(j202_soc_core_memory0_ram_dout0[153]), 
        .B(n20456), .Y(n16203) );
  sky130_fd_sc_hd__nand2_1 U23279 ( .A(j202_soc_core_memory0_ram_dout0[121]), 
        .B(n20460), .Y(n16202) );
  sky130_fd_sc_hd__nand2_1 U23280 ( .A(j202_soc_core_memory0_ram_dout0[185]), 
        .B(n20459), .Y(n16201) );
  sky130_fd_sc_hd__nand2_1 U23281 ( .A(n16206), .B(n16207), .Y(n16815) );
  sky130_fd_sc_hd__nand2_1 U23282 ( .A(n21074), .B(n20485), .Y(n20515) );
  sky130_fd_sc_hd__nand2b_1 U23283 ( .A_N(n20515), .B(n16205), .Y(n16270) );
  sky130_fd_sc_hd__o22ai_1 U23284 ( .A1(n16207), .A2(n16857), .B1(n16206), 
        .B2(n16270), .Y(n16208) );
  sky130_fd_sc_hd__a21oi_1 U23285 ( .A1(n16209), .A2(n16815), .B1(n16208), .Y(
        n16210) );
  sky130_fd_sc_hd__o211ai_1 U23286 ( .A1(n16211), .A2(n17102), .B1(n16210), 
        .C1(n16870), .Y(n16212) );
  sky130_fd_sc_hd__o21ai_1 U23287 ( .A1(n16213), .A2(n16212), .B1(n16871), .Y(
        n16287) );
  sky130_fd_sc_hd__nand3_1 U23288 ( .A(n16215), .B(n16751), .C(n16214), .Y(
        n16225) );
  sky130_fd_sc_hd__nor3_1 U23289 ( .A(n16217), .B(n16216), .C(n16225), .Y(
        n16218) );
  sky130_fd_sc_hd__nand2_1 U23290 ( .A(n16774), .B(n16218), .Y(n16219) );
  sky130_fd_sc_hd__nand2_1 U23291 ( .A(n16219), .B(n20385), .Y(n16236) );
  sky130_fd_sc_hd__o21ai_1 U23292 ( .A1(n16790), .A2(n16220), .B1(n20374), .Y(
        n16235) );
  sky130_fd_sc_hd__nand2_1 U23293 ( .A(n17101), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n16222) );
  sky130_fd_sc_hd__nand3_1 U23294 ( .A(n16222), .B(n16789), .C(n16221), .Y(
        n16224) );
  sky130_fd_sc_hd__o21ai_1 U23295 ( .A1(n16224), .A2(n16223), .B1(n20393), .Y(
        n16234) );
  sky130_fd_sc_hd__nand2_1 U23296 ( .A(n16226), .B(n19130), .Y(n16805) );
  sky130_fd_sc_hd__nand3_1 U23297 ( .A(n16805), .B(n16785), .C(n16778), .Y(
        n16830) );
  sky130_fd_sc_hd__nor2_1 U23298 ( .A(n16830), .B(n16228), .Y(n16230) );
  sky130_fd_sc_hd__nand4_1 U23299 ( .A(n16231), .B(n16230), .C(n16229), .D(
        n16818), .Y(n16232) );
  sky130_fd_sc_hd__nand2_1 U23300 ( .A(n16232), .B(n20368), .Y(n16233) );
  sky130_fd_sc_hd__nand4_1 U23301 ( .A(n16236), .B(n16235), .C(n16234), .D(
        n16233), .Y(n16237) );
  sky130_fd_sc_hd__nand2_1 U23302 ( .A(n16237), .B(n16801), .Y(n16286) );
  sky130_fd_sc_hd__o31a_1 U23303 ( .A1(n16240), .A2(n16239), .A3(n16238), .B1(
        n20374), .X(n16257) );
  sky130_fd_sc_hd__nor2_1 U23304 ( .A(n16831), .B(n16241), .Y(n16254) );
  sky130_fd_sc_hd__nor2b_1 U23305 ( .B_N(n16242), .A(n16780), .Y(n16244) );
  sky130_fd_sc_hd__nand4_1 U23306 ( .A(n16249), .B(n16244), .C(n16792), .D(
        n16243), .Y(n16245) );
  sky130_fd_sc_hd__nand2_1 U23307 ( .A(n16245), .B(n20368), .Y(n16253) );
  sky130_fd_sc_hd__nor3_1 U23308 ( .A(n16808), .B(n16804), .C(n16832), .Y(
        n16250) );
  sky130_fd_sc_hd__nand2_1 U23309 ( .A(n16826), .B(n16246), .Y(n16806) );
  sky130_fd_sc_hd__nor2_1 U23310 ( .A(n16247), .B(n16806), .Y(n16248) );
  sky130_fd_sc_hd__nand4_1 U23311 ( .A(n16250), .B(n16817), .C(n16249), .D(
        n16248), .Y(n16251) );
  sky130_fd_sc_hd__nand2_1 U23312 ( .A(n16251), .B(n20385), .Y(n16252) );
  sky130_fd_sc_hd__o211ai_1 U23313 ( .A1(n16254), .A2(n17102), .B1(n16253), 
        .C1(n16252), .Y(n16256) );
  sky130_fd_sc_hd__nand4_1 U23315 ( .A(n16260), .B(n16259), .C(n16258), .D(
        n16751), .Y(n16261) );
  sky130_fd_sc_hd__nand2_1 U23316 ( .A(n16261), .B(n20385), .Y(n16282) );
  sky130_fd_sc_hd__nand4_1 U23317 ( .A(n16264), .B(n16263), .C(n16754), .D(
        n16262), .Y(n16265) );
  sky130_fd_sc_hd__nand2_1 U23318 ( .A(n16265), .B(n20393), .Y(n16281) );
  sky130_fd_sc_hd__and3_1 U23320 ( .A(n16268), .B(n16267), .C(n16266), .X(
        n16269) );
  sky130_fd_sc_hd__o211ai_1 U23321 ( .A1(n16271), .A2(n16819), .B1(n16270), 
        .C1(n16269), .Y(n16753) );
  sky130_fd_sc_hd__o21ai_1 U23322 ( .A1(n16272), .A2(n16753), .B1(n20374), .Y(
        n16280) );
  sky130_fd_sc_hd__nand3_1 U23323 ( .A(n16276), .B(n16275), .C(n16274), .Y(
        n16278) );
  sky130_fd_sc_hd__nand4_1 U23325 ( .A(n16282), .B(n16281), .C(n16280), .D(
        n16279), .Y(n16283) );
  sky130_fd_sc_hd__nand2_1 U23326 ( .A(n16283), .B(n16770), .Y(n16284) );
  sky130_fd_sc_hd__nand4_1 U23327 ( .A(n16287), .B(n16286), .C(n16285), .D(
        n16284), .Y(n16288) );
  sky130_fd_sc_hd__nand2_1 U23328 ( .A(n16288), .B(n21629), .Y(n16291) );
  sky130_fd_sc_hd__a22oi_1 U23329 ( .A1(n21516), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[25]), .B1(n20540), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[57]), .Y(n16290) );
  sky130_fd_sc_hd__a22oi_1 U23330 ( .A1(n20759), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[89]), .B1(n21513), .B2(
        j202_soc_core_uart_div0[1]), .Y(n16289) );
  sky130_fd_sc_hd__nand3_1 U23331 ( .A(n16291), .B(n16290), .C(n16289), .Y(
        n16292) );
  sky130_fd_sc_hd__a21oi_1 U23332 ( .A1(j202_soc_core_memory0_ram_dout0[505]), 
        .A2(n11207), .B1(n16292), .Y(n16293) );
  sky130_fd_sc_hd__nor2_1 U23333 ( .A(n16296), .B(n17030), .Y(n16298) );
  sky130_fd_sc_hd__o21ai_1 U23334 ( .A1(n16296), .A2(n17036), .B1(n16295), .Y(
        n16297) );
  sky130_fd_sc_hd__a21oi_1 U23335 ( .A1(n17040), .A2(n16298), .B1(n16297), .Y(
        n16301) );
  sky130_fd_sc_hd__nand2_1 U23336 ( .A(n16895), .B(n16893), .Y(n16300) );
  sky130_fd_sc_hd__xor2_1 U23337 ( .A(n16301), .B(n16300), .X(n25288) );
  sky130_fd_sc_hd__nand2_1 U23338 ( .A(n25288), .B(n17225), .Y(n16307) );
  sky130_fd_sc_hd__ha_1 U23339 ( .A(n16302), .B(j202_soc_core_j22_cpu_pc[25]), 
        .COUT(n16888), .SUM(n16303) );
  sky130_fd_sc_hd__o22ai_1 U23340 ( .A1(n25286), .A2(n13365), .B1(n27796), 
        .B2(n11186), .Y(n16304) );
  sky130_fd_sc_hd__a21oi_1 U23341 ( .A1(n22701), .A2(n28475), .B1(n16304), .Y(
        n16306) );
  sky130_fd_sc_hd__nor2_1 U23342 ( .A(n16587), .B(n16679), .Y(n16964) );
  sky130_fd_sc_hd__nand2_1 U23343 ( .A(n16964), .B(n16308), .Y(n16312) );
  sky130_fd_sc_hd__nor2_1 U23344 ( .A(n16310), .B(n16309), .Y(n16941) );
  sky130_fd_sc_hd__nand2_1 U23345 ( .A(n16941), .B(n16311), .Y(n16675) );
  sky130_fd_sc_hd__o21ai_1 U23346 ( .A1(n16312), .A2(n16675), .B1(n17099), .Y(
        n16331) );
  sky130_fd_sc_hd__and4_1 U23347 ( .A(n16578), .B(n16632), .C(n16346), .D(
        n17288), .X(n16313) );
  sky130_fd_sc_hd__nand3_1 U23348 ( .A(n16314), .B(n16313), .C(n16655), .Y(
        n16967) );
  sky130_fd_sc_hd__nand4_1 U23349 ( .A(n16959), .B(n16672), .C(n16576), .D(
        n16334), .Y(n16316) );
  sky130_fd_sc_hd__nand2_1 U23350 ( .A(n17003), .B(n16617), .Y(n16315) );
  sky130_fd_sc_hd__nor2_1 U23351 ( .A(n16316), .B(n16315), .Y(n16317) );
  sky130_fd_sc_hd__nand3_1 U23352 ( .A(n16318), .B(n16317), .C(n16663), .Y(
        n16319) );
  sky130_fd_sc_hd__nand2_1 U23353 ( .A(n16319), .B(n16992), .Y(n16330) );
  sky130_fd_sc_hd__nand4_1 U23354 ( .A(n17003), .B(n16578), .C(n16577), .D(
        n16632), .Y(n16320) );
  sky130_fd_sc_hd__nand2_1 U23356 ( .A(n16321), .B(n16610), .Y(n16322) );
  sky130_fd_sc_hd__nor2_1 U23357 ( .A(n16322), .B(n16660), .Y(n16592) );
  sky130_fd_sc_hd__nand2_1 U23358 ( .A(n16989), .B(n16960), .Y(n16323) );
  sky130_fd_sc_hd__nor2_1 U23359 ( .A(n16323), .B(n16945), .Y(n16325) );
  sky130_fd_sc_hd__nor2_1 U23360 ( .A(n16976), .B(n16943), .Y(n16324) );
  sky130_fd_sc_hd__nand4_1 U23361 ( .A(n16592), .B(n16326), .C(n16325), .D(
        n16324), .Y(n16327) );
  sky130_fd_sc_hd__nand2_1 U23362 ( .A(n16327), .B(n16994), .Y(n16328) );
  sky130_fd_sc_hd__nand4_1 U23363 ( .A(n16331), .B(n16330), .C(n16329), .D(
        n16328), .Y(n16332) );
  sky130_fd_sc_hd__nand2_1 U23364 ( .A(n21629), .B(n20505), .Y(n16667) );
  sky130_fd_sc_hd__nand2_1 U23365 ( .A(n16332), .B(n20643), .Y(n16395) );
  sky130_fd_sc_hd__a2bb2oi_1 U23366 ( .B1(j202_soc_core_uart_div0[7]), .B2(
        n21513), .A1_N(n21512), .A2_N(n16333), .Y(n16389) );
  sky130_fd_sc_hd__nand2b_1 U23367 ( .A_N(n21515), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[63]), .Y(n16388) );
  sky130_fd_sc_hd__nand2_1 U23368 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[31]), .Y(n16387) );
  sky130_fd_sc_hd__nand4_1 U23369 ( .A(n16389), .B(n21768), .C(n16388), .D(
        n16387), .Y(n16344) );
  sky130_fd_sc_hd__nor2_1 U23370 ( .A(n16680), .B(n16335), .Y(n16961) );
  sky130_fd_sc_hd__nand4b_1 U23371 ( .A_N(n16336), .B(n16663), .C(n16961), .D(
        n20656), .Y(n16337) );
  sky130_fd_sc_hd__nand2_1 U23372 ( .A(n16337), .B(n17099), .Y(n16343) );
  sky130_fd_sc_hd__nand2_1 U23373 ( .A(n16338), .B(n16980), .Y(n16339) );
  sky130_fd_sc_hd__o22ai_1 U23374 ( .A1(n16356), .A2(n16339), .B1(n17001), 
        .B2(n16678), .Y(n16340) );
  sky130_fd_sc_hd__a21oi_1 U23375 ( .A1(n16992), .A2(n16341), .B1(n16340), .Y(
        n16342) );
  sky130_fd_sc_hd__nand2_1 U23376 ( .A(n21629), .B(n20508), .Y(n17146) );
  sky130_fd_sc_hd__a21oi_1 U23377 ( .A1(n16343), .A2(n16342), .B1(n17146), .Y(
        n16390) );
  sky130_fd_sc_hd__nor2_1 U23378 ( .A(n16344), .B(n16390), .Y(n16383) );
  sky130_fd_sc_hd__nor2_1 U23379 ( .A(n21359), .B(n16356), .Y(n21083) );
  sky130_fd_sc_hd__nor2_1 U23380 ( .A(n16345), .B(n21083), .Y(n16940) );
  sky130_fd_sc_hd__nand4_1 U23381 ( .A(n16623), .B(n16940), .C(n16347), .D(
        n16346), .Y(n16348) );
  sky130_fd_sc_hd__nand2_1 U23382 ( .A(n16348), .B(n17099), .Y(n16365) );
  sky130_fd_sc_hd__nand4_1 U23383 ( .A(n16618), .B(n16349), .C(n19203), .D(
        n16677), .Y(n16351) );
  sky130_fd_sc_hd__nand3_1 U23384 ( .A(n16350), .B(n16977), .C(n16632), .Y(
        n16650) );
  sky130_fd_sc_hd__nor3_1 U23385 ( .A(n16351), .B(n16650), .C(n16575), .Y(
        n16352) );
  sky130_fd_sc_hd__nand2_1 U23386 ( .A(n16623), .B(n16352), .Y(n16353) );
  sky130_fd_sc_hd__nand2_1 U23387 ( .A(n16353), .B(n16994), .Y(n16364) );
  sky130_fd_sc_hd__nand3_1 U23388 ( .A(n16988), .B(n16977), .C(n16367), .Y(
        n16598) );
  sky130_fd_sc_hd__nand4b_1 U23389 ( .A_N(n16598), .B(n16990), .C(n16959), .D(
        n16686), .Y(n16355) );
  sky130_fd_sc_hd__nand4_1 U23390 ( .A(n16605), .B(n16655), .C(n16648), .D(
        n16663), .Y(n16354) );
  sky130_fd_sc_hd__o21ai_1 U23391 ( .A1(n16355), .A2(n16354), .B1(n16980), .Y(
        n16363) );
  sky130_fd_sc_hd__nor2_1 U23392 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .B(n16356), .Y(n16670) );
  sky130_fd_sc_hd__nor2_1 U23393 ( .A(n16670), .B(n16357), .Y(n17006) );
  sky130_fd_sc_hd__nand3_1 U23394 ( .A(n16689), .B(n16678), .C(n16977), .Y(
        n16358) );
  sky130_fd_sc_hd__nor2_1 U23395 ( .A(n16358), .B(n16943), .Y(n16360) );
  sky130_fd_sc_hd__nand3_1 U23396 ( .A(n16989), .B(n16694), .C(n16672), .Y(
        n16630) );
  sky130_fd_sc_hd__nor2_1 U23397 ( .A(n16630), .B(n16575), .Y(n16359) );
  sky130_fd_sc_hd__nand3_1 U23398 ( .A(n17006), .B(n16360), .C(n16359), .Y(
        n16361) );
  sky130_fd_sc_hd__nand2_1 U23399 ( .A(n16361), .B(n16992), .Y(n16362) );
  sky130_fd_sc_hd__nand4_1 U23400 ( .A(n16365), .B(n16364), .C(n16363), .D(
        n16362), .Y(n16366) );
  sky130_fd_sc_hd__nand2_1 U23401 ( .A(n16366), .B(n20784), .Y(n16393) );
  sky130_fd_sc_hd__nand4_1 U23402 ( .A(n16368), .B(n16989), .C(n17002), .D(
        n16367), .Y(n16369) );
  sky130_fd_sc_hd__nand2_1 U23403 ( .A(n16369), .B(n16992), .Y(n16381) );
  sky130_fd_sc_hd__nand2_1 U23404 ( .A(n16577), .B(n16573), .Y(n16602) );
  sky130_fd_sc_hd__nand4b_1 U23405 ( .A_N(n16602), .B(n16977), .C(n16959), .D(
        n16619), .Y(n16370) );
  sky130_fd_sc_hd__o21ai_1 U23406 ( .A1(n16370), .A2(n16976), .B1(n16994), .Y(
        n16380) );
  sky130_fd_sc_hd__nand2_1 U23407 ( .A(n17241), .B(n20374), .Y(n16371) );
  sky130_fd_sc_hd__nand4_1 U23408 ( .A(n16618), .B(n16372), .C(n16632), .D(
        n16371), .Y(n16373) );
  sky130_fd_sc_hd__and3_1 U23410 ( .A(n16672), .B(n16374), .C(n16960), .X(
        n16978) );
  sky130_fd_sc_hd__nor2_1 U23411 ( .A(n16376), .B(n16375), .Y(n16377) );
  sky130_fd_sc_hd__nand4_1 U23412 ( .A(n16978), .B(n16377), .C(n16648), .D(
        n16689), .Y(n16586) );
  sky130_fd_sc_hd__nand2_1 U23413 ( .A(n16586), .B(n17099), .Y(n16378) );
  sky130_fd_sc_hd__nand4_1 U23414 ( .A(n16381), .B(n16380), .C(n16379), .D(
        n16378), .Y(n16382) );
  sky130_fd_sc_hd__nand2_1 U23415 ( .A(n16382), .B(n20757), .Y(n16392) );
  sky130_fd_sc_hd__nand4_1 U23416 ( .A(n16395), .B(n16383), .C(n16393), .D(
        n16392), .Y(n16384) );
  sky130_fd_sc_hd__a21oi_1 U23417 ( .A1(j202_soc_core_memory0_ram_dout0[95]), 
        .A2(n21642), .B1(n16384), .Y(n16386) );
  sky130_fd_sc_hd__nand2_1 U23418 ( .A(j202_soc_core_memory0_ram_dout0[159]), 
        .B(n21489), .Y(n16385) );
  sky130_fd_sc_hd__nand2_1 U23419 ( .A(j202_soc_core_memory0_ram_dout0[511]), 
        .B(n21650), .Y(n16397) );
  sky130_fd_sc_hd__nand4_1 U23420 ( .A(n16389), .B(n21653), .C(n16388), .D(
        n16387), .Y(n16391) );
  sky130_fd_sc_hd__nor2_1 U23421 ( .A(n16391), .B(n16390), .Y(n16394) );
  sky130_fd_sc_hd__and3_1 U23422 ( .A(n16394), .B(n16393), .C(n16392), .X(
        n16396) );
  sky130_fd_sc_hd__nand3_1 U23423 ( .A(n16397), .B(n16396), .C(n16395), .Y(
        n19851) );
  sky130_fd_sc_hd__nand2_1 U23424 ( .A(n14828), .B(
        j202_soc_core_j22_cpu_rf_gpr[350]), .Y(n16403) );
  sky130_fd_sc_hd__nand2_1 U23425 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_rf_gpr[223]), .Y(n16402) );
  sky130_fd_sc_hd__nand2_1 U23426 ( .A(n16398), .B(
        j202_soc_core_j22_cpu_rf_gpr[127]), .Y(n16401) );
  sky130_fd_sc_hd__nand2_1 U23427 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[287]), .Y(n16400) );
  sky130_fd_sc_hd__nand4_1 U23428 ( .A(n16403), .B(n16402), .C(n16401), .D(
        n16400), .Y(n16409) );
  sky130_fd_sc_hd__nand2_1 U23429 ( .A(n16425), .B(
        j202_soc_core_j22_cpu_rf_gpr[159]), .Y(n16407) );
  sky130_fd_sc_hd__nand2_1 U23430 ( .A(n16043), .B(
        j202_soc_core_j22_cpu_rf_gpr[255]), .Y(n16406) );
  sky130_fd_sc_hd__nand2_1 U23431 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[95]), .Y(n16405) );
  sky130_fd_sc_hd__nand2_1 U23432 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_rf_gpr[63]), .Y(n16404) );
  sky130_fd_sc_hd__nand4_1 U23433 ( .A(n16407), .B(n16406), .C(n16405), .D(
        n16404), .Y(n16408) );
  sky130_fd_sc_hd__nor2_1 U23434 ( .A(n16409), .B(n16408), .Y(n16423) );
  sky130_fd_sc_hd__nand2_1 U23435 ( .A(n11194), .B(
        j202_soc_core_j22_cpu_rf_gpr[318]), .Y(n16414) );
  sky130_fd_sc_hd__nand2_1 U23436 ( .A(n16410), .B(
        j202_soc_core_j22_cpu_rf_gpr[191]), .Y(n16413) );
  sky130_fd_sc_hd__nand2_1 U23437 ( .A(n15937), .B(
        j202_soc_core_j22_cpu_rf_gpr[414]), .Y(n16412) );
  sky130_fd_sc_hd__nand2_1 U23438 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[446]), .Y(n16411) );
  sky130_fd_sc_hd__and4_1 U23439 ( .A(n16414), .B(n16413), .C(n16412), .D(
        n16411), .X(n16422) );
  sky130_fd_sc_hd__nor2_1 U23440 ( .A(n16489), .B(n13537), .Y(n16420) );
  sky130_fd_sc_hd__a21oi_1 U23441 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[31]), .B1(n14743), .Y(n16418) );
  sky130_fd_sc_hd__nand2_1 U23442 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[510]), .Y(n16417) );
  sky130_fd_sc_hd__nand2_1 U23443 ( .A(n11124), .B(
        j202_soc_core_j22_cpu_rf_gpr[382]), .Y(n16416) );
  sky130_fd_sc_hd__nand2_1 U23444 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[478]), .Y(n16415) );
  sky130_fd_sc_hd__nand4_1 U23445 ( .A(n16418), .B(n16417), .C(n16416), .D(
        n16415), .Y(n16419) );
  sky130_fd_sc_hd__nor2_1 U23446 ( .A(n16420), .B(n16419), .Y(n16421) );
  sky130_fd_sc_hd__nand3_1 U23447 ( .A(n16423), .B(n16422), .C(n16421), .Y(
        n26416) );
  sky130_fd_sc_hd__nand2_1 U23448 ( .A(n26416), .B(n16424), .Y(n16459) );
  sky130_fd_sc_hd__nand2_1 U23449 ( .A(n16425), .B(
        j202_soc_core_j22_cpu_rf_gpr[158]), .Y(n16431) );
  sky130_fd_sc_hd__nand2_1 U23450 ( .A(n16426), .B(
        j202_soc_core_j22_cpu_rf_gpr[254]), .Y(n16430) );
  sky130_fd_sc_hd__nand2_1 U23451 ( .A(n11195), .B(
        j202_soc_core_j22_cpu_rf_gpr[413]), .Y(n16429) );
  sky130_fd_sc_hd__nand2_1 U23452 ( .A(n16427), .B(
        j202_soc_core_j22_cpu_rf_gpr[94]), .Y(n16428) );
  sky130_fd_sc_hd__nand4_1 U23453 ( .A(n16431), .B(n16430), .C(n16429), .D(
        n16428), .Y(n16439) );
  sky130_fd_sc_hd__nand2_1 U23454 ( .A(n16432), .B(
        j202_soc_core_j22_cpu_rf_gpr[349]), .Y(n16437) );
  sky130_fd_sc_hd__nand2_1 U23455 ( .A(n16433), .B(
        j202_soc_core_j22_cpu_rf_gpr[222]), .Y(n16436) );
  sky130_fd_sc_hd__nand2_1 U23456 ( .A(n16399), .B(
        j202_soc_core_j22_cpu_rf_gpr[286]), .Y(n16435) );
  sky130_fd_sc_hd__nand2_1 U23457 ( .A(n15783), .B(
        j202_soc_core_j22_cpu_rf_gpr[126]), .Y(n16434) );
  sky130_fd_sc_hd__nand4_1 U23458 ( .A(n16437), .B(n16436), .C(n16435), .D(
        n16434), .Y(n16438) );
  sky130_fd_sc_hd__nor2_1 U23459 ( .A(n16439), .B(n16438), .Y(n16456) );
  sky130_fd_sc_hd__nand2_1 U23460 ( .A(n11125), .B(
        j202_soc_core_j22_cpu_rf_gpr[317]), .Y(n16443) );
  sky130_fd_sc_hd__nand2_1 U23461 ( .A(n16410), .B(
        j202_soc_core_j22_cpu_rf_gpr[190]), .Y(n16442) );
  sky130_fd_sc_hd__nand2_1 U23462 ( .A(n11196), .B(
        j202_soc_core_j22_cpu_rf_gpr[381]), .Y(n16441) );
  sky130_fd_sc_hd__nand2_1 U23463 ( .A(n14821), .B(
        j202_soc_core_j22_cpu_rf_gpr[477]), .Y(n16440) );
  sky130_fd_sc_hd__nor2_1 U23464 ( .A(n16445), .B(n16444), .Y(n16454) );
  sky130_fd_sc_hd__a21oi_1 U23465 ( .A1(n13053), .A2(
        j202_soc_core_j22_cpu_rf_tmp[30]), .B1(n14743), .Y(n16452) );
  sky130_fd_sc_hd__nand2_1 U23466 ( .A(n16446), .B(
        j202_soc_core_j22_cpu_rf_gpr[62]), .Y(n16451) );
  sky130_fd_sc_hd__nand2_1 U23467 ( .A(n16447), .B(
        j202_soc_core_j22_cpu_rf_gpr[509]), .Y(n16450) );
  sky130_fd_sc_hd__nand2_1 U23468 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[445]), .Y(n16449) );
  sky130_fd_sc_hd__nand4_1 U23469 ( .A(n16452), .B(n16451), .C(n16450), .D(
        n16449), .Y(n16453) );
  sky130_fd_sc_hd__nor2_1 U23470 ( .A(n16454), .B(n16453), .Y(n16455) );
  sky130_fd_sc_hd__nand3_1 U23471 ( .A(n16456), .B(n13063), .C(n16455), .Y(
        n26330) );
  sky130_fd_sc_hd__nand2_1 U23472 ( .A(n26330), .B(n16457), .Y(n16458) );
  sky130_fd_sc_hd__nand2_1 U23473 ( .A(n16459), .B(n16458), .Y(n25803) );
  sky130_fd_sc_hd__nand2_1 U23474 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[223]), .Y(n16465) );
  sky130_fd_sc_hd__nand2_1 U23475 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[478]), .Y(n16464) );
  sky130_fd_sc_hd__nand2_1 U23476 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[510]), .Y(n16463) );
  sky130_fd_sc_hd__nand2_1 U23477 ( .A(n16461), .B(
        j202_soc_core_j22_cpu_rf_gpr[255]), .Y(n16462) );
  sky130_fd_sc_hd__nand4_1 U23478 ( .A(n16465), .B(n16464), .C(n16463), .D(
        n16462), .Y(n16472) );
  sky130_fd_sc_hd__nand2_1 U23479 ( .A(n23500), .B(
        j202_soc_core_j22_cpu_rf_gpr[31]), .Y(n16470) );
  sky130_fd_sc_hd__nand2_1 U23480 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[95]), .Y(n16469) );
  sky130_fd_sc_hd__nand2_1 U23481 ( .A(n16466), .B(
        j202_soc_core_j22_cpu_rf_gpr[414]), .Y(n16468) );
  sky130_fd_sc_hd__nand2_1 U23482 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[159]), .Y(n16467) );
  sky130_fd_sc_hd__nand4_1 U23483 ( .A(n16470), .B(n16469), .C(n16468), .D(
        n16467), .Y(n16471) );
  sky130_fd_sc_hd__nor2_1 U23484 ( .A(n16472), .B(n16471), .Y(n16483) );
  sky130_fd_sc_hd__nand2_1 U23485 ( .A(n14275), .B(
        j202_soc_core_j22_cpu_rf_gpr[287]), .Y(n16476) );
  sky130_fd_sc_hd__nand2_1 U23486 ( .A(n13566), .B(
        j202_soc_core_j22_cpu_rf_gpr[63]), .Y(n16475) );
  sky130_fd_sc_hd__nand2_1 U23487 ( .A(n23776), .B(
        j202_soc_core_j22_cpu_rf_gpr[382]), .Y(n16474) );
  sky130_fd_sc_hd__nand2_1 U23488 ( .A(n16064), .B(
        j202_soc_core_j22_cpu_rf_gpr[350]), .Y(n16473) );
  sky130_fd_sc_hd__and4_1 U23489 ( .A(n16476), .B(n16475), .C(n16474), .D(
        n16473), .X(n16482) );
  sky130_fd_sc_hd__nand2_1 U23490 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[318]), .Y(n16480) );
  sky130_fd_sc_hd__nand2_1 U23491 ( .A(n23823), .B(
        j202_soc_core_j22_cpu_rf_gpr[446]), .Y(n16479) );
  sky130_fd_sc_hd__nand2_1 U23492 ( .A(n11199), .B(
        j202_soc_core_j22_cpu_rf_gpr[191]), .Y(n16478) );
  sky130_fd_sc_hd__nand2_1 U23493 ( .A(n15992), .B(
        j202_soc_core_j22_cpu_rf_gpr[127]), .Y(n16477) );
  sky130_fd_sc_hd__and4_1 U23494 ( .A(n16480), .B(n16479), .C(n16478), .D(
        n16477), .X(n16481) );
  sky130_fd_sc_hd__nand3_1 U23495 ( .A(n16483), .B(n16482), .C(n16481), .Y(
        n22466) );
  sky130_fd_sc_hd__o22a_1 U23496 ( .A1(n16486), .A2(n16077), .B1(n16485), .B2(
        n14342), .X(n16497) );
  sky130_fd_sc_hd__o22a_1 U23497 ( .A1(n16489), .A2(n16488), .B1(n16487), .B2(
        n22463), .X(n16496) );
  sky130_fd_sc_hd__o22a_1 U23498 ( .A1(n16492), .A2(n16491), .B1(n16490), .B2(
        n22462), .X(n16495) );
  sky130_fd_sc_hd__a21oi_1 U23499 ( .A1(n11201), .A2(
        j202_soc_core_j22_cpu_rf_gpr[510]), .B1(n16493), .Y(n16494) );
  sky130_fd_sc_hd__nand4_1 U23500 ( .A(n16497), .B(n16496), .C(n16495), .D(
        n16494), .Y(n16498) );
  sky130_fd_sc_hd__a21oi_1 U23501 ( .A1(n22466), .A2(n16523), .B1(n16498), .Y(
        n26408) );
  sky130_fd_sc_hd__nand2_1 U23502 ( .A(n26408), .B(n16543), .Y(n16499) );
  sky130_fd_sc_hd__o21a_1 U23503 ( .A1(n26408), .A2(n16541), .B1(n16499), .X(
        n25804) );
  sky130_fd_sc_hd__xnor2_1 U23504 ( .A(n25803), .B(n25804), .Y(n26206) );
  sky130_fd_sc_hd__o22ai_1 U23505 ( .A1(n16501), .A2(n26435), .B1(n26296), 
        .B2(n16500), .Y(n16546) );
  sky130_fd_sc_hd__nand2_1 U23506 ( .A(n23792), .B(
        j202_soc_core_j22_cpu_rf_gpr[222]), .Y(n16505) );
  sky130_fd_sc_hd__nand2_1 U23507 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[477]), .Y(n16504) );
  sky130_fd_sc_hd__nand2_1 U23508 ( .A(n13820), .B(
        j202_soc_core_j22_cpu_rf_gpr[509]), .Y(n16503) );
  sky130_fd_sc_hd__nand2_1 U23509 ( .A(n23754), .B(
        j202_soc_core_j22_cpu_rf_gpr[254]), .Y(n16502) );
  sky130_fd_sc_hd__nand4_1 U23510 ( .A(n16505), .B(n16504), .C(n16503), .D(
        n16502), .Y(n16513) );
  sky130_fd_sc_hd__nand2_1 U23511 ( .A(n16506), .B(
        j202_soc_core_j22_cpu_rf_gpr[30]), .Y(n16511) );
  sky130_fd_sc_hd__nand2_1 U23512 ( .A(n16507), .B(
        j202_soc_core_j22_cpu_rf_gpr[94]), .Y(n16510) );
  sky130_fd_sc_hd__nand2_1 U23513 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_rf_gpr[413]), .Y(n16509) );
  sky130_fd_sc_hd__nand2_1 U23514 ( .A(n15951), .B(
        j202_soc_core_j22_cpu_rf_gpr[158]), .Y(n16508) );
  sky130_fd_sc_hd__nand4_1 U23515 ( .A(n16511), .B(n16510), .C(n16509), .D(
        n16508), .Y(n16512) );
  sky130_fd_sc_hd__nor2_1 U23516 ( .A(n16513), .B(n16512), .Y(n16522) );
  sky130_fd_sc_hd__a22oi_1 U23517 ( .A1(n23776), .A2(
        j202_soc_core_j22_cpu_rf_gpr[381]), .B1(n14275), .B2(
        j202_soc_core_j22_cpu_rf_gpr[286]), .Y(n16521) );
  sky130_fd_sc_hd__a22oi_1 U23518 ( .A1(n13566), .A2(
        j202_soc_core_j22_cpu_rf_gpr[62]), .B1(n15017), .B2(
        j202_soc_core_j22_cpu_rf_gpr[349]), .Y(n16520) );
  sky130_fd_sc_hd__nand2_1 U23519 ( .A(n23781), .B(
        j202_soc_core_j22_cpu_rf_gpr[317]), .Y(n16518) );
  sky130_fd_sc_hd__nand2_1 U23520 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_gpr[445]), .Y(n16517) );
  sky130_fd_sc_hd__nand2_1 U23521 ( .A(n23802), .B(
        j202_soc_core_j22_cpu_rf_gpr[190]), .Y(n16516) );
  sky130_fd_sc_hd__nand2_1 U23522 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[126]), .Y(n16515) );
  sky130_fd_sc_hd__and4_1 U23523 ( .A(n16518), .B(n16517), .C(n16516), .D(
        n16515), .X(n16519) );
  sky130_fd_sc_hd__nand4_1 U23524 ( .A(n16522), .B(n16521), .C(n16520), .D(
        n16519), .Y(n22585) );
  sky130_fd_sc_hd__nand2_1 U23525 ( .A(n22585), .B(n16523), .Y(n16540) );
  sky130_fd_sc_hd__o22ai_1 U23527 ( .A1(n16528), .A2(n11202), .B1(n16527), 
        .B2(n14342), .Y(n16529) );
  sky130_fd_sc_hd__nor2_1 U23528 ( .A(n16530), .B(n16529), .Y(n16539) );
  sky130_fd_sc_hd__nand2_1 U23529 ( .A(n16531), .B(
        j202_soc_core_j22_cpu_rf_gpr[30]), .Y(n16538) );
  sky130_fd_sc_hd__nand2_1 U23530 ( .A(n16532), .B(
        j202_soc_core_j22_cpu_rf_pr[30]), .Y(n16537) );
  sky130_fd_sc_hd__nand2_1 U23531 ( .A(n16533), .B(
        j202_soc_core_j22_cpu_pc[30]), .Y(n16536) );
  sky130_fd_sc_hd__nand2_1 U23532 ( .A(n16534), .B(
        j202_soc_core_j22_cpu_rf_gbr[30]), .Y(n16535) );
  sky130_fd_sc_hd__nand3_1 U23533 ( .A(n16540), .B(n16539), .C(n13108), .Y(
        n28446) );
  sky130_fd_sc_hd__nand2_1 U23534 ( .A(n28446), .B(n16541), .Y(n16542) );
  sky130_fd_sc_hd__nor2_1 U23536 ( .A(n16546), .B(n16547), .Y(n16730) );
  sky130_fd_sc_hd__nor2_1 U23537 ( .A(n16730), .B(n16723), .Y(n16549) );
  sky130_fd_sc_hd__nand2_1 U23538 ( .A(n16549), .B(n16718), .Y(n16552) );
  sky130_fd_sc_hd__nor2_1 U23539 ( .A(n16552), .B(n16544), .Y(n16554) );
  sky130_fd_sc_hd__nand2_1 U23540 ( .A(n16545), .B(n16554), .Y(n16558) );
  sky130_fd_sc_hd__nand2_1 U23541 ( .A(n16547), .B(n16546), .Y(n16731) );
  sky130_fd_sc_hd__o21ai_1 U23542 ( .A1(n16721), .A2(n16730), .B1(n16731), .Y(
        n16548) );
  sky130_fd_sc_hd__a21oi_1 U23543 ( .A1(n16549), .A2(n16720), .B1(n16548), .Y(
        n16550) );
  sky130_fd_sc_hd__a21oi_1 U23545 ( .A1(n16555), .A2(n16554), .B1(n16553), .Y(
        n16556) );
  sky130_fd_sc_hd__nand2_1 U23546 ( .A(n21925), .B(n26416), .Y(n16562) );
  sky130_fd_sc_hd__ha_1 U23547 ( .A(n16559), .B(j202_soc_core_j22_cpu_pc[29]), 
        .COUT(n16735), .SUM(n25465) );
  sky130_fd_sc_hd__xor2_1 U23548 ( .A(j202_soc_core_j22_cpu_pc[31]), .B(n16560), .X(n27587) );
  sky130_fd_sc_hd__nand2_1 U23549 ( .A(n27587), .B(n21322), .Y(n16561) );
  sky130_fd_sc_hd__o211ai_1 U23550 ( .A1(n26408), .A2(n22745), .B1(n16562), 
        .C1(n16561), .Y(n16563) );
  sky130_fd_sc_hd__nand2_1 U23551 ( .A(n27587), .B(n17048), .Y(n16565) );
  sky130_fd_sc_hd__nand2_1 U23552 ( .A(n22701), .B(n28431), .Y(n16564) );
  sky130_fd_sc_hd__nand2_1 U23553 ( .A(n16565), .B(n16564), .Y(n17059) );
  sky130_fd_sc_hd__inv_1 U23554 ( .A(n21045), .Y(n17056) );
  sky130_fd_sc_hd__nand2_1 U23555 ( .A(n16654), .B(n16573), .Y(n16574) );
  sky130_fd_sc_hd__nor2_1 U23556 ( .A(n16574), .B(n16660), .Y(n16581) );
  sky130_fd_sc_hd__nor2_1 U23557 ( .A(n16598), .B(n16575), .Y(n16580) );
  sky130_fd_sc_hd__nand4_1 U23558 ( .A(n17003), .B(n16578), .C(n16577), .D(
        n16576), .Y(n17005) );
  sky130_fd_sc_hd__nor2_1 U23559 ( .A(n16976), .B(n17005), .Y(n16579) );
  sky130_fd_sc_hd__nand4_1 U23560 ( .A(n17006), .B(n16581), .C(n16580), .D(
        n16579), .Y(n16585) );
  sky130_fd_sc_hd__nand3_1 U23561 ( .A(n17002), .B(n16960), .C(n17288), .Y(
        n16653) );
  sky130_fd_sc_hd__nor3_1 U23562 ( .A(n16603), .B(n16653), .C(n17005), .Y(
        n16583) );
  sky130_fd_sc_hd__nand3_1 U23563 ( .A(n16583), .B(n16965), .C(n16582), .Y(
        n16584) );
  sky130_fd_sc_hd__a22o_1 U23564 ( .A1(n16992), .A2(n16585), .B1(n16584), .B2(
        n16994), .X(n16596) );
  sky130_fd_sc_hd__nor2_1 U23565 ( .A(n16587), .B(n16968), .Y(n16588) );
  sky130_fd_sc_hd__nand4_1 U23566 ( .A(n16588), .B(n16989), .C(n16694), .D(
        n16619), .Y(n16589) );
  sky130_fd_sc_hd__nor2_1 U23567 ( .A(n16589), .B(n16942), .Y(n16590) );
  sky130_fd_sc_hd__nand3_1 U23568 ( .A(n16592), .B(n16591), .C(n16590), .Y(
        n16593) );
  sky130_fd_sc_hd__o2bb2ai_1 U23569 ( .B1(n17007), .B2(n16594), .A1_N(n16980), 
        .A2_N(n16593), .Y(n16595) );
  sky130_fd_sc_hd__nor2_1 U23570 ( .A(n16596), .B(n16595), .Y(n16629) );
  sky130_fd_sc_hd__nor2_1 U23571 ( .A(n16598), .B(n16597), .Y(n16684) );
  sky130_fd_sc_hd__a21oi_1 U23572 ( .A1(n19124), .A2(n19148), .B1(n16599), .Y(
        n16600) );
  sky130_fd_sc_hd__nand3_1 U23573 ( .A(n16684), .B(n16651), .C(n16600), .Y(
        n16607) );
  sky130_fd_sc_hd__nor3_1 U23574 ( .A(n16603), .B(n16602), .C(n16601), .Y(
        n16604) );
  sky130_fd_sc_hd__nand4_1 U23575 ( .A(n16623), .B(n17006), .C(n16605), .D(
        n16604), .Y(n16606) );
  sky130_fd_sc_hd__a22oi_1 U23576 ( .A1(n16607), .A2(n16980), .B1(n16606), 
        .B2(n16992), .Y(n16627) );
  sky130_fd_sc_hd__nor2_1 U23577 ( .A(n16612), .B(n16611), .Y(n16613) );
  sky130_fd_sc_hd__nand4_1 U23578 ( .A(n16615), .B(n16614), .C(n16613), .D(
        n16618), .Y(n16616) );
  sky130_fd_sc_hd__nand2_1 U23579 ( .A(n16616), .B(n17099), .Y(n16626) );
  sky130_fd_sc_hd__nor2_1 U23580 ( .A(n16631), .B(n16620), .Y(n16621) );
  sky130_fd_sc_hd__nand4_1 U23581 ( .A(n16623), .B(n16622), .C(n16682), .D(
        n16621), .Y(n16624) );
  sky130_fd_sc_hd__nand2_1 U23582 ( .A(n16624), .B(n16994), .Y(n16625) );
  sky130_fd_sc_hd__nand3_1 U23583 ( .A(n16627), .B(n16626), .C(n16625), .Y(
        n16628) );
  sky130_fd_sc_hd__o2bb2ai_1 U23584 ( .B1(n20823), .B2(n16629), .A1_N(n16996), 
        .A2_N(n16628), .Y(n16716) );
  sky130_fd_sc_hd__nor2_1 U23585 ( .A(n16631), .B(n16630), .Y(n17004) );
  sky130_fd_sc_hd__nor2_1 U23586 ( .A(n16634), .B(n16633), .Y(n16635) );
  sky130_fd_sc_hd__nand4_1 U23587 ( .A(n17004), .B(n16636), .C(n16635), .D(
        n16987), .Y(n16647) );
  sky130_fd_sc_hd__a21oi_1 U23588 ( .A1(n16638), .A2(n21088), .B1(n16637), .Y(
        n16640) );
  sky130_fd_sc_hd__nand4b_1 U23589 ( .A_N(n16943), .B(n16640), .C(n16639), .D(
        n16686), .Y(n16969) );
  sky130_fd_sc_hd__nor2_1 U23590 ( .A(n16642), .B(n16641), .Y(n16643) );
  sky130_fd_sc_hd__nand4_1 U23591 ( .A(n16645), .B(n16644), .C(n16643), .D(
        n17003), .Y(n16646) );
  sky130_fd_sc_hd__a22oi_1 U23592 ( .A1(n16647), .A2(n16980), .B1(n16646), 
        .B2(n16994), .Y(n16669) );
  sky130_fd_sc_hd__nand3_1 U23593 ( .A(n16648), .B(n16686), .C(n16963), .Y(
        n16649) );
  sky130_fd_sc_hd__nor2_1 U23594 ( .A(n16650), .B(n16649), .Y(n16652) );
  sky130_fd_sc_hd__nand4_1 U23595 ( .A(n16652), .B(n16651), .C(n17003), .D(
        n16689), .Y(n16666) );
  sky130_fd_sc_hd__nand3_1 U23596 ( .A(n16656), .B(n16655), .C(n16654), .Y(
        n16659) );
  sky130_fd_sc_hd__nor2_1 U23597 ( .A(n16659), .B(n16658), .Y(n16664) );
  sky130_fd_sc_hd__nand4_1 U23598 ( .A(n16664), .B(n16704), .C(n16663), .D(
        n16662), .Y(n16665) );
  sky130_fd_sc_hd__a22oi_1 U23599 ( .A1(n16666), .A2(n17099), .B1(n16665), 
        .B2(n16992), .Y(n16668) );
  sky130_fd_sc_hd__a21oi_1 U23600 ( .A1(n16669), .A2(n16668), .B1(n16667), .Y(
        n16714) );
  sky130_fd_sc_hd__nand4b_1 U23601 ( .A_N(n16674), .B(n16673), .C(n16672), .D(
        n16671), .Y(n16676) );
  sky130_fd_sc_hd__nand3_1 U23603 ( .A(n16678), .B(n17002), .C(n16677), .Y(
        n16687) );
  sky130_fd_sc_hd__nor2_1 U23604 ( .A(n16680), .B(n16679), .Y(n16681) );
  sky130_fd_sc_hd__nand4_1 U23605 ( .A(n16684), .B(n16683), .C(n16682), .D(
        n16681), .Y(n16685) );
  sky130_fd_sc_hd__nand2_1 U23606 ( .A(n16685), .B(n16994), .Y(n16708) );
  sky130_fd_sc_hd__nand2_1 U23607 ( .A(n16686), .B(n20656), .Y(n16688) );
  sky130_fd_sc_hd__nor2_1 U23608 ( .A(n16688), .B(n16687), .Y(n16951) );
  sky130_fd_sc_hd__nand4_1 U23609 ( .A(n16692), .B(n16951), .C(n16691), .D(
        n16690), .Y(n16693) );
  sky130_fd_sc_hd__nand2_1 U23610 ( .A(n16693), .B(n16992), .Y(n16707) );
  sky130_fd_sc_hd__nand3_1 U23611 ( .A(n16959), .B(n16977), .C(n16694), .Y(
        n16695) );
  sky130_fd_sc_hd__nor3_1 U23612 ( .A(n16697), .B(n16696), .C(n16695), .Y(
        n16949) );
  sky130_fd_sc_hd__nor2_1 U23613 ( .A(n16700), .B(n16699), .Y(n16703) );
  sky130_fd_sc_hd__nor2_1 U23614 ( .A(n16945), .B(n16701), .Y(n16702) );
  sky130_fd_sc_hd__nand4_1 U23615 ( .A(n16949), .B(n16704), .C(n16703), .D(
        n16702), .Y(n16705) );
  sky130_fd_sc_hd__nand2_1 U23616 ( .A(n16705), .B(n16980), .Y(n16706) );
  sky130_fd_sc_hd__nand4_1 U23617 ( .A(n16709), .B(n16708), .C(n16707), .D(
        n16706), .Y(n16710) );
  sky130_fd_sc_hd__nand2_1 U23618 ( .A(n16710), .B(n20784), .Y(n16713) );
  sky130_fd_sc_hd__a22oi_1 U23619 ( .A1(n21516), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[30]), .B1(n20540), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[62]), .Y(n16712) );
  sky130_fd_sc_hd__a22oi_1 U23620 ( .A1(n20759), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[94]), .B1(n21513), .B2(
        j202_soc_core_uart_div0[6]), .Y(n16711) );
  sky130_fd_sc_hd__nand4b_1 U23621 ( .A_N(n16714), .B(n16713), .C(n16712), .D(
        n16711), .Y(n16715) );
  sky130_fd_sc_hd__a21o_1 U23622 ( .A1(n16716), .A2(n21629), .B1(n16715), .X(
        n16717) );
  sky130_fd_sc_hd__a21oi_1 U23623 ( .A1(j202_soc_core_memory0_ram_dout0[510]), 
        .A2(n11207), .B1(n16717), .Y(n20091) );
  sky130_fd_sc_hd__nand2_1 U23624 ( .A(n26168), .B(n22739), .Y(n17067) );
  sky130_fd_sc_hd__nor2_1 U23625 ( .A(n16723), .B(n16719), .Y(n16725) );
  sky130_fd_sc_hd__nand2_1 U23626 ( .A(n16725), .B(n17029), .Y(n16727) );
  sky130_fd_sc_hd__nor2_1 U23627 ( .A(n16727), .B(n17030), .Y(n16729) );
  sky130_fd_sc_hd__o21ai_1 U23628 ( .A1(n16723), .A2(n16722), .B1(n16721), .Y(
        n16724) );
  sky130_fd_sc_hd__a21oi_1 U23629 ( .A1(n17034), .A2(n16725), .B1(n16724), .Y(
        n16726) );
  sky130_fd_sc_hd__o21ai_1 U23630 ( .A1(n16727), .A2(n17036), .B1(n16726), .Y(
        n16728) );
  sky130_fd_sc_hd__nand2_1 U23632 ( .A(n16732), .B(n16731), .Y(n16733) );
  sky130_fd_sc_hd__xor2_1 U23633 ( .A(n16734), .B(n16733), .X(n25141) );
  sky130_fd_sc_hd__ha_1 U23634 ( .A(n16735), .B(j202_soc_core_j22_cpu_pc[30]), 
        .COUT(n16560), .SUM(n25138) );
  sky130_fd_sc_hd__nand2_1 U23635 ( .A(n25138), .B(n21322), .Y(n16737) );
  sky130_fd_sc_hd__nand2_1 U23636 ( .A(n25138), .B(n17048), .Y(n16736) );
  sky130_fd_sc_hd__o211ai_1 U23637 ( .A1(n26435), .A2(n11186), .B1(n16737), 
        .C1(n16736), .Y(n17060) );
  sky130_fd_sc_hd__nand3_1 U23638 ( .A(n16742), .B(n16741), .C(n16740), .Y(
        n16744) );
  sky130_fd_sc_hd__o21ai_1 U23639 ( .A1(n16744), .A2(n16743), .B1(n20393), .Y(
        n16769) );
  sky130_fd_sc_hd__nor2_1 U23640 ( .A(n16762), .B(n16849), .Y(n16750) );
  sky130_fd_sc_hd__nand4_1 U23642 ( .A(n16751), .B(n16750), .C(n16749), .D(
        n16748), .Y(n16752) );
  sky130_fd_sc_hd__o21ai_1 U23643 ( .A1(n16753), .A2(n16752), .B1(n20374), .Y(
        n16768) );
  sky130_fd_sc_hd__nand4_1 U23644 ( .A(n16858), .B(n16756), .C(n16755), .D(
        n16754), .Y(n16760) );
  sky130_fd_sc_hd__nand2_1 U23645 ( .A(n16757), .B(n16851), .Y(n16758) );
  sky130_fd_sc_hd__nand2_1 U23646 ( .A(n16759), .B(n16758), .Y(n16843) );
  sky130_fd_sc_hd__o21ai_1 U23647 ( .A1(n16760), .A2(n16843), .B1(n20368), .Y(
        n16767) );
  sky130_fd_sc_hd__a211o_1 U23648 ( .A1(n16764), .A2(n16763), .B1(n16762), 
        .C1(n16761), .X(n16765) );
  sky130_fd_sc_hd__nand2_1 U23649 ( .A(n16765), .B(n20385), .Y(n16766) );
  sky130_fd_sc_hd__nand4_1 U23650 ( .A(n16769), .B(n16768), .C(n16767), .D(
        n16766), .Y(n16771) );
  sky130_fd_sc_hd__nand2_1 U23651 ( .A(n16771), .B(n16770), .Y(n16876) );
  sky130_fd_sc_hd__nand2_1 U23652 ( .A(n16774), .B(n16773), .Y(n16800) );
  sky130_fd_sc_hd__nand2_1 U23653 ( .A(n16776), .B(n16775), .Y(n16781) );
  sky130_fd_sc_hd__nand2_1 U23654 ( .A(n16778), .B(n16777), .Y(n16779) );
  sky130_fd_sc_hd__nor3_1 U23655 ( .A(n16781), .B(n16780), .C(n16779), .Y(
        n16798) );
  sky130_fd_sc_hd__nor2_1 U23656 ( .A(n16782), .B(n16804), .Y(n16783) );
  sky130_fd_sc_hd__nand4_1 U23657 ( .A(n16785), .B(n16823), .C(n16784), .D(
        n16783), .Y(n16787) );
  sky130_fd_sc_hd__o21ai_1 U23658 ( .A1(n16787), .A2(n16786), .B1(n20368), .Y(
        n16797) );
  sky130_fd_sc_hd__nor2_1 U23659 ( .A(n16791), .B(n16790), .Y(n16793) );
  sky130_fd_sc_hd__nand4_1 U23660 ( .A(n16794), .B(n16793), .C(n16792), .D(
        n16809), .Y(n16795) );
  sky130_fd_sc_hd__o211ai_1 U23662 ( .A1(n16798), .A2(n17102), .B1(n16797), 
        .C1(n16796), .Y(n16799) );
  sky130_fd_sc_hd__a21o_1 U23663 ( .A1(n16800), .A2(n20385), .B1(n16799), .X(
        n16802) );
  sky130_fd_sc_hd__nand2_1 U23664 ( .A(n16802), .B(n16801), .Y(n16875) );
  sky130_fd_sc_hd__nor2_1 U23665 ( .A(n16804), .B(n16803), .Y(n16812) );
  sky130_fd_sc_hd__nor2_1 U23666 ( .A(n16807), .B(n16806), .Y(n16811) );
  sky130_fd_sc_hd__nand4_1 U23667 ( .A(n16812), .B(n16811), .C(n16810), .D(
        n16809), .Y(n16813) );
  sky130_fd_sc_hd__o21ai_0 U23668 ( .A1(n16814), .A2(n16813), .B1(n20368), .Y(
        n16839) );
  sky130_fd_sc_hd__nand2_1 U23669 ( .A(n16817), .B(n16816), .Y(n16825) );
  sky130_fd_sc_hd__nand2_1 U23671 ( .A(n16821), .B(n20393), .Y(n16822) );
  sky130_fd_sc_hd__o21ai_1 U23672 ( .A1(n19394), .A2(n16823), .B1(n16822), .Y(
        n16824) );
  sky130_fd_sc_hd__a21oi_1 U23673 ( .A1(n16848), .A2(n16825), .B1(n16824), .Y(
        n16838) );
  sky130_fd_sc_hd__nand3_1 U23674 ( .A(n16828), .B(n16827), .C(n16826), .Y(
        n16829) );
  sky130_fd_sc_hd__o21ai_1 U23675 ( .A1(n16830), .A2(n16829), .B1(n20374), .Y(
        n16837) );
  sky130_fd_sc_hd__nor2_1 U23676 ( .A(n16832), .B(n16831), .Y(n16833) );
  sky130_fd_sc_hd__nand2_1 U23677 ( .A(n16834), .B(n16833), .Y(n16835) );
  sky130_fd_sc_hd__nand2_1 U23678 ( .A(n16835), .B(n20385), .Y(n16836) );
  sky130_fd_sc_hd__nand4_1 U23679 ( .A(n16839), .B(n16838), .C(n16837), .D(
        n16836), .Y(n16841) );
  sky130_fd_sc_hd__nand2_1 U23680 ( .A(n16841), .B(n16840), .Y(n16874) );
  sky130_fd_sc_hd__nand3_1 U23682 ( .A(n16846), .B(n16864), .C(n16845), .Y(
        n16847) );
  sky130_fd_sc_hd__nand2_1 U23683 ( .A(n16847), .B(n20393), .Y(n16854) );
  sky130_fd_sc_hd__nand2_1 U23684 ( .A(n16849), .B(n16848), .Y(n16853) );
  sky130_fd_sc_hd__nand3_1 U23685 ( .A(n16851), .B(n20374), .C(n16850), .Y(
        n16852) );
  sky130_fd_sc_hd__nand4_1 U23686 ( .A(n16855), .B(n16854), .C(n16853), .D(
        n16852), .Y(n16863) );
  sky130_fd_sc_hd__nand4_1 U23687 ( .A(n16859), .B(n16865), .C(n16858), .D(
        n16857), .Y(n16860) );
  sky130_fd_sc_hd__o21a_1 U23688 ( .A1(n16861), .A2(n16860), .B1(n20385), .X(
        n16862) );
  sky130_fd_sc_hd__nor2_1 U23689 ( .A(n16863), .B(n16862), .Y(n16869) );
  sky130_fd_sc_hd__nand3_1 U23690 ( .A(n16866), .B(n16865), .C(n16864), .Y(
        n16867) );
  sky130_fd_sc_hd__nand2_1 U23691 ( .A(n16867), .B(n20368), .Y(n16868) );
  sky130_fd_sc_hd__nand3_1 U23692 ( .A(n16870), .B(n16869), .C(n16868), .Y(
        n16872) );
  sky130_fd_sc_hd__nand2_1 U23693 ( .A(n16872), .B(n16871), .Y(n16873) );
  sky130_fd_sc_hd__nand4_1 U23694 ( .A(n16876), .B(n16875), .C(n16874), .D(
        n16873), .Y(n16877) );
  sky130_fd_sc_hd__nand2_1 U23695 ( .A(n16877), .B(n21629), .Y(n16880) );
  sky130_fd_sc_hd__a22oi_1 U23696 ( .A1(n21516), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[26]), .B1(n20540), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[58]), .Y(n16879) );
  sky130_fd_sc_hd__a22oi_1 U23697 ( .A1(n20759), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[90]), .B1(n21513), .B2(
        j202_soc_core_uart_div0[2]), .Y(n16878) );
  sky130_fd_sc_hd__nand3_1 U23698 ( .A(n16880), .B(n16879), .C(n16878), .Y(
        n16881) );
  sky130_fd_sc_hd__a21oi_1 U23699 ( .A1(j202_soc_core_memory0_ram_dout0[506]), 
        .A2(n11207), .B1(n16881), .Y(n16887) );
  sky130_fd_sc_hd__a22oi_1 U23700 ( .A1(j202_soc_core_memory0_ram_dout0[250]), 
        .A2(j202_soc_core_memory0_ram_dout0_sel[7]), .B1(n20455), .B2(
        j202_soc_core_memory0_ram_dout0[218]), .Y(n16885) );
  sky130_fd_sc_hd__nand2_1 U23701 ( .A(j202_soc_core_memory0_ram_dout0[90]), 
        .B(n20458), .Y(n16883) );
  sky130_fd_sc_hd__ha_1 U23702 ( .A(n16888), .B(j202_soc_core_j22_cpu_pc[26]), 
        .COUT(n16190), .SUM(n27863) );
  sky130_fd_sc_hd__o22ai_1 U23703 ( .A1(n27849), .A2(n13365), .B1(n27825), 
        .B2(n11186), .Y(n16889) );
  sky130_fd_sc_hd__a21oi_1 U23704 ( .A1(n22701), .A2(n28471), .B1(n16889), .Y(
        n16891) );
  sky130_fd_sc_hd__nand2_1 U23705 ( .A(n22702), .B(n28471), .Y(n16890) );
  sky130_fd_sc_hd__nand2_1 U23706 ( .A(n16892), .B(n16895), .Y(n16898) );
  sky130_fd_sc_hd__nor2_1 U23707 ( .A(n16898), .B(n17030), .Y(n16900) );
  sky130_fd_sc_hd__a21oi_1 U23708 ( .A1(n16896), .A2(n16895), .B1(n16894), .Y(
        n16897) );
  sky130_fd_sc_hd__a21oi_1 U23710 ( .A1(n17040), .A2(n16900), .B1(n16899), .Y(
        n16905) );
  sky130_fd_sc_hd__nand2_1 U23711 ( .A(n16903), .B(n16902), .Y(n16904) );
  sky130_fd_sc_hd__xor2_1 U23712 ( .A(n16905), .B(n16904), .X(n27853) );
  sky130_fd_sc_hd__nand2_1 U23713 ( .A(n27853), .B(n17225), .Y(n16906) );
  sky130_fd_sc_hd__nand3_2 U23714 ( .A(n16907), .B(n13055), .C(n16906), .Y(
        n21042) );
  sky130_fd_sc_hd__a22oi_1 U23715 ( .A1(n16909), .A2(
        j202_soc_core_j22_cpu_rfuo_sr__i__3_), .B1(
        j202_soc_core_j22_cpu_rfuo_sr__i__2_), .B2(n16908), .Y(n16916) );
  sky130_fd_sc_hd__nand2_1 U23716 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__1_), 
        .B(n16910), .Y(n16911) );
  sky130_fd_sc_hd__nand3_1 U23717 ( .A(n16911), .B(n21801), .C(
        j202_soc_core_intr_level__0_), .Y(n16914) );
  sky130_fd_sc_hd__nand2_1 U23718 ( .A(n22154), .B(
        j202_soc_core_intr_level__2_), .Y(n16913) );
  sky130_fd_sc_hd__nand2_1 U23719 ( .A(n22287), .B(
        j202_soc_core_intr_level__1_), .Y(n16912) );
  sky130_fd_sc_hd__nand3_1 U23720 ( .A(n16914), .B(n16913), .C(n16912), .Y(
        n16915) );
  sky130_fd_sc_hd__nand2_1 U23721 ( .A(n16916), .B(n16915), .Y(n16918) );
  sky130_fd_sc_hd__a21oi_1 U23722 ( .A1(n18866), .A2(
        j202_soc_core_intr_level__3_), .B1(j202_soc_core_intr_level__4_), .Y(
        n16917) );
  sky130_fd_sc_hd__a21oi_1 U23723 ( .A1(n16918), .A2(n16917), .B1(n28376), .Y(
        n28106) );
  sky130_fd_sc_hd__nand2_1 U23724 ( .A(n28109), .B(n28106), .Y(n28084) );
  sky130_fd_sc_hd__nand3_1 U23725 ( .A(n28084), .B(
        j202_soc_core_j22_cpu_ifetchl), .C(n24792), .Y(n21055) );
  sky130_fd_sc_hd__nor2_1 U23726 ( .A(n16919), .B(n29484), .Y(n16924) );
  sky130_fd_sc_hd__nand2_1 U23727 ( .A(n28109), .B(n19539), .Y(n24541) );
  sky130_fd_sc_hd__nand2_1 U23728 ( .A(n24541), .B(
        j202_soc_core_j22_cpu_id_opn_v_), .Y(n16920) );
  sky130_fd_sc_hd__nand2_1 U23729 ( .A(n16924), .B(n16920), .Y(n16923) );
  sky130_fd_sc_hd__mux2i_1 U23730 ( .A0(n16923), .A1(n16922), .S(n24302), .Y(
        n16932) );
  sky130_fd_sc_hd__nand2_1 U23731 ( .A(n28109), .B(n16933), .Y(n16929) );
  sky130_fd_sc_hd__nor2_1 U23732 ( .A(j202_soc_core_j22_cpu_ifetchl), .B(
        n29746), .Y(n24707) );
  sky130_fd_sc_hd__nor2_1 U23733 ( .A(n29088), .B(n24707), .Y(n16926) );
  sky130_fd_sc_hd__nand3_1 U23734 ( .A(n23643), .B(n19539), .C(n19429), .Y(
        n16925) );
  sky130_fd_sc_hd__and3_1 U23735 ( .A(n28084), .B(n16926), .C(n16925), .X(
        n16927) );
  sky130_fd_sc_hd__o21a_1 U23736 ( .A1(n16929), .A2(n16928), .B1(n16927), .X(
        n24710) );
  sky130_fd_sc_hd__nand2_1 U23737 ( .A(n29746), .B(n29745), .Y(n24588) );
  sky130_fd_sc_hd__nor3_1 U23738 ( .A(n16930), .B(n28340), .C(n24588), .Y(
        n16931) );
  sky130_fd_sc_hd__nand3_1 U23739 ( .A(n16932), .B(n24710), .C(n16931), .Y(
        n24589) );
  sky130_fd_sc_hd__nand2_1 U23740 ( .A(n24589), .B(n16934), .Y(n28384) );
  sky130_fd_sc_hd__nand2_1 U23741 ( .A(j202_soc_core_memory0_ram_dout0[156]), 
        .B(n21489), .Y(n16937) );
  sky130_fd_sc_hd__nand2_1 U23742 ( .A(j202_soc_core_memory0_ram_dout0[124]), 
        .B(n21488), .Y(n16936) );
  sky130_fd_sc_hd__nand2_1 U23743 ( .A(j202_soc_core_memory0_ram_dout0[92]), 
        .B(n21642), .Y(n16935) );
  sky130_fd_sc_hd__o31a_1 U23744 ( .A1(n19130), .A2(n18700), .A3(n19185), .B1(
        n16938), .X(n16939) );
  sky130_fd_sc_hd__nand4_1 U23745 ( .A(n16941), .B(n16940), .C(n16939), .D(
        n16963), .Y(n16954) );
  sky130_fd_sc_hd__nor2_1 U23746 ( .A(n16943), .B(n16942), .Y(n16948) );
  sky130_fd_sc_hd__a31oi_1 U23747 ( .A1(n16948), .A2(n16947), .A3(n16946), 
        .B1(n17009), .Y(n16953) );
  sky130_fd_sc_hd__o22ai_1 U23748 ( .A1(n17001), .A2(n16951), .B1(n16950), 
        .B2(n16949), .Y(n16952) );
  sky130_fd_sc_hd__a211o_1 U23749 ( .A1(n16954), .A2(n17099), .B1(n16953), 
        .C1(n16952), .X(n16955) );
  sky130_fd_sc_hd__nand2_1 U23750 ( .A(n16955), .B(n20784), .Y(n17024) );
  sky130_fd_sc_hd__nand2_1 U23751 ( .A(n20759), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[92]), .Y(n17019) );
  sky130_fd_sc_hd__nand2_1 U23752 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[28]), .Y(n17018) );
  sky130_fd_sc_hd__nand3_1 U23753 ( .A(n17019), .B(n21768), .C(n17018), .Y(
        n16958) );
  sky130_fd_sc_hd__nand2_1 U23754 ( .A(n20540), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[60]), .Y(n16957) );
  sky130_fd_sc_hd__nand2_1 U23755 ( .A(n21513), .B(j202_soc_core_uart_div0[4]), 
        .Y(n16956) );
  sky130_fd_sc_hd__nand2_1 U23756 ( .A(n16957), .B(n16956), .Y(n17020) );
  sky130_fd_sc_hd__nor2_1 U23757 ( .A(n16958), .B(n17020), .Y(n16975) );
  sky130_fd_sc_hd__nand4_1 U23758 ( .A(n16961), .B(n16960), .C(n17002), .D(
        n16959), .Y(n16962) );
  sky130_fd_sc_hd__o21ai_1 U23759 ( .A1(n16962), .A2(n16981), .B1(n16992), .Y(
        n16973) );
  sky130_fd_sc_hd__nand3_1 U23760 ( .A(n16965), .B(n16964), .C(n16963), .Y(
        n16966) );
  sky130_fd_sc_hd__nand2_1 U23761 ( .A(n16966), .B(n17099), .Y(n16972) );
  sky130_fd_sc_hd__nand2_1 U23763 ( .A(n16969), .B(n16994), .Y(n16970) );
  sky130_fd_sc_hd__nand4_1 U23764 ( .A(n16973), .B(n16972), .C(n16971), .D(
        n16970), .Y(n16974) );
  sky130_fd_sc_hd__nand2_1 U23765 ( .A(n16974), .B(n20643), .Y(n17022) );
  sky130_fd_sc_hd__nand3_1 U23766 ( .A(n17024), .B(n16975), .C(n17022), .Y(
        n17016) );
  sky130_fd_sc_hd__nand3_1 U23767 ( .A(n16979), .B(n16978), .C(n16977), .Y(
        n16982) );
  sky130_fd_sc_hd__o211ai_1 U23769 ( .A1(n16986), .A2(n16985), .B1(n16989), 
        .C1(n16984), .Y(n16993) );
  sky130_fd_sc_hd__nand4_1 U23770 ( .A(n16990), .B(n16989), .C(n16988), .D(
        n16987), .Y(n16991) );
  sky130_fd_sc_hd__a22oi_1 U23771 ( .A1(n16993), .A2(n16992), .B1(n16991), 
        .B2(n17099), .Y(n16999) );
  sky130_fd_sc_hd__nand2_1 U23772 ( .A(n16995), .B(n16994), .Y(n16998) );
  sky130_fd_sc_hd__a31oi_1 U23773 ( .A1(n17000), .A2(n16999), .A3(n16998), 
        .B1(n16997), .Y(n17015) );
  sky130_fd_sc_hd__a31oi_1 U23774 ( .A1(n17004), .A2(n17003), .A3(n17002), 
        .B1(n17001), .Y(n17013) );
  sky130_fd_sc_hd__o22ai_1 U23775 ( .A1(n17009), .A2(n17008), .B1(n17007), 
        .B2(n17006), .Y(n17012) );
  sky130_fd_sc_hd__o31a_1 U23776 ( .A1(n17013), .A2(n17012), .A3(n17011), .B1(
        n20508), .X(n17014) );
  sky130_fd_sc_hd__o21a_1 U23777 ( .A1(n17015), .A2(n17014), .B1(n21629), .X(
        n17025) );
  sky130_fd_sc_hd__nor2_1 U23778 ( .A(n17016), .B(n17025), .Y(n17017) );
  sky130_fd_sc_hd__nand2_1 U23779 ( .A(j202_soc_core_memory0_ram_dout0[508]), 
        .B(n21650), .Y(n17028) );
  sky130_fd_sc_hd__nand3_1 U23780 ( .A(n17019), .B(n17018), .C(n21653), .Y(
        n17021) );
  sky130_fd_sc_hd__nor2_1 U23781 ( .A(n17021), .B(n17020), .Y(n17023) );
  sky130_fd_sc_hd__nand3_1 U23782 ( .A(n17024), .B(n17023), .C(n17022), .Y(
        n17026) );
  sky130_fd_sc_hd__nor2_1 U23783 ( .A(n17026), .B(n17025), .Y(n17027) );
  sky130_fd_sc_hd__nand2_1 U23784 ( .A(n17028), .B(n17027), .Y(n20089) );
  sky130_fd_sc_hd__nand2_1 U23785 ( .A(n20090), .B(n20089), .Y(n26166) );
  sky130_fd_sc_hd__nand2_1 U23786 ( .A(n17029), .B(n17033), .Y(n17037) );
  sky130_fd_sc_hd__nor2_1 U23787 ( .A(n17037), .B(n17030), .Y(n17039) );
  sky130_fd_sc_hd__a21oi_1 U23788 ( .A1(n17034), .A2(n17033), .B1(n17032), .Y(
        n17035) );
  sky130_fd_sc_hd__o21ai_1 U23789 ( .A1(n17037), .A2(n17036), .B1(n17035), .Y(
        n17038) );
  sky130_fd_sc_hd__a21oi_1 U23790 ( .A1(n17040), .A2(n17039), .B1(n17038), .Y(
        n17045) );
  sky130_fd_sc_hd__nand2_1 U23791 ( .A(n17043), .B(n17042), .Y(n17044) );
  sky130_fd_sc_hd__xor2_1 U23792 ( .A(n17045), .B(n17044), .X(n25864) );
  sky130_fd_sc_hd__ha_1 U23793 ( .A(n17046), .B(j202_soc_core_j22_cpu_pc[28]), 
        .COUT(n16559), .SUM(n17047) );
  sky130_fd_sc_hd__a2bb2oi_1 U23794 ( .B1(n17048), .B2(n17047), .A1_N(n27026), 
        .A2_N(n11186), .Y(n17050) );
  sky130_fd_sc_hd__nand2_1 U23795 ( .A(n21924), .B(n25825), .Y(n17049) );
  sky130_fd_sc_hd__o211ai_1 U23796 ( .A1(n22705), .A2(n25862), .B1(n17050), 
        .C1(n17049), .Y(n17051) );
  sky130_fd_sc_hd__a21oi_1 U23797 ( .A1(n25864), .A2(n17225), .B1(n17051), .Y(
        n17052) );
  sky130_fd_sc_hd__nor2_1 U23798 ( .A(n17054), .B(n17095), .Y(n17055) );
  sky130_fd_sc_hd__nand3_1 U23799 ( .A(n17056), .B(n30029), .C(n17055), .Y(
        n28385) );
  sky130_fd_sc_hd__nor3_1 U23802 ( .A(n17061), .B(n17060), .C(n17059), .Y(
        n17062) );
  sky130_fd_sc_hd__nand4_1 U23803 ( .A(n17068), .B(n11103), .C(n17067), .D(
        n17066), .Y(n17076) );
  sky130_fd_sc_hd__nand2_1 U23805 ( .A(n17095), .B(n21042), .Y(n20894) );
  sky130_fd_sc_hd__nand2_1 U23806 ( .A(n20894), .B(n28384), .Y(n17073) );
  sky130_fd_sc_hd__nor2_2 U23807 ( .A(n17073), .B(n29436), .Y(n21188) );
  sky130_fd_sc_hd__nand3_1 U23808 ( .A(n20892), .B(n17074), .C(n12293), .Y(
        n17075) );
  sky130_fd_sc_hd__nor2_1 U23809 ( .A(n17076), .B(n17075), .Y(n17079) );
  sky130_fd_sc_hd__nor3_1 U23810 ( .A(n12334), .B(n12353), .C(n29479), .Y(
        n17077) );
  sky130_fd_sc_hd__nand4_1 U23811 ( .A(n20895), .B(n17079), .C(n17078), .D(
        n17077), .Y(n17092) );
  sky130_fd_sc_hd__nand2_1 U23812 ( .A(n12353), .B(n21042), .Y(n17081) );
  sky130_fd_sc_hd__inv_1 U23813 ( .A(n17095), .Y(n24143) );
  sky130_fd_sc_hd__nor2_1 U23814 ( .A(n17081), .B(n17080), .Y(n17089) );
  sky130_fd_sc_hd__and4_1 U23815 ( .A(n17084), .B(n17083), .C(n11208), .D(
        n17082), .X(n17086) );
  sky130_fd_sc_hd__nand3_1 U23816 ( .A(n17087), .B(n17086), .C(n17085), .Y(
        n17088) );
  sky130_fd_sc_hd__nor2_1 U23817 ( .A(n17092), .B(n30066), .Y(n24146) );
  sky130_fd_sc_hd__nor2_1 U23818 ( .A(io_in[14]), .B(n17093), .Y(n20889) );
  sky130_fd_sc_hd__nand2b_1 U23819 ( .A_N(n20889), .B(n17094), .Y(n17098) );
  sky130_fd_sc_hd__nand2_1 U23820 ( .A(n17095), .B(n17098), .Y(n17097) );
  sky130_fd_sc_hd__nand2_1 U23821 ( .A(n24143), .B(n12421), .Y(n17096) );
  sky130_fd_sc_hd__o211a_2 U23822 ( .A1(n17098), .A2(n12421), .B1(n17097), 
        .C1(n17096), .X(n24145) );
  sky130_fd_sc_hd__nand3_1 U23823 ( .A(n19143), .B(n19140), .C(n20673), .Y(
        n20371) );
  sky130_fd_sc_hd__nor2_1 U23824 ( .A(n13179), .B(n19145), .Y(n19136) );
  sky130_fd_sc_hd__nor2_1 U23825 ( .A(n19140), .B(n11150), .Y(n17160) );
  sky130_fd_sc_hd__nand2_1 U23826 ( .A(n19136), .B(n17160), .Y(n19562) );
  sky130_fd_sc_hd__nand2_1 U23827 ( .A(n18706), .B(n21359), .Y(n17123) );
  sky130_fd_sc_hd__nor2_1 U23828 ( .A(n20485), .B(n19125), .Y(n19159) );
  sky130_fd_sc_hd__nand2b_1 U23829 ( .A_N(n17123), .B(n19159), .Y(n20306) );
  sky130_fd_sc_hd__nand2_1 U23830 ( .A(n19562), .B(n20306), .Y(n20345) );
  sky130_fd_sc_hd__nor2_1 U23831 ( .A(n19608), .B(n20345), .Y(n19402) );
  sky130_fd_sc_hd__nand2_1 U23832 ( .A(n19159), .B(n18727), .Y(n19397) );
  sky130_fd_sc_hd__nor2_1 U23833 ( .A(n13179), .B(n19397), .Y(n20296) );
  sky130_fd_sc_hd__nand2_1 U23834 ( .A(n18706), .B(n13179), .Y(n20301) );
  sky130_fd_sc_hd__nor2_1 U23835 ( .A(n17243), .B(n20301), .Y(n19561) );
  sky130_fd_sc_hd__nand2_1 U23836 ( .A(n19561), .B(n20485), .Y(n20387) );
  sky130_fd_sc_hd__nand2b_1 U23837 ( .A_N(n17100), .B(n17099), .Y(n20293) );
  sky130_fd_sc_hd__nand3_1 U23838 ( .A(n20338), .B(n20387), .C(n20293), .Y(
        n20327) );
  sky130_fd_sc_hd__nor2_1 U23839 ( .A(n17104), .B(n19145), .Y(n19584) );
  sky130_fd_sc_hd__nand2_1 U23840 ( .A(n19584), .B(n21359), .Y(n20310) );
  sky130_fd_sc_hd__nand2_1 U23841 ( .A(n17101), .B(n11150), .Y(n19641) );
  sky130_fd_sc_hd__nand2_1 U23842 ( .A(n20310), .B(n19641), .Y(n19654) );
  sky130_fd_sc_hd__a31oi_1 U23843 ( .A1(n19402), .A2(n17103), .A3(n20317), 
        .B1(n17102), .Y(n17119) );
  sky130_fd_sc_hd__nor2_1 U23844 ( .A(n21359), .B(n19397), .Y(n19581) );
  sky130_fd_sc_hd__nor2_1 U23845 ( .A(n17104), .B(n20515), .Y(n20376) );
  sky130_fd_sc_hd__nand2_1 U23846 ( .A(n20376), .B(n21359), .Y(n20307) );
  sky130_fd_sc_hd__nor2_1 U23847 ( .A(n19581), .B(n17105), .Y(n17134) );
  sky130_fd_sc_hd__nand2_1 U23848 ( .A(n19143), .B(n18706), .Y(n20343) );
  sky130_fd_sc_hd__nand2b_1 U23849 ( .A_N(n20343), .B(n13179), .Y(n20360) );
  sky130_fd_sc_hd__nor2_1 U23850 ( .A(n13179), .B(n20515), .Y(n17150) );
  sky130_fd_sc_hd__nand2_1 U23851 ( .A(n17150), .B(n17160), .Y(n19575) );
  sky130_fd_sc_hd__nand3_1 U23852 ( .A(n19143), .B(n18727), .C(n13179), .Y(
        n20268) );
  sky130_fd_sc_hd__nand3_1 U23853 ( .A(n19132), .B(n21359), .C(n17160), .Y(
        n20348) );
  sky130_fd_sc_hd__and3_1 U23854 ( .A(n20360), .B(n19575), .C(n17106), .X(
        n19623) );
  sky130_fd_sc_hd__nand2_1 U23855 ( .A(n17160), .B(n13179), .Y(n17110) );
  sky130_fd_sc_hd__nor2_1 U23856 ( .A(n21595), .B(n17110), .Y(n17112) );
  sky130_fd_sc_hd__nor2_1 U23857 ( .A(n17112), .B(n17107), .Y(n17109) );
  sky130_fd_sc_hd__nand2_1 U23858 ( .A(n17251), .B(n13199), .Y(n19180) );
  sky130_fd_sc_hd__nor2_1 U23859 ( .A(n17108), .B(n19180), .Y(n20490) );
  sky130_fd_sc_hd__nand2_1 U23860 ( .A(n20490), .B(n19140), .Y(n20326) );
  sky130_fd_sc_hd__nand4_1 U23861 ( .A(n17134), .B(n19623), .C(n17109), .D(
        n20326), .Y(n17115) );
  sky130_fd_sc_hd__nand2_1 U23862 ( .A(n20809), .B(n17160), .Y(n19329) );
  sky130_fd_sc_hd__nand2_1 U23863 ( .A(n20360), .B(n19329), .Y(n19665) );
  sky130_fd_sc_hd__nor2_1 U23864 ( .A(n13182), .B(n19180), .Y(n19206) );
  sky130_fd_sc_hd__nand2_1 U23865 ( .A(n19206), .B(n19140), .Y(n19656) );
  sky130_fd_sc_hd__nor2_1 U23866 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n19656), .Y(n20381) );
  sky130_fd_sc_hd__nor2_1 U23867 ( .A(n19665), .B(n20381), .Y(n19350) );
  sky130_fd_sc_hd__nand2b_1 U23868 ( .A_N(n17110), .B(n21074), .Y(n20377) );
  sky130_fd_sc_hd__nor2_1 U23869 ( .A(n13199), .B(n20377), .Y(n19615) );
  sky130_fd_sc_hd__nand2_1 U23870 ( .A(n19132), .B(n18695), .Y(n19549) );
  sky130_fd_sc_hd__nand2b_1 U23871 ( .A_N(n19549), .B(n13179), .Y(n20389) );
  sky130_fd_sc_hd__nor2_1 U23872 ( .A(n19615), .B(n17111), .Y(n17113) );
  sky130_fd_sc_hd__nand2b_1 U23873 ( .A_N(n20301), .B(n19159), .Y(n19369) );
  sky130_fd_sc_hd__nand2_1 U23874 ( .A(n17112), .B(n13199), .Y(n19612) );
  sky130_fd_sc_hd__nand4_1 U23875 ( .A(n19350), .B(n17113), .C(n19369), .D(
        n19612), .Y(n17114) );
  sky130_fd_sc_hd__a22oi_1 U23876 ( .A1(n17115), .A2(n20368), .B1(n17114), 
        .B2(n20385), .Y(n17118) );
  sky130_fd_sc_hd__nand2_1 U23877 ( .A(n20303), .B(n20673), .Y(n20560) );
  sky130_fd_sc_hd__nand2b_1 U23878 ( .A_N(n19549), .B(n21359), .Y(n17162) );
  sky130_fd_sc_hd__nand2_1 U23879 ( .A(n20349), .B(n17162), .Y(n19664) );
  sky130_fd_sc_hd__nand3_1 U23880 ( .A(n20335), .B(n20317), .C(n20387), .Y(
        n17116) );
  sky130_fd_sc_hd__nand2_1 U23881 ( .A(n20277), .B(n20343), .Y(n20395) );
  sky130_fd_sc_hd__nor2_1 U23882 ( .A(n17148), .B(n19613), .Y(n20366) );
  sky130_fd_sc_hd__nand2b_1 U23883 ( .A_N(n20395), .B(n20366), .Y(n19317) );
  sky130_fd_sc_hd__nand3b_1 U23885 ( .A_N(n17119), .B(n17118), .C(n17117), .Y(
        n17120) );
  sky130_fd_sc_hd__nand2_1 U23886 ( .A(n17120), .B(n20757), .Y(n17185) );
  sky130_fd_sc_hd__nand2_1 U23887 ( .A(n20303), .B(n18727), .Y(n19348) );
  sky130_fd_sc_hd__nor2_1 U23888 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n19348), .Y(n19319) );
  sky130_fd_sc_hd__nand3_1 U23889 ( .A(n20809), .B(n18695), .C(n13179), .Y(
        n20339) );
  sky130_fd_sc_hd__nand3_1 U23890 ( .A(n20363), .B(n20339), .C(n20307), .Y(
        n17121) );
  sky130_fd_sc_hd__nor2_1 U23891 ( .A(n17121), .B(n20395), .Y(n17171) );
  sky130_fd_sc_hd__nand2b_1 U23892 ( .A_N(n17123), .B(n17122), .Y(n20372) );
  sky130_fd_sc_hd__nand2_1 U23893 ( .A(n20372), .B(n20306), .Y(n19555) );
  sky130_fd_sc_hd__nor2_1 U23894 ( .A(n19555), .B(n19392), .Y(n19585) );
  sky130_fd_sc_hd__nand2b_1 U23895 ( .A_N(n19329), .B(n21359), .Y(n20289) );
  sky130_fd_sc_hd__nand2_1 U23896 ( .A(n20289), .B(n20377), .Y(n17124) );
  sky130_fd_sc_hd__nor2_1 U23897 ( .A(n17124), .B(n19664), .Y(n17125) );
  sky130_fd_sc_hd__nand4_1 U23898 ( .A(n17171), .B(n19585), .C(n17125), .D(
        n20338), .Y(n17126) );
  sky130_fd_sc_hd__nand2_1 U23899 ( .A(n17126), .B(n20374), .Y(n17145) );
  sky130_fd_sc_hd__nor2_1 U23900 ( .A(n20376), .B(n17127), .Y(n17128) );
  sky130_fd_sc_hd__nand3_1 U23901 ( .A(n17128), .B(n20310), .C(n20344), .Y(
        n19373) );
  sky130_fd_sc_hd__nand3_1 U23902 ( .A(n20360), .B(n20387), .C(n20268), .Y(
        n17131) );
  sky130_fd_sc_hd__nand2_1 U23903 ( .A(n18695), .B(n21359), .Y(n20388) );
  sky130_fd_sc_hd__nand2b_1 U23904 ( .A_N(n20388), .B(n20809), .Y(n20364) );
  sky130_fd_sc_hd__nand2_1 U23905 ( .A(n19369), .B(n20364), .Y(n17129) );
  sky130_fd_sc_hd__nor2_1 U23906 ( .A(n17129), .B(n19615), .Y(n17130) );
  sky130_fd_sc_hd__nand4b_1 U23907 ( .A_N(n17131), .B(n17130), .C(n20326), .D(
        n20389), .Y(n17132) );
  sky130_fd_sc_hd__o21ai_0 U23908 ( .A1(n19373), .A2(n17132), .B1(n20368), .Y(
        n17144) );
  sky130_fd_sc_hd__nand3_1 U23909 ( .A(n20347), .B(n17133), .C(n20306), .Y(
        n19322) );
  sky130_fd_sc_hd__nor2_1 U23910 ( .A(n19322), .B(n17135), .Y(n19652) );
  sky130_fd_sc_hd__nand2b_1 U23911 ( .A_N(n19329), .B(n13179), .Y(n19571) );
  sky130_fd_sc_hd__nand2_1 U23912 ( .A(n19571), .B(n20364), .Y(n20291) );
  sky130_fd_sc_hd__nor2_1 U23913 ( .A(n13179), .B(n20343), .Y(n19370) );
  sky130_fd_sc_hd__nor2_1 U23914 ( .A(n20485), .B(n20377), .Y(n19574) );
  sky130_fd_sc_hd__nand2b_1 U23915 ( .A_N(n19574), .B(n20349), .Y(n19579) );
  sky130_fd_sc_hd__nor2_1 U23916 ( .A(n19370), .B(n19579), .Y(n17136) );
  sky130_fd_sc_hd__nand4_1 U23917 ( .A(n19652), .B(n20317), .C(n19544), .D(
        n17136), .Y(n17137) );
  sky130_fd_sc_hd__nand2_1 U23918 ( .A(n17137), .B(n20385), .Y(n17143) );
  sky130_fd_sc_hd__nand2_1 U23919 ( .A(n19549), .B(n20339), .Y(n20362) );
  sky130_fd_sc_hd__nand4b_1 U23920 ( .A_N(n20296), .B(n20326), .C(n19571), .D(
        n20307), .Y(n19643) );
  sky130_fd_sc_hd__nor2_1 U23921 ( .A(n20362), .B(n19643), .Y(n19377) );
  sky130_fd_sc_hd__nor2_1 U23922 ( .A(n19584), .B(n19559), .Y(n17140) );
  sky130_fd_sc_hd__nor2_1 U23923 ( .A(n19574), .B(n17138), .Y(n17139) );
  sky130_fd_sc_hd__nand4_1 U23924 ( .A(n19377), .B(n19585), .C(n17140), .D(
        n17139), .Y(n17141) );
  sky130_fd_sc_hd__nand2_1 U23925 ( .A(n17141), .B(n20393), .Y(n17142) );
  sky130_fd_sc_hd__nand4_1 U23926 ( .A(n17145), .B(n17144), .C(n17143), .D(
        n17142), .Y(n17147) );
  sky130_fd_sc_hd__nand2_1 U23927 ( .A(n17147), .B(n20617), .Y(n17184) );
  sky130_fd_sc_hd__nand2_1 U23928 ( .A(n20326), .B(n20348), .Y(n20314) );
  sky130_fd_sc_hd__nor2_1 U23929 ( .A(n17148), .B(n20314), .Y(n20280) );
  sky130_fd_sc_hd__nand4_1 U23930 ( .A(n20280), .B(n19575), .C(n19622), .D(
        n20277), .Y(n19374) );
  sky130_fd_sc_hd__nand2_1 U23931 ( .A(n19584), .B(n13179), .Y(n19649) );
  sky130_fd_sc_hd__nand2_1 U23932 ( .A(n19649), .B(n19612), .Y(n20297) );
  sky130_fd_sc_hd__nor2_1 U23933 ( .A(n19574), .B(n20297), .Y(n19565) );
  sky130_fd_sc_hd__nor2_1 U23934 ( .A(n19615), .B(n19319), .Y(n17149) );
  sky130_fd_sc_hd__nand2_1 U23935 ( .A(n20376), .B(n13179), .Y(n20390) );
  sky130_fd_sc_hd__nand3_1 U23936 ( .A(n19565), .B(n17149), .C(n20390), .Y(
        n20272) );
  sky130_fd_sc_hd__o21ai_1 U23937 ( .A1(n19374), .A2(n20272), .B1(n20374), .Y(
        n17169) );
  sky130_fd_sc_hd__nor2_1 U23938 ( .A(n19559), .B(n19370), .Y(n20316) );
  sky130_fd_sc_hd__nor2_1 U23939 ( .A(n20043), .B(n17151), .Y(n20315) );
  sky130_fd_sc_hd__nor2_1 U23940 ( .A(n17152), .B(n20315), .Y(n19405) );
  sky130_fd_sc_hd__and4_1 U23941 ( .A(n19405), .B(n20366), .C(n20326), .D(
        n20363), .X(n17153) );
  sky130_fd_sc_hd__nand3_1 U23942 ( .A(n19617), .B(n17153), .C(n19565), .Y(
        n17154) );
  sky130_fd_sc_hd__nand2_1 U23943 ( .A(n17154), .B(n20368), .Y(n17168) );
  sky130_fd_sc_hd__nand4b_1 U23944 ( .A_N(n19615), .B(n20349), .C(n20307), .D(
        n19649), .Y(n17155) );
  sky130_fd_sc_hd__nand2_1 U23945 ( .A(n19561), .B(n13199), .Y(n20379) );
  sky130_fd_sc_hd__nand2_1 U23946 ( .A(n17156), .B(n20673), .Y(n17157) );
  sky130_fd_sc_hd__nand2_1 U23947 ( .A(n20379), .B(n17157), .Y(n19398) );
  sky130_fd_sc_hd__nand3_1 U23948 ( .A(n19402), .B(n19371), .C(n17158), .Y(
        n17159) );
  sky130_fd_sc_hd__nand2_1 U23949 ( .A(n17159), .B(n20385), .Y(n17167) );
  sky130_fd_sc_hd__nand2_1 U23951 ( .A(n20326), .B(n17162), .Y(n19344) );
  sky130_fd_sc_hd__nor3_1 U23952 ( .A(n20296), .B(n17163), .C(n19344), .Y(
        n17164) );
  sky130_fd_sc_hd__nand2_1 U23953 ( .A(n19565), .B(n17164), .Y(n17165) );
  sky130_fd_sc_hd__nand2_1 U23954 ( .A(n17165), .B(n20393), .Y(n17166) );
  sky130_fd_sc_hd__nand4_1 U23955 ( .A(n17169), .B(n17168), .C(n17167), .D(
        n17166), .Y(n17170) );
  sky130_fd_sc_hd__nand2_1 U23956 ( .A(n17170), .B(n20784), .Y(n17183) );
  sky130_fd_sc_hd__nand2_1 U23957 ( .A(n20310), .B(n20339), .Y(n19580) );
  sky130_fd_sc_hd__o21ai_0 U23958 ( .A1(n19580), .A2(n19317), .B1(n20374), .Y(
        n17180) );
  sky130_fd_sc_hd__and3_1 U23959 ( .A(n20379), .B(n20389), .C(n20371), .X(
        n19345) );
  sky130_fd_sc_hd__nand4_1 U23960 ( .A(n17171), .B(n19345), .C(n19571), .D(
        n19575), .Y(n17172) );
  sky130_fd_sc_hd__nand2_1 U23961 ( .A(n17172), .B(n20368), .Y(n17179) );
  sky130_fd_sc_hd__nand3_1 U23962 ( .A(n19544), .B(n20390), .C(n20306), .Y(
        n19576) );
  sky130_fd_sc_hd__nand2_1 U23963 ( .A(n20387), .B(n19575), .Y(n19651) );
  sky130_fd_sc_hd__nor2_1 U23964 ( .A(n19651), .B(n20381), .Y(n20367) );
  sky130_fd_sc_hd__nand2_1 U23965 ( .A(n20310), .B(n20389), .Y(n20350) );
  sky130_fd_sc_hd__nand4_1 U23966 ( .A(n19552), .B(n20367), .C(n20334), .D(
        n19562), .Y(n17173) );
  sky130_fd_sc_hd__nand2_1 U23967 ( .A(n17173), .B(n20393), .Y(n17178) );
  sky130_fd_sc_hd__nand2_1 U23968 ( .A(n19562), .B(n20289), .Y(n19321) );
  sky130_fd_sc_hd__nor2_1 U23969 ( .A(n19554), .B(n19321), .Y(n19346) );
  sky130_fd_sc_hd__nand3_1 U23970 ( .A(n20360), .B(n20326), .C(n20377), .Y(
        n17174) );
  sky130_fd_sc_hd__nor2_1 U23971 ( .A(n17174), .B(n20350), .Y(n17175) );
  sky130_fd_sc_hd__nand2_1 U23972 ( .A(n19346), .B(n17175), .Y(n17176) );
  sky130_fd_sc_hd__nand2_1 U23973 ( .A(n17176), .B(n20385), .Y(n17177) );
  sky130_fd_sc_hd__nand4_1 U23974 ( .A(n17180), .B(n17179), .C(n17178), .D(
        n17177), .Y(n17181) );
  sky130_fd_sc_hd__nand2_1 U23975 ( .A(n17181), .B(n20643), .Y(n17182) );
  sky130_fd_sc_hd__nand4_1 U23976 ( .A(n17185), .B(n17184), .C(n17183), .D(
        n17182), .Y(n17213) );
  sky130_fd_sc_hd__nor2_1 U23977 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[1]), 
        .B(n27957), .Y(n24720) );
  sky130_fd_sc_hd__a22oi_1 U23978 ( .A1(n24720), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[18]), .B1(n21505), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[2]), .Y(n17187) );
  sky130_fd_sc_hd__nor2_1 U23979 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[0]), 
        .B(n24722), .Y(n21504) );
  sky130_fd_sc_hd__nor2_1 U23980 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[0]), 
        .B(j202_soc_core_uart_TOP_rx_fifo_rp[1]), .Y(n21506) );
  sky130_fd_sc_hd__a22oi_1 U23981 ( .A1(n21504), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[10]), .B1(n21506), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[26]), .Y(n17186) );
  sky130_fd_sc_hd__nand2_1 U23982 ( .A(n17187), .B(n17186), .Y(n17188) );
  sky130_fd_sc_hd__nand2_1 U23983 ( .A(n21513), .B(n17188), .Y(n17194) );
  sky130_fd_sc_hd__nor2_1 U23984 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[2]), .B(n17189), .Y(n17191) );
  sky130_fd_sc_hd__nand3_1 U23985 ( .A(n17192), .B(n17191), .C(n17190), .Y(
        n21519) );
  sky130_fd_sc_hd__nand2_1 U23986 ( .A(n21446), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[98]), .Y(n17193) );
  sky130_fd_sc_hd__nand2_1 U23987 ( .A(n17194), .B(n17193), .Y(n17206) );
  sky130_fd_sc_hd__nand2_1 U23988 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[2]), .Y(n17195) );
  sky130_fd_sc_hd__o21a_1 U23989 ( .A1(n17196), .A2(n21512), .B1(n17195), .X(
        n17208) );
  sky130_fd_sc_hd__nand2b_1 U23990 ( .A_N(n21515), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[34]), .Y(n17207) );
  sky130_fd_sc_hd__nand3_1 U23991 ( .A(n17208), .B(n17207), .C(n21768), .Y(
        n17197) );
  sky130_fd_sc_hd__nor2_1 U23992 ( .A(n17206), .B(n17197), .Y(n17204) );
  sky130_fd_sc_hd__mux2_2 U23993 ( .A0(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[2]), .A1(
        j202_soc_core_aquc_ADR__2_), .S(n29435), .X(n28203) );
  sky130_fd_sc_hd__or4_1 U23994 ( .A(n29435), .B(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[7]), .C(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[5]), .D(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[6]), .X(n17199) );
  sky130_fd_sc_hd__a21oi_1 U23995 ( .A1(n17200), .A2(n17199), .B1(n17198), .Y(
        n28202) );
  sky130_fd_sc_hd__and3_1 U23996 ( .A(n29435), .B(n28202), .C(
        j202_soc_core_aquc_ADR__3_), .X(n17201) );
  sky130_fd_sc_hd__nand3_1 U23997 ( .A(n28164), .B(n28203), .C(n17201), .Y(
        n19595) );
  sky130_fd_sc_hd__nand3_1 U23998 ( .A(n19598), .B(j202_soc_core_aquc_ADR__3_), 
        .C(n28164), .Y(n19600) );
  sky130_fd_sc_hd__o22ai_1 U23999 ( .A1(n29119), .A2(n19595), .B1(n17202), 
        .B2(n19600), .Y(n17203) );
  sky130_fd_sc_hd__nand2_1 U24000 ( .A(n17203), .B(n19605), .Y(n17214) );
  sky130_fd_sc_hd__nand2_1 U24001 ( .A(n20786), .B(
        j202_soc_core_bldc_core_00_pwm_period[2]), .Y(n17210) );
  sky130_fd_sc_hd__nand4b_1 U24002 ( .A_N(n17213), .B(n17204), .C(n17214), .D(
        n17210), .Y(n17205) );
  sky130_fd_sc_hd__nand2_1 U24003 ( .A(j202_soc_core_memory0_ram_dout0[482]), 
        .B(n21650), .Y(n17217) );
  sky130_fd_sc_hd__nand4_1 U24004 ( .A(n17209), .B(n17208), .C(n21653), .D(
        n17207), .Y(n17212) );
  sky130_fd_sc_hd__nor2_1 U24005 ( .A(n17212), .B(n17211), .Y(n17216) );
  sky130_fd_sc_hd__nand4_1 U24006 ( .A(n17217), .B(n17216), .C(n17215), .D(
        n17214), .Y(n17218) );
  sky130_fd_sc_hd__nand2_1 U24007 ( .A(n20255), .B(n22739), .Y(n17231) );
  sky130_fd_sc_hd__xnor2_1 U24008 ( .A(j202_soc_core_j22_cpu_pc[1]), .B(n13913), .Y(n27125) );
  sky130_fd_sc_hd__nand2_1 U24009 ( .A(n17221), .B(n17220), .Y(n17224) );
  sky130_fd_sc_hd__o21ai_0 U24010 ( .A1(n20431), .A2(n20435), .B1(n20432), .Y(
        n17223) );
  sky130_fd_sc_hd__xnor2_1 U24011 ( .A(n17224), .B(n17223), .Y(n24048) );
  sky130_fd_sc_hd__a22oi_1 U24012 ( .A1(n21322), .A2(n27125), .B1(n24048), 
        .B2(n17225), .Y(n17230) );
  sky130_fd_sc_hd__nand2_1 U24013 ( .A(n22701), .B(n28521), .Y(n17227) );
  sky130_fd_sc_hd__o211a_2 U24014 ( .A1(n26937), .A2(n22745), .B1(n17228), 
        .C1(n17227), .X(n17229) );
  sky130_fd_sc_hd__nand3_1 U24015 ( .A(n17231), .B(n17230), .C(n17229), .Y(
        n29557) );
  sky130_fd_sc_hd__nor2_1 U24016 ( .A(n19148), .B(n13179), .Y(n18724) );
  sky130_fd_sc_hd__nand2_1 U24017 ( .A(n18715), .B(n18724), .Y(n21097) );
  sky130_fd_sc_hd__nand2b_1 U24018 ( .A_N(n21097), .B(n19130), .Y(n21380) );
  sky130_fd_sc_hd__nand2_1 U24019 ( .A(n18715), .B(n21075), .Y(n20058) );
  sky130_fd_sc_hd__nand2_1 U24020 ( .A(n18715), .B(n17237), .Y(n21527) );
  sky130_fd_sc_hd__nand2b_1 U24021 ( .A_N(n21527), .B(n13179), .Y(n21572) );
  sky130_fd_sc_hd__nand3_1 U24022 ( .A(n18715), .B(n21359), .C(n19804), .Y(
        n21364) );
  sky130_fd_sc_hd__nand2_1 U24023 ( .A(n21572), .B(n21364), .Y(n21137) );
  sky130_fd_sc_hd__nand2_1 U24024 ( .A(n17242), .B(n13182), .Y(n17238) );
  sky130_fd_sc_hd__nor2_1 U24025 ( .A(n17238), .B(n21132), .Y(n21142) );
  sky130_fd_sc_hd__nand2_1 U24026 ( .A(n21142), .B(n19148), .Y(n21362) );
  sky130_fd_sc_hd__nor2_1 U24027 ( .A(n21595), .B(n17238), .Y(n21613) );
  sky130_fd_sc_hd__nand2_1 U24028 ( .A(n21613), .B(n19148), .Y(n21574) );
  sky130_fd_sc_hd__nand2_1 U24029 ( .A(n21362), .B(n21574), .Y(n17282) );
  sky130_fd_sc_hd__nor2_1 U24030 ( .A(n21137), .B(n17282), .Y(n21098) );
  sky130_fd_sc_hd__o22ai_1 U24031 ( .A1(n21412), .A2(n21386), .B1(n21395), 
        .B2(n21098), .Y(n17249) );
  sky130_fd_sc_hd__nor3_1 U24032 ( .A(n11150), .B(n21595), .C(n17239), .Y(
        n17285) );
  sky130_fd_sc_hd__nand3_1 U24033 ( .A(n21104), .B(n17251), .C(n17240), .Y(
        n21575) );
  sky130_fd_sc_hd__nand3_1 U24034 ( .A(n17241), .B(n21104), .C(n21103), .Y(
        n21567) );
  sky130_fd_sc_hd__nand3b_1 U24035 ( .A_N(n17285), .B(n21575), .C(n21567), .Y(
        n17245) );
  sky130_fd_sc_hd__nand2_1 U24036 ( .A(n17242), .B(n11150), .Y(n17254) );
  sky130_fd_sc_hd__nor2_1 U24037 ( .A(n17243), .B(n17254), .Y(n17272) );
  sky130_fd_sc_hd__nor2_1 U24038 ( .A(n19148), .B(n11150), .Y(n17244) );
  sky130_fd_sc_hd__nand3_1 U24039 ( .A(n21104), .B(n21074), .C(n17244), .Y(
        n21415) );
  sky130_fd_sc_hd__nand3_1 U24040 ( .A(n21554), .B(n21415), .C(n21527), .Y(
        n21401) );
  sky130_fd_sc_hd__nor3_1 U24041 ( .A(n17245), .B(n21401), .C(n17282), .Y(
        n17247) );
  sky130_fd_sc_hd__nor2_1 U24042 ( .A(n13179), .B(n21527), .Y(n21556) );
  sky130_fd_sc_hd__nand3_1 U24043 ( .A(n21104), .B(n19148), .C(n17250), .Y(
        n21583) );
  sky130_fd_sc_hd__nand3b_1 U24044 ( .A_N(n17282), .B(n17259), .C(n21583), .Y(
        n21522) );
  sky130_fd_sc_hd__o21ai_1 U24045 ( .A1(n21389), .A2(n21522), .B1(n21610), .Y(
        n17246) );
  sky130_fd_sc_hd__o21ai_1 U24046 ( .A1(n17247), .A2(n21150), .B1(n17246), .Y(
        n17248) );
  sky130_fd_sc_hd__nor2_1 U24047 ( .A(n17249), .B(n17248), .Y(n17304) );
  sky130_fd_sc_hd__nand2_1 U24048 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .B(n19140), .Y(n21405) );
  sky130_fd_sc_hd__nor2_1 U24049 ( .A(n17265), .B(n19125), .Y(n17281) );
  sky130_fd_sc_hd__nand2_1 U24050 ( .A(n17281), .B(n18752), .Y(n21550) );
  sky130_fd_sc_hd__nand3_1 U24051 ( .A(n21104), .B(n17250), .C(n19804), .Y(
        n21573) );
  sky130_fd_sc_hd__nand2_1 U24052 ( .A(n21550), .B(n21573), .Y(n21530) );
  sky130_fd_sc_hd__nor2_1 U24053 ( .A(n13182), .B(n17269), .Y(n17255) );
  sky130_fd_sc_hd__nand2_1 U24054 ( .A(n17255), .B(n21101), .Y(n21096) );
  sky130_fd_sc_hd__nand2_1 U24055 ( .A(n18742), .B(n17251), .Y(n17267) );
  sky130_fd_sc_hd__nand3_1 U24056 ( .A(n21096), .B(n21575), .C(n21593), .Y(
        n17252) );
  sky130_fd_sc_hd__nor2_1 U24057 ( .A(n21530), .B(n17252), .Y(n21376) );
  sky130_fd_sc_hd__nand2_1 U24058 ( .A(n21376), .B(n21574), .Y(n17253) );
  sky130_fd_sc_hd__nand2_1 U24059 ( .A(n17253), .B(n21603), .Y(n17263) );
  sky130_fd_sc_hd__nand3_1 U24060 ( .A(n21399), .B(n21415), .C(n21536), .Y(
        n17257) );
  sky130_fd_sc_hd__nor2_1 U24061 ( .A(n17272), .B(n21082), .Y(n17256) );
  sky130_fd_sc_hd__nand2_1 U24062 ( .A(n17255), .B(n21104), .Y(n21616) );
  sky130_fd_sc_hd__nand4b_1 U24063 ( .A_N(n17257), .B(n17256), .C(n21616), .D(
        n21572), .Y(n17258) );
  sky130_fd_sc_hd__nand2_1 U24064 ( .A(n17258), .B(n21617), .Y(n17262) );
  sky130_fd_sc_hd__nand2_1 U24065 ( .A(n18715), .B(n21103), .Y(n21375) );
  sky130_fd_sc_hd__nand2_1 U24066 ( .A(n17259), .B(n21375), .Y(n21107) );
  sky130_fd_sc_hd__nor2_1 U24068 ( .A(n21145), .B(n21571), .Y(n21127) );
  sky130_fd_sc_hd__o21a_1 U24069 ( .A1(n21127), .A2(n21532), .B1(n21610), .X(
        n21124) );
  sky130_fd_sc_hd__nand4_1 U24070 ( .A(n17263), .B(n17262), .C(n17261), .D(
        n17290), .Y(n17280) );
  sky130_fd_sc_hd__nor2_1 U24071 ( .A(n19140), .B(n17264), .Y(n21624) );
  sky130_fd_sc_hd__nand2_1 U24072 ( .A(n18724), .B(n18712), .Y(n18707) );
  sky130_fd_sc_hd__nor2_1 U24073 ( .A(n17265), .B(n18707), .Y(n18716) );
  sky130_fd_sc_hd__nand3_1 U24074 ( .A(n21616), .B(n20166), .C(n21574), .Y(
        n17266) );
  sky130_fd_sc_hd__nor2_1 U24075 ( .A(n17265), .B(n17269), .Y(n17291) );
  sky130_fd_sc_hd__nand2_1 U24076 ( .A(n17291), .B(n21359), .Y(n21568) );
  sky130_fd_sc_hd__nand2_1 U24077 ( .A(n21568), .B(n21364), .Y(n21148) );
  sky130_fd_sc_hd__nor2_1 U24078 ( .A(n17266), .B(n21148), .Y(n21547) );
  sky130_fd_sc_hd__nor2_1 U24079 ( .A(n18731), .B(n17267), .Y(n21525) );
  sky130_fd_sc_hd__nand2b_1 U24080 ( .A_N(n17269), .B(n17268), .Y(n21606) );
  sky130_fd_sc_hd__nand4_1 U24081 ( .A(n21547), .B(n21570), .C(n21399), .D(
        n21606), .Y(n17270) );
  sky130_fd_sc_hd__nand2_1 U24082 ( .A(n17270), .B(n21598), .Y(n17278) );
  sky130_fd_sc_hd__nand2_1 U24083 ( .A(n21362), .B(n21567), .Y(n21139) );
  sky130_fd_sc_hd__nor2_1 U24084 ( .A(n21146), .B(n21122), .Y(n17273) );
  sky130_fd_sc_hd__nand2_1 U24085 ( .A(n17271), .B(n21075), .Y(n21384) );
  sky130_fd_sc_hd__nand2_1 U24086 ( .A(n17291), .B(n13179), .Y(n21365) );
  sky130_fd_sc_hd__nand4_1 U24087 ( .A(n17273), .B(n21384), .C(n21615), .D(
        n21365), .Y(n17274) );
  sky130_fd_sc_hd__a22oi_1 U24088 ( .A1(n21139), .A2(n21617), .B1(n17274), 
        .B2(n21603), .Y(n17277) );
  sky130_fd_sc_hd__nor2_1 U24089 ( .A(n21101), .B(n21571), .Y(n21426) );
  sky130_fd_sc_hd__nand3_1 U24090 ( .A(n21521), .B(n17287), .C(n21567), .Y(
        n21552) );
  sky130_fd_sc_hd__nand4_1 U24091 ( .A(n21538), .B(n21125), .C(n17288), .D(
        n21575), .Y(n17275) );
  sky130_fd_sc_hd__nand2_1 U24092 ( .A(n17275), .B(n21610), .Y(n17276) );
  sky130_fd_sc_hd__nand3_1 U24093 ( .A(n17278), .B(n17277), .C(n17276), .Y(
        n17279) );
  sky130_fd_sc_hd__nor2_1 U24094 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .B(n18744), .Y(n21591) );
  sky130_fd_sc_hd__a22oi_1 U24095 ( .A1(n17280), .A2(n21624), .B1(n17279), 
        .B2(n21591), .Y(n17303) );
  sky130_fd_sc_hd__nand2_1 U24096 ( .A(n17281), .B(n18724), .Y(n21607) );
  sky130_fd_sc_hd__nand2_1 U24097 ( .A(n21607), .B(n21573), .Y(n17289) );
  sky130_fd_sc_hd__nand3_1 U24098 ( .A(n18752), .B(n21360), .C(n21074), .Y(
        n21421) );
  sky130_fd_sc_hd__nand2_1 U24099 ( .A(n21413), .B(n21428), .Y(n17283) );
  sky130_fd_sc_hd__nor3_1 U24100 ( .A(n17284), .B(n17289), .C(n17283), .Y(
        n17300) );
  sky130_fd_sc_hd__nand2_1 U24101 ( .A(n21607), .B(n21421), .Y(n17286) );
  sky130_fd_sc_hd__nand2_1 U24102 ( .A(n17285), .B(n19148), .Y(n21110) );
  sky130_fd_sc_hd__nand2_1 U24103 ( .A(n21110), .B(n21384), .Y(n21353) );
  sky130_fd_sc_hd__nor2_1 U24104 ( .A(n17286), .B(n21353), .Y(n21569) );
  sky130_fd_sc_hd__nand2_1 U24105 ( .A(n21554), .B(n21570), .Y(n21599) );
  sky130_fd_sc_hd__a31oi_1 U24106 ( .A1(n21569), .A2(n17287), .A3(n21423), 
        .B1(n21150), .Y(n17298) );
  sky130_fd_sc_hd__nand2_1 U24107 ( .A(n21572), .B(n17293), .Y(n21349) );
  sky130_fd_sc_hd__nor2_1 U24108 ( .A(n17289), .B(n21349), .Y(n21419) );
  sky130_fd_sc_hd__nand2_1 U24110 ( .A(n21600), .B(n13179), .Y(n21388) );
  sky130_fd_sc_hd__nand2_1 U24111 ( .A(n21380), .B(n21388), .Y(n17295) );
  sky130_fd_sc_hd__nand3_1 U24112 ( .A(n21384), .B(n21355), .C(n21550), .Y(
        n21605) );
  sky130_fd_sc_hd__nor2_1 U24113 ( .A(n21525), .B(n21605), .Y(n21597) );
  sky130_fd_sc_hd__nand2_1 U24114 ( .A(n21102), .B(n21104), .Y(n17292) );
  sky130_fd_sc_hd__nand2_1 U24115 ( .A(n21597), .B(n17292), .Y(n21565) );
  sky130_fd_sc_hd__nand2_1 U24116 ( .A(n17293), .B(n21575), .Y(n21141) );
  sky130_fd_sc_hd__nor2_1 U24117 ( .A(n17294), .B(n21141), .Y(n21584) );
  sky130_fd_sc_hd__nand2b_1 U24118 ( .A_N(n21565), .B(n21584), .Y(n21099) );
  sky130_fd_sc_hd__o21a_1 U24119 ( .A1(n17295), .A2(n21099), .B1(n21603), .X(
        n17296) );
  sky130_fd_sc_hd__nor3_1 U24120 ( .A(n17298), .B(n17297), .C(n17296), .Y(
        n17299) );
  sky130_fd_sc_hd__nor2_1 U24122 ( .A(n19140), .B(
        j202_soc_core_bootrom_00_address_w[8]), .Y(n21589) );
  sky130_fd_sc_hd__nand2_1 U24123 ( .A(n17301), .B(n21589), .Y(n17302) );
  sky130_fd_sc_hd__o211ai_1 U24124 ( .A1(n17304), .A2(n21405), .B1(n17303), 
        .C1(n17302), .Y(n17305) );
  sky130_fd_sc_hd__nand2_1 U24125 ( .A(n17305), .B(n21629), .Y(n17330) );
  sky130_fd_sc_hd__nand2b_1 U24126 ( .A_N(n21515), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[39]), .Y(n17324) );
  sky130_fd_sc_hd__nand2_1 U24127 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[7]), .Y(n17323) );
  sky130_fd_sc_hd__nand3_1 U24128 ( .A(n17324), .B(n21768), .C(n17323), .Y(
        n17314) );
  sky130_fd_sc_hd__o22a_1 U24129 ( .A1(n17307), .A2(n21512), .B1(n17306), .B2(
        n21519), .X(n17322) );
  sky130_fd_sc_hd__nand2_1 U24130 ( .A(n21504), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[15]), .Y(n17311) );
  sky130_fd_sc_hd__nand2_1 U24131 ( .A(n24720), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[23]), .Y(n17310) );
  sky130_fd_sc_hd__nand2_1 U24132 ( .A(n21505), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[7]), .Y(n17309) );
  sky130_fd_sc_hd__nand2_1 U24133 ( .A(n21506), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[31]), .Y(n17308) );
  sky130_fd_sc_hd__nand4_1 U24134 ( .A(n17311), .B(n17310), .C(n17309), .D(
        n17308), .Y(n17312) );
  sky130_fd_sc_hd__nand2_1 U24135 ( .A(n21513), .B(n17312), .Y(n17325) );
  sky130_fd_sc_hd__nand2_1 U24136 ( .A(n17322), .B(n17325), .Y(n17313) );
  sky130_fd_sc_hd__nor2_1 U24137 ( .A(n17314), .B(n17313), .Y(n17315) );
  sky130_fd_sc_hd__nand2_1 U24138 ( .A(n20786), .B(
        j202_soc_core_bldc_core_00_pwm_period[7]), .Y(n17326) );
  sky130_fd_sc_hd__nand3_1 U24139 ( .A(n17330), .B(n17315), .C(n17326), .Y(
        n17316) );
  sky130_fd_sc_hd__a21oi_1 U24140 ( .A1(j202_soc_core_memory0_ram_dout0[455]), 
        .A2(j202_soc_core_memory0_ram_dout0_sel[14]), .B1(n17316), .Y(n17318)
         );
  sky130_fd_sc_hd__nand4_1 U24141 ( .A(n17320), .B(n17319), .C(n17318), .D(
        n17317), .Y(n17321) );
  sky130_fd_sc_hd__nand2_1 U24142 ( .A(j202_soc_core_memory0_ram_dout0[487]), 
        .B(n21650), .Y(n17332) );
  sky130_fd_sc_hd__nand4_1 U24143 ( .A(n17325), .B(n17324), .C(n21653), .D(
        n17323), .Y(n17328) );
  sky130_fd_sc_hd__nor3_1 U24144 ( .A(n17329), .B(n17328), .C(n17327), .Y(
        n17331) );
  sky130_fd_sc_hd__buf_2 U24145 ( .A(n23507), .X(n29439) );
  sky130_fd_sc_hd__xnor2_1 U24146 ( .A(j202_soc_core_j22_cpu_ml_bufa[22]), .B(
        j202_soc_core_j22_cpu_ml_bufa[21]), .Y(n17334) );
  sky130_fd_sc_hd__xnor2_1 U24147 ( .A(n18966), .B(n22087), .Y(n17345) );
  sky130_fd_sc_hd__xnor2_1 U24148 ( .A(n18994), .B(n22087), .Y(n17416) );
  sky130_fd_sc_hd__xor2_1 U24149 ( .A(j202_soc_core_j22_cpu_ml_bufa[23]), .B(
        n25627), .X(n17335) );
  sky130_fd_sc_hd__o22ai_1 U24150 ( .A1(n18474), .A2(n17345), .B1(n17416), 
        .B2(n18471), .Y(n17427) );
  sky130_fd_sc_hd__xnor2_1 U24151 ( .A(n18377), .B(n22023), .Y(n17336) );
  sky130_fd_sc_hd__xnor2_1 U24152 ( .A(j202_soc_core_j22_cpu_ml_bufa[20]), .B(
        j202_soc_core_j22_cpu_ml_bufa[19]), .Y(n17337) );
  sky130_fd_sc_hd__xnor2_1 U24153 ( .A(n22024), .B(n22299), .Y(n17365) );
  sky130_fd_sc_hd__xnor2_1 U24154 ( .A(n18925), .B(n22299), .Y(n17413) );
  sky130_fd_sc_hd__xor2_1 U24155 ( .A(j202_soc_core_j22_cpu_ml_bufa[20]), .B(
        j202_soc_core_j22_cpu_ml_bufa[21]), .X(n17338) );
  sky130_fd_sc_hd__o22ai_1 U24156 ( .A1(n18533), .A2(n17365), .B1(n17413), 
        .B2(n18530), .Y(n17402) );
  sky130_fd_sc_hd__xnor2_1 U24157 ( .A(j202_soc_core_j22_cpu_ml_bufa[26]), .B(
        j202_soc_core_j22_cpu_ml_bufa[25]), .Y(n17339) );
  sky130_fd_sc_hd__xnor2_1 U24158 ( .A(n18962), .B(n23571), .Y(n17372) );
  sky130_fd_sc_hd__xnor2_1 U24159 ( .A(n18999), .B(n23571), .Y(n17417) );
  sky130_fd_sc_hd__inv_1 U24160 ( .A(j202_soc_core_j22_cpu_ml_bufa[27]), .Y(
        n22526) );
  sky130_fd_sc_hd__o22ai_1 U24161 ( .A1(n18989), .A2(n17372), .B1(n17417), 
        .B2(n12044), .Y(n17421) );
  sky130_fd_sc_hd__xnor2_1 U24162 ( .A(j202_soc_core_j22_cpu_ml_bufa[30]), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .Y(n17341) );
  sky130_fd_sc_hd__xnor2_1 U24164 ( .A(n18367), .B(n25777), .Y(n17346) );
  sky130_fd_sc_hd__xnor2_1 U24165 ( .A(n18387), .B(n25777), .Y(n17414) );
  sky130_fd_sc_hd__xor2_1 U24166 ( .A(j202_soc_core_j22_cpu_ml_bufa[31]), .B(
        n12425), .X(n17342) );
  sky130_fd_sc_hd__nand2_4 U24167 ( .A(n17342), .B(n18993), .Y(n18990) );
  sky130_fd_sc_hd__o22ai_1 U24168 ( .A1(n18993), .A2(n17346), .B1(n17414), 
        .B2(n18990), .Y(n17420) );
  sky130_fd_sc_hd__xnor2_1 U24169 ( .A(j202_soc_core_j22_cpu_ml_bufa[28]), .B(
        j202_soc_core_j22_cpu_ml_bufa[27]), .Y(n17343) );
  sky130_fd_sc_hd__buf_4 U24170 ( .A(n17343), .X(n19023) );
  sky130_fd_sc_hd__xnor2_1 U24171 ( .A(n18964), .B(n25389), .Y(n17347) );
  sky130_fd_sc_hd__xnor2_1 U24172 ( .A(n18366), .B(n25389), .Y(n17418) );
  sky130_fd_sc_hd__buf_2 U24173 ( .A(j202_soc_core_j22_cpu_ml_bufa[28]), .X(
        n23582) );
  sky130_fd_sc_hd__xor2_1 U24174 ( .A(j202_soc_core_j22_cpu_ml_bufa[29]), .B(
        n23582), .X(n17344) );
  sky130_fd_sc_hd__nand2_4 U24175 ( .A(n17344), .B(n19023), .Y(n19020) );
  sky130_fd_sc_hd__o22ai_1 U24176 ( .A1(n19023), .A2(n17347), .B1(n17418), 
        .B2(n19020), .Y(n17419) );
  sky130_fd_sc_hd__xnor2_1 U24177 ( .A(n18925), .B(n22087), .Y(n17367) );
  sky130_fd_sc_hd__o22ai_1 U24178 ( .A1(n18474), .A2(n17367), .B1(n17345), 
        .B2(n18471), .Y(n17363) );
  sky130_fd_sc_hd__xnor2_1 U24179 ( .A(n18366), .B(n25777), .Y(n17371) );
  sky130_fd_sc_hd__o22ai_1 U24180 ( .A1(n18993), .A2(n17371), .B1(n17346), 
        .B2(n18990), .Y(n17362) );
  sky130_fd_sc_hd__xnor2_1 U24181 ( .A(n18999), .B(n25389), .Y(n17370) );
  sky130_fd_sc_hd__o22ai_1 U24182 ( .A1(n19023), .A2(n17370), .B1(n17347), 
        .B2(n19020), .Y(n17361) );
  sky130_fd_sc_hd__o21ai_1 U24183 ( .A1(n28435), .A2(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[4]), .B1(n24674), .Y(n17349) );
  sky130_fd_sc_hd__nor2_1 U24184 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .B(j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]), .Y(n17348) );
  sky130_fd_sc_hd__nand2_1 U24185 ( .A(n17349), .B(n17348), .Y(n17354) );
  sky130_fd_sc_hd__nand4_1 U24186 ( .A(n17351), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]), .C(n24674), .D(n17350), .Y(
        n17353) );
  sky130_fd_sc_hd__nand2_1 U24187 ( .A(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[4]), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]), .Y(n17352) );
  sky130_fd_sc_hd__nand2_1 U24188 ( .A(n23492), .B(n17355), .Y(n17964) );
  sky130_fd_sc_hd__nand3_2 U24189 ( .A(n17357), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[0]), .C(n18831), .Y(n22845) );
  sky130_fd_sc_hd__nand3_1 U24190 ( .A(n18834), .B(n17359), .C(n22845), .Y(
        n17358) );
  sky130_fd_sc_hd__nand2_4 U24191 ( .A(n17965), .B(n11478), .Y(n24854) );
  sky130_fd_sc_hd__a21oi_1 U24192 ( .A1(j202_soc_core_j22_cpu_ml_mach[22]), 
        .A2(n25679), .B1(n13087), .Y(n17360) );
  sky130_fd_sc_hd__o21ai_1 U24193 ( .A1(n22112), .A2(n11145), .B1(n17360), .Y(
        n17386) );
  sky130_fd_sc_hd__xnor2_1 U24194 ( .A(n18387), .B(n22023), .Y(n17364) );
  sky130_fd_sc_hd__xnor2_1 U24195 ( .A(n18971), .B(n23571), .Y(n17379) );
  sky130_fd_sc_hd__xnor2_1 U24196 ( .A(n18941), .B(n23571), .Y(n17373) );
  sky130_fd_sc_hd__o22ai_1 U24197 ( .A1(n18989), .A2(n17379), .B1(n17373), 
        .B2(n12044), .Y(n17391) );
  sky130_fd_sc_hd__xnor2_1 U24198 ( .A(n18367), .B(n22023), .Y(n17366) );
  sky130_fd_sc_hd__xnor2_1 U24199 ( .A(n22024), .B(n22087), .Y(n17383) );
  sky130_fd_sc_hd__o22ai_1 U24200 ( .A1(n18474), .A2(n17383), .B1(n17367), 
        .B2(n18471), .Y(n18958) );
  sky130_fd_sc_hd__xnor2_1 U24201 ( .A(j202_soc_core_j22_cpu_ml_bufa[24]), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .Y(n17368) );
  sky130_fd_sc_hd__buf_6 U24202 ( .A(j202_soc_core_j22_cpu_ml_bufa[25]), .X(
        n17635) );
  sky130_fd_sc_hd__buf_6 U24203 ( .A(n17635), .X(n23567) );
  sky130_fd_sc_hd__xnor2_1 U24204 ( .A(n18966), .B(n23567), .Y(n17381) );
  sky130_fd_sc_hd__xnor2_1 U24205 ( .A(n18994), .B(n23567), .Y(n17374) );
  sky130_fd_sc_hd__xor2_1 U24206 ( .A(n17635), .B(
        j202_soc_core_j22_cpu_ml_bufa[24]), .X(n17369) );
  sky130_fd_sc_hd__xnor2_1 U24207 ( .A(n18962), .B(n25389), .Y(n17387) );
  sky130_fd_sc_hd__o22ai_1 U24208 ( .A1(n19023), .A2(n17387), .B1(n17370), 
        .B2(n19020), .Y(n17377) );
  sky130_fd_sc_hd__xnor2_1 U24209 ( .A(n18964), .B(n25777), .Y(n17380) );
  sky130_fd_sc_hd__o22ai_1 U24210 ( .A1(n18993), .A2(n17380), .B1(n17371), 
        .B2(n18990), .Y(n17376) );
  sky130_fd_sc_hd__o22ai_1 U24211 ( .A1(n18989), .A2(n17373), .B1(n17372), 
        .B2(n12044), .Y(n17405) );
  sky130_fd_sc_hd__xnor2_1 U24212 ( .A(n18971), .B(n23567), .Y(n17406) );
  sky130_fd_sc_hd__a21oi_1 U24213 ( .A1(j202_soc_core_j22_cpu_ml_mach[21]), 
        .A2(n25679), .B1(n13087), .Y(n17375) );
  sky130_fd_sc_hd__fah_1 U24215 ( .A(n17378), .B(n17377), .CI(n17376), .COUT(
        n18980), .SUM(n17393) );
  sky130_fd_sc_hd__xnor2_1 U24216 ( .A(n18994), .B(n23571), .Y(n18967) );
  sky130_fd_sc_hd__o22ai_1 U24217 ( .A1(n18989), .A2(n18967), .B1(n17379), 
        .B2(n18986), .Y(n18961) );
  sky130_fd_sc_hd__xnor2_1 U24218 ( .A(n18999), .B(n25777), .Y(n18963) );
  sky130_fd_sc_hd__o22ai_1 U24219 ( .A1(n18993), .A2(n18963), .B1(n17380), 
        .B2(n18990), .Y(n18960) );
  sky130_fd_sc_hd__xnor2_1 U24220 ( .A(n18925), .B(n23567), .Y(n18973) );
  sky130_fd_sc_hd__xnor2_1 U24221 ( .A(n18366), .B(n22023), .Y(n17382) );
  sky130_fd_sc_hd__fah_1 U24222 ( .A(n17386), .B(n17385), .CI(n17384), .COUT(
        n18970), .SUM(n17398) );
  sky130_fd_sc_hd__xnor2_1 U24223 ( .A(n18941), .B(n25389), .Y(n18972) );
  sky130_fd_sc_hd__o22ai_1 U24224 ( .A1(n19023), .A2(n18972), .B1(n17387), 
        .B2(n19020), .Y(n18977) );
  sky130_fd_sc_hd__a21oi_1 U24225 ( .A1(j202_soc_core_j22_cpu_ml_mach[23]), 
        .A2(n25679), .B1(n13087), .Y(n17388) );
  sky130_fd_sc_hd__o21ai_1 U24226 ( .A1(n17488), .A2(n11145), .B1(n17388), .Y(
        n18976) );
  sky130_fd_sc_hd__fah_1 U24227 ( .A(n17391), .B(n17390), .CI(n17389), .COUT(
        n18975), .SUM(n17394) );
  sky130_fd_sc_hd__fah_1 U24228 ( .A(n17394), .B(n17393), .CI(n17392), .COUT(
        n18968), .SUM(n17397) );
  sky130_fd_sc_hd__xnor2_1 U24229 ( .A(n17395), .B(n19009), .Y(n17396) );
  sky130_fd_sc_hd__xor2_1 U24230 ( .A(n19011), .B(n17396), .X(n17441) );
  sky130_fd_sc_hd__fah_1 U24231 ( .A(n17397), .B(n17398), .CI(n17399), .COUT(
        n19011), .SUM(n18646) );
  sky130_fd_sc_hd__fa_1 U24232 ( .A(n17402), .B(n17401), .CIN(n17400), .COUT(
        n17384), .SUM(n18459) );
  sky130_fd_sc_hd__fah_1 U24233 ( .A(n17405), .B(n17404), .CI(n17403), .COUT(
        n17392), .SUM(n18458) );
  sky130_fd_sc_hd__xnor2_1 U24234 ( .A(n18941), .B(n23567), .Y(n17415) );
  sky130_fd_sc_hd__a21oi_1 U24235 ( .A1(j202_soc_core_j22_cpu_ml_mach[20]), 
        .A2(n22940), .B1(n13087), .Y(n17407) );
  sky130_fd_sc_hd__o21ai_1 U24236 ( .A1(n17720), .A2(n11145), .B1(n17407), .Y(
        n17435) );
  sky130_fd_sc_hd__xnor2_1 U24237 ( .A(n22024), .B(n22811), .Y(n17412) );
  sky130_fd_sc_hd__xnor2_1 U24238 ( .A(n18925), .B(n22811), .Y(n18341) );
  sky130_fd_sc_hd__xnor2_1 U24239 ( .A(n17408), .B(
        j202_soc_core_j22_cpu_ml_bufa[19]), .Y(n17409) );
  sky130_fd_sc_hd__xnor2_1 U24241 ( .A(n18371), .B(n22023), .Y(n17411) );
  sky130_fd_sc_hd__a21o_1 U24242 ( .A1(n17410), .A2(n18496), .B1(n17412), .X(
        n18414) );
  sky130_fd_sc_hd__xnor2_1 U24243 ( .A(n18966), .B(n22299), .Y(n17431) );
  sky130_fd_sc_hd__o22ai_1 U24244 ( .A1(n18533), .A2(n17413), .B1(n17431), 
        .B2(n18530), .Y(n18419) );
  sky130_fd_sc_hd__xnor2_1 U24245 ( .A(n18377), .B(n25777), .Y(n17432) );
  sky130_fd_sc_hd__o22ai_1 U24246 ( .A1(n18993), .A2(n17414), .B1(n17432), 
        .B2(n18990), .Y(n18418) );
  sky130_fd_sc_hd__xnor2_1 U24247 ( .A(n18962), .B(n23567), .Y(n17433) );
  sky130_fd_sc_hd__xnor2_1 U24248 ( .A(n18971), .B(n22087), .Y(n17429) );
  sky130_fd_sc_hd__xnor2_1 U24250 ( .A(n18964), .B(n23571), .Y(n18402) );
  sky130_fd_sc_hd__o22ai_1 U24251 ( .A1(n18989), .A2(n17417), .B1(n18402), 
        .B2(n12044), .Y(n18412) );
  sky130_fd_sc_hd__xnor2_1 U24252 ( .A(n18367), .B(n25389), .Y(n18404) );
  sky130_fd_sc_hd__o22ai_1 U24253 ( .A1(n19023), .A2(n17418), .B1(n18404), 
        .B2(n19020), .Y(n18411) );
  sky130_fd_sc_hd__fah_1 U24254 ( .A(n17421), .B(n17420), .CI(n17419), .COUT(
        n17423), .SUM(n18437) );
  sky130_fd_sc_hd__fah_1 U24255 ( .A(n17424), .B(n17423), .CI(n17422), .COUT(
        n17399), .SUM(n18453) );
  sky130_fd_sc_hd__fah_1 U24256 ( .A(n17427), .B(n17426), .CI(n17425), .COUT(
        n17424), .SUM(n18447) );
  sky130_fd_sc_hd__a21oi_1 U24257 ( .A1(j202_soc_core_j22_cpu_ml_mach[19]), 
        .A2(n22940), .B1(n13087), .Y(n17428) );
  sky130_fd_sc_hd__o21ai_1 U24258 ( .A1(n17710), .A2(n11145), .B1(n17428), .Y(
        n18391) );
  sky130_fd_sc_hd__xnor2_1 U24259 ( .A(n18941), .B(n22087), .Y(n18356) );
  sky130_fd_sc_hd__xnor2_1 U24260 ( .A(n18372), .B(n22023), .Y(n17430) );
  sky130_fd_sc_hd__xnor2_1 U24261 ( .A(n18994), .B(n22299), .Y(n18384) );
  sky130_fd_sc_hd__o22ai_1 U24262 ( .A1(n18533), .A2(n17431), .B1(n18384), 
        .B2(n18530), .Y(n18353) );
  sky130_fd_sc_hd__xnor2_1 U24263 ( .A(n18371), .B(
        j202_soc_core_j22_cpu_ml_bufa[31]), .Y(n18342) );
  sky130_fd_sc_hd__o22ai_1 U24264 ( .A1(n18993), .A2(n17432), .B1(n18342), 
        .B2(n18990), .Y(n18352) );
  sky130_fd_sc_hd__xnor2_1 U24265 ( .A(n18999), .B(n23567), .Y(n18386) );
  sky130_fd_sc_hd__fah_1 U24266 ( .A(n17436), .B(n17435), .CI(n17434), .COUT(
        n18457), .SUM(n18445) );
  sky130_fd_sc_hd__o21ai_1 U24267 ( .A1(n18646), .A2(n18647), .B1(n13059), .Y(
        n17439) );
  sky130_fd_sc_hd__nand2_1 U24268 ( .A(n18646), .B(n18647), .Y(n17438) );
  sky130_fd_sc_hd__nand2_1 U24269 ( .A(n17439), .B(n17438), .Y(n17442) );
  sky130_fd_sc_hd__nor2_1 U24270 ( .A(n17441), .B(n17442), .Y(n17440) );
  sky130_fd_sc_hd__nand2_1 U24271 ( .A(n17442), .B(n17441), .Y(n19059) );
  sky130_fd_sc_hd__nand2_1 U24272 ( .A(n19061), .B(n19059), .Y(n18677) );
  sky130_fd_sc_hd__xnor2_1 U24273 ( .A(j202_soc_core_j22_cpu_ml_bufa[16]), .B(
        j202_soc_core_j22_cpu_ml_bufa[15]), .Y(n17443) );
  sky130_fd_sc_hd__xnor2_1 U24274 ( .A(n18999), .B(n25761), .Y(n17536) );
  sky130_fd_sc_hd__xnor2_1 U24275 ( .A(n18964), .B(n25761), .Y(n17445) );
  sky130_fd_sc_hd__xor2_1 U24276 ( .A(j202_soc_core_j22_cpu_ml_bufa[17]), .B(
        n24829), .X(n17444) );
  sky130_fd_sc_hd__o22ai_1 U24277 ( .A1(n18486), .A2(n17536), .B1(n17445), 
        .B2(n18483), .Y(n17568) );
  sky130_fd_sc_hd__nor2b_1 U24278 ( .B_N(n18470), .A(n19002), .Y(n17523) );
  sky130_fd_sc_hd__xnor2_1 U24279 ( .A(n18366), .B(n25761), .Y(n17447) );
  sky130_fd_sc_hd__o22ai_1 U24280 ( .A1(n18486), .A2(n17445), .B1(n17447), 
        .B2(n18483), .Y(n17522) );
  sky130_fd_sc_hd__o22ai_1 U24281 ( .A1(n24854), .A2(n18982), .B1(n22889), 
        .B2(n18224), .Y(n17566) );
  sky130_fd_sc_hd__xnor2_1 U24282 ( .A(n18367), .B(n25761), .Y(n17478) );
  sky130_fd_sc_hd__xnor2_1 U24283 ( .A(n18363), .B(n22087), .Y(n17466) );
  sky130_fd_sc_hd__xnor2_1 U24284 ( .A(n22087), .B(n18470), .Y(n17448) );
  sky130_fd_sc_hd__o22ai_1 U24285 ( .A1(n18474), .A2(n17466), .B1(n17448), 
        .B2(n18471), .Y(n17476) );
  sky130_fd_sc_hd__inv_2 U24286 ( .A(j202_soc_core_j22_cpu_ml_bufa[6]), .Y(
        n17449) );
  sky130_fd_sc_hd__xnor2_1 U24287 ( .A(n17449), .B(
        j202_soc_core_j22_cpu_ml_bufa[7]), .Y(n17450) );
  sky130_fd_sc_hd__buf_4 U24288 ( .A(n30022), .X(n18192) );
  sky130_fd_sc_hd__xnor2_1 U24289 ( .A(n22024), .B(n27618), .Y(n17508) );
  sky130_fd_sc_hd__buf_6 U24290 ( .A(n11350), .X(n24345) );
  sky130_fd_sc_hd__xnor2_1 U24291 ( .A(n18941), .B(n24345), .Y(n17467) );
  sky130_fd_sc_hd__xnor2_1 U24292 ( .A(n18962), .B(n24345), .Y(n17504) );
  sky130_fd_sc_hd__o22ai_1 U24293 ( .A1(n18027), .A2(n17467), .B1(n17504), 
        .B2(n11119), .Y(n17511) );
  sky130_fd_sc_hd__nand2b_1 U24294 ( .A_N(n18470), .B(n22087), .Y(n17456) );
  sky130_fd_sc_hd__o22ai_1 U24295 ( .A1(n18474), .A2(n17456), .B1(n17455), 
        .B2(n18471), .Y(n17510) );
  sky130_fd_sc_hd__xnor2_1 U24296 ( .A(j202_soc_core_j22_cpu_ml_bufa[14]), .B(
        j202_soc_core_j22_cpu_ml_bufa[13]), .Y(n17457) );
  sky130_fd_sc_hd__buf_4 U24297 ( .A(n17457), .X(n18492) );
  sky130_fd_sc_hd__xnor2_1 U24298 ( .A(n18999), .B(n18887), .Y(n17468) );
  sky130_fd_sc_hd__xnor2_1 U24299 ( .A(n18964), .B(n18887), .Y(n17506) );
  sky130_fd_sc_hd__xnor2_1 U24300 ( .A(n11417), .B(n24454), .Y(n17458) );
  sky130_fd_sc_hd__nand2b_4 U24301 ( .A_N(n17458), .B(n18492), .Y(n18489) );
  sky130_fd_sc_hd__o22ai_1 U24302 ( .A1(n18492), .A2(n17468), .B1(n17506), 
        .B2(n18489), .Y(n17509) );
  sky130_fd_sc_hd__xnor2_1 U24303 ( .A(n18387), .B(n22811), .Y(n17463) );
  sky130_fd_sc_hd__xnor2_1 U24304 ( .A(n18377), .B(n22811), .Y(n17498) );
  sky130_fd_sc_hd__o22ai_1 U24305 ( .A1(n18496), .A2(n17463), .B1(n17498), 
        .B2(n17410), .Y(n17474) );
  sky130_fd_sc_hd__xnor2_2 U24306 ( .A(j202_soc_core_j22_cpu_ml_bufa[10]), .B(
        n12050), .Y(n17460) );
  sky130_fd_sc_hd__buf_4 U24308 ( .A(j202_soc_core_j22_cpu_ml_bufa[11]), .X(
        n21280) );
  sky130_fd_sc_hd__xnor2_1 U24309 ( .A(n18994), .B(n21280), .Y(n17464) );
  sky130_fd_sc_hd__xnor2_1 U24310 ( .A(n18971), .B(n21280), .Y(n17502) );
  sky130_fd_sc_hd__xor2_1 U24311 ( .A(j202_soc_core_j22_cpu_ml_bufa[11]), .B(
        j202_soc_core_j22_cpu_ml_bufa[10]), .X(n17459) );
  sky130_fd_sc_hd__o22ai_1 U24313 ( .A1(n18079), .A2(n17464), .B1(n17502), 
        .B2(n18036), .Y(n17473) );
  sky130_fd_sc_hd__xnor2_1 U24314 ( .A(j202_soc_core_j22_cpu_ml_bufa[8]), .B(
        j202_soc_core_j22_cpu_ml_bufa[7]), .Y(n17461) );
  sky130_fd_sc_hd__buf_6 U24315 ( .A(n12050), .X(n24799) );
  sky130_fd_sc_hd__xnor2_1 U24316 ( .A(n18925), .B(n24799), .Y(n17465) );
  sky130_fd_sc_hd__xnor2_1 U24317 ( .A(n18966), .B(n24799), .Y(n17500) );
  sky130_fd_sc_hd__xor2_1 U24318 ( .A(n12050), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n17462) );
  sky130_fd_sc_hd__xnor2_1 U24319 ( .A(n18367), .B(n22811), .Y(n17517) );
  sky130_fd_sc_hd__o22ai_1 U24320 ( .A1(n18496), .A2(n17517), .B1(n17463), 
        .B2(n17410), .Y(n17484) );
  sky130_fd_sc_hd__xnor2_1 U24321 ( .A(n18966), .B(n21280), .Y(n17516) );
  sky130_fd_sc_hd__o22ai_1 U24322 ( .A1(n18079), .A2(n17516), .B1(n17464), 
        .B2(n18036), .Y(n17483) );
  sky130_fd_sc_hd__xnor2_1 U24323 ( .A(n22024), .B(n24799), .Y(n17519) );
  sky130_fd_sc_hd__xnor2_1 U24324 ( .A(n18372), .B(n22087), .Y(n17469) );
  sky130_fd_sc_hd__o22ai_1 U24325 ( .A1(n18474), .A2(n17469), .B1(n17466), 
        .B2(n18471), .Y(n17481) );
  sky130_fd_sc_hd__xnor2_1 U24326 ( .A(n18971), .B(n24345), .Y(n17470) );
  sky130_fd_sc_hd__o22ai_1 U24327 ( .A1(n18027), .A2(n17470), .B1(n17467), 
        .B2(n11119), .Y(n17480) );
  sky130_fd_sc_hd__xnor2_1 U24328 ( .A(n18962), .B(n18887), .Y(n17471) );
  sky130_fd_sc_hd__o22ai_1 U24329 ( .A1(n18492), .A2(n17471), .B1(n17468), 
        .B2(n18489), .Y(n17479) );
  sky130_fd_sc_hd__xnor2_1 U24330 ( .A(n18371), .B(n22087), .Y(n17561) );
  sky130_fd_sc_hd__o22ai_1 U24331 ( .A1(n18474), .A2(n17561), .B1(n17469), 
        .B2(n18471), .Y(n17546) );
  sky130_fd_sc_hd__xnor2_1 U24332 ( .A(n18994), .B(n24345), .Y(n17560) );
  sky130_fd_sc_hd__o22ai_1 U24333 ( .A1(n18027), .A2(n17560), .B1(n17470), 
        .B2(n11119), .Y(n17545) );
  sky130_fd_sc_hd__xnor2_1 U24334 ( .A(n18941), .B(n18887), .Y(n17562) );
  sky130_fd_sc_hd__o22ai_1 U24335 ( .A1(n18492), .A2(n17562), .B1(n17471), 
        .B2(n18489), .Y(n17544) );
  sky130_fd_sc_hd__xnor2_1 U24337 ( .A(n18372), .B(n22299), .Y(n17485) );
  sky130_fd_sc_hd__xnor2_1 U24338 ( .A(n18363), .B(n22299), .Y(n17493) );
  sky130_fd_sc_hd__o22ai_1 U24339 ( .A1(n18533), .A2(n17485), .B1(n17493), 
        .B2(n18530), .Y(n17691) );
  sky130_fd_sc_hd__xnor2_1 U24340 ( .A(n18387), .B(n25761), .Y(n17496) );
  sky130_fd_sc_hd__xnor2_1 U24341 ( .A(n17487), .B(n17486), .Y(n17690) );
  sky130_fd_sc_hd__fah_1 U24342 ( .A(n17484), .B(n17483), .CI(n17482), .COUT(
        n17540), .SUM(n17513) );
  sky130_fd_sc_hd__xnor2_1 U24343 ( .A(n18371), .B(n22299), .Y(n17520) );
  sky130_fd_sc_hd__o22ai_1 U24344 ( .A1(n18533), .A2(n17520), .B1(n17485), 
        .B2(n18530), .Y(n17491) );
  sky130_fd_sc_hd__o22ai_1 U24345 ( .A1(n24854), .A2(n17488), .B1(n22081), 
        .B2(n18536), .Y(n17489) );
  sky130_fd_sc_hd__fah_1 U24346 ( .A(n17491), .B(n17490), .CI(n17489), .COUT(
        n17512), .SUM(n17815) );
  sky130_fd_sc_hd__xnor2_1 U24347 ( .A(n18371), .B(n22811), .Y(n17497) );
  sky130_fd_sc_hd__xnor2_1 U24348 ( .A(n18372), .B(n22811), .Y(n17695) );
  sky130_fd_sc_hd__o22ai_1 U24349 ( .A1(n18496), .A2(n17497), .B1(n17695), 
        .B2(n17410), .Y(n17716) );
  sky130_fd_sc_hd__buf_2 U24350 ( .A(j202_soc_core_j22_cpu_ml_bufb[0]), .X(
        n18210) );
  sky130_fd_sc_hd__xnor2_1 U24351 ( .A(n22299), .B(n18210), .Y(n17492) );
  sky130_fd_sc_hd__o22ai_1 U24352 ( .A1(n18533), .A2(n17493), .B1(n17492), 
        .B2(n18530), .Y(n17715) );
  sky130_fd_sc_hd__xor2_1 U24353 ( .A(j202_soc_core_j22_cpu_ml_bufa[5]), .B(
        j202_soc_core_j22_cpu_ml_bufa[4]), .X(n17494) );
  sky130_fd_sc_hd__xnor2_1 U24354 ( .A(j202_soc_core_j22_cpu_ml_bufa[4]), .B(
        j202_soc_core_j22_cpu_ml_bufa[3]), .Y(n17495) );
  sky130_fd_sc_hd__buf_4 U24355 ( .A(n17495), .X(n18205) );
  sky130_fd_sc_hd__xnor2_1 U24356 ( .A(n22024), .B(n24366), .Y(n17718) );
  sky130_fd_sc_hd__xnor2_1 U24357 ( .A(n18999), .B(n24345), .Y(n17503) );
  sky130_fd_sc_hd__xnor2_1 U24358 ( .A(n18964), .B(n24345), .Y(n17719) );
  sky130_fd_sc_hd__o22ai_1 U24359 ( .A1(n18027), .A2(n17503), .B1(n17719), 
        .B2(n11119), .Y(n17700) );
  sky130_fd_sc_hd__xnor2_1 U24360 ( .A(n18366), .B(n18887), .Y(n17505) );
  sky130_fd_sc_hd__xnor2_1 U24361 ( .A(n18367), .B(n18887), .Y(n17696) );
  sky130_fd_sc_hd__o22ai_1 U24362 ( .A1(n18492), .A2(n17505), .B1(n17696), 
        .B2(n18489), .Y(n17699) );
  sky130_fd_sc_hd__xnor2_1 U24363 ( .A(n18925), .B(n27618), .Y(n17507) );
  sky130_fd_sc_hd__xnor2_1 U24364 ( .A(n18966), .B(n27618), .Y(n17693) );
  sky130_fd_sc_hd__o22ai_1 U24365 ( .A1(n18192), .A2(n17507), .B1(n17693), 
        .B2(n18189), .Y(n17698) );
  sky130_fd_sc_hd__xnor2_1 U24366 ( .A(n18377), .B(n25761), .Y(n17692) );
  sky130_fd_sc_hd__o22ai_1 U24367 ( .A1(n18486), .A2(n17496), .B1(n17692), 
        .B2(n18483), .Y(n17713) );
  sky130_fd_sc_hd__xnor2_1 U24368 ( .A(n18941), .B(n21280), .Y(n17501) );
  sky130_fd_sc_hd__xnor2_1 U24369 ( .A(n18962), .B(n21280), .Y(n17697) );
  sky130_fd_sc_hd__o22ai_1 U24370 ( .A1(n18079), .A2(n17501), .B1(n17697), 
        .B2(n18036), .Y(n17712) );
  sky130_fd_sc_hd__xnor2_1 U24371 ( .A(n18994), .B(n24799), .Y(n17499) );
  sky130_fd_sc_hd__xnor2_1 U24372 ( .A(n18971), .B(n24799), .Y(n17694) );
  sky130_fd_sc_hd__o22ai_1 U24373 ( .A1(n18496), .A2(n17498), .B1(n17497), 
        .B2(n17410), .Y(n17757) );
  sky130_fd_sc_hd__o22ai_1 U24374 ( .A1(n18079), .A2(n17502), .B1(n17501), 
        .B2(n18036), .Y(n17755) );
  sky130_fd_sc_hd__o22ai_1 U24375 ( .A1(n18027), .A2(n17504), .B1(n17503), 
        .B2(n11119), .Y(n17754) );
  sky130_fd_sc_hd__o22ai_1 U24376 ( .A1(n18492), .A2(n17506), .B1(n17505), 
        .B2(n18489), .Y(n17753) );
  sky130_fd_sc_hd__o22ai_1 U24377 ( .A1(n18192), .A2(n17508), .B1(n17507), 
        .B2(n18189), .Y(n17752) );
  sky130_fd_sc_hd__fah_1 U24379 ( .A(n17514), .B(n17513), .CI(n17512), .COUT(
        n17553), .SUM(n17845) );
  sky130_fd_sc_hd__xnor2_1 U24380 ( .A(n18387), .B(n22299), .Y(n17563) );
  sky130_fd_sc_hd__xnor2_1 U24381 ( .A(n18377), .B(n22299), .Y(n17521) );
  sky130_fd_sc_hd__o22ai_1 U24382 ( .A1(n18533), .A2(n17563), .B1(n17521), 
        .B2(n18530), .Y(n17549) );
  sky130_fd_sc_hd__nand2b_1 U24383 ( .A_N(n18470), .B(n23567), .Y(n17515) );
  sky130_fd_sc_hd__xnor2_1 U24384 ( .A(n18925), .B(n21280), .Y(n17565) );
  sky130_fd_sc_hd__o22ai_1 U24385 ( .A1(n18079), .A2(n17565), .B1(n17516), 
        .B2(n18036), .Y(n17547) );
  sky130_fd_sc_hd__xnor2_1 U24386 ( .A(n18366), .B(n22811), .Y(n17537) );
  sky130_fd_sc_hd__o22ai_1 U24387 ( .A1(n18496), .A2(n17537), .B1(n17517), 
        .B2(n17410), .Y(n17543) );
  sky130_fd_sc_hd__xnor2_1 U24388 ( .A(n18363), .B(n23567), .Y(n17564) );
  sky130_fd_sc_hd__xnor2_1 U24389 ( .A(n23567), .B(n18210), .Y(n17518) );
  sky130_fd_sc_hd__o22ai_1 U24390 ( .A1(n18533), .A2(n17521), .B1(n17520), 
        .B2(n18530), .Y(n17526) );
  sky130_fd_sc_hd__xnor2_1 U24391 ( .A(n17523), .B(n17522), .Y(n17525) );
  sky130_fd_sc_hd__xnor2_1 U24392 ( .A(n17553), .B(n17554), .Y(n17533) );
  sky130_fd_sc_hd__o21ai_1 U24394 ( .A1(n17850), .A2(n17854), .B1(n17851), .Y(
        n17535) );
  sky130_fd_sc_hd__nand2_1 U24395 ( .A(n17854), .B(n17850), .Y(n17534) );
  sky130_fd_sc_hd__nand2_1 U24396 ( .A(n17535), .B(n17534), .Y(n17859) );
  sky130_fd_sc_hd__xnor2_1 U24397 ( .A(n18962), .B(n25761), .Y(n17588) );
  sky130_fd_sc_hd__o22ai_1 U24398 ( .A1(n18486), .A2(n17588), .B1(n17536), 
        .B2(n18483), .Y(n17600) );
  sky130_fd_sc_hd__nor2b_1 U24399 ( .B_N(n18470), .A(n18989), .Y(n17577) );
  sky130_fd_sc_hd__xnor2_1 U24400 ( .A(n18964), .B(n22811), .Y(n17575) );
  sky130_fd_sc_hd__o22ai_1 U24401 ( .A1(n18496), .A2(n17575), .B1(n17537), 
        .B2(n17410), .Y(n17576) );
  sky130_fd_sc_hd__xnor2_1 U24402 ( .A(n17577), .B(n17576), .Y(n17599) );
  sky130_fd_sc_hd__inv_2 U24403 ( .A(n24854), .Y(n25679) );
  sky130_fd_sc_hd__fah_1 U24404 ( .A(n17540), .B(n17539), .CI(n17538), .COUT(
        n17602), .SUM(n17569) );
  sky130_fd_sc_hd__fah_1 U24405 ( .A(n17543), .B(n17542), .CI(n17541), .COUT(
        n17580), .SUM(n17558) );
  sky130_fd_sc_hd__nand2b_1 U24407 ( .A_N(n17554), .B(n17550), .Y(n17551) );
  sky130_fd_sc_hd__nand2_1 U24408 ( .A(n17552), .B(n17551), .Y(n17556) );
  sky130_fd_sc_hd__nand2_1 U24409 ( .A(n17554), .B(n17553), .Y(n17555) );
  sky130_fd_sc_hd__nand2_1 U24410 ( .A(n17556), .B(n17555), .Y(n17573) );
  sky130_fd_sc_hd__fah_1 U24411 ( .A(n17559), .B(n17558), .CI(n17557), .COUT(
        n17607), .SUM(n17554) );
  sky130_fd_sc_hd__xnor2_1 U24412 ( .A(n18966), .B(n24345), .Y(n17592) );
  sky130_fd_sc_hd__o22ai_1 U24413 ( .A1(n18027), .A2(n17592), .B1(n17560), 
        .B2(n11119), .Y(n17585) );
  sky130_fd_sc_hd__xnor2_1 U24414 ( .A(n18377), .B(n22087), .Y(n17586) );
  sky130_fd_sc_hd__xnor2_1 U24416 ( .A(n18971), .B(n18887), .Y(n17594) );
  sky130_fd_sc_hd__o22ai_1 U24417 ( .A1(n18492), .A2(n17594), .B1(n17562), 
        .B2(n18489), .Y(n17583) );
  sky130_fd_sc_hd__xnor2_1 U24418 ( .A(n18367), .B(n22299), .Y(n17595) );
  sky130_fd_sc_hd__o22ai_1 U24419 ( .A1(n18533), .A2(n17595), .B1(n17563), 
        .B2(n18530), .Y(n17582) );
  sky130_fd_sc_hd__xnor2_1 U24420 ( .A(n18372), .B(n23567), .Y(n17593) );
  sky130_fd_sc_hd__xnor2_1 U24421 ( .A(n22024), .B(n21280), .Y(n17597) );
  sky130_fd_sc_hd__o22ai_1 U24422 ( .A1(n18079), .A2(n17597), .B1(n17565), 
        .B2(n18036), .Y(n17581) );
  sky130_fd_sc_hd__fah_1 U24423 ( .A(n17571), .B(n17570), .CI(n17569), .COUT(
        n17605), .SUM(n17850) );
  sky130_fd_sc_hd__nor2_1 U24424 ( .A(n17859), .B(n17860), .Y(n19303) );
  sky130_fd_sc_hd__xnor2_1 U24425 ( .A(n18999), .B(n22811), .Y(n17619) );
  sky130_fd_sc_hd__o22ai_1 U24426 ( .A1(n18496), .A2(n17619), .B1(n17575), 
        .B2(n17410), .Y(n17638) );
  sky130_fd_sc_hd__fah_1 U24427 ( .A(n17580), .B(n17579), .CI(n17578), .COUT(
        n17640), .SUM(n17601) );
  sky130_fd_sc_hd__xnor2_1 U24429 ( .A(n18387), .B(n22087), .Y(n17633) );
  sky130_fd_sc_hd__nand2b_1 U24430 ( .A_N(n18470), .B(n23571), .Y(n17587) );
  sky130_fd_sc_hd__o22ai_1 U24431 ( .A1(n18989), .A2(n17587), .B1(n22526), 
        .B2(n12044), .Y(n17612) );
  sky130_fd_sc_hd__xnor2_1 U24432 ( .A(n18941), .B(n25761), .Y(n17632) );
  sky130_fd_sc_hd__o22ai_1 U24433 ( .A1(n18486), .A2(n17632), .B1(n17588), 
        .B2(n18483), .Y(n17611) );
  sky130_fd_sc_hd__fah_1 U24434 ( .A(n17591), .B(n17590), .CI(n17589), .COUT(
        n17623), .SUM(n17606) );
  sky130_fd_sc_hd__xnor2_1 U24435 ( .A(n18925), .B(n24345), .Y(n17620) );
  sky130_fd_sc_hd__o22ai_1 U24436 ( .A1(n18027), .A2(n17620), .B1(n17592), 
        .B2(n11119), .Y(n17615) );
  sky130_fd_sc_hd__xnor2_1 U24437 ( .A(n18371), .B(n17635), .Y(n17636) );
  sky130_fd_sc_hd__xnor2_1 U24438 ( .A(n18994), .B(n18887), .Y(n17634) );
  sky130_fd_sc_hd__o22ai_1 U24439 ( .A1(n18492), .A2(n17634), .B1(n17594), 
        .B2(n18489), .Y(n17613) );
  sky130_fd_sc_hd__xnor2_1 U24440 ( .A(n18366), .B(n22299), .Y(n17630) );
  sky130_fd_sc_hd__xnor2_1 U24441 ( .A(n18363), .B(n23571), .Y(n17631) );
  sky130_fd_sc_hd__xnor2_1 U24442 ( .A(n23571), .B(n18470), .Y(n17596) );
  sky130_fd_sc_hd__o22ai_1 U24443 ( .A1(n18989), .A2(n17631), .B1(n17596), 
        .B2(n18986), .Y(n17609) );
  sky130_fd_sc_hd__a21o_1 U24444 ( .A1(n18036), .A2(n18079), .B1(n17597), .X(
        n17608) );
  sky130_fd_sc_hd__xnor2_1 U24445 ( .A(n17623), .B(n17624), .Y(n17604) );
  sky130_fd_sc_hd__fah_1 U24446 ( .A(n17603), .B(n17602), .CI(n17601), .COUT(
        n17622), .SUM(n17574) );
  sky130_fd_sc_hd__xnor2_1 U24447 ( .A(n17604), .B(n17622), .Y(n17684) );
  sky130_fd_sc_hd__fa_1 U24448 ( .A(n17610), .B(n17609), .CIN(n17608), .COUT(
        n17654), .SUM(n17628) );
  sky130_fd_sc_hd__fa_1 U24449 ( .A(n17615), .B(n17614), .CIN(n17613), .COUT(
        n17652), .SUM(n17629) );
  sky130_fd_sc_hd__fah_1 U24450 ( .A(n17618), .B(n17617), .CI(n17616), .COUT(
        n17666), .SUM(n17639) );
  sky130_fd_sc_hd__xnor2_1 U24451 ( .A(n18962), .B(n22811), .Y(n17651) );
  sky130_fd_sc_hd__o22ai_1 U24452 ( .A1(n18496), .A2(n17651), .B1(n17619), 
        .B2(n17410), .Y(n17681) );
  sky130_fd_sc_hd__nor2b_1 U24453 ( .B_N(n18470), .A(n19023), .Y(n17657) );
  sky130_fd_sc_hd__xnor2_1 U24454 ( .A(n22024), .B(n24345), .Y(n17678) );
  sky130_fd_sc_hd__o22ai_1 U24455 ( .A1(n18027), .A2(n17678), .B1(n17620), 
        .B2(n11119), .Y(n17656) );
  sky130_fd_sc_hd__xnor2_1 U24456 ( .A(n17657), .B(n17656), .Y(n17680) );
  sky130_fd_sc_hd__xnor2_1 U24457 ( .A(n17666), .B(n17665), .Y(n17621) );
  sky130_fd_sc_hd__xnor2_1 U24458 ( .A(n17664), .B(n17621), .Y(n17688) );
  sky130_fd_sc_hd__nand2_1 U24460 ( .A(n17624), .B(n17623), .Y(n17625) );
  sky130_fd_sc_hd__nand2_1 U24461 ( .A(n17626), .B(n17625), .Y(n17687) );
  sky130_fd_sc_hd__fah_1 U24462 ( .A(n17629), .B(n17628), .CI(n17627), .COUT(
        n17661), .SUM(n17624) );
  sky130_fd_sc_hd__xnor2_1 U24463 ( .A(n18964), .B(n22299), .Y(n17655) );
  sky130_fd_sc_hd__o22ai_1 U24464 ( .A1(n18533), .A2(n17655), .B1(n17630), 
        .B2(n18530), .Y(n17648) );
  sky130_fd_sc_hd__xnor2_1 U24465 ( .A(n18372), .B(n23571), .Y(n17650) );
  sky130_fd_sc_hd__o22ai_1 U24466 ( .A1(n18989), .A2(n17650), .B1(n17631), 
        .B2(n12044), .Y(n17647) );
  sky130_fd_sc_hd__xnor2_1 U24467 ( .A(n18971), .B(n25761), .Y(n17672) );
  sky130_fd_sc_hd__o22ai_1 U24468 ( .A1(n18486), .A2(n17672), .B1(n17632), 
        .B2(n18483), .Y(n17646) );
  sky130_fd_sc_hd__xnor2_1 U24469 ( .A(n18367), .B(n22087), .Y(n17676) );
  sky130_fd_sc_hd__o22ai_1 U24470 ( .A1(n18474), .A2(n17676), .B1(n17633), 
        .B2(n18471), .Y(n17645) );
  sky130_fd_sc_hd__xnor2_1 U24471 ( .A(n18966), .B(n18887), .Y(n17649) );
  sky130_fd_sc_hd__o22ai_1 U24472 ( .A1(n18492), .A2(n17649), .B1(n17634), 
        .B2(n18489), .Y(n17644) );
  sky130_fd_sc_hd__xnor2_1 U24473 ( .A(n18377), .B(n17635), .Y(n17675) );
  sky130_fd_sc_hd__xnor2_1 U24474 ( .A(n17661), .B(n17662), .Y(n17642) );
  sky130_fd_sc_hd__xnor2_1 U24475 ( .A(n17642), .B(n17660), .Y(n17686) );
  sky130_fd_sc_hd__xnor2_1 U24476 ( .A(n18925), .B(n18887), .Y(n18490) );
  sky130_fd_sc_hd__o22ai_1 U24477 ( .A1(n18492), .A2(n18490), .B1(n17649), 
        .B2(n18489), .Y(n18551) );
  sky130_fd_sc_hd__xnor2_1 U24478 ( .A(n18371), .B(n23571), .Y(n18497) );
  sky130_fd_sc_hd__o22ai_1 U24479 ( .A1(n18989), .A2(n18497), .B1(n17650), 
        .B2(n12044), .Y(n18550) );
  sky130_fd_sc_hd__xnor2_1 U24480 ( .A(n18941), .B(n22811), .Y(n18494) );
  sky130_fd_sc_hd__o22ai_1 U24481 ( .A1(n18496), .A2(n18494), .B1(n17651), 
        .B2(n17410), .Y(n18549) );
  sky130_fd_sc_hd__fah_1 U24482 ( .A(n17654), .B(n17653), .CI(n17652), .COUT(
        n18593), .SUM(n17664) );
  sky130_fd_sc_hd__xnor2_1 U24483 ( .A(n18999), .B(n22299), .Y(n18531) );
  sky130_fd_sc_hd__o22ai_1 U24484 ( .A1(n18533), .A2(n18531), .B1(n17655), 
        .B2(n18530), .Y(n18590) );
  sky130_fd_sc_hd__or2_1 U24485 ( .A(n17657), .B(n17656), .X(n18589) );
  sky130_fd_sc_hd__o22ai_1 U24486 ( .A1(n24854), .A2(n24440), .B1(n18026), 
        .B2(n18536), .Y(n18588) );
  sky130_fd_sc_hd__nand2b_1 U24487 ( .A_N(n17662), .B(n17658), .Y(n17659) );
  sky130_fd_sc_hd__nand2_1 U24488 ( .A(n17662), .B(n17661), .Y(n17663) );
  sky130_fd_sc_hd__o21ai_1 U24489 ( .A1(n17666), .A2(n17665), .B1(n17664), .Y(
        n17668) );
  sky130_fd_sc_hd__nand2_1 U24490 ( .A(n17666), .B(n17665), .Y(n17667) );
  sky130_fd_sc_hd__nand2_1 U24491 ( .A(n17668), .B(n17667), .Y(n18575) );
  sky130_fd_sc_hd__fah_1 U24492 ( .A(n17671), .B(n17670), .CI(n17669), .COUT(
        n18576), .SUM(n17662) );
  sky130_fd_sc_hd__xnor2_1 U24493 ( .A(n18994), .B(n25761), .Y(n18484) );
  sky130_fd_sc_hd__o22ai_1 U24494 ( .A1(n18486), .A2(n18484), .B1(n17672), 
        .B2(n18483), .Y(n18554) );
  sky130_fd_sc_hd__nand2b_1 U24495 ( .A_N(n18470), .B(n25389), .Y(n17674) );
  sky130_fd_sc_hd__o22ai_1 U24496 ( .A1(n19023), .A2(n17674), .B1(n17673), 
        .B2(n19020), .Y(n18553) );
  sky130_fd_sc_hd__xnor2_1 U24497 ( .A(n18387), .B(n23567), .Y(n18499) );
  sky130_fd_sc_hd__xnor2_1 U24498 ( .A(n18366), .B(n22087), .Y(n18472) );
  sky130_fd_sc_hd__o22ai_1 U24499 ( .A1(n18474), .A2(n18472), .B1(n17676), 
        .B2(n18471), .Y(n18548) );
  sky130_fd_sc_hd__xnor2_1 U24500 ( .A(n18363), .B(n25389), .Y(n18487) );
  sky130_fd_sc_hd__xnor2_1 U24501 ( .A(n25389), .B(n18210), .Y(n17677) );
  sky130_fd_sc_hd__o22ai_1 U24502 ( .A1(n19023), .A2(n18487), .B1(n17677), 
        .B2(n19020), .Y(n18547) );
  sky130_fd_sc_hd__a21o_1 U24503 ( .A1(n11119), .A2(n18027), .B1(n17678), .X(
        n18546) );
  sky130_fd_sc_hd__fa_1 U24504 ( .A(n17681), .B(n17680), .CIN(n17679), .COUT(
        n18579), .SUM(n17665) );
  sky130_fd_sc_hd__xnor2_1 U24505 ( .A(n18576), .B(n18577), .Y(n17682) );
  sky130_fd_sc_hd__xnor2_1 U24506 ( .A(n18575), .B(n17682), .Y(n18614) );
  sky130_fd_sc_hd__fah_1 U24507 ( .A(n17685), .B(n17683), .CI(n17684), .COUT(
        n17863), .SUM(n17862) );
  sky130_fd_sc_hd__fah_1 U24508 ( .A(n17688), .B(n17687), .CI(n17686), .COUT(
        n17865), .SUM(n17864) );
  sky130_fd_sc_hd__nand2_1 U24509 ( .A(n22956), .B(n17868), .Y(n18335) );
  sky130_fd_sc_hd__xnor2_1 U24510 ( .A(n18371), .B(n25761), .Y(n17745) );
  sky130_fd_sc_hd__xnor2_1 U24511 ( .A(n18994), .B(n27618), .Y(n17746) );
  sky130_fd_sc_hd__o22ai_1 U24512 ( .A1(n18192), .A2(n17693), .B1(n17746), 
        .B2(n18189), .Y(n17708) );
  sky130_fd_sc_hd__xnor2_1 U24513 ( .A(n18941), .B(n24799), .Y(n17743) );
  sky130_fd_sc_hd__xnor2_1 U24514 ( .A(n18363), .B(n22811), .Y(n17737) );
  sky130_fd_sc_hd__o22ai_1 U24515 ( .A1(n18496), .A2(n17695), .B1(n17737), 
        .B2(n17410), .Y(n17706) );
  sky130_fd_sc_hd__xnor2_1 U24516 ( .A(n18387), .B(n18887), .Y(n17731) );
  sky130_fd_sc_hd__o22ai_1 U24517 ( .A1(n18492), .A2(n17696), .B1(n17731), 
        .B2(n18489), .Y(n17705) );
  sky130_fd_sc_hd__xnor2_1 U24518 ( .A(n18999), .B(n21280), .Y(n17733) );
  sky130_fd_sc_hd__o22ai_1 U24519 ( .A1(n18079), .A2(n17697), .B1(n17733), 
        .B2(n18036), .Y(n17704) );
  sky130_fd_sc_hd__fah_1 U24520 ( .A(n17703), .B(n17702), .CI(n17701), .COUT(
        n17814), .SUM(n17822) );
  sky130_fd_sc_hd__fah_1 U24521 ( .A(n17709), .B(n17708), .CI(n17707), .COUT(
        n17771), .SUM(n17776) );
  sky130_fd_sc_hd__xnor2_1 U24522 ( .A(n18925), .B(n24366), .Y(n17717) );
  sky130_fd_sc_hd__xnor2_1 U24523 ( .A(n18966), .B(n24366), .Y(n17726) );
  sky130_fd_sc_hd__o22ai_1 U24524 ( .A1(n18205), .A2(n17717), .B1(n17726), 
        .B2(n12048), .Y(n17792) );
  sky130_fd_sc_hd__nor2b_1 U24525 ( .B_N(n18210), .A(n18496), .Y(n17789) );
  sky130_fd_sc_hd__xnor2_1 U24526 ( .A(n18372), .B(n25761), .Y(n17744) );
  sky130_fd_sc_hd__o22ai_1 U24528 ( .A1(n18486), .A2(n17744), .B1(n17795), 
        .B2(n18483), .Y(n17788) );
  sky130_fd_sc_hd__o22ai_1 U24529 ( .A1(n24854), .A2(n17710), .B1(n22815), 
        .B2(n18224), .Y(n17790) );
  sky130_fd_sc_hd__fah_1 U24530 ( .A(n17713), .B(n17712), .CI(n17711), .COUT(
        n17701), .SUM(n17751) );
  sky130_fd_sc_hd__o22ai_1 U24531 ( .A1(n18205), .A2(n17718), .B1(n17717), 
        .B2(n12048), .Y(n17723) );
  sky130_fd_sc_hd__nor2b_1 U24532 ( .B_N(n18470), .A(n18533), .Y(n17761) );
  sky130_fd_sc_hd__xnor2_1 U24533 ( .A(n18366), .B(n24345), .Y(n17735) );
  sky130_fd_sc_hd__o22ai_1 U24534 ( .A1(n18027), .A2(n17719), .B1(n17735), 
        .B2(n11119), .Y(n17760) );
  sky130_fd_sc_hd__xnor2_1 U24535 ( .A(n17761), .B(n17760), .Y(n17722) );
  sky130_fd_sc_hd__o22ai_1 U24536 ( .A1(n24854), .A2(n17720), .B1(n22318), 
        .B2(n11561), .Y(n17721) );
  sky130_fd_sc_hd__nor2_1 U24537 ( .A(n17807), .B(n17806), .Y(n17748) );
  sky130_fd_sc_hd__fah_1 U24538 ( .A(n17723), .B(n17722), .CI(n17721), .COUT(
        n17749), .SUM(n17873) );
  sky130_fd_sc_hd__xnor2_1 U24539 ( .A(n18367), .B(n24345), .Y(n17734) );
  sky130_fd_sc_hd__xnor2_1 U24540 ( .A(n18387), .B(n24345), .Y(n17787) );
  sky130_fd_sc_hd__o22ai_1 U24541 ( .A1(n18027), .A2(n17734), .B1(n17787), 
        .B2(n11119), .Y(n17894) );
  sky130_fd_sc_hd__xnor2_1 U24542 ( .A(n18377), .B(n18887), .Y(n17730) );
  sky130_fd_sc_hd__xnor2_1 U24543 ( .A(n18371), .B(n18887), .Y(n17798) );
  sky130_fd_sc_hd__o22ai_1 U24544 ( .A1(n18492), .A2(n17730), .B1(n17798), 
        .B2(n18489), .Y(n17893) );
  sky130_fd_sc_hd__xnor2_1 U24545 ( .A(j202_soc_core_j22_cpu_ml_bufa[2]), .B(
        j202_soc_core_j22_cpu_ml_bufa[1]), .Y(n17724) );
  sky130_fd_sc_hd__xnor2_1 U24546 ( .A(n22024), .B(n21219), .Y(n17738) );
  sky130_fd_sc_hd__xnor2_1 U24547 ( .A(n18925), .B(n21219), .Y(n17796) );
  sky130_fd_sc_hd__xor2_1 U24548 ( .A(j202_soc_core_j22_cpu_ml_bufa[3]), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n17725) );
  sky130_fd_sc_hd__nand2_2 U24549 ( .A(n17725), .B(n17724), .Y(n18206) );
  sky130_fd_sc_hd__o22ai_1 U24550 ( .A1(n18209), .A2(n17738), .B1(n17796), 
        .B2(n18206), .Y(n17892) );
  sky130_fd_sc_hd__xnor2_1 U24551 ( .A(n18994), .B(n24366), .Y(n17898) );
  sky130_fd_sc_hd__o22ai_1 U24552 ( .A1(n18205), .A2(n17726), .B1(n17898), 
        .B2(n18202), .Y(n17897) );
  sky130_fd_sc_hd__xnor2_1 U24553 ( .A(n18964), .B(n21280), .Y(n17732) );
  sky130_fd_sc_hd__xnor2_1 U24554 ( .A(n18366), .B(n21280), .Y(n17797) );
  sky130_fd_sc_hd__o22ai_1 U24555 ( .A1(n18079), .A2(n17732), .B1(n17797), 
        .B2(n18036), .Y(n17896) );
  sky130_fd_sc_hd__xnor2_1 U24556 ( .A(n18962), .B(n24799), .Y(n17742) );
  sky130_fd_sc_hd__xnor2_1 U24557 ( .A(n18999), .B(n24799), .Y(n17793) );
  sky130_fd_sc_hd__nand2b_1 U24558 ( .A_N(n18470), .B(n22811), .Y(n17728) );
  sky130_fd_sc_hd__o22ai_1 U24559 ( .A1(n18496), .A2(n17728), .B1(n17727), 
        .B2(n17410), .Y(n17741) );
  sky130_fd_sc_hd__o22ai_1 U24560 ( .A1(n18079), .A2(n17733), .B1(n17732), 
        .B2(n18036), .Y(n17739) );
  sky130_fd_sc_hd__o22ai_1 U24561 ( .A1(n18027), .A2(n17735), .B1(n17734), 
        .B2(n11119), .Y(n17783) );
  sky130_fd_sc_hd__xnor2_1 U24562 ( .A(n22811), .B(n18210), .Y(n17736) );
  sky130_fd_sc_hd__o22ai_1 U24563 ( .A1(n18496), .A2(n17737), .B1(n17736), 
        .B2(n17410), .Y(n17782) );
  sky130_fd_sc_hd__a21o_1 U24564 ( .A1(n18206), .A2(n18209), .B1(n17738), .X(
        n17781) );
  sky130_fd_sc_hd__o22ai_1 U24565 ( .A1(n18486), .A2(n17745), .B1(n17744), 
        .B2(n18483), .Y(n17779) );
  sky130_fd_sc_hd__xnor2_1 U24566 ( .A(n18971), .B(n27618), .Y(n17784) );
  sky130_fd_sc_hd__o22ai_1 U24567 ( .A1(n18192), .A2(n17746), .B1(n17784), 
        .B2(n18189), .Y(n17778) );
  sky130_fd_sc_hd__fah_1 U24568 ( .A(n17751), .B(n17750), .CI(n17749), .COUT(
        n17827), .SUM(n17806) );
  sky130_fd_sc_hd__nand2b_1 U24570 ( .A_N(n18470), .B(n22299), .Y(n17759) );
  sky130_fd_sc_hd__o22ai_1 U24571 ( .A1(n18533), .A2(n17759), .B1(n17758), 
        .B2(n18530), .Y(n17765) );
  sky130_fd_sc_hd__o22ai_1 U24573 ( .A1(n24854), .A2(n17762), .B1(n22279), 
        .B2(n18536), .Y(n17763) );
  sky130_fd_sc_hd__fah_1 U24574 ( .A(n17765), .B(n17764), .CI(n17763), .COUT(
        n17816), .SUM(n17774) );
  sky130_fd_sc_hd__fah_1 U24575 ( .A(n17769), .B(n17770), .CI(n17771), .COUT(
        n17823), .SUM(n17772) );
  sky130_fd_sc_hd__fah_1 U24576 ( .A(n17774), .B(n17773), .CI(n17772), .COUT(
        n17825), .SUM(n17909) );
  sky130_fd_sc_hd__fah_1 U24577 ( .A(n17783), .B(n17782), .CI(n17781), .COUT(
        n17768), .SUM(n17890) );
  sky130_fd_sc_hd__xnor2_1 U24578 ( .A(n18941), .B(n27618), .Y(n17899) );
  sky130_fd_sc_hd__o22ai_1 U24579 ( .A1(n18192), .A2(n17784), .B1(n17899), 
        .B2(n18189), .Y(n17880) );
  sky130_fd_sc_hd__nand2b_1 U24580 ( .A_N(n18470), .B(n25761), .Y(n17786) );
  sky130_fd_sc_hd__o22ai_1 U24581 ( .A1(n18486), .A2(n17786), .B1(n17785), 
        .B2(n18483), .Y(n17901) );
  sky130_fd_sc_hd__xnor2_1 U24582 ( .A(n18377), .B(n24345), .Y(n17884) );
  sky130_fd_sc_hd__o22ai_1 U24583 ( .A1(n18027), .A2(n17787), .B1(n17884), 
        .B2(n11119), .Y(n17900) );
  sky130_fd_sc_hd__or2_1 U24584 ( .A(n17901), .B(n17900), .X(n17879) );
  sky130_fd_sc_hd__xnor2_1 U24585 ( .A(n17789), .B(n17788), .Y(n17878) );
  sky130_fd_sc_hd__xnor2_1 U24586 ( .A(n18964), .B(n24799), .Y(n17883) );
  sky130_fd_sc_hd__xnor2_1 U24587 ( .A(n25761), .B(n18210), .Y(n17794) );
  sky130_fd_sc_hd__o22ai_1 U24588 ( .A1(n18486), .A2(n17795), .B1(n17794), 
        .B2(n18483), .Y(n17919) );
  sky130_fd_sc_hd__inv_4 U24589 ( .A(j202_soc_core_j22_cpu_ml_bufa[0]), .Y(
        n18188) );
  sky130_fd_sc_hd__nand2_2 U24590 ( .A(n21943), .B(n18188), .Y(n18185) );
  sky130_fd_sc_hd__buf_6 U24591 ( .A(j202_soc_core_j22_cpu_ml_bufa[1]), .X(
        n21943) );
  sky130_fd_sc_hd__xnor2_1 U24592 ( .A(n22024), .B(n21943), .Y(n17881) );
  sky130_fd_sc_hd__a21o_1 U24593 ( .A1(n18185), .A2(n18188), .B1(n17881), .X(
        n17918) );
  sky130_fd_sc_hd__o22ai_1 U24594 ( .A1(n24854), .A2(n18406), .B1(n22366), 
        .B2(n11561), .Y(n17887) );
  sky130_fd_sc_hd__xnor2_1 U24595 ( .A(n18966), .B(n21219), .Y(n17913) );
  sky130_fd_sc_hd__o22ai_1 U24596 ( .A1(n18209), .A2(n17796), .B1(n17913), 
        .B2(n18206), .Y(n17917) );
  sky130_fd_sc_hd__xnor2_1 U24597 ( .A(n18367), .B(n21280), .Y(n17882) );
  sky130_fd_sc_hd__o22ai_1 U24598 ( .A1(n18079), .A2(n17797), .B1(n17882), 
        .B2(n18036), .Y(n17916) );
  sky130_fd_sc_hd__xnor2_1 U24599 ( .A(n18372), .B(n18887), .Y(n17885) );
  sky130_fd_sc_hd__o21ai_1 U24600 ( .A1(n17911), .A2(n17910), .B1(n17912), .Y(
        n17803) );
  sky130_fd_sc_hd__nand2_1 U24601 ( .A(n17910), .B(n17911), .Y(n17802) );
  sky130_fd_sc_hd__nand2_1 U24602 ( .A(n17803), .B(n17802), .Y(n17877) );
  sky130_fd_sc_hd__nand2_1 U24604 ( .A(n17875), .B(n17874), .Y(n17804) );
  sky130_fd_sc_hd__nand2_1 U24605 ( .A(n17805), .B(n17804), .Y(n17908) );
  sky130_fd_sc_hd__xnor2_1 U24606 ( .A(n17807), .B(n17806), .Y(n17808) );
  sky130_fd_sc_hd__xnor2_1 U24607 ( .A(n17809), .B(n17808), .Y(n17907) );
  sky130_fd_sc_hd__fah_1 U24608 ( .A(n17812), .B(n17811), .CI(n17810), .COUT(
        n17828), .SUM(n18332) );
  sky130_fd_sc_hd__fah_1 U24609 ( .A(n17818), .B(n17817), .CI(n17816), .COUT(
        n17840), .SUM(n17826) );
  sky130_fd_sc_hd__fah_1 U24610 ( .A(n17821), .B(n17820), .CI(n17819), .COUT(
        n17846), .SUM(n17841) );
  sky130_fd_sc_hd__fah_1 U24611 ( .A(n17827), .B(n17826), .CI(n17825), .COUT(
        n17831), .SUM(n17810) );
  sky130_fd_sc_hd__o21ai_1 U24612 ( .A1(n17830), .A2(n17831), .B1(n17829), .Y(
        n17833) );
  sky130_fd_sc_hd__nand2_1 U24613 ( .A(n17831), .B(n17830), .Y(n17832) );
  sky130_fd_sc_hd__nand2_1 U24614 ( .A(n17833), .B(n17832), .Y(n17855) );
  sky130_fd_sc_hd__fah_1 U24615 ( .A(n17836), .B(n17835), .CI(n17834), .COUT(
        n17552), .SUM(n17849) );
  sky130_fd_sc_hd__nand2b_1 U24616 ( .A_N(n17841), .B(n17837), .Y(n17838) );
  sky130_fd_sc_hd__nand2_1 U24617 ( .A(n17839), .B(n17838), .Y(n17843) );
  sky130_fd_sc_hd__nand2_1 U24618 ( .A(n17841), .B(n17840), .Y(n17842) );
  sky130_fd_sc_hd__nand2_1 U24619 ( .A(n17843), .B(n17842), .Y(n17848) );
  sky130_fd_sc_hd__fah_1 U24620 ( .A(n17846), .B(n17845), .CI(n17844), .COUT(
        n17854), .SUM(n17847) );
  sky130_fd_sc_hd__nor2_1 U24621 ( .A(n17855), .B(n17856), .Y(n21752) );
  sky130_fd_sc_hd__xnor2_1 U24622 ( .A(n17852), .B(n17851), .Y(n17853) );
  sky130_fd_sc_hd__nand2_1 U24623 ( .A(n17856), .B(n17855), .Y(n22873) );
  sky130_fd_sc_hd__o21ai_1 U24624 ( .A1(n22873), .A2(n22869), .B1(n22870), .Y(
        n17858) );
  sky130_fd_sc_hd__a21oi_2 U24625 ( .A1(n21753), .A2(n18334), .B1(n17858), .Y(
        n19304) );
  sky130_fd_sc_hd__nand2_1 U24626 ( .A(n17860), .B(n17859), .Y(n21273) );
  sky130_fd_sc_hd__nand2_1 U24627 ( .A(n17862), .B(n17861), .Y(n21269) );
  sky130_fd_sc_hd__nand2_1 U24628 ( .A(n17864), .B(n17863), .Y(n22960) );
  sky130_fd_sc_hd__nand2_1 U24629 ( .A(n17866), .B(n17865), .Y(n22954) );
  sky130_fd_sc_hd__o21ai_1 U24630 ( .A1(n22960), .A2(n22953), .B1(n22954), .Y(
        n17867) );
  sky130_fd_sc_hd__o21ai_1 U24631 ( .A1(n18335), .A2(n19304), .B1(n17869), .Y(
        n17870) );
  sky130_fd_sc_hd__fah_1 U24632 ( .A(n17873), .B(n17872), .CI(n17871), .COUT(
        n17809), .SUM(n17948) );
  sky130_fd_sc_hd__xnor2_1 U24633 ( .A(n17875), .B(n17874), .Y(n17876) );
  sky130_fd_sc_hd__fah_1 U24634 ( .A(n17880), .B(n17879), .CI(n17878), .COUT(
        n17889), .SUM(n17998) );
  sky130_fd_sc_hd__xnor2_1 U24635 ( .A(n18925), .B(n21943), .Y(n17924) );
  sky130_fd_sc_hd__o22ai_1 U24636 ( .A1(n18188), .A2(n17881), .B1(n17924), 
        .B2(n18185), .Y(n17975) );
  sky130_fd_sc_hd__xnor2_1 U24637 ( .A(n18387), .B(n21280), .Y(n17926) );
  sky130_fd_sc_hd__o22ai_1 U24638 ( .A1(n18079), .A2(n17882), .B1(n17926), 
        .B2(n18036), .Y(n17974) );
  sky130_fd_sc_hd__xnor2_1 U24639 ( .A(n18366), .B(n24799), .Y(n17935) );
  sky130_fd_sc_hd__xnor2_1 U24640 ( .A(n18371), .B(n24345), .Y(n17925) );
  sky130_fd_sc_hd__o22ai_1 U24641 ( .A1(n18027), .A2(n17884), .B1(n17925), 
        .B2(n11119), .Y(n17938) );
  sky130_fd_sc_hd__xnor2_1 U24642 ( .A(n18363), .B(n18887), .Y(n17929) );
  sky130_fd_sc_hd__o22ai_1 U24643 ( .A1(n18492), .A2(n17885), .B1(n17929), 
        .B2(n18489), .Y(n17937) );
  sky130_fd_sc_hd__o22ai_1 U24644 ( .A1(n24854), .A2(n18360), .B1(n22844), 
        .B2(n18536), .Y(n17967) );
  sky130_fd_sc_hd__fah_1 U24645 ( .A(n17891), .B(n17890), .CI(n17889), .COUT(
        n17875), .SUM(n17943) );
  sky130_fd_sc_hd__fah_1 U24646 ( .A(n17897), .B(n17896), .CI(n17895), .COUT(
        n17800), .SUM(n17922) );
  sky130_fd_sc_hd__xnor2_1 U24647 ( .A(n18971), .B(n24366), .Y(n17915) );
  sky130_fd_sc_hd__o22ai_1 U24648 ( .A1(n18205), .A2(n17898), .B1(n17915), 
        .B2(n12048), .Y(n17932) );
  sky130_fd_sc_hd__xnor2_1 U24649 ( .A(n18962), .B(n27618), .Y(n17914) );
  sky130_fd_sc_hd__o22ai_1 U24650 ( .A1(n18192), .A2(n17899), .B1(n17914), 
        .B2(n18189), .Y(n17931) );
  sky130_fd_sc_hd__xnor2_1 U24651 ( .A(n17901), .B(n17900), .Y(n17930) );
  sky130_fd_sc_hd__nand2_1 U24652 ( .A(n17903), .B(n17902), .Y(n17904) );
  sky130_fd_sc_hd__nand2_1 U24653 ( .A(n17946), .B(n17904), .Y(n17906) );
  sky130_fd_sc_hd__nand2_1 U24654 ( .A(n17943), .B(n17944), .Y(n17905) );
  sky130_fd_sc_hd__fah_1 U24655 ( .A(n17909), .B(n17908), .CI(n17907), .COUT(
        n18333), .SUM(n18327) );
  sky130_fd_sc_hd__nor2_2 U24656 ( .A(n18326), .B(n18327), .Y(n22215) );
  sky130_fd_sc_hd__xnor2_1 U24657 ( .A(n18994), .B(n21219), .Y(n17927) );
  sky130_fd_sc_hd__o22ai_1 U24658 ( .A1(n18209), .A2(n17913), .B1(n17927), 
        .B2(n18206), .Y(n17942) );
  sky130_fd_sc_hd__xnor2_1 U24659 ( .A(n18999), .B(n27618), .Y(n17936) );
  sky130_fd_sc_hd__o22ai_1 U24660 ( .A1(n18192), .A2(n17914), .B1(n17936), 
        .B2(n18189), .Y(n17941) );
  sky130_fd_sc_hd__xnor2_1 U24661 ( .A(n18941), .B(n24366), .Y(n17976) );
  sky130_fd_sc_hd__o22ai_1 U24662 ( .A1(n18205), .A2(n17915), .B1(n17976), 
        .B2(n12048), .Y(n17940) );
  sky130_fd_sc_hd__fah_1 U24663 ( .A(n17923), .B(n17922), .CI(n17921), .COUT(
        n17944), .SUM(n18003) );
  sky130_fd_sc_hd__xnor2_1 U24664 ( .A(n18966), .B(n21943), .Y(n17983) );
  sky130_fd_sc_hd__o22ai_1 U24665 ( .A1(n18188), .A2(n17924), .B1(n17983), 
        .B2(n18185), .Y(n17978) );
  sky130_fd_sc_hd__xnor2_1 U24666 ( .A(n18372), .B(n24345), .Y(n17980) );
  sky130_fd_sc_hd__o22ai_1 U24667 ( .A1(n18027), .A2(n17925), .B1(n17980), 
        .B2(n11119), .Y(n17977) );
  sky130_fd_sc_hd__xnor2_1 U24668 ( .A(n18377), .B(n21280), .Y(n17982) );
  sky130_fd_sc_hd__o22ai_1 U24669 ( .A1(n18079), .A2(n17926), .B1(n17982), 
        .B2(n18036), .Y(n17963) );
  sky130_fd_sc_hd__xnor2_1 U24670 ( .A(n18971), .B(n21219), .Y(n17989) );
  sky130_fd_sc_hd__o22ai_1 U24671 ( .A1(n18209), .A2(n17927), .B1(n17989), 
        .B2(n18206), .Y(n17962) );
  sky130_fd_sc_hd__xnor2_1 U24672 ( .A(n18887), .B(n18210), .Y(n17928) );
  sky130_fd_sc_hd__o22ai_1 U24673 ( .A1(n18492), .A2(n17929), .B1(n17928), 
        .B2(n18489), .Y(n17961) );
  sky130_fd_sc_hd__nand2b_1 U24674 ( .A_N(n18470), .B(n18887), .Y(n17934) );
  sky130_fd_sc_hd__o22ai_1 U24675 ( .A1(n18492), .A2(n17934), .B1(n17933), 
        .B2(n18489), .Y(n17960) );
  sky130_fd_sc_hd__xnor2_1 U24676 ( .A(n18367), .B(n24799), .Y(n17987) );
  sky130_fd_sc_hd__xnor2_1 U24677 ( .A(n18964), .B(n27618), .Y(n17985) );
  sky130_fd_sc_hd__o22ai_1 U24678 ( .A1(n18192), .A2(n17936), .B1(n17985), 
        .B2(n18189), .Y(n17958) );
  sky130_fd_sc_hd__fah_1 U24679 ( .A(n17939), .B(n17938), .CI(n17937), .COUT(
        n17968), .SUM(n17956) );
  sky130_fd_sc_hd__fa_1 U24680 ( .A(n17942), .B(n17941), .CIN(n17940), .COUT(
        n17972), .SUM(n17955) );
  sky130_fd_sc_hd__xnor2_1 U24681 ( .A(n17944), .B(n17943), .Y(n17945) );
  sky130_fd_sc_hd__xnor2_1 U24682 ( .A(n17946), .B(n17945), .Y(n18008) );
  sky130_fd_sc_hd__fah_1 U24683 ( .A(n17951), .B(n17950), .CI(n17949), .COUT(
        n18002), .SUM(n18313) );
  sky130_fd_sc_hd__fah_1 U24684 ( .A(n17954), .B(n17953), .CI(n17952), .COUT(
        n17951), .SUM(n18307) );
  sky130_fd_sc_hd__fah_1 U24685 ( .A(n17957), .B(n17956), .CI(n17955), .COUT(
        n17949), .SUM(n18306) );
  sky130_fd_sc_hd__o22ai_1 U24686 ( .A1(n22365), .A2(n22561), .B1(n24464), 
        .B2(n11561), .Y(n18046) );
  sky130_fd_sc_hd__xnor2_1 U24687 ( .A(n18387), .B(n24799), .Y(n17986) );
  sky130_fd_sc_hd__xnor2_1 U24688 ( .A(n18377), .B(n24799), .Y(n18020) );
  sky130_fd_sc_hd__xnor2_1 U24689 ( .A(n18941), .B(n21219), .Y(n17988) );
  sky130_fd_sc_hd__xnor2_1 U24690 ( .A(n18962), .B(n21219), .Y(n18029) );
  sky130_fd_sc_hd__o22ai_1 U24691 ( .A1(n18209), .A2(n17988), .B1(n18029), 
        .B2(n18206), .Y(n18054) );
  sky130_fd_sc_hd__xnor2_1 U24692 ( .A(n18363), .B(n24345), .Y(n17979) );
  sky130_fd_sc_hd__xnor2_1 U24693 ( .A(n24345), .B(n18210), .Y(n17966) );
  sky130_fd_sc_hd__o22ai_1 U24694 ( .A1(n18027), .A2(n17979), .B1(n17966), 
        .B2(n11119), .Y(n18053) );
  sky130_fd_sc_hd__xnor2_1 U24695 ( .A(n18999), .B(n24366), .Y(n17990) );
  sky130_fd_sc_hd__xnor2_1 U24696 ( .A(n18964), .B(n24366), .Y(n18035) );
  sky130_fd_sc_hd__o22ai_1 U24697 ( .A1(n18205), .A2(n17990), .B1(n18035), 
        .B2(n12048), .Y(n18052) );
  sky130_fd_sc_hd__xnor2_1 U24698 ( .A(n18371), .B(n21280), .Y(n17981) );
  sky130_fd_sc_hd__xnor2_1 U24699 ( .A(n18372), .B(n21280), .Y(n18038) );
  sky130_fd_sc_hd__o22ai_1 U24700 ( .A1(n18079), .A2(n17981), .B1(n18038), 
        .B2(n18036), .Y(n18051) );
  sky130_fd_sc_hd__xnor2_1 U24701 ( .A(n18366), .B(n27618), .Y(n17984) );
  sky130_fd_sc_hd__xnor2_1 U24702 ( .A(n18367), .B(n27618), .Y(n18040) );
  sky130_fd_sc_hd__o22ai_1 U24703 ( .A1(n18192), .A2(n17984), .B1(n18040), 
        .B2(n18189), .Y(n18050) );
  sky130_fd_sc_hd__fa_2 U24704 ( .A(n17969), .B(n17968), .CIN(n17967), .COUT(
        n17997), .SUM(n18001) );
  sky130_fd_sc_hd__fah_1 U24705 ( .A(n17972), .B(n17971), .CI(n17970), .COUT(
        n18004), .SUM(n18000) );
  sky130_fd_sc_hd__fah_1 U24706 ( .A(n17975), .B(n17974), .CI(n17973), .COUT(
        n17969), .SUM(n18301) );
  sky130_fd_sc_hd__xnor2_1 U24707 ( .A(n18962), .B(n24366), .Y(n17991) );
  sky130_fd_sc_hd__o22ai_1 U24708 ( .A1(n18205), .A2(n17976), .B1(n17991), 
        .B2(n12048), .Y(n18064) );
  sky130_fd_sc_hd__ha_1 U24709 ( .A(n17978), .B(n17977), .COUT(n17954), .SUM(
        n18063) );
  sky130_fd_sc_hd__o22ai_1 U24710 ( .A1(n22365), .A2(n18475), .B1(n18888), 
        .B2(n18536), .Y(n18062) );
  sky130_fd_sc_hd__nor2b_1 U24711 ( .B_N(n18470), .A(n18492), .Y(n18013) );
  sky130_fd_sc_hd__o22ai_1 U24712 ( .A1(n18027), .A2(n17980), .B1(n17979), 
        .B2(n11119), .Y(n18012) );
  sky130_fd_sc_hd__o22ai_1 U24713 ( .A1(n18079), .A2(n17982), .B1(n17981), 
        .B2(n18036), .Y(n18011) );
  sky130_fd_sc_hd__xnor2_1 U24714 ( .A(n18994), .B(n21943), .Y(n17992) );
  sky130_fd_sc_hd__o22ai_1 U24715 ( .A1(n18188), .A2(n17983), .B1(n17992), 
        .B2(n18185), .Y(n18016) );
  sky130_fd_sc_hd__o22ai_1 U24716 ( .A1(n18192), .A2(n17985), .B1(n17984), 
        .B2(n18189), .Y(n18015) );
  sky130_fd_sc_hd__o22ai_1 U24717 ( .A1(n18209), .A2(n17989), .B1(n17988), 
        .B2(n18206), .Y(n18019) );
  sky130_fd_sc_hd__o22ai_1 U24718 ( .A1(n18205), .A2(n17991), .B1(n17990), 
        .B2(n12048), .Y(n18018) );
  sky130_fd_sc_hd__xnor2_1 U24719 ( .A(n18971), .B(n21943), .Y(n18028) );
  sky130_fd_sc_hd__o22ai_1 U24720 ( .A1(n18188), .A2(n17992), .B1(n18028), 
        .B2(n18185), .Y(n18025) );
  sky130_fd_sc_hd__nand2b_1 U24721 ( .A_N(n18470), .B(n24345), .Y(n17995) );
  sky130_fd_sc_hd__o22ai_1 U24722 ( .A1(n18027), .A2(n17995), .B1(n17994), 
        .B2(n11119), .Y(n18024) );
  sky130_fd_sc_hd__nor2_1 U24723 ( .A(n18320), .B(n18321), .Y(n19109) );
  sky130_fd_sc_hd__fah_1 U24724 ( .A(n18007), .B(n18006), .CI(n18005), .COUT(
        n18322), .SUM(n18321) );
  sky130_fd_sc_hd__fah_1 U24725 ( .A(n18010), .B(n18009), .CI(n18008), .COUT(
        n18324), .SUM(n18323) );
  sky130_fd_sc_hd__nand2_1 U24727 ( .A(n18329), .B(n22207), .Y(n18331) );
  sky130_fd_sc_hd__fah_1 U24728 ( .A(n18013), .B(n18012), .CI(n18011), .COUT(
        n18070), .SUM(n18067) );
  sky130_fd_sc_hd__xnor2_1 U24729 ( .A(n18371), .B(n24799), .Y(n18021) );
  sky130_fd_sc_hd__xnor2_1 U24730 ( .A(n18372), .B(n24799), .Y(n18081) );
  sky130_fd_sc_hd__nand2b_1 U24731 ( .A_N(n18470), .B(n21280), .Y(n18023) );
  sky130_fd_sc_hd__o22ai_1 U24732 ( .A1(n18079), .A2(n18023), .B1(n18022), 
        .B2(n18036), .Y(n18076) );
  sky130_fd_sc_hd__o22ai_1 U24733 ( .A1(n22365), .A2(n22630), .B1(n21883), 
        .B2(n18536), .Y(n18085) );
  sky130_fd_sc_hd__o22ai_1 U24734 ( .A1(n22365), .A2(n18026), .B1(n24445), 
        .B2(n11561), .Y(n18042) );
  sky130_fd_sc_hd__nor2b_1 U24735 ( .B_N(n18470), .A(n18027), .Y(n18034) );
  sky130_fd_sc_hd__xnor2_1 U24736 ( .A(n18941), .B(n21943), .Y(n18030) );
  sky130_fd_sc_hd__o22ai_1 U24737 ( .A1(n18188), .A2(n18028), .B1(n18030), 
        .B2(n18185), .Y(n18033) );
  sky130_fd_sc_hd__xnor2_1 U24738 ( .A(n18999), .B(n21219), .Y(n18074) );
  sky130_fd_sc_hd__xnor2_1 U24739 ( .A(n18387), .B(n27618), .Y(n18039) );
  sky130_fd_sc_hd__xnor2_1 U24740 ( .A(n18377), .B(n27618), .Y(n18083) );
  sky130_fd_sc_hd__o22ai_1 U24741 ( .A1(n18192), .A2(n18039), .B1(n18083), 
        .B2(n18189), .Y(n18247) );
  sky130_fd_sc_hd__xnor2_1 U24742 ( .A(n18962), .B(n21943), .Y(n18080) );
  sky130_fd_sc_hd__o22ai_1 U24743 ( .A1(n18188), .A2(n18030), .B1(n18080), 
        .B2(n18185), .Y(n18246) );
  sky130_fd_sc_hd__xnor2_1 U24744 ( .A(n18363), .B(n21280), .Y(n18037) );
  sky130_fd_sc_hd__xnor2_1 U24745 ( .A(n21280), .B(n18210), .Y(n18031) );
  sky130_fd_sc_hd__o22ai_1 U24746 ( .A1(n18079), .A2(n18037), .B1(n18031), 
        .B2(n18036), .Y(n18245) );
  sky130_fd_sc_hd__fa_1 U24747 ( .A(n18034), .B(n18033), .CIN(n18032), .COUT(
        n18041), .SUM(n18270) );
  sky130_fd_sc_hd__xnor2_1 U24748 ( .A(n18366), .B(n24366), .Y(n18075) );
  sky130_fd_sc_hd__o22ai_1 U24749 ( .A1(n18205), .A2(n18035), .B1(n18075), 
        .B2(n12048), .Y(n18049) );
  sky130_fd_sc_hd__o22ai_1 U24750 ( .A1(n18079), .A2(n18038), .B1(n18037), 
        .B2(n18036), .Y(n18048) );
  sky130_fd_sc_hd__o22ai_1 U24751 ( .A1(n18192), .A2(n18040), .B1(n18039), 
        .B2(n18189), .Y(n18047) );
  sky130_fd_sc_hd__fah_1 U24752 ( .A(n18052), .B(n18051), .CI(n18050), .COUT(
        n18044), .SUM(n18072) );
  sky130_fd_sc_hd__fah_1 U24753 ( .A(n18058), .B(n18057), .CI(n18056), .COUT(
        n18305), .SUM(n18298) );
  sky130_fd_sc_hd__fah_1 U24754 ( .A(n18061), .B(n18060), .CI(n18059), .COUT(
        n18297), .SUM(n18091) );
  sky130_fd_sc_hd__nor2_1 U24755 ( .A(n18291), .B(n18292), .Y(n18293) );
  sky130_fd_sc_hd__fa_1 U24756 ( .A(n18073), .B(n18072), .CIN(n18071), .COUT(
        n18059), .SUM(n18283) );
  sky130_fd_sc_hd__xnor2_1 U24757 ( .A(n18964), .B(n21219), .Y(n18082) );
  sky130_fd_sc_hd__o22ai_1 U24758 ( .A1(n18209), .A2(n18074), .B1(n18082), 
        .B2(n18206), .Y(n18250) );
  sky130_fd_sc_hd__xnor2_1 U24759 ( .A(n18367), .B(n24366), .Y(n18084) );
  sky130_fd_sc_hd__o22ai_1 U24760 ( .A1(n18205), .A2(n18075), .B1(n18084), 
        .B2(n12048), .Y(n18249) );
  sky130_fd_sc_hd__ha_1 U24761 ( .A(n18077), .B(n18076), .COUT(n18086), .SUM(
        n18248) );
  sky130_fd_sc_hd__o22ai_1 U24762 ( .A1(n22365), .A2(n22522), .B1(n18078), 
        .B2(n11561), .Y(n18241) );
  sky130_fd_sc_hd__nor2b_1 U24763 ( .B_N(n18470), .A(n18079), .Y(n18233) );
  sky130_fd_sc_hd__xnor2_1 U24764 ( .A(n18999), .B(n21943), .Y(n18187) );
  sky130_fd_sc_hd__o22ai_1 U24765 ( .A1(n18188), .A2(n18080), .B1(n18187), 
        .B2(n18185), .Y(n18232) );
  sky130_fd_sc_hd__xnor2_1 U24766 ( .A(n18363), .B(n24799), .Y(n18212) );
  sky130_fd_sc_hd__xnor2_1 U24767 ( .A(n18366), .B(n21219), .Y(n18208) );
  sky130_fd_sc_hd__xnor2_1 U24768 ( .A(n18371), .B(n27618), .Y(n18191) );
  sky130_fd_sc_hd__o22ai_1 U24769 ( .A1(n18192), .A2(n18083), .B1(n18191), 
        .B2(n18189), .Y(n18235) );
  sky130_fd_sc_hd__xnor2_1 U24770 ( .A(n18387), .B(n24366), .Y(n18204) );
  sky130_fd_sc_hd__o22ai_1 U24771 ( .A1(n18205), .A2(n18084), .B1(n18204), 
        .B2(n12048), .Y(n18234) );
  sky130_fd_sc_hd__fa_1 U24772 ( .A(n18087), .B(n18086), .CIN(n18085), .COUT(
        n18090), .SUM(n18275) );
  sky130_fd_sc_hd__fah_1 U24773 ( .A(n18093), .B(n18092), .CI(n18091), .COUT(
        n18291), .SUM(n18290) );
  sky130_fd_sc_hd__nor2_1 U24774 ( .A(n18289), .B(n18290), .Y(n18094) );
  sky130_fd_sc_hd__nand2_1 U24775 ( .A(n18884), .B(n22567), .Y(n18295) );
  sky130_fd_sc_hd__xnor2_1 U24776 ( .A(n18377), .B(n21219), .Y(n18104) );
  sky130_fd_sc_hd__xnor2_1 U24777 ( .A(n18371), .B(n21219), .Y(n18095) );
  sky130_fd_sc_hd__o22ai_1 U24778 ( .A1(n18209), .A2(n18104), .B1(n18095), 
        .B2(n18206), .Y(n18113) );
  sky130_fd_sc_hd__xnor2_1 U24779 ( .A(n18372), .B(n24366), .Y(n18109) );
  sky130_fd_sc_hd__xnor2_1 U24780 ( .A(n18363), .B(n24366), .Y(n18097) );
  sky130_fd_sc_hd__o22ai_1 U24781 ( .A1(n18205), .A2(n18109), .B1(n18097), 
        .B2(n12048), .Y(n18112) );
  sky130_fd_sc_hd__xnor2_1 U24782 ( .A(n18372), .B(n21219), .Y(n18117) );
  sky130_fd_sc_hd__o22ai_1 U24783 ( .A1(n18209), .A2(n18095), .B1(n18117), 
        .B2(n18206), .Y(n18125) );
  sky130_fd_sc_hd__xnor2_1 U24784 ( .A(n24366), .B(n18210), .Y(n18096) );
  sky130_fd_sc_hd__o22ai_1 U24785 ( .A1(n18205), .A2(n18097), .B1(n18096), 
        .B2(n12048), .Y(n18124) );
  sky130_fd_sc_hd__nand2b_1 U24786 ( .A_N(n18470), .B(n24366), .Y(n18099) );
  sky130_fd_sc_hd__o22ai_1 U24787 ( .A1(n18205), .A2(n18099), .B1(n18098), 
        .B2(n12048), .Y(n18102) );
  sky130_fd_sc_hd__xnor2_1 U24788 ( .A(n18387), .B(n21943), .Y(n18100) );
  sky130_fd_sc_hd__xnor2_1 U24789 ( .A(n18377), .B(n21943), .Y(n18119) );
  sky130_fd_sc_hd__o22ai_1 U24790 ( .A1(n18188), .A2(n18100), .B1(n18119), 
        .B2(n18185), .Y(n18101) );
  sky130_fd_sc_hd__xnor2_1 U24791 ( .A(n18367), .B(n21943), .Y(n18103) );
  sky130_fd_sc_hd__o22ai_1 U24792 ( .A1(n18188), .A2(n18103), .B1(n18100), 
        .B2(n18185), .Y(n18108) );
  sky130_fd_sc_hd__ha_1 U24793 ( .A(n18102), .B(n18101), .COUT(n18107), .SUM(
        n18123) );
  sky130_fd_sc_hd__o22ai_1 U24794 ( .A1(n22365), .A2(n22148), .B1(n22131), 
        .B2(n11561), .Y(n18106) );
  sky130_fd_sc_hd__xnor2_1 U24795 ( .A(n18366), .B(n21943), .Y(n18180) );
  sky130_fd_sc_hd__o22ai_1 U24796 ( .A1(n18188), .A2(n18180), .B1(n18103), 
        .B2(n18185), .Y(n18178) );
  sky130_fd_sc_hd__xnor2_1 U24797 ( .A(n18387), .B(n21219), .Y(n18181) );
  sky130_fd_sc_hd__o22ai_1 U24798 ( .A1(n18209), .A2(n18181), .B1(n18104), 
        .B2(n18206), .Y(n18177) );
  sky130_fd_sc_hd__xnor2_1 U24799 ( .A(n18363), .B(n27618), .Y(n18170) );
  sky130_fd_sc_hd__xnor2_1 U24800 ( .A(n27618), .B(n18210), .Y(n18105) );
  sky130_fd_sc_hd__o22ai_1 U24801 ( .A1(n18192), .A2(n18170), .B1(n18105), 
        .B2(n18189), .Y(n18176) );
  sky130_fd_sc_hd__fah_1 U24802 ( .A(n18108), .B(n18107), .CI(n18106), .COUT(
        n18167), .SUM(n18158) );
  sky130_fd_sc_hd__xnor2_1 U24803 ( .A(n18371), .B(n24366), .Y(n18169) );
  sky130_fd_sc_hd__o22ai_1 U24804 ( .A1(n18205), .A2(n18169), .B1(n18109), 
        .B2(n12048), .Y(n18172) );
  sky130_fd_sc_hd__nand2b_1 U24805 ( .A_N(n18470), .B(n27618), .Y(n18111) );
  sky130_fd_sc_hd__o22ai_1 U24806 ( .A1(n18192), .A2(n18111), .B1(n18110), 
        .B2(n18189), .Y(n18171) );
  sky130_fd_sc_hd__xnor2_1 U24807 ( .A(n18371), .B(n21943), .Y(n18118) );
  sky130_fd_sc_hd__xnor2_1 U24808 ( .A(n18372), .B(n21943), .Y(n18126) );
  sky130_fd_sc_hd__o22ai_1 U24809 ( .A1(n18188), .A2(n18118), .B1(n18126), 
        .B2(n18185), .Y(n18132) );
  sky130_fd_sc_hd__nand2b_1 U24810 ( .A_N(n18470), .B(n21219), .Y(n18116) );
  sky130_fd_sc_hd__o22ai_1 U24811 ( .A1(n18209), .A2(n18116), .B1(n18115), 
        .B2(n18206), .Y(n18131) );
  sky130_fd_sc_hd__o22ai_1 U24812 ( .A1(n22365), .A2(n22318), .B1(n21849), 
        .B2(n11561), .Y(n18144) );
  sky130_fd_sc_hd__nor2b_1 U24813 ( .B_N(n18470), .A(n18205), .Y(n18122) );
  sky130_fd_sc_hd__xnor2_1 U24814 ( .A(n18363), .B(n21219), .Y(n18130) );
  sky130_fd_sc_hd__o22ai_1 U24815 ( .A1(n18209), .A2(n18117), .B1(n18130), 
        .B2(n18206), .Y(n18121) );
  sky130_fd_sc_hd__o22ai_1 U24816 ( .A1(n18188), .A2(n18119), .B1(n18118), 
        .B2(n18185), .Y(n18120) );
  sky130_fd_sc_hd__o22ai_1 U24817 ( .A1(n22365), .A2(n22279), .B1(n22245), 
        .B2(n18224), .Y(n18157) );
  sky130_fd_sc_hd__fah_1 U24818 ( .A(n18122), .B(n18121), .CI(n18120), .COUT(
        n18156), .SUM(n18143) );
  sky130_fd_sc_hd__fah_1 U24819 ( .A(n18125), .B(n18124), .CI(n18123), .COUT(
        n18159), .SUM(n18155) );
  sky130_fd_sc_hd__nor2_1 U24820 ( .A(n18153), .B(n18154), .Y(n22238) );
  sky130_fd_sc_hd__nor2b_1 U24821 ( .B_N(n18470), .A(n18209), .Y(n18135) );
  sky130_fd_sc_hd__xnor2_1 U24822 ( .A(n18363), .B(n21943), .Y(n18127) );
  sky130_fd_sc_hd__o22ai_1 U24823 ( .A1(n18188), .A2(n18126), .B1(n18127), 
        .B2(n18185), .Y(n18134) );
  sky130_fd_sc_hd__o22ai_1 U24824 ( .A1(n18188), .A2(n18127), .B1(n18210), 
        .B2(n18185), .Y(n18137) );
  sky130_fd_sc_hd__nand2b_1 U24825 ( .A_N(n18470), .B(n21943), .Y(n18128) );
  sky130_fd_sc_hd__nand2_1 U24826 ( .A(n18185), .B(n18128), .Y(n18136) );
  sky130_fd_sc_hd__xnor2_1 U24827 ( .A(n21219), .B(n18210), .Y(n18129) );
  sky130_fd_sc_hd__o22ai_1 U24828 ( .A1(n18209), .A2(n18130), .B1(n18129), 
        .B2(n18206), .Y(n18148) );
  sky130_fd_sc_hd__ha_1 U24829 ( .A(n18132), .B(n18131), .COUT(n18145), .SUM(
        n18147) );
  sky130_fd_sc_hd__o22ai_1 U24830 ( .A1(n22365), .A2(n22815), .B1(n21221), 
        .B2(n11561), .Y(n18146) );
  sky130_fd_sc_hd__o22ai_1 U24831 ( .A1(n22365), .A2(n22366), .B1(n19244), 
        .B2(n18536), .Y(n19239) );
  sky130_fd_sc_hd__fah_1 U24832 ( .A(n18135), .B(n18134), .CI(n18133), .COUT(
        n18141), .SUM(n19238) );
  sky130_fd_sc_hd__ha_1 U24833 ( .A(n18137), .B(n18136), .COUT(n18133), .SUM(
        n18139) );
  sky130_fd_sc_hd__o2bb2ai_1 U24834 ( .B1(n21942), .B2(n11561), .A1_N(n22979), 
        .A2_N(j202_soc_core_j22_cpu_ml_macl[17]), .Y(n18140) );
  sky130_fd_sc_hd__nor2_1 U24835 ( .A(n18139), .B(n18140), .Y(n18138) );
  sky130_fd_sc_hd__nor2b_1 U24837 ( .B_N(n18470), .A(n18188), .Y(n21704) );
  sky130_fd_sc_hd__nand2_1 U24838 ( .A(n21703), .B(n21704), .Y(n21705) );
  sky130_fd_sc_hd__nand2_1 U24839 ( .A(n18140), .B(n18139), .Y(n21938) );
  sky130_fd_sc_hd__nand2_1 U24840 ( .A(n19238), .B(n19239), .Y(n19240) );
  sky130_fd_sc_hd__nand2_1 U24841 ( .A(n18142), .B(n18141), .Y(n21215) );
  sky130_fd_sc_hd__o21ai_2 U24842 ( .A1(n21214), .A2(n21217), .B1(n21215), .Y(
        n21846) );
  sky130_fd_sc_hd__fah_1 U24843 ( .A(n18145), .B(n18144), .CI(n18143), .COUT(
        n18153), .SUM(n18152) );
  sky130_fd_sc_hd__fah_1 U24844 ( .A(n18148), .B(n18147), .CI(n18146), .COUT(
        n18151), .SUM(n18142) );
  sky130_fd_sc_hd__nand2_1 U24845 ( .A(n18150), .B(n18149), .Y(n21844) );
  sky130_fd_sc_hd__nand2_1 U24846 ( .A(n18152), .B(n18151), .Y(n21843) );
  sky130_fd_sc_hd__nand2_1 U24847 ( .A(n18154), .B(n18153), .Y(n22239) );
  sky130_fd_sc_hd__fah_1 U24848 ( .A(n18157), .B(n18156), .CI(n18155), .COUT(
        n18162), .SUM(n18154) );
  sky130_fd_sc_hd__fah_1 U24849 ( .A(n18160), .B(n18159), .CI(n18158), .COUT(
        n18164), .SUM(n18163) );
  sky130_fd_sc_hd__nor2_1 U24850 ( .A(n18162), .B(n18163), .Y(n18161) );
  sky130_fd_sc_hd__inv_1 U24851 ( .A(n18161), .Y(n22126) );
  sky130_fd_sc_hd__nand2_1 U24852 ( .A(n18163), .B(n18162), .Y(n22125) );
  sky130_fd_sc_hd__nand2_1 U24853 ( .A(n18165), .B(n18164), .Y(n18812) );
  sky130_fd_sc_hd__xnor2_1 U24855 ( .A(n18377), .B(n24366), .Y(n18203) );
  sky130_fd_sc_hd__o22ai_1 U24856 ( .A1(n18205), .A2(n18203), .B1(n18169), 
        .B2(n12048), .Y(n18216) );
  sky130_fd_sc_hd__xnor2_1 U24857 ( .A(n18372), .B(n27618), .Y(n18190) );
  sky130_fd_sc_hd__o22ai_1 U24858 ( .A1(n18192), .A2(n18190), .B1(n18170), 
        .B2(n18189), .Y(n18215) );
  sky130_fd_sc_hd__ha_1 U24859 ( .A(n18172), .B(n18171), .COUT(n18214), .SUM(
        n18175) );
  sky130_fd_sc_hd__fah_1 U24860 ( .A(n18178), .B(n18177), .CI(n18176), .COUT(
        n18198), .SUM(n18168) );
  sky130_fd_sc_hd__o22ai_1 U24861 ( .A1(n22365), .A2(n18179), .B1(n21733), 
        .B2(n18536), .Y(n18197) );
  sky130_fd_sc_hd__xnor2_1 U24862 ( .A(n18964), .B(n21943), .Y(n18186) );
  sky130_fd_sc_hd__o22ai_1 U24863 ( .A1(n18188), .A2(n18186), .B1(n18180), 
        .B2(n18185), .Y(n18200) );
  sky130_fd_sc_hd__xnor2_1 U24864 ( .A(n18367), .B(n21219), .Y(n18207) );
  sky130_fd_sc_hd__o22ai_1 U24865 ( .A1(n18209), .A2(n18207), .B1(n18181), 
        .B2(n18206), .Y(n18199) );
  sky130_fd_sc_hd__fah_1 U24866 ( .A(n18184), .B(n18183), .CI(n18182), .COUT(
        n18219), .SUM(n18218) );
  sky130_fd_sc_hd__o22ai_1 U24867 ( .A1(n18188), .A2(n18187), .B1(n18186), 
        .B2(n18185), .Y(n18238) );
  sky130_fd_sc_hd__o22ai_1 U24868 ( .A1(n18192), .A2(n18191), .B1(n18190), 
        .B2(n18189), .Y(n18223) );
  sky130_fd_sc_hd__nand2b_1 U24869 ( .A_N(n18470), .B(n24799), .Y(n18194) );
  sky130_fd_sc_hd__o22ai_1 U24870 ( .A1(n22365), .A2(n22889), .B1(n18195), 
        .B2(n18536), .Y(n18236) );
  sky130_fd_sc_hd__fah_1 U24871 ( .A(n18201), .B(n18200), .CI(n18199), .COUT(
        n18230), .SUM(n18196) );
  sky130_fd_sc_hd__o22ai_1 U24872 ( .A1(n18205), .A2(n18204), .B1(n18203), 
        .B2(n12048), .Y(n18227) );
  sky130_fd_sc_hd__o22ai_1 U24873 ( .A1(n18209), .A2(n18208), .B1(n18207), 
        .B2(n18206), .Y(n18226) );
  sky130_fd_sc_hd__xnor2_1 U24874 ( .A(n24799), .B(n18210), .Y(n18211) );
  sky130_fd_sc_hd__fah_1 U24875 ( .A(n18216), .B(n18215), .CI(n18214), .COUT(
        n18228), .SUM(n18184) );
  sky130_fd_sc_hd__nor2_1 U24876 ( .A(n22885), .B(n22880), .Y(n18222) );
  sky130_fd_sc_hd__nand2_1 U24877 ( .A(n18218), .B(n18217), .Y(n22883) );
  sky130_fd_sc_hd__nand2_1 U24878 ( .A(n18220), .B(n18219), .Y(n22881) );
  sky130_fd_sc_hd__o21ai_1 U24879 ( .A1(n22883), .A2(n22880), .B1(n22881), .Y(
        n18221) );
  sky130_fd_sc_hd__fah_1 U24880 ( .A(n18227), .B(n18226), .CI(n18225), .COUT(
        n18251), .SUM(n18229) );
  sky130_fd_sc_hd__fah_1 U24881 ( .A(n18230), .B(n18229), .CI(n18228), .COUT(
        n18257), .SUM(n18253) );
  sky130_fd_sc_hd__fah_1 U24882 ( .A(n18233), .B(n18232), .CI(n18231), .COUT(
        n18240), .SUM(n18244) );
  sky130_fd_sc_hd__fah_1 U24883 ( .A(n18238), .B(n18237), .CI(n18236), .COUT(
        n18242), .SUM(n18255) );
  sky130_fd_sc_hd__fah_1 U24884 ( .A(n18241), .B(n18240), .CI(n18239), .COUT(
        n18276), .SUM(n18268) );
  sky130_fd_sc_hd__fa_1 U24885 ( .A(n18247), .B(n18246), .CIN(n18245), .COUT(
        n18271), .SUM(n18274) );
  sky130_fd_sc_hd__fah_1 U24886 ( .A(n12117), .B(n18252), .CI(n18251), .COUT(
        n18272), .SUM(n18258) );
  sky130_fd_sc_hd__fah_1 U24887 ( .A(n18255), .B(n18254), .CI(n18253), .COUT(
        n18259), .SUM(n18220) );
  sky130_fd_sc_hd__fah_1 U24888 ( .A(n18258), .B(n18257), .CI(n18256), .COUT(
        n18261), .SUM(n18260) );
  sky130_fd_sc_hd__nand2_1 U24889 ( .A(n21286), .B(n13076), .Y(n18265) );
  sky130_fd_sc_hd__nand2_1 U24890 ( .A(n18260), .B(n18259), .Y(n19278) );
  sky130_fd_sc_hd__nand2_1 U24891 ( .A(n18262), .B(n18261), .Y(n21285) );
  sky130_fd_sc_hd__a21oi_1 U24892 ( .A1(n21286), .A2(n21283), .B1(n18263), .Y(
        n18264) );
  sky130_fd_sc_hd__fah_1 U24893 ( .A(n18271), .B(n18270), .CI(n18269), .COUT(
        n18088), .SUM(n18280) );
  sky130_fd_sc_hd__fah_1 U24894 ( .A(n18274), .B(n18273), .CI(n18272), .COUT(
        n18279), .SUM(n18266) );
  sky130_fd_sc_hd__fah_1 U24895 ( .A(n18280), .B(n18279), .CI(n18278), .COUT(
        n18286), .SUM(n18285) );
  sky130_fd_sc_hd__nand2_1 U24896 ( .A(n18285), .B(n18284), .Y(n22974) );
  sky130_fd_sc_hd__nand2_1 U24897 ( .A(n18287), .B(n18286), .Y(n22972) );
  sky130_fd_sc_hd__o21ai_1 U24898 ( .A1(n22974), .A2(n22971), .B1(n22972), .Y(
        n18288) );
  sky130_fd_sc_hd__nand2_1 U24899 ( .A(n18290), .B(n18289), .Y(n22566) );
  sky130_fd_sc_hd__nand2_1 U24900 ( .A(n18292), .B(n18291), .Y(n18883) );
  sky130_fd_sc_hd__o21a_1 U24901 ( .A1(n18293), .A2(n22566), .B1(n18883), .X(
        n18294) );
  sky130_fd_sc_hd__o21ai_2 U24902 ( .A1(n18295), .A2(n18881), .B1(n18294), .Y(
        n21684) );
  sky130_fd_sc_hd__fah_1 U24903 ( .A(n18298), .B(n18297), .CI(n18296), .COUT(
        n18314), .SUM(n18292) );
  sky130_fd_sc_hd__fah_1 U24905 ( .A(n18304), .B(n18303), .CI(n18302), .COUT(
        n18309), .SUM(n18296) );
  sky130_fd_sc_hd__nor2_1 U24907 ( .A(n18314), .B(n18315), .Y(n21974) );
  sky130_fd_sc_hd__fah_1 U24908 ( .A(n18310), .B(n18309), .CI(n18308), .COUT(
        n18316), .SUM(n18315) );
  sky130_fd_sc_hd__nor2_1 U24911 ( .A(n21974), .B(n21969), .Y(n18319) );
  sky130_fd_sc_hd__nand2_1 U24912 ( .A(n18315), .B(n18314), .Y(n21972) );
  sky130_fd_sc_hd__nand2_1 U24913 ( .A(n18317), .B(n18316), .Y(n21970) );
  sky130_fd_sc_hd__o21ai_1 U24914 ( .A1(n21972), .A2(n21969), .B1(n21970), .Y(
        n18318) );
  sky130_fd_sc_hd__a21oi_2 U24915 ( .A1(n21684), .A2(n18319), .B1(n18318), .Y(
        n19110) );
  sky130_fd_sc_hd__nand2_1 U24916 ( .A(n18321), .B(n18320), .Y(n21232) );
  sky130_fd_sc_hd__nand2_1 U24917 ( .A(n18323), .B(n18322), .Y(n21236) );
  sky130_fd_sc_hd__nand2_1 U24918 ( .A(n18325), .B(n18324), .Y(n22209) );
  sky130_fd_sc_hd__nand2_1 U24919 ( .A(n18327), .B(n18326), .Y(n22216) );
  sky130_fd_sc_hd__o21ai_1 U24920 ( .A1(n22209), .A2(n22215), .B1(n22216), .Y(
        n18328) );
  sky130_fd_sc_hd__a21oi_1 U24921 ( .A1(n21866), .A2(n18329), .B1(n18328), .Y(
        n18330) );
  sky130_fd_sc_hd__nor2_1 U24922 ( .A(n18333), .B(n18332), .Y(n22108) );
  sky130_fd_sc_hd__nor2_1 U24923 ( .A(n18683), .B(n22108), .Y(n22872) );
  sky130_fd_sc_hd__xnor2_1 U24924 ( .A(n18971), .B(n22299), .Y(n18383) );
  sky130_fd_sc_hd__xnor2_1 U24925 ( .A(n18941), .B(n22299), .Y(n18365) );
  sky130_fd_sc_hd__o22ai_1 U24926 ( .A1(n18533), .A2(n18383), .B1(n18365), 
        .B2(n18530), .Y(n18482) );
  sky130_fd_sc_hd__a21oi_1 U24927 ( .A1(j202_soc_core_j22_cpu_ml_mach[16]), 
        .A2(n25679), .B1(n13087), .Y(n18339) );
  sky130_fd_sc_hd__xnor2_1 U24929 ( .A(n22024), .B(n25761), .Y(n18345) );
  sky130_fd_sc_hd__xnor2_1 U24930 ( .A(n18925), .B(n25761), .Y(n18368) );
  sky130_fd_sc_hd__o22ai_1 U24931 ( .A1(n18486), .A2(n18345), .B1(n18368), 
        .B2(n18483), .Y(n18357) );
  sky130_fd_sc_hd__xnor2_1 U24932 ( .A(n18358), .B(n18357), .Y(n18480) );
  sky130_fd_sc_hd__xnor2_1 U24933 ( .A(n18966), .B(n22811), .Y(n18380) );
  sky130_fd_sc_hd__o22ai_1 U24934 ( .A1(n18496), .A2(n18341), .B1(n18380), 
        .B2(n17410), .Y(n18400) );
  sky130_fd_sc_hd__xnor2_1 U24935 ( .A(n18372), .B(n25777), .Y(n18376) );
  sky130_fd_sc_hd__o22ai_1 U24936 ( .A1(n18993), .A2(n18342), .B1(n18376), 
        .B2(n18990), .Y(n18399) );
  sky130_fd_sc_hd__nand2b_1 U24937 ( .A_N(n18470), .B(n22023), .Y(n18343) );
  sky130_fd_sc_hd__xnor2_1 U24938 ( .A(n18366), .B(n23571), .Y(n18401) );
  sky130_fd_sc_hd__xnor2_1 U24939 ( .A(n18367), .B(n23571), .Y(n18374) );
  sky130_fd_sc_hd__o22ai_1 U24940 ( .A1(n18989), .A2(n18401), .B1(n18374), 
        .B2(n12044), .Y(n18394) );
  sky130_fd_sc_hd__xnor2_1 U24941 ( .A(n18363), .B(n22023), .Y(n18344) );
  sky130_fd_sc_hd__nand2_1 U24942 ( .A(n18347), .B(n18346), .Y(n18348) );
  sky130_fd_sc_hd__nand2_1 U24943 ( .A(n18478), .B(n18348), .Y(n18350) );
  sky130_fd_sc_hd__nand2_1 U24944 ( .A(n18476), .B(n18477), .Y(n18349) );
  sky130_fd_sc_hd__nand2_1 U24945 ( .A(n18350), .B(n18349), .Y(n18514) );
  sky130_fd_sc_hd__fah_1 U24946 ( .A(n18353), .B(n18352), .CI(n18351), .COUT(
        n18389), .SUM(n18410) );
  sky130_fd_sc_hd__xnor2_1 U24947 ( .A(n18962), .B(n22087), .Y(n18381) );
  sky130_fd_sc_hd__o22ai_1 U24948 ( .A1(n18474), .A2(n18356), .B1(n18381), 
        .B2(n18471), .Y(n18362) );
  sky130_fd_sc_hd__a21oi_1 U24949 ( .A1(j202_soc_core_j22_cpu_ml_mach[17]), 
        .A2(n22940), .B1(n13087), .Y(n18359) );
  sky130_fd_sc_hd__o21ai_1 U24950 ( .A1(n18360), .A2(n11145), .B1(n18359), .Y(
        n18361) );
  sky130_fd_sc_hd__xnor2_1 U24951 ( .A(n18994), .B(n22811), .Y(n18379) );
  sky130_fd_sc_hd__xnor2_1 U24952 ( .A(n18971), .B(n22811), .Y(n18495) );
  sky130_fd_sc_hd__o22ai_1 U24953 ( .A1(n18496), .A2(n18379), .B1(n18495), 
        .B2(n17410), .Y(n18529) );
  sky130_fd_sc_hd__xnor2_1 U24954 ( .A(n18363), .B(n25777), .Y(n18375) );
  sky130_fd_sc_hd__xnor2_1 U24955 ( .A(n25777), .B(n18470), .Y(n18364) );
  sky130_fd_sc_hd__o22ai_1 U24956 ( .A1(n18993), .A2(n18375), .B1(n18364), 
        .B2(n18990), .Y(n18528) );
  sky130_fd_sc_hd__xnor2_1 U24957 ( .A(n22024), .B(n18887), .Y(n18491) );
  sky130_fd_sc_hd__a21o_1 U24958 ( .A1(n18489), .A2(n18492), .B1(n18491), .X(
        n18527) );
  sky130_fd_sc_hd__xnor2_1 U24959 ( .A(n18962), .B(n22299), .Y(n18532) );
  sky130_fd_sc_hd__xnor2_1 U24961 ( .A(n18387), .B(n23571), .Y(n18373) );
  sky130_fd_sc_hd__xnor2_1 U24962 ( .A(n18377), .B(n23571), .Y(n18498) );
  sky130_fd_sc_hd__o22ai_1 U24963 ( .A1(n18989), .A2(n18373), .B1(n18498), 
        .B2(n12044), .Y(n18502) );
  sky130_fd_sc_hd__xnor2_1 U24964 ( .A(n18366), .B(n23567), .Y(n18382) );
  sky130_fd_sc_hd__xnor2_1 U24965 ( .A(n18367), .B(n23567), .Y(n18500) );
  sky130_fd_sc_hd__xnor2_1 U24966 ( .A(n18966), .B(n25761), .Y(n18485) );
  sky130_fd_sc_hd__o22ai_1 U24967 ( .A1(n18486), .A2(n18368), .B1(n18485), 
        .B2(n18483), .Y(n18526) );
  sky130_fd_sc_hd__nand2b_1 U24968 ( .A_N(n18470), .B(n25777), .Y(n18370) );
  sky130_fd_sc_hd__o22ai_1 U24969 ( .A1(n18993), .A2(n18370), .B1(n13026), 
        .B2(n18990), .Y(n18525) );
  sky130_fd_sc_hd__xnor2_1 U24970 ( .A(n18371), .B(n25389), .Y(n18378) );
  sky130_fd_sc_hd__xnor2_1 U24971 ( .A(n18372), .B(n25389), .Y(n18488) );
  sky130_fd_sc_hd__o22ai_1 U24972 ( .A1(n19023), .A2(n18378), .B1(n18488), 
        .B2(n19020), .Y(n18524) );
  sky130_fd_sc_hd__o22ai_1 U24973 ( .A1(n18989), .A2(n18374), .B1(n18373), 
        .B2(n12044), .Y(n18468) );
  sky130_fd_sc_hd__xnor2_1 U24974 ( .A(n18377), .B(n25389), .Y(n18388) );
  sky130_fd_sc_hd__o22ai_1 U24975 ( .A1(n19023), .A2(n18388), .B1(n18378), 
        .B2(n19020), .Y(n18467) );
  sky130_fd_sc_hd__o22ai_1 U24976 ( .A1(n18496), .A2(n18380), .B1(n18379), 
        .B2(n17410), .Y(n18466) );
  sky130_fd_sc_hd__xnor2_1 U24977 ( .A(n18999), .B(n22087), .Y(n18469) );
  sky130_fd_sc_hd__o22ai_1 U24978 ( .A1(n18474), .A2(n18381), .B1(n18469), 
        .B2(n18471), .Y(n18465) );
  sky130_fd_sc_hd__xnor2_1 U24979 ( .A(n18964), .B(n23567), .Y(n18385) );
  sky130_fd_sc_hd__o22ai_1 U24980 ( .A1(n18533), .A2(n18384), .B1(n18383), 
        .B2(n18530), .Y(n18397) );
  sky130_fd_sc_hd__xnor2_1 U24981 ( .A(n18387), .B(n25389), .Y(n18403) );
  sky130_fd_sc_hd__o22ai_1 U24982 ( .A1(n19023), .A2(n18403), .B1(n18388), 
        .B2(n19020), .Y(n18395) );
  sky130_fd_sc_hd__fah_1 U24983 ( .A(n18394), .B(n18393), .CI(n18392), .COUT(
        n18428), .SUM(n18477) );
  sky130_fd_sc_hd__o22ai_1 U24984 ( .A1(n18989), .A2(n18402), .B1(n18401), 
        .B2(n12044), .Y(n18422) );
  sky130_fd_sc_hd__o22ai_1 U24985 ( .A1(n19023), .A2(n18404), .B1(n18403), 
        .B2(n19020), .Y(n18421) );
  sky130_fd_sc_hd__a21oi_1 U24986 ( .A1(j202_soc_core_j22_cpu_ml_mach[18]), 
        .A2(n22940), .B1(n13087), .Y(n18405) );
  sky130_fd_sc_hd__o21ai_1 U24987 ( .A1(n18406), .A2(n11145), .B1(n18405), .Y(
        n18420) );
  sky130_fd_sc_hd__xnor2_1 U24988 ( .A(n18442), .B(n18441), .Y(n18407) );
  sky130_fd_sc_hd__xnor2_1 U24989 ( .A(n18440), .B(n18407), .Y(n18518) );
  sky130_fd_sc_hd__fah_1 U24990 ( .A(n18410), .B(n18409), .CI(n18408), .COUT(
        n18433), .SUM(n18513) );
  sky130_fd_sc_hd__fah_1 U24991 ( .A(n18416), .B(n18415), .CI(n18414), .COUT(
        n17434), .SUM(n18435) );
  sky130_fd_sc_hd__fah_1 U24992 ( .A(n18422), .B(n18421), .CI(n18420), .COUT(
        n18441), .SUM(n18509) );
  sky130_fd_sc_hd__nand2_1 U24993 ( .A(n18511), .B(n18509), .Y(n18429) );
  sky130_fd_sc_hd__o21ai_1 U24994 ( .A1(n18520), .A2(n18518), .B1(n18517), .Y(
        n18431) );
  sky130_fd_sc_hd__nand2_1 U24995 ( .A(n18520), .B(n18518), .Y(n18430) );
  sky130_fd_sc_hd__nand2_1 U24996 ( .A(n18431), .B(n18430), .Y(n18663) );
  sky130_fd_sc_hd__fah_1 U24997 ( .A(n18436), .B(n18435), .CI(n18434), .COUT(
        n18462), .SUM(n18432) );
  sky130_fd_sc_hd__fa_1 U24998 ( .A(n18439), .B(n18438), .CIN(n18437), .COUT(
        n18454), .SUM(n18461) );
  sky130_fd_sc_hd__o21ai_1 U24999 ( .A1(n18442), .A2(n18441), .B1(n18440), .Y(
        n18444) );
  sky130_fd_sc_hd__nand2_1 U25000 ( .A(n18442), .B(n18441), .Y(n18443) );
  sky130_fd_sc_hd__nand2_1 U25001 ( .A(n18444), .B(n18443), .Y(n18460) );
  sky130_fd_sc_hd__o21ai_1 U25002 ( .A1(n18449), .A2(n18450), .B1(n18448), .Y(
        n18452) );
  sky130_fd_sc_hd__nand2_1 U25003 ( .A(n18450), .B(n18449), .Y(n18451) );
  sky130_fd_sc_hd__nand2_1 U25004 ( .A(n18452), .B(n18451), .Y(n18665) );
  sky130_fd_sc_hd__xnor2_1 U25005 ( .A(n18454), .B(n18453), .Y(n18455) );
  sky130_fd_sc_hd__xnor2_1 U25006 ( .A(n18456), .B(n18455), .Y(n18643) );
  sky130_fd_sc_hd__fa_1 U25007 ( .A(n18459), .B(n18458), .CIN(n18457), .COUT(
        n18647), .SUM(n18642) );
  sky130_fd_sc_hd__xnor2_1 U25010 ( .A(n18643), .B(n18463), .Y(n18666) );
  sky130_fd_sc_hd__xnor2_1 U25011 ( .A(n18964), .B(n22087), .Y(n18473) );
  sky130_fd_sc_hd__o22ai_1 U25012 ( .A1(n18474), .A2(n18469), .B1(n18473), 
        .B2(n18471), .Y(n18542) );
  sky130_fd_sc_hd__nor2b_1 U25013 ( .B_N(n18470), .A(n18993), .Y(n18535) );
  sky130_fd_sc_hd__o22ai_1 U25014 ( .A1(n24854), .A2(n19092), .B1(n18475), 
        .B2(n18536), .Y(n18540) );
  sky130_fd_sc_hd__xnor2_1 U25015 ( .A(n18477), .B(n18476), .Y(n18479) );
  sky130_fd_sc_hd__xnor2_1 U25016 ( .A(n18479), .B(n18478), .Y(n18556) );
  sky130_fd_sc_hd__fah_1 U25017 ( .A(n18482), .B(n18481), .CI(n18480), .COUT(
        n18478), .SUM(n18619) );
  sky130_fd_sc_hd__o22ai_1 U25018 ( .A1(n18486), .A2(n18485), .B1(n18484), 
        .B2(n18483), .Y(n18587) );
  sky130_fd_sc_hd__o22ai_1 U25019 ( .A1(n19023), .A2(n18488), .B1(n18487), 
        .B2(n19020), .Y(n18586) );
  sky130_fd_sc_hd__o22ai_1 U25020 ( .A1(n18492), .A2(n18491), .B1(n18490), 
        .B2(n18489), .Y(n18585) );
  sky130_fd_sc_hd__o22ai_1 U25021 ( .A1(n18496), .A2(n18495), .B1(n18494), 
        .B2(n17410), .Y(n18584) );
  sky130_fd_sc_hd__o22ai_1 U25022 ( .A1(n18989), .A2(n18498), .B1(n18497), 
        .B2(n12044), .Y(n18583) );
  sky130_fd_sc_hd__nand2_1 U25025 ( .A(n18623), .B(n18619), .Y(n18506) );
  sky130_fd_sc_hd__nand2_1 U25026 ( .A(n18507), .B(n18506), .Y(n18555) );
  sky130_fd_sc_hd__fah_1 U25029 ( .A(n18514), .B(n18513), .CI(n18512), .COUT(
        n18520), .SUM(n18560) );
  sky130_fd_sc_hd__o21ai_1 U25030 ( .A1(n18562), .A2(n18561), .B1(n18560), .Y(
        n18516) );
  sky130_fd_sc_hd__nand2_1 U25031 ( .A(n18562), .B(n18561), .Y(n18515) );
  sky130_fd_sc_hd__nand2_1 U25032 ( .A(n18516), .B(n18515), .Y(n18661) );
  sky130_fd_sc_hd__xnor2_1 U25033 ( .A(n18518), .B(n18517), .Y(n18519) );
  sky130_fd_sc_hd__xnor2_1 U25034 ( .A(n18520), .B(n18519), .Y(n18662) );
  sky130_fd_sc_hd__fah_1 U25035 ( .A(n18523), .B(n18522), .CI(n18521), .COUT(
        n18512), .SUM(n18630) );
  sky130_fd_sc_hd__fah_1 U25036 ( .A(n18526), .B(n18525), .CI(n18524), .COUT(
        n18504), .SUM(n18607) );
  sky130_fd_sc_hd__o22ai_1 U25037 ( .A1(n18533), .A2(n18532), .B1(n18531), 
        .B2(n18530), .Y(n18571) );
  sky130_fd_sc_hd__xnor2_1 U25038 ( .A(n18535), .B(n18534), .Y(n18570) );
  sky130_fd_sc_hd__o22ai_1 U25039 ( .A1(n24854), .A2(n24455), .B1(n22561), 
        .B2(n18536), .Y(n18569) );
  sky130_fd_sc_hd__fah_1 U25040 ( .A(n18539), .B(n18538), .CI(n18537), .COUT(
        n18557), .SUM(n18627) );
  sky130_fd_sc_hd__fah_1 U25041 ( .A(n18542), .B(n18541), .CI(n18540), .COUT(
        n18537), .SUM(n18601) );
  sky130_fd_sc_hd__fah_1 U25042 ( .A(n18545), .B(n18544), .CI(n18543), .COUT(
        n18623), .SUM(n18600) );
  sky130_fd_sc_hd__nand2_1 U25044 ( .A(n18632), .B(n18630), .Y(n18558) );
  sky130_fd_sc_hd__nand2_1 U25045 ( .A(n18559), .B(n18558), .Y(n18659) );
  sky130_fd_sc_hd__nor2_1 U25046 ( .A(n18659), .B(n18660), .Y(n19105) );
  sky130_fd_sc_hd__fah_1 U25047 ( .A(n18565), .B(n18564), .CI(n18563), .COUT(
        n18599), .SUM(n18608) );
  sky130_fd_sc_hd__fah_1 U25048 ( .A(n18568), .B(n18567), .CI(n18566), .COUT(
        n18610), .SUM(n18591) );
  sky130_fd_sc_hd__fah_1 U25049 ( .A(n18571), .B(n18570), .CI(n18569), .COUT(
        n18605), .SUM(n18609) );
  sky130_fd_sc_hd__xnor2_1 U25050 ( .A(n18610), .B(n18609), .Y(n18572) );
  sky130_fd_sc_hd__xnor2_1 U25051 ( .A(n18608), .B(n18572), .Y(n18618) );
  sky130_fd_sc_hd__nand2b_1 U25052 ( .A_N(n18577), .B(n18573), .Y(n18574) );
  sky130_fd_sc_hd__nand2_1 U25053 ( .A(n18577), .B(n18576), .Y(n18578) );
  sky130_fd_sc_hd__fah_1 U25054 ( .A(n18581), .B(n18580), .CI(n18579), .COUT(
        n18598), .SUM(n18577) );
  sky130_fd_sc_hd__fah_1 U25055 ( .A(n18587), .B(n18586), .CI(n18585), .COUT(
        n18545), .SUM(n18603) );
  sky130_fd_sc_hd__fah_1 U25056 ( .A(n18590), .B(n18589), .CI(n18588), .COUT(
        n18602), .SUM(n18592) );
  sky130_fd_sc_hd__nand2_1 U25057 ( .A(n18593), .B(n18592), .Y(n18594) );
  sky130_fd_sc_hd__nand2_1 U25058 ( .A(n18595), .B(n18594), .Y(n18596) );
  sky130_fd_sc_hd__fah_1 U25059 ( .A(n18598), .B(n18597), .CI(n18596), .COUT(
        n18635), .SUM(n18616) );
  sky130_fd_sc_hd__fah_1 U25060 ( .A(n18604), .B(n18603), .CI(n18602), .COUT(
        n18625), .SUM(n18597) );
  sky130_fd_sc_hd__fah_1 U25061 ( .A(n18607), .B(n18606), .CI(n18605), .COUT(
        n18628), .SUM(n18624) );
  sky130_fd_sc_hd__o21ai_1 U25062 ( .A1(n18610), .A2(n18609), .B1(n18608), .Y(
        n18612) );
  sky130_fd_sc_hd__nand2_1 U25063 ( .A(n18610), .B(n18609), .Y(n18611) );
  sky130_fd_sc_hd__xnor2_1 U25064 ( .A(n18634), .B(n18633), .Y(n18613) );
  sky130_fd_sc_hd__xnor2_1 U25065 ( .A(n18635), .B(n18613), .Y(n18652) );
  sky130_fd_sc_hd__nor2_2 U25066 ( .A(n18651), .B(n18652), .Y(n19087) );
  sky130_fd_sc_hd__fah_1 U25067 ( .A(n18618), .B(n18617), .CI(n18616), .COUT(
        n18651), .SUM(n18650) );
  sky130_fd_sc_hd__nor2_1 U25068 ( .A(n18649), .B(n18650), .Y(n22562) );
  sky130_fd_sc_hd__xnor2_1 U25069 ( .A(n18621), .B(n18620), .Y(n18622) );
  sky130_fd_sc_hd__xor2_1 U25070 ( .A(n18623), .B(n18622), .X(n18640) );
  sky130_fd_sc_hd__fah_1 U25071 ( .A(n18628), .B(n18627), .CI(n18626), .COUT(
        n18632), .SUM(n18638) );
  sky130_fd_sc_hd__xnor2_1 U25072 ( .A(n18630), .B(n18629), .Y(n18631) );
  sky130_fd_sc_hd__xnor2_1 U25073 ( .A(n18632), .B(n18631), .Y(n18656) );
  sky130_fd_sc_hd__o21ai_1 U25074 ( .A1(n18634), .A2(n18635), .B1(n18633), .Y(
        n18637) );
  sky130_fd_sc_hd__nand2_1 U25075 ( .A(n18635), .B(n18634), .Y(n18636) );
  sky130_fd_sc_hd__nand2_1 U25076 ( .A(n18637), .B(n18636), .Y(n18653) );
  sky130_fd_sc_hd__fah_1 U25077 ( .A(n18640), .B(n18639), .CI(n18638), .COUT(
        n18655), .SUM(n18654) );
  sky130_fd_sc_hd__nor2_1 U25078 ( .A(n18653), .B(n18654), .Y(n21681) );
  sky130_fd_sc_hd__o21ai_1 U25079 ( .A1(n18643), .A2(n18642), .B1(n18641), .Y(
        n18645) );
  sky130_fd_sc_hd__nand2_1 U25080 ( .A(n18643), .B(n18642), .Y(n18644) );
  sky130_fd_sc_hd__nand2_1 U25081 ( .A(n18645), .B(n18644), .Y(n18672) );
  sky130_fd_sc_hd__xnor2_1 U25082 ( .A(n18647), .B(n18646), .Y(n18648) );
  sky130_fd_sc_hd__xnor2_1 U25083 ( .A(n13059), .B(n18648), .Y(n18673) );
  sky130_fd_sc_hd__nand2_1 U25084 ( .A(n23030), .B(n13086), .Y(n18675) );
  sky130_fd_sc_hd__nand2_1 U25085 ( .A(n18650), .B(n18649), .Y(n22563) );
  sky130_fd_sc_hd__nand2_1 U25086 ( .A(n18652), .B(n18651), .Y(n19088) );
  sky130_fd_sc_hd__nand2_1 U25087 ( .A(n18654), .B(n18653), .Y(n21961) );
  sky130_fd_sc_hd__nand2_1 U25088 ( .A(n18656), .B(n18655), .Y(n21958) );
  sky130_fd_sc_hd__nand2_1 U25090 ( .A(n18662), .B(n18661), .Y(n21190) );
  sky130_fd_sc_hd__nand2_1 U25091 ( .A(n18664), .B(n18663), .Y(n22197) );
  sky130_fd_sc_hd__nand2_1 U25092 ( .A(n18666), .B(n18665), .Y(n22191) );
  sky130_fd_sc_hd__o21ai_1 U25093 ( .A1(n22197), .A2(n22190), .B1(n22191), .Y(
        n18667) );
  sky130_fd_sc_hd__a21oi_1 U25094 ( .A1(n18668), .A2(n22196), .B1(n18667), .Y(
        n18669) );
  sky130_fd_sc_hd__buf_6 U25095 ( .A(n18671), .X(n23036) );
  sky130_fd_sc_hd__nand2_1 U25096 ( .A(n18673), .B(n18672), .Y(n22105) );
  sky130_fd_sc_hd__o21ai_2 U25097 ( .A1(n12349), .A2(n18675), .B1(n18674), .Y(
        n18676) );
  sky130_fd_sc_hd__xnor2_2 U25098 ( .A(n18677), .B(n18676), .Y(n23478) );
  sky130_fd_sc_hd__nand2_1 U25099 ( .A(n18681), .B(n18680), .Y(n18682) );
  sky130_fd_sc_hd__nand2_1 U25100 ( .A(n28045), .B(n18682), .Y(n24852) );
  sky130_fd_sc_hd__nand2_1 U25101 ( .A(n18685), .B(n18684), .Y(n18688) );
  sky130_fd_sc_hd__o21ai_0 U25102 ( .A1(n22108), .A2(n22967), .B1(n22109), .Y(
        n18687) );
  sky130_fd_sc_hd__xnor2_1 U25103 ( .A(n18688), .B(n18687), .Y(n22083) );
  sky130_fd_sc_hd__nand2_1 U25104 ( .A(n22083), .B(n25679), .Y(n22381) );
  sky130_fd_sc_hd__nand2_1 U25105 ( .A(j202_soc_core_j22_cpu_ma_M_address[0]), 
        .B(j202_soc_core_j22_cpu_ma_M_MEM[1]), .Y(n18794) );
  sky130_fd_sc_hd__nor2_1 U25106 ( .A(n23511), .B(n18794), .Y(n23506) );
  sky130_fd_sc_hd__nor2_1 U25107 ( .A(j202_soc_core_j22_cpu_ma_M_address[0]), 
        .B(n18689), .Y(n23502) );
  sky130_fd_sc_hd__nand2b_1 U25108 ( .A_N(n21515), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[47]), .Y(n18786) );
  sky130_fd_sc_hd__nand2_1 U25109 ( .A(n18786), .B(n21768), .Y(n18693) );
  sky130_fd_sc_hd__nand2_1 U25110 ( .A(n20759), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[79]), .Y(n18692) );
  sky130_fd_sc_hd__nand2_1 U25111 ( .A(n21446), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[111]), .Y(n18691) );
  sky130_fd_sc_hd__nand2_1 U25112 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[15]), .Y(n18690) );
  sky130_fd_sc_hd__nand3_1 U25113 ( .A(n18692), .B(n18691), .C(n18690), .Y(
        n18785) );
  sky130_fd_sc_hd__nor2_1 U25114 ( .A(n18693), .B(n18785), .Y(n18784) );
  sky130_fd_sc_hd__nand2b_1 U25115 ( .A_N(n20058), .B(n18744), .Y(n20167) );
  sky130_fd_sc_hd__nor2_1 U25116 ( .A(n18711), .B(n18694), .Y(n19904) );
  sky130_fd_sc_hd__nand2_1 U25117 ( .A(n19904), .B(n21101), .Y(n20215) );
  sky130_fd_sc_hd__nand2_1 U25118 ( .A(n20167), .B(n20215), .Y(n20037) );
  sky130_fd_sc_hd__nand2_1 U25119 ( .A(n20199), .B(n18752), .Y(n19876) );
  sky130_fd_sc_hd__nand2_1 U25120 ( .A(n19865), .B(n18695), .Y(n18696) );
  sky130_fd_sc_hd__nand2b_1 U25121 ( .A_N(n18696), .B(n21104), .Y(n20113) );
  sky130_fd_sc_hd__nand2_1 U25122 ( .A(n19876), .B(n20113), .Y(n20024) );
  sky130_fd_sc_hd__nand2b_1 U25123 ( .A_N(n20034), .B(n13179), .Y(n20137) );
  sky130_fd_sc_hd__nor2_1 U25124 ( .A(n18697), .B(n18696), .Y(n20100) );
  sky130_fd_sc_hd__nand2_1 U25125 ( .A(n18753), .B(n21359), .Y(n20129) );
  sky130_fd_sc_hd__nand2_1 U25126 ( .A(n20152), .B(n20129), .Y(n20213) );
  sky130_fd_sc_hd__nor2_1 U25127 ( .A(n18768), .B(n20213), .Y(n18701) );
  sky130_fd_sc_hd__nor2_1 U25128 ( .A(n18731), .B(n20034), .Y(n20060) );
  sky130_fd_sc_hd__nor2_1 U25129 ( .A(n18764), .B(n18731), .Y(n18743) );
  sky130_fd_sc_hd__nor2_1 U25130 ( .A(n18698), .B(n18699), .Y(n20055) );
  sky130_fd_sc_hd__nor2_1 U25131 ( .A(n20060), .B(n20055), .Y(n20014) );
  sky130_fd_sc_hd__nand2_1 U25132 ( .A(n18716), .B(n18744), .Y(n20128) );
  sky130_fd_sc_hd__nor2_1 U25133 ( .A(n18700), .B(n18699), .Y(n20029) );
  sky130_fd_sc_hd__nand2_1 U25134 ( .A(n20029), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n20102) );
  sky130_fd_sc_hd__nand4_1 U25135 ( .A(n18701), .B(n20014), .C(n20128), .D(
        n20102), .Y(n18702) );
  sky130_fd_sc_hd__nor3_1 U25136 ( .A(n20037), .B(n20024), .C(n18702), .Y(
        n18721) );
  sky130_fd_sc_hd__nor2_1 U25137 ( .A(n21088), .B(n19119), .Y(n20225) );
  sky130_fd_sc_hd__nand2b_1 U25138 ( .A_N(n21097), .B(n19140), .Y(n20023) );
  sky130_fd_sc_hd__nor2_1 U25139 ( .A(n20213), .B(n18728), .Y(n20162) );
  sky130_fd_sc_hd__nand3_1 U25140 ( .A(n18715), .B(n19140), .C(n18763), .Y(
        n20138) );
  sky130_fd_sc_hd__nand2_1 U25141 ( .A(n18703), .B(n18752), .Y(n19951) );
  sky130_fd_sc_hd__nand2_1 U25142 ( .A(n20138), .B(n19951), .Y(n20036) );
  sky130_fd_sc_hd__nor2_1 U25143 ( .A(n18730), .B(n18704), .Y(n20013) );
  sky130_fd_sc_hd__nand4_1 U25144 ( .A(n20162), .B(n20118), .C(n20052), .D(
        n19876), .Y(n18710) );
  sky130_fd_sc_hd__nor2_1 U25145 ( .A(n21088), .B(
        j202_soc_core_bootrom_00_address_w[4]), .Y(n20227) );
  sky130_fd_sc_hd__nor2_1 U25146 ( .A(n18764), .B(n21101), .Y(n18705) );
  sky130_fd_sc_hd__nand3_1 U25147 ( .A(n18706), .B(n21075), .C(n18705), .Y(
        n19949) );
  sky130_fd_sc_hd__nand2b_1 U25148 ( .A_N(n20034), .B(n18752), .Y(n20182) );
  sky130_fd_sc_hd__nor2_1 U25149 ( .A(n18741), .B(n18723), .Y(n19965) );
  sky130_fd_sc_hd__nor2_1 U25150 ( .A(n18713), .B(n18707), .Y(n19981) );
  sky130_fd_sc_hd__nand2_1 U25151 ( .A(n19981), .B(n21101), .Y(n20216) );
  sky130_fd_sc_hd__nand3_1 U25152 ( .A(n18742), .B(n21359), .C(n18712), .Y(
        n18708) );
  sky130_fd_sc_hd__nand3_1 U25153 ( .A(n19965), .B(n20216), .C(n18708), .Y(
        n18709) );
  sky130_fd_sc_hd__nor2_1 U25154 ( .A(n20024), .B(n18709), .Y(n20008) );
  sky130_fd_sc_hd__a2bb2oi_1 U25155 ( .B1(n20210), .B2(n18710), .A1_N(n20038), 
        .A2_N(n20008), .Y(n18719) );
  sky130_fd_sc_hd__nand2_1 U25156 ( .A(n20199), .B(n18724), .Y(n20047) );
  sky130_fd_sc_hd__nor2_1 U25157 ( .A(n18711), .B(n20034), .Y(n20046) );
  sky130_fd_sc_hd__nand3_1 U25158 ( .A(n20148), .B(n20047), .C(n19895), .Y(
        n18717) );
  sky130_fd_sc_hd__nand2_1 U25159 ( .A(n21075), .B(n18712), .Y(n20044) );
  sky130_fd_sc_hd__nor2_1 U25160 ( .A(n18713), .B(n20044), .Y(n19874) );
  sky130_fd_sc_hd__nand2_1 U25161 ( .A(n19874), .B(n21101), .Y(n20173) );
  sky130_fd_sc_hd__nand2_1 U25162 ( .A(n19866), .B(n19865), .Y(n20001) );
  sky130_fd_sc_hd__nand2b_1 U25163 ( .A_N(n20001), .B(n13179), .Y(n19937) );
  sky130_fd_sc_hd__nand2_1 U25164 ( .A(n19937), .B(n20052), .Y(n20146) );
  sky130_fd_sc_hd__nor2_1 U25165 ( .A(n18714), .B(n20146), .Y(n19996) );
  sky130_fd_sc_hd__nand2_1 U25166 ( .A(n18715), .B(n18752), .Y(n19942) );
  sky130_fd_sc_hd__nor2_1 U25167 ( .A(n18744), .B(n19942), .Y(n19956) );
  sky130_fd_sc_hd__nand2_1 U25168 ( .A(n18716), .B(n19140), .Y(n20183) );
  sky130_fd_sc_hd__nand3_1 U25169 ( .A(n19996), .B(n20006), .C(n20183), .Y(
        n20212) );
  sky130_fd_sc_hd__o21ai_1 U25170 ( .A1(n18717), .A2(n20212), .B1(n20179), .Y(
        n18718) );
  sky130_fd_sc_hd__o211ai_1 U25171 ( .A1(n18721), .A2(n18720), .B1(n18719), 
        .C1(n18718), .Y(n18722) );
  sky130_fd_sc_hd__nand2_1 U25172 ( .A(n18722), .B(n20126), .Y(n18782) );
  sky130_fd_sc_hd__nor2_1 U25173 ( .A(n20060), .B(n18723), .Y(n20205) );
  sky130_fd_sc_hd__nand2_1 U25174 ( .A(n20199), .B(n21075), .Y(n20153) );
  sky130_fd_sc_hd__nand2_1 U25175 ( .A(n20205), .B(n20153), .Y(n19993) );
  sky130_fd_sc_hd__nor2_1 U25176 ( .A(n20037), .B(n19993), .Y(n18726) );
  sky130_fd_sc_hd__nor2_1 U25177 ( .A(n18725), .B(n20034), .Y(n18755) );
  sky130_fd_sc_hd__nand2_1 U25178 ( .A(n19999), .B(n21097), .Y(n20175) );
  sky130_fd_sc_hd__nand3_1 U25179 ( .A(n18743), .B(n11150), .C(n21101), .Y(
        n19966) );
  sky130_fd_sc_hd__nand4_1 U25180 ( .A(n18726), .B(n20130), .C(n19966), .D(
        n19937), .Y(n18739) );
  sky130_fd_sc_hd__nand2_1 U25181 ( .A(n18743), .B(n18727), .Y(n20002) );
  sky130_fd_sc_hd__nor2_1 U25182 ( .A(n18729), .B(n18728), .Y(n20187) );
  sky130_fd_sc_hd__nand2_1 U25183 ( .A(n20199), .B(n18730), .Y(n19971) );
  sky130_fd_sc_hd__nand2b_1 U25184 ( .A_N(n19971), .B(n18731), .Y(n19905) );
  sky130_fd_sc_hd__a31oi_1 U25185 ( .A1(n20187), .A2(n20006), .A3(n19905), 
        .B1(n20200), .Y(n18738) );
  sky130_fd_sc_hd__nand2_1 U25186 ( .A(n20023), .B(n19966), .Y(n18732) );
  sky130_fd_sc_hd__nand3_1 U25187 ( .A(n20167), .B(n20173), .C(n19895), .Y(
        n19881) );
  sky130_fd_sc_hd__nor2_1 U25188 ( .A(n18732), .B(n19881), .Y(n20223) );
  sky130_fd_sc_hd__nor2_1 U25189 ( .A(n20046), .B(n20055), .Y(n18733) );
  sky130_fd_sc_hd__nand4_1 U25190 ( .A(n18733), .B(n20216), .C(n20173), .D(
        n19876), .Y(n18735) );
  sky130_fd_sc_hd__nand2_1 U25191 ( .A(n20205), .B(n20023), .Y(n18734) );
  sky130_fd_sc_hd__o21ai_1 U25193 ( .A1(n19910), .A2(n20223), .B1(n18736), .Y(
        n18737) );
  sky130_fd_sc_hd__a211o_1 U25194 ( .A1(n18739), .A2(n20227), .B1(n18738), 
        .C1(n18737), .X(n18740) );
  sky130_fd_sc_hd__nand2_1 U25195 ( .A(n18740), .B(n20196), .Y(n18781) );
  sky130_fd_sc_hd__nor2_1 U25196 ( .A(n18741), .B(n20100), .Y(n20020) );
  sky130_fd_sc_hd__nand2_1 U25197 ( .A(n18743), .B(n18742), .Y(n21121) );
  sky130_fd_sc_hd__nand2b_1 U25198 ( .A_N(n21121), .B(n18744), .Y(n20139) );
  sky130_fd_sc_hd__nand3_1 U25199 ( .A(n20020), .B(n20139), .C(n20023), .Y(
        n19970) );
  sky130_fd_sc_hd__nand2_1 U25200 ( .A(n20216), .B(n20137), .Y(n19976) );
  sky130_fd_sc_hd__nor2_1 U25201 ( .A(n18744), .B(n21121), .Y(n19903) );
  sky130_fd_sc_hd__nor2_1 U25202 ( .A(n18745), .B(n19903), .Y(n19935) );
  sky130_fd_sc_hd__nand2b_1 U25203 ( .A_N(n19976), .B(n19935), .Y(n18746) );
  sky130_fd_sc_hd__nand3_1 U25205 ( .A(n19937), .B(n20215), .C(n19895), .Y(
        n20132) );
  sky130_fd_sc_hd__nand2_1 U25206 ( .A(n20172), .B(n20113), .Y(n20015) );
  sky130_fd_sc_hd__nor3_1 U25207 ( .A(n18755), .B(n20100), .C(n20036), .Y(
        n18747) );
  sky130_fd_sc_hd__nand3b_1 U25208 ( .A_N(n20132), .B(n19889), .C(n18747), .Y(
        n18748) );
  sky130_fd_sc_hd__nand2_1 U25209 ( .A(n18748), .B(n20227), .Y(n18760) );
  sky130_fd_sc_hd__nand2b_1 U25210 ( .A_N(n20058), .B(n19140), .Y(n20214) );
  sky130_fd_sc_hd__nand3_1 U25211 ( .A(n20167), .B(n20214), .C(n19897), .Y(
        n18770) );
  sky130_fd_sc_hd__nand2_1 U25212 ( .A(n19874), .B(n21145), .Y(n20000) );
  sky130_fd_sc_hd__nand2_1 U25213 ( .A(n20000), .B(n20129), .Y(n18749) );
  sky130_fd_sc_hd__nor2_1 U25214 ( .A(n19946), .B(n18768), .Y(n19877) );
  sky130_fd_sc_hd__nand4b_1 U25215 ( .A_N(n18749), .B(n19877), .C(n20139), .D(
        n19937), .Y(n18750) );
  sky130_fd_sc_hd__o21ai_1 U25216 ( .A1(n18770), .A2(n18750), .B1(n20179), .Y(
        n18759) );
  sky130_fd_sc_hd__nand2_1 U25217 ( .A(n18751), .B(n18763), .Y(n20181) );
  sky130_fd_sc_hd__nand2_1 U25218 ( .A(n18753), .B(n18752), .Y(n20033) );
  sky130_fd_sc_hd__and3_1 U25219 ( .A(n20033), .B(n19951), .C(n21121), .X(
        n18754) );
  sky130_fd_sc_hd__nand3_1 U25220 ( .A(n20181), .B(n18754), .C(n20172), .Y(
        n18757) );
  sky130_fd_sc_hd__nor2_1 U25221 ( .A(n18755), .B(n20046), .Y(n18756) );
  sky130_fd_sc_hd__nand4_1 U25222 ( .A(n18756), .B(n20216), .C(n19876), .D(
        n20167), .Y(n20206) );
  sky130_fd_sc_hd__nand4_1 U25224 ( .A(n18761), .B(n18760), .C(n18759), .D(
        n18758), .Y(n18762) );
  sky130_fd_sc_hd__nand2_1 U25225 ( .A(n18762), .B(n20235), .Y(n18780) );
  sky130_fd_sc_hd__nand3_1 U25226 ( .A(n19866), .B(n18764), .C(n18763), .Y(
        n20103) );
  sky130_fd_sc_hd__nand2_1 U25227 ( .A(n20216), .B(n20103), .Y(n19943) );
  sky130_fd_sc_hd__nand4_1 U25228 ( .A(n19892), .B(n18765), .C(n19877), .D(
        n20167), .Y(n18767) );
  sky130_fd_sc_hd__nand3_1 U25229 ( .A(n20173), .B(n20216), .C(n20182), .Y(
        n18766) );
  sky130_fd_sc_hd__nand2_1 U25230 ( .A(n19876), .B(n20103), .Y(n20056) );
  sky130_fd_sc_hd__nor2_1 U25231 ( .A(n18766), .B(n20056), .Y(n20115) );
  sky130_fd_sc_hd__a2bb2oi_1 U25232 ( .B1(n20210), .B2(n18767), .A1_N(n20200), 
        .A2_N(n20115), .Y(n18777) );
  sky130_fd_sc_hd__nor2_1 U25233 ( .A(n20100), .B(n18768), .Y(n19891) );
  sky130_fd_sc_hd__nand3_1 U25234 ( .A(n19891), .B(n19889), .C(n20128), .Y(
        n18769) );
  sky130_fd_sc_hd__nor2_1 U25235 ( .A(n18770), .B(n18769), .Y(n18771) );
  sky130_fd_sc_hd__nand2_1 U25236 ( .A(n18771), .B(n19996), .Y(n18772) );
  sky130_fd_sc_hd__nand2_1 U25237 ( .A(n18772), .B(n20227), .Y(n18776) );
  sky130_fd_sc_hd__nor2_1 U25238 ( .A(n18773), .B(n19956), .Y(n20186) );
  sky130_fd_sc_hd__nand2_1 U25239 ( .A(n20216), .B(n19951), .Y(n19879) );
  sky130_fd_sc_hd__nand4_1 U25240 ( .A(n20186), .B(n19959), .C(n20130), .D(
        n20182), .Y(n18774) );
  sky130_fd_sc_hd__nand2_1 U25241 ( .A(n18774), .B(n20225), .Y(n18775) );
  sky130_fd_sc_hd__nand3_1 U25242 ( .A(n18777), .B(n18776), .C(n18775), .Y(
        n18778) );
  sky130_fd_sc_hd__nand2_1 U25243 ( .A(n18778), .B(n20194), .Y(n18779) );
  sky130_fd_sc_hd__nand4_1 U25244 ( .A(n18782), .B(n18781), .C(n18780), .D(
        n18779), .Y(n18783) );
  sky130_fd_sc_hd__nand2_1 U25245 ( .A(n18783), .B(n21629), .Y(n18791) );
  sky130_fd_sc_hd__nand2_1 U25246 ( .A(n20786), .B(
        j202_soc_core_bldc_core_00_pwm_duty[3]), .Y(n18788) );
  sky130_fd_sc_hd__nand2_1 U25247 ( .A(j202_soc_core_memory0_ram_dout0[495]), 
        .B(n21650), .Y(n18793) );
  sky130_fd_sc_hd__nand3_1 U25248 ( .A(n18787), .B(n21653), .C(n18786), .Y(
        n18790) );
  sky130_fd_sc_hd__nor2_1 U25249 ( .A(n18790), .B(n18789), .Y(n18792) );
  sky130_fd_sc_hd__nand2_1 U25250 ( .A(n18795), .B(n23511), .Y(n19235) );
  sky130_fd_sc_hd__nor2_1 U25251 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[0]), .B(
        n23511), .Y(n18798) );
  sky130_fd_sc_hd__nor2_1 U25252 ( .A(n18798), .B(n26189), .Y(n25940) );
  sky130_fd_sc_hd__nand2_1 U25253 ( .A(n18799), .B(n23511), .Y(n24069) );
  sky130_fd_sc_hd__nand2_1 U25254 ( .A(n10971), .B(n25938), .Y(n18800) );
  sky130_fd_sc_hd__nand3_1 U25255 ( .A(n26345), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .C(n26142), .Y(n25263) );
  sky130_fd_sc_hd__nand2_1 U25256 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[0]), .Y(n26264) );
  sky130_fd_sc_hd__nand2_1 U25257 ( .A(n25263), .B(n26264), .Y(n25830) );
  sky130_fd_sc_hd__nand2_1 U25258 ( .A(n26208), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n18802) );
  sky130_fd_sc_hd__nand2_1 U25259 ( .A(n18802), .B(n26341), .Y(n18804) );
  sky130_fd_sc_hd__mux2i_1 U25260 ( .A0(j202_soc_core_j22_cpu_exuop_EXU_[5]), 
        .A1(j202_soc_core_j22_cpu_exuop_EXU_[3]), .S(
        j202_soc_core_j22_cpu_exuop_EXU_[0]), .Y(n18803) );
  sky130_fd_sc_hd__nand2_1 U25261 ( .A(n18804), .B(n18803), .Y(n18818) );
  sky130_fd_sc_hd__nand2b_1 U25262 ( .A_N(n26208), .B(n22117), .Y(n18805) );
  sky130_fd_sc_hd__nand2_1 U25263 ( .A(n26295), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[5]), .Y(n26340) );
  sky130_fd_sc_hd__nand2_1 U25264 ( .A(n24879), .B(n25263), .Y(n18808) );
  sky130_fd_sc_hd__nand2_1 U25265 ( .A(n18808), .B(n27786), .Y(n18811) );
  sky130_fd_sc_hd__nand3_1 U25266 ( .A(n26426), .B(n26295), .C(n18809), .Y(
        n25397) );
  sky130_fd_sc_hd__nand2_1 U25267 ( .A(n24879), .B(n27785), .Y(n18810) );
  sky130_fd_sc_hd__nand2_1 U25268 ( .A(n18811), .B(n18810), .Y(n18853) );
  sky130_fd_sc_hd__nand2_1 U25269 ( .A(n12141), .B(n18812), .Y(n18813) );
  sky130_fd_sc_hd__xor2_1 U25270 ( .A(n18814), .B(n18813), .X(n24324) );
  sky130_fd_sc_hd__nand2_1 U25271 ( .A(n24324), .B(n24461), .Y(n22387) );
  sky130_fd_sc_hd__nand2_1 U25272 ( .A(n18816), .B(n22751), .Y(n18817) );
  sky130_fd_sc_hd__xor2_1 U25273 ( .A(n22752), .B(n18817), .X(n24086) );
  sky130_fd_sc_hd__nor2_1 U25274 ( .A(n26340), .B(n28541), .Y(n25999) );
  sky130_fd_sc_hd__nand2_1 U25275 ( .A(n26937), .B(n28515), .Y(n18819) );
  sky130_fd_sc_hd__nand2_1 U25276 ( .A(n25999), .B(n18819), .Y(n27795) );
  sky130_fd_sc_hd__nand2_1 U25277 ( .A(n28541), .B(n26419), .Y(n18844) );
  sky130_fd_sc_hd__nand2b_1 U25278 ( .A_N(n18844), .B(n28509), .Y(n26943) );
  sky130_fd_sc_hd__o22ai_1 U25279 ( .A1(n11191), .A2(n27795), .B1(n26430), 
        .B2(n26943), .Y(n18824) );
  sky130_fd_sc_hd__nand2b_1 U25280 ( .A_N(n18844), .B(n18819), .Y(n27803) );
  sky130_fd_sc_hd__nand2_1 U25281 ( .A(n28515), .B(n28502), .Y(n23523) );
  sky130_fd_sc_hd__nand2_1 U25282 ( .A(n18821), .B(n18820), .Y(n25996) );
  sky130_fd_sc_hd__o22ai_1 U25283 ( .A1(n26317), .A2(n27803), .B1(n26431), 
        .B2(n25996), .Y(n18823) );
  sky130_fd_sc_hd__nand2_1 U25284 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[5]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[3]), .Y(n26268) );
  sky130_fd_sc_hd__nor2_1 U25285 ( .A(n26268), .B(n26377), .Y(n23520) );
  sky130_fd_sc_hd__nand2_1 U25286 ( .A(n23520), .B(n27147), .Y(n23531) );
  sky130_fd_sc_hd__nand2b_1 U25287 ( .A_N(n23531), .B(n26426), .Y(n26936) );
  sky130_fd_sc_hd__nand2_1 U25288 ( .A(n26377), .B(n18828), .Y(n26425) );
  sky130_fd_sc_hd__nand2_1 U25289 ( .A(n27147), .B(n26284), .Y(n26332) );
  sky130_fd_sc_hd__nor2_1 U25290 ( .A(n26425), .B(n26332), .Y(n23533) );
  sky130_fd_sc_hd__nand2_1 U25291 ( .A(n23533), .B(n26426), .Y(n26932) );
  sky130_fd_sc_hd__o22ai_1 U25292 ( .A1(n26311), .A2(n26936), .B1(n28487), 
        .B2(n26932), .Y(n18822) );
  sky130_fd_sc_hd__nor3_1 U25293 ( .A(n18824), .B(n18823), .C(n18822), .Y(
        n18849) );
  sky130_fd_sc_hd__nand2b_1 U25294 ( .A_N(n26048), .B(n18825), .Y(n27793) );
  sky130_fd_sc_hd__nand2_1 U25295 ( .A(n26375), .B(n26377), .Y(n23519) );
  sky130_fd_sc_hd__nand2_1 U25296 ( .A(n23519), .B(n27147), .Y(n18829) );
  sky130_fd_sc_hd__nand2_1 U25297 ( .A(n18826), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[1]), .Y(n26144) );
  sky130_fd_sc_hd__nand2_1 U25298 ( .A(n26144), .B(n18827), .Y(n23530) );
  sky130_fd_sc_hd__a21oi_1 U25299 ( .A1(n18829), .A2(n18828), .B1(n23530), .Y(
        n21210) );
  sky130_fd_sc_hd__nand2b_1 U25300 ( .A_N(n21210), .B(n26426), .Y(n22251) );
  sky130_fd_sc_hd__mux2_2 U25301 ( .A0(n27793), .A1(n22251), .S(n28489), .X(
        n18848) );
  sky130_fd_sc_hd__nand2_1 U25302 ( .A(n26149), .B(n28104), .Y(n21206) );
  sky130_fd_sc_hd__nor2_1 U25303 ( .A(n26144), .B(n26048), .Y(n25109) );
  sky130_fd_sc_hd__a21oi_1 U25304 ( .A1(n28489), .A2(n27791), .B1(n25109), .Y(
        n18843) );
  sky130_fd_sc_hd__nand2_1 U25306 ( .A(n24677), .B(n18831), .Y(n18833) );
  sky130_fd_sc_hd__nand2_1 U25307 ( .A(n22980), .B(n22365), .Y(n23587) );
  sky130_fd_sc_hd__nor2_1 U25308 ( .A(n18836), .B(n24463), .Y(n22383) );
  sky130_fd_sc_hd__nand2b_1 U25309 ( .A_N(n22845), .B(n27052), .Y(n26001) );
  sky130_fd_sc_hd__nand2_1 U25310 ( .A(n28056), .B(n27828), .Y(n22850) );
  sky130_fd_sc_hd__nand2_1 U25311 ( .A(n23004), .B(n27618), .Y(n22385) );
  sky130_fd_sc_hd__nand2_1 U25312 ( .A(n18837), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n21200) );
  sky130_fd_sc_hd__nand2b_1 U25313 ( .A_N(n26048), .B(n18838), .Y(n27787) );
  sky130_fd_sc_hd__nor2_1 U25314 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[3]), 
        .B(n26374), .Y(n23532) );
  sky130_fd_sc_hd__nand2b_1 U25315 ( .A_N(n26048), .B(n23532), .Y(n21707) );
  sky130_fd_sc_hd__nand2_1 U25316 ( .A(n25271), .B(n26003), .Y(n18839) );
  sky130_fd_sc_hd__o211ai_1 U25317 ( .A1(n26926), .A2(n22385), .B1(n27787), 
        .C1(n18839), .Y(n18840) );
  sky130_fd_sc_hd__a21oi_1 U25318 ( .A1(n22383), .A2(n26414), .B1(n18840), .Y(
        n18842) );
  sky130_fd_sc_hd__xor2_1 U25319 ( .A(n28489), .B(n24879), .X(n26249) );
  sky130_fd_sc_hd__nor2_1 U25320 ( .A(n21201), .B(n26048), .Y(n27806) );
  sky130_fd_sc_hd__nand2_1 U25321 ( .A(n26249), .B(n27806), .Y(n18841) );
  sky130_fd_sc_hd__nand3_1 U25322 ( .A(n26421), .B(n26240), .C(n28515), .Y(
        n18845) );
  sky130_fd_sc_hd__a22oi_1 U25323 ( .A1(n27810), .A2(n25916), .B1(n27808), 
        .B2(n22260), .Y(n18847) );
  sky130_fd_sc_hd__nand4_1 U25324 ( .A(n18849), .B(n18848), .C(n12116), .D(
        n18847), .Y(n18850) );
  sky130_fd_sc_hd__a21oi_1 U25325 ( .A1(n24086), .A2(n27789), .B1(n18850), .Y(
        n18851) );
  sky130_fd_sc_hd__a21oi_1 U25327 ( .A1(n26195), .A2(n18853), .B1(n18852), .Y(
        n18854) );
  sky130_fd_sc_hd__nand2b_1 U25328 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[7]), .Y(n22380) );
  sky130_fd_sc_hd__nand2_1 U25329 ( .A(n24682), .B(n27355), .Y(n18856) );
  sky130_fd_sc_hd__nor2_1 U25330 ( .A(n12041), .B(n18855), .Y(n22266) );
  sky130_fd_sc_hd__nand2_1 U25331 ( .A(n18858), .B(n22996), .Y(n18879) );
  sky130_fd_sc_hd__nand3_1 U25332 ( .A(n11094), .B(n18860), .C(n18859), .Y(
        n18861) );
  sky130_fd_sc_hd__nor2_1 U25333 ( .A(n18869), .B(n18861), .Y(n22988) );
  sky130_fd_sc_hd__nand2_1 U25334 ( .A(n22988), .B(j202_soc_core_j22_cpu_pc[7]), .Y(n18863) );
  sky130_fd_sc_hd__nand2_1 U25335 ( .A(n22987), .B(
        j202_soc_core_j22_cpu_rf_gbr[7]), .Y(n18862) );
  sky130_fd_sc_hd__o211a_2 U25336 ( .A1(n18864), .A2(n22084), .B1(n18863), 
        .C1(n18862), .X(n18878) );
  sky130_fd_sc_hd__nand2_1 U25337 ( .A(n18865), .B(n11094), .Y(n22897) );
  sky130_fd_sc_hd__o22ai_1 U25338 ( .A1(n18867), .A2(n22897), .B1(n18866), 
        .B2(n22894), .Y(n18876) );
  sky130_fd_sc_hd__nand2_1 U25339 ( .A(n18868), .B(n11094), .Y(n22285) );
  sky130_fd_sc_hd__nand3_1 U25340 ( .A(n18870), .B(n11094), .C(n18869), .Y(
        n22982) );
  sky130_fd_sc_hd__a2bb2oi_1 U25341 ( .B1(j202_soc_core_j22_cpu_rf_pr[7]), 
        .B2(n18872), .A1_N(n22982), .A2_N(n18871), .Y(n18873) );
  sky130_fd_sc_hd__o21ai_1 U25342 ( .A1(n22285), .A2(n18874), .B1(n18873), .Y(
        n18875) );
  sky130_fd_sc_hd__nor2_1 U25343 ( .A(n18876), .B(n18875), .Y(n18877) );
  sky130_fd_sc_hd__nand3_1 U25344 ( .A(n18879), .B(n18878), .C(n18877), .Y(
        n22384) );
  sky130_fd_sc_hd__nor2_1 U25345 ( .A(j202_soc_core_j22_cpu_memop_MEM__0_), 
        .B(n22779), .Y(n22950) );
  sky130_fd_sc_hd__nand2_1 U25346 ( .A(n22384), .B(n22950), .Y(n18880) );
  sky130_fd_sc_hd__inv_1 U25347 ( .A(n18881), .Y(n22568) );
  sky130_fd_sc_hd__a21oi_1 U25348 ( .A1(n22568), .A2(n22567), .B1(n18882), .Y(
        n18886) );
  sky130_fd_sc_hd__nand2_1 U25349 ( .A(n18884), .B(n18883), .Y(n18885) );
  sky130_fd_sc_hd__xor2_1 U25350 ( .A(n18886), .B(n18885), .X(n24337) );
  sky130_fd_sc_hd__nand2_1 U25351 ( .A(n24337), .B(n24461), .Y(n26061) );
  sky130_fd_sc_hd__o22a_1 U25352 ( .A1(n17933), .A2(n26001), .B1(n18888), .B2(
        n24463), .X(n26044) );
  sky130_fd_sc_hd__nand2_1 U25353 ( .A(n18889), .B(n22996), .Y(n18901) );
  sky130_fd_sc_hd__o22ai_1 U25354 ( .A1(n18891), .A2(n22983), .B1(n22982), 
        .B2(n18890), .Y(n18892) );
  sky130_fd_sc_hd__a21oi_1 U25355 ( .A1(n22986), .A2(
        j202_soc_core_j22_cpu_rf_gpr[15]), .B1(n18892), .Y(n18900) );
  sky130_fd_sc_hd__nand2_1 U25356 ( .A(n22988), .B(
        j202_soc_core_j22_cpu_pc[15]), .Y(n18894) );
  sky130_fd_sc_hd__nand2_1 U25357 ( .A(n22987), .B(
        j202_soc_core_j22_cpu_rf_gbr[15]), .Y(n18893) );
  sky130_fd_sc_hd__nand2_1 U25358 ( .A(n18894), .B(n18893), .Y(n18898) );
  sky130_fd_sc_hd__o22ai_1 U25359 ( .A1(n18896), .A2(n22897), .B1(n18895), 
        .B2(n22285), .Y(n18897) );
  sky130_fd_sc_hd__nor2_1 U25360 ( .A(n18898), .B(n18897), .Y(n18899) );
  sky130_fd_sc_hd__nand3_1 U25361 ( .A(n18901), .B(n18900), .C(n18899), .Y(
        n22472) );
  sky130_fd_sc_hd__nor2_1 U25362 ( .A(n24587), .B(n22779), .Y(n23973) );
  sky130_fd_sc_hd__nand2b_1 U25363 ( .A_N(n23973), .B(n24304), .Y(n24450) );
  sky130_fd_sc_hd__nand2_1 U25364 ( .A(n22472), .B(n24450), .Y(n18902) );
  sky130_fd_sc_hd__nand3_1 U25365 ( .A(n26061), .B(n26044), .C(n18902), .Y(
        n18904) );
  sky130_fd_sc_hd__nand2_1 U25366 ( .A(n18902), .B(n24467), .Y(n18903) );
  sky130_fd_sc_hd__nand2_1 U25367 ( .A(n18904), .B(n18903), .Y(n19097) );
  sky130_fd_sc_hd__a21oi_1 U25368 ( .A1(j202_soc_core_j22_cpu_ml_mach[31]), 
        .A2(n25679), .B1(n13087), .Y(n22026) );
  sky130_fd_sc_hd__o21ai_1 U25369 ( .A1(n19092), .A2(n11145), .B1(n22026), .Y(
        n22033) );
  sky130_fd_sc_hd__xnor2_1 U25370 ( .A(n22024), .B(n25777), .Y(n18906) );
  sky130_fd_sc_hd__xnor2_1 U25371 ( .A(n18925), .B(n25777), .Y(n18914) );
  sky130_fd_sc_hd__o22ai_1 U25372 ( .A1(n18993), .A2(n18906), .B1(n18914), 
        .B2(n18990), .Y(n22030) );
  sky130_fd_sc_hd__xnor2_1 U25373 ( .A(n18925), .B(n22023), .Y(n18905) );
  sky130_fd_sc_hd__a21o_1 U25374 ( .A1(n18990), .A2(n18993), .B1(n18906), .X(
        n22028) );
  sky130_fd_sc_hd__xnor2_1 U25375 ( .A(n18966), .B(n22023), .Y(n18907) );
  sky130_fd_sc_hd__a21oi_1 U25376 ( .A1(j202_soc_core_j22_cpu_ml_mach[30]), 
        .A2(n22940), .B1(n13087), .Y(n18908) );
  sky130_fd_sc_hd__o21ai_1 U25377 ( .A1(n24455), .A2(n11145), .B1(n18908), .Y(
        n18911) );
  sky130_fd_sc_hd__xnor2_1 U25378 ( .A(n22024), .B(n25389), .Y(n18910) );
  sky130_fd_sc_hd__xnor2_1 U25379 ( .A(n18925), .B(n25389), .Y(n18934) );
  sky130_fd_sc_hd__xnor2_1 U25380 ( .A(n18994), .B(n22023), .Y(n18909) );
  sky130_fd_sc_hd__a21o_1 U25381 ( .A1(n19020), .A2(n19023), .B1(n18910), .X(
        n18921) );
  sky130_fd_sc_hd__fa_1 U25382 ( .A(n18913), .B(n18912), .CIN(n18911), .COUT(
        n22031), .SUM(n18951) );
  sky130_fd_sc_hd__xnor2_1 U25383 ( .A(n18966), .B(n25777), .Y(n18916) );
  sky130_fd_sc_hd__o22ai_1 U25384 ( .A1(n18993), .A2(n18914), .B1(n18916), 
        .B2(n18990), .Y(n18933) );
  sky130_fd_sc_hd__a21oi_1 U25385 ( .A1(j202_soc_core_j22_cpu_ml_mach[29]), 
        .A2(n25679), .B1(n13087), .Y(n18915) );
  sky130_fd_sc_hd__o21ai_1 U25386 ( .A1(n24440), .A2(n11145), .B1(n18915), .Y(
        n18932) );
  sky130_fd_sc_hd__xnor2_1 U25387 ( .A(n18994), .B(n25777), .Y(n18935) );
  sky130_fd_sc_hd__o22ai_1 U25388 ( .A1(n18993), .A2(n18916), .B1(n18935), 
        .B2(n18990), .Y(n18930) );
  sky130_fd_sc_hd__xnor2_1 U25389 ( .A(n18971), .B(n22023), .Y(n18917) );
  sky130_fd_sc_hd__nor2_1 U25390 ( .A(n18918), .B(n18919), .Y(n22786) );
  sky130_fd_sc_hd__nand2_1 U25391 ( .A(n18919), .B(n18918), .Y(n22784) );
  sky130_fd_sc_hd__fa_1 U25392 ( .A(n11402), .B(n18922), .CIN(n18921), .COUT(
        n18952), .SUM(n18955) );
  sky130_fd_sc_hd__a21oi_1 U25393 ( .A1(j202_soc_core_j22_cpu_ml_mach[28]), 
        .A2(n25679), .B1(n13087), .Y(n18924) );
  sky130_fd_sc_hd__o21ai_1 U25394 ( .A1(n21893), .A2(n11145), .B1(n18924), .Y(
        n18940) );
  sky130_fd_sc_hd__xnor2_1 U25395 ( .A(n22024), .B(n23571), .Y(n18927) );
  sky130_fd_sc_hd__xnor2_1 U25396 ( .A(n18925), .B(n23571), .Y(n18988) );
  sky130_fd_sc_hd__o22ai_1 U25397 ( .A1(n18989), .A2(n18927), .B1(n18988), 
        .B2(n12044), .Y(n18946) );
  sky130_fd_sc_hd__xnor2_1 U25398 ( .A(n18941), .B(n22023), .Y(n18926) );
  sky130_fd_sc_hd__fah_1 U25399 ( .A(n18930), .B(n18929), .CI(n18928), .COUT(
        n18931), .SUM(n18938) );
  sky130_fd_sc_hd__fa_1 U25400 ( .A(n18933), .B(n18932), .CIN(n18931), .COUT(
        n18950), .SUM(n18953) );
  sky130_fd_sc_hd__xnor2_1 U25401 ( .A(n18966), .B(n25389), .Y(n19022) );
  sky130_fd_sc_hd__o22ai_1 U25402 ( .A1(n19023), .A2(n18934), .B1(n19022), 
        .B2(n19020), .Y(n18949) );
  sky130_fd_sc_hd__xnor2_1 U25403 ( .A(n18971), .B(n25777), .Y(n18942) );
  sky130_fd_sc_hd__o22ai_1 U25404 ( .A1(n18993), .A2(n18935), .B1(n18942), 
        .B2(n18990), .Y(n18948) );
  sky130_fd_sc_hd__a21oi_1 U25405 ( .A1(j202_soc_core_j22_cpu_ml_mach[27]), 
        .A2(n25679), .B1(n13087), .Y(n18936) );
  sky130_fd_sc_hd__o21ai_1 U25406 ( .A1(n18937), .A2(n11145), .B1(n18936), .Y(
        n18947) );
  sky130_fd_sc_hd__xnor2_1 U25407 ( .A(n18941), .B(n25777), .Y(n18992) );
  sky130_fd_sc_hd__o22ai_1 U25408 ( .A1(n18993), .A2(n18942), .B1(n18992), 
        .B2(n18990), .Y(n19036) );
  sky130_fd_sc_hd__xnor2_1 U25409 ( .A(n18962), .B(n22023), .Y(n18943) );
  sky130_fd_sc_hd__nor2_1 U25410 ( .A(n19081), .B(n19082), .Y(n22593) );
  sky130_fd_sc_hd__fah_1 U25411 ( .A(n18952), .B(n18951), .CI(n18950), .COUT(
        n18919), .SUM(n19083) );
  sky130_fd_sc_hd__fah_1 U25412 ( .A(n18955), .B(n18954), .CI(n18953), .COUT(
        n19084), .SUM(n19081) );
  sky130_fd_sc_hd__nand2_1 U25413 ( .A(n23020), .B(n12098), .Y(n22783) );
  sky130_fd_sc_hd__fah_1 U25414 ( .A(n18961), .B(n18960), .CI(n18959), .COUT(
        n19007), .SUM(n18979) );
  sky130_fd_sc_hd__xnor2_1 U25415 ( .A(n18962), .B(n25777), .Y(n18991) );
  sky130_fd_sc_hd__o22ai_1 U25416 ( .A1(n18993), .A2(n18991), .B1(n18963), 
        .B2(n18990), .Y(n18985) );
  sky130_fd_sc_hd__xnor2_1 U25417 ( .A(n18964), .B(n22023), .Y(n18965) );
  sky130_fd_sc_hd__xnor2_1 U25418 ( .A(n18966), .B(n23571), .Y(n18987) );
  sky130_fd_sc_hd__inv_2 U25419 ( .A(n19027), .Y(n18983) );
  sky130_fd_sc_hd__xnor2_1 U25420 ( .A(n18971), .B(n25389), .Y(n18995) );
  sky130_fd_sc_hd__o22ai_1 U25421 ( .A1(n19023), .A2(n18995), .B1(n18972), 
        .B2(n19020), .Y(n19005) );
  sky130_fd_sc_hd__xnor2_1 U25422 ( .A(n22024), .B(n23567), .Y(n19001) );
  sky130_fd_sc_hd__a21oi_1 U25423 ( .A1(j202_soc_core_j22_cpu_ml_mach[24]), 
        .A2(n25679), .B1(n13087), .Y(n18974) );
  sky130_fd_sc_hd__fah_1 U25425 ( .A(n18977), .B(n18976), .CI(n18975), .COUT(
        n18997), .SUM(n18969) );
  sky130_fd_sc_hd__fah_1 U25426 ( .A(n18980), .B(n18979), .CI(n18978), .COUT(
        n18996), .SUM(n19010) );
  sky130_fd_sc_hd__a21oi_1 U25427 ( .A1(j202_soc_core_j22_cpu_ml_mach[25]), 
        .A2(n22940), .B1(n13087), .Y(n18981) );
  sky130_fd_sc_hd__o22ai_1 U25429 ( .A1(n18989), .A2(n18988), .B1(n18987), 
        .B2(n12044), .Y(n19033) );
  sky130_fd_sc_hd__o22ai_1 U25430 ( .A1(n18993), .A2(n18992), .B1(n18991), 
        .B2(n18990), .Y(n19032) );
  sky130_fd_sc_hd__xnor2_1 U25431 ( .A(n18994), .B(n25389), .Y(n19021) );
  sky130_fd_sc_hd__o22ai_1 U25432 ( .A1(n19023), .A2(n19021), .B1(n18995), 
        .B2(n19020), .Y(n19031) );
  sky130_fd_sc_hd__fa_1 U25433 ( .A(n18998), .B(n18997), .CIN(n18996), .COUT(
        n19018), .SUM(n19014) );
  sky130_fd_sc_hd__xnor2_1 U25434 ( .A(n18999), .B(n22023), .Y(n19000) );
  sky130_fd_sc_hd__fah_1 U25435 ( .A(n19005), .B(n19004), .CI(n19003), .COUT(
        n19029), .SUM(n18998) );
  sky130_fd_sc_hd__o21ai_1 U25436 ( .A1(n19010), .A2(n19011), .B1(n19009), .Y(
        n19013) );
  sky130_fd_sc_hd__nand2_1 U25437 ( .A(n19011), .B(n19010), .Y(n19012) );
  sky130_fd_sc_hd__nand2_1 U25438 ( .A(n19013), .B(n19012), .Y(n19063) );
  sky130_fd_sc_hd__fah_1 U25439 ( .A(n19016), .B(n19015), .CI(n19014), .COUT(
        n19065), .SUM(n19064) );
  sky130_fd_sc_hd__nor2_1 U25440 ( .A(n22915), .B(n22920), .Y(n19295) );
  sky130_fd_sc_hd__o22ai_1 U25441 ( .A1(n19023), .A2(n19022), .B1(n19021), 
        .B2(n19020), .Y(n19045) );
  sky130_fd_sc_hd__a21oi_1 U25442 ( .A1(j202_soc_core_j22_cpu_ml_mach[26]), 
        .A2(n22940), .B1(n13087), .Y(n19024) );
  sky130_fd_sc_hd__o21ai_1 U25443 ( .A1(n19307), .A2(n11145), .B1(n19024), .Y(
        n19044) );
  sky130_fd_sc_hd__fah_1 U25444 ( .A(n19030), .B(n19029), .CI(n19028), .COUT(
        n19041), .SUM(n19017) );
  sky130_fd_sc_hd__fa_1 U25445 ( .A(n19033), .B(n19032), .CIN(n19031), .COUT(
        n19051), .SUM(n19037) );
  sky130_fd_sc_hd__fa_1 U25446 ( .A(n19036), .B(n19035), .CIN(n19034), .COUT(
        n19048), .SUM(n19050) );
  sky130_fd_sc_hd__fah_1 U25447 ( .A(n19039), .B(n19038), .CI(n19037), .COUT(
        n19049), .SUM(n19019) );
  sky130_fd_sc_hd__fah_1 U25448 ( .A(n19042), .B(n19041), .CI(n19040), .COUT(
        n19069), .SUM(n19068) );
  sky130_fd_sc_hd__fa_1 U25449 ( .A(n19045), .B(n19044), .CIN(n19043), .COUT(
        n19057), .SUM(n19042) );
  sky130_fd_sc_hd__fah_1 U25450 ( .A(n19051), .B(n19050), .CI(n19049), .COUT(
        n19055), .SUM(n19040) );
  sky130_fd_sc_hd__inv_1 U25451 ( .A(n21907), .Y(n21256) );
  sky130_fd_sc_hd__fah_1 U25452 ( .A(n19054), .B(n19053), .CI(n19052), .COUT(
        n19082), .SUM(n19071) );
  sky130_fd_sc_hd__fah_1 U25453 ( .A(n19057), .B(n19056), .CI(n19055), .COUT(
        n19072), .SUM(n19070) );
  sky130_fd_sc_hd__nor2_1 U25454 ( .A(n19071), .B(n19072), .Y(n19058) );
  sky130_fd_sc_hd__nand2_1 U25456 ( .A(n21256), .B(n21903), .Y(n19076) );
  sky130_fd_sc_hd__nor2_4 U25457 ( .A(n19080), .B(n22918), .Y(n22017) );
  sky130_fd_sc_hd__nand2_1 U25458 ( .A(n19064), .B(n19063), .Y(n22919) );
  sky130_fd_sc_hd__nand2_1 U25459 ( .A(n19066), .B(n19065), .Y(n22916) );
  sky130_fd_sc_hd__o21ai_1 U25460 ( .A1(n22919), .A2(n22915), .B1(n22916), .Y(
        n19296) );
  sky130_fd_sc_hd__nand2_1 U25461 ( .A(n19068), .B(n19067), .Y(n21258) );
  sky130_fd_sc_hd__nand2_1 U25462 ( .A(n19070), .B(n19069), .Y(n21905) );
  sky130_fd_sc_hd__inv_1 U25463 ( .A(n21905), .Y(n19074) );
  sky130_fd_sc_hd__nand2_1 U25464 ( .A(n19072), .B(n19071), .Y(n21902) );
  sky130_fd_sc_hd__a21oi_1 U25465 ( .A1(n19074), .A2(n21903), .B1(n19073), .Y(
        n19075) );
  sky130_fd_sc_hd__o21ai_1 U25466 ( .A1(n21258), .A2(n19076), .B1(n19075), .Y(
        n19077) );
  sky130_fd_sc_hd__a21oi_1 U25467 ( .A1(n19078), .A2(n19296), .B1(n19077), .Y(
        n19079) );
  sky130_fd_sc_hd__o21ai_2 U25468 ( .A1(n19080), .A2(n22921), .B1(n19079), .Y(
        n22789) );
  sky130_fd_sc_hd__nand2_1 U25469 ( .A(n19082), .B(n19081), .Y(n23019) );
  sky130_fd_sc_hd__nand2_1 U25470 ( .A(n19084), .B(n19083), .Y(n22592) );
  sky130_fd_sc_hd__a21oi_1 U25471 ( .A1(n19085), .A2(n12098), .B1(n22049), .Y(
        n22785) );
  sky130_fd_sc_hd__nand2_1 U25472 ( .A(n19089), .B(n19088), .Y(n19091) );
  sky130_fd_sc_hd__o21ai_2 U25473 ( .A1(n22562), .A2(n11866), .B1(n22563), .Y(
        n19090) );
  sky130_fd_sc_hd__xnor2_2 U25474 ( .A(n19091), .B(n19090), .Y(n26032) );
  sky130_fd_sc_hd__nand2_1 U25475 ( .A(n28056), .B(n18887), .Y(n26035) );
  sky130_fd_sc_hd__o21ai_1 U25476 ( .A1(n19092), .A2(n28045), .B1(n26035), .Y(
        n19093) );
  sky130_fd_sc_hd__a21oi_1 U25477 ( .A1(n26032), .A2(n25679), .B1(n19093), .Y(
        n19094) );
  sky130_fd_sc_hd__nand2_1 U25478 ( .A(n19095), .B(n19094), .Y(n26076) );
  sky130_fd_sc_hd__nand2_1 U25479 ( .A(n27717), .B(n27828), .Y(n22309) );
  sky130_fd_sc_hd__nand2_1 U25480 ( .A(n26076), .B(n23044), .Y(n19096) );
  sky130_fd_sc_hd__nand2_1 U25481 ( .A(j202_soc_core_qspi_wb_wdat[15]), .B(
        n29830), .Y(n29154) );
  sky130_fd_sc_hd__nand2_1 U25482 ( .A(n29439), .B(n22739), .Y(n19104) );
  sky130_fd_sc_hd__nor2_1 U25483 ( .A(n19099), .B(n21660), .Y(n22740) );
  sky130_fd_sc_hd__xnor2_1 U25484 ( .A(n14285), .B(n22740), .Y(n24713) );
  sky130_fd_sc_hd__o22a_1 U25485 ( .A1(n27616), .A2(n11186), .B1(n26309), .B2(
        n22743), .X(n19100) );
  sky130_fd_sc_hd__a21oi_1 U25487 ( .A1(n24713), .A2(n22747), .B1(n19101), .Y(
        n19103) );
  sky130_fd_sc_hd__nand2_1 U25488 ( .A(n24086), .B(n17225), .Y(n19102) );
  sky130_fd_sc_hd__nand3_1 U25489 ( .A(n19104), .B(n19103), .C(n19102), .Y(
        n29556) );
  sky130_fd_sc_hd__o21ai_2 U25490 ( .A1(n21192), .A2(n11866), .B1(n21193), .Y(
        n19107) );
  sky130_fd_sc_hd__xnor2_2 U25491 ( .A(n19108), .B(n19107), .Y(n25890) );
  sky130_fd_sc_hd__nand2_1 U25492 ( .A(n21234), .B(n21232), .Y(n19111) );
  sky130_fd_sc_hd__inv_1 U25493 ( .A(n19110), .Y(n22213) );
  sky130_fd_sc_hd__xnor2_1 U25494 ( .A(n19111), .B(n22213), .Y(n22368) );
  sky130_fd_sc_hd__nand2_1 U25495 ( .A(n22368), .B(n25679), .Y(n19114) );
  sky130_fd_sc_hd__nand2b_1 U25496 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[2]), .Y(n19113) );
  sky130_fd_sc_hd__nand2_1 U25497 ( .A(n28056), .B(n12436), .Y(n19112) );
  sky130_fd_sc_hd__nand3_1 U25499 ( .A(n19115), .B(
        j202_soc_core_j22_cpu_ma_M_MEM[1]), .C(n23511), .Y(n22229) );
  sky130_fd_sc_hd__nand2_1 U25500 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[1]), .B(
        j202_soc_core_j22_cpu_ma_M_address[1]), .Y(n19116) );
  sky130_fd_sc_hd__nor2_1 U25501 ( .A(j202_soc_core_j22_cpu_ma_M_address[0]), 
        .B(n19116), .Y(n22114) );
  sky130_fd_sc_hd__nand2_1 U25502 ( .A(j202_soc_core_memory0_ram_dout0[330]), 
        .B(n21490), .Y(n19118) );
  sky130_fd_sc_hd__nand2_1 U25503 ( .A(j202_soc_core_memory0_ram_dout0[426]), 
        .B(n12156), .Y(n19117) );
  sky130_fd_sc_hd__nand2_1 U25504 ( .A(n20742), .B(n20837), .Y(n19141) );
  sky130_fd_sc_hd__nand2_1 U25505 ( .A(n21088), .B(n13199), .Y(n19121) );
  sky130_fd_sc_hd__nor2_1 U25506 ( .A(n19121), .B(n19120), .Y(n20634) );
  sky130_fd_sc_hd__nand2_1 U25507 ( .A(n19129), .B(n11150), .Y(n20516) );
  sky130_fd_sc_hd__nand2_1 U25508 ( .A(n19122), .B(n20303), .Y(n20841) );
  sky130_fd_sc_hd__nor2_1 U25509 ( .A(n20634), .B(n20677), .Y(n20472) );
  sky130_fd_sc_hd__nand2b_1 U25510 ( .A_N(n20516), .B(n19143), .Y(n20675) );
  sky130_fd_sc_hd__nand2_1 U25511 ( .A(n19124), .B(n19123), .Y(n20775) );
  sky130_fd_sc_hd__nor2_1 U25512 ( .A(n19125), .B(n19185), .Y(n20828) );
  sky130_fd_sc_hd__nand4_1 U25513 ( .A(n20472), .B(n20675), .C(n20775), .D(
        n19126), .Y(n19127) );
  sky130_fd_sc_hd__nand2b_1 U25514 ( .A_N(n20467), .B(n20485), .Y(n20817) );
  sky130_fd_sc_hd__nand2b_1 U25515 ( .A_N(n20814), .B(n13199), .Y(n20852) );
  sky130_fd_sc_hd__nand2_1 U25516 ( .A(n19712), .B(n19159), .Y(n20687) );
  sky130_fd_sc_hd__nand3_1 U25517 ( .A(n20817), .B(n20852), .C(n20687), .Y(
        n20625) );
  sky130_fd_sc_hd__nor3_1 U25518 ( .A(n19141), .B(n19127), .C(n20625), .Y(
        n19135) );
  sky130_fd_sc_hd__nor2_1 U25519 ( .A(n19140), .B(n19148), .Y(n20804) );
  sky130_fd_sc_hd__nor2_1 U25520 ( .A(n19128), .B(n20515), .Y(n20731) );
  sky130_fd_sc_hd__nand2_1 U25521 ( .A(n20731), .B(n21359), .Y(n20793) );
  sky130_fd_sc_hd__nand2_1 U25522 ( .A(n19129), .B(n13182), .Y(n19183) );
  sky130_fd_sc_hd__nor2_1 U25523 ( .A(n19183), .B(n21132), .Y(n20486) );
  sky130_fd_sc_hd__nand3_1 U25524 ( .A(n20852), .B(n20793), .C(n20466), .Y(
        n19158) );
  sky130_fd_sc_hd__nand2b_1 U25525 ( .A_N(n20467), .B(n13199), .Y(n20635) );
  sky130_fd_sc_hd__nand2_1 U25526 ( .A(n19131), .B(n19130), .Y(n20829) );
  sky130_fd_sc_hd__nand2_1 U25527 ( .A(n20635), .B(n20829), .Y(n20499) );
  sky130_fd_sc_hd__nor2_1 U25528 ( .A(n20485), .B(n19203), .Y(n20474) );
  sky130_fd_sc_hd__nor2_1 U25529 ( .A(n20827), .B(n20474), .Y(n20838) );
  sky130_fd_sc_hd__nand2b_1 U25530 ( .A_N(n19185), .B(n19143), .Y(n20767) );
  sky130_fd_sc_hd__nand2b_1 U25531 ( .A_N(n19183), .B(n19132), .Y(n20528) );
  sky130_fd_sc_hd__nand4_1 U25532 ( .A(n20838), .B(n20767), .C(n20742), .D(
        n20528), .Y(n19133) );
  sky130_fd_sc_hd__nor3_1 U25533 ( .A(n19158), .B(n20499), .C(n19133), .Y(
        n19134) );
  sky130_fd_sc_hd__o22ai_1 U25534 ( .A1(n20632), .A2(n19135), .B1(n20846), 
        .B2(n19134), .Y(n19152) );
  sky130_fd_sc_hd__nand2b_1 U25535 ( .A_N(n19145), .B(n19146), .Y(n19193) );
  sky130_fd_sc_hd__nor2_1 U25536 ( .A(n21359), .B(n19193), .Y(n20765) );
  sky130_fd_sc_hd__nor2_1 U25537 ( .A(n21088), .B(n20603), .Y(n20743) );
  sky130_fd_sc_hd__nor2_1 U25538 ( .A(n20765), .B(n20743), .Y(n20798) );
  sky130_fd_sc_hd__nand2_1 U25539 ( .A(n20798), .B(n20841), .Y(n20821) );
  sky130_fd_sc_hd__nand2_1 U25540 ( .A(n19136), .B(n19146), .Y(n20762) );
  sky130_fd_sc_hd__nand2b_1 U25541 ( .A_N(n20515), .B(n19144), .Y(n20836) );
  sky130_fd_sc_hd__nand2_1 U25542 ( .A(n20762), .B(n20836), .Y(n20633) );
  sky130_fd_sc_hd__nand2_1 U25543 ( .A(n19162), .B(n20817), .Y(n19139) );
  sky130_fd_sc_hd__nand2_1 U25544 ( .A(n20467), .B(n19203), .Y(n19137) );
  sky130_fd_sc_hd__nand2_1 U25545 ( .A(n19137), .B(n13199), .Y(n20746) );
  sky130_fd_sc_hd__nand4_1 U25546 ( .A(n20746), .B(n20656), .C(n20852), .D(
        n20793), .Y(n19138) );
  sky130_fd_sc_hd__or3_1 U25547 ( .A(n20821), .B(n19139), .C(n19138), .X(
        n20834) );
  sky130_fd_sc_hd__nand2_1 U25548 ( .A(n19148), .B(n19140), .Y(n20684) );
  sky130_fd_sc_hd__nand2_1 U25549 ( .A(n20834), .B(n20856), .Y(n19151) );
  sky130_fd_sc_hd__nand2_1 U25550 ( .A(n20532), .B(n21598), .Y(n20790) );
  sky130_fd_sc_hd__nand2b_1 U25551 ( .A_N(n20490), .B(n20790), .Y(n20598) );
  sky130_fd_sc_hd__nand3_1 U25552 ( .A(n20740), .B(n19142), .C(n20843), .Y(
        n19149) );
  sky130_fd_sc_hd__nand3_1 U25553 ( .A(n19143), .B(
        j202_soc_core_bootrom_00_address_w[4]), .C(n11150), .Y(n20831) );
  sky130_fd_sc_hd__nor2_1 U25554 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n20831), .Y(n20815) );
  sky130_fd_sc_hd__nand2_1 U25555 ( .A(n20766), .B(n20675), .Y(n20744) );
  sky130_fd_sc_hd__nand2b_1 U25556 ( .A_N(n20656), .B(n20485), .Y(n20774) );
  sky130_fd_sc_hd__nand2b_1 U25557 ( .A_N(n20731), .B(n20774), .Y(n20595) );
  sky130_fd_sc_hd__nand2b_1 U25558 ( .A_N(n19145), .B(n19144), .Y(n20799) );
  sky130_fd_sc_hd__nand2_1 U25559 ( .A(n20809), .B(n19146), .Y(n20559) );
  sky130_fd_sc_hd__nand2b_1 U25560 ( .A_N(n20559), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n20736) );
  sky130_fd_sc_hd__nand4_1 U25561 ( .A(n19147), .B(n20471), .C(n20799), .D(
        n20736), .Y(n19175) );
  sky130_fd_sc_hd__nor2_1 U25562 ( .A(n19148), .B(n18744), .Y(n20850) );
  sky130_fd_sc_hd__o21ai_1 U25563 ( .A1(n19149), .A2(n19175), .B1(n20850), .Y(
        n19150) );
  sky130_fd_sc_hd__nand3b_1 U25564 ( .A_N(n19152), .B(n19151), .C(n19150), .Y(
        n19153) );
  sky130_fd_sc_hd__nand2_1 U25565 ( .A(n19153), .B(n20508), .Y(n19173) );
  sky130_fd_sc_hd__nand2b_1 U25566 ( .A_N(n20559), .B(n13179), .Y(n20792) );
  sky130_fd_sc_hd__nand4_1 U25567 ( .A(n20837), .B(n20829), .C(n20792), .D(
        n20799), .Y(n19154) );
  sky130_fd_sc_hd__nor2_1 U25568 ( .A(n19154), .B(n20625), .Y(n20638) );
  sky130_fd_sc_hd__nand2b_1 U25569 ( .A_N(n19185), .B(n19159), .Y(n20623) );
  sky130_fd_sc_hd__nand2_1 U25570 ( .A(n20623), .B(n20841), .Y(n19155) );
  sky130_fd_sc_hd__nor3_1 U25571 ( .A(n19155), .B(n20765), .C(n20744), .Y(
        n19156) );
  sky130_fd_sc_hd__nand2_1 U25572 ( .A(n20638), .B(n19156), .Y(n19170) );
  sky130_fd_sc_hd__nor2_1 U25573 ( .A(n19157), .B(n20743), .Y(n20530) );
  sky130_fd_sc_hd__nand2b_1 U25574 ( .A_N(n20516), .B(n19159), .Y(n20741) );
  sky130_fd_sc_hd__nand2_1 U25575 ( .A(n20741), .B(n20559), .Y(n19160) );
  sky130_fd_sc_hd__nand2_1 U25576 ( .A(n20762), .B(n20623), .Y(n20561) );
  sky130_fd_sc_hd__nor3_1 U25577 ( .A(n19160), .B(n20598), .C(n20561), .Y(
        n19161) );
  sky130_fd_sc_hd__a31oi_1 U25578 ( .A1(n20530), .A2(n20664), .A3(n19161), 
        .B1(n20846), .Y(n19169) );
  sky130_fd_sc_hd__nand2_1 U25579 ( .A(n20830), .B(n20767), .Y(n20737) );
  sky130_fd_sc_hd__nand2_1 U25580 ( .A(n20742), .B(n20774), .Y(n20844) );
  sky130_fd_sc_hd__nand3_1 U25581 ( .A(n19162), .B(n20521), .C(n20680), .Y(
        n19163) );
  sky130_fd_sc_hd__nor3_1 U25582 ( .A(n20737), .B(n20844), .C(n19163), .Y(
        n19167) );
  sky130_fd_sc_hd__nand3_1 U25583 ( .A(n20739), .B(n20831), .C(n20830), .Y(
        n20626) );
  sky130_fd_sc_hd__nor2_1 U25584 ( .A(n21595), .B(n19183), .Y(n19164) );
  sky130_fd_sc_hd__nor2_1 U25585 ( .A(n19164), .B(n20474), .Y(n20523) );
  sky130_fd_sc_hd__nand2_1 U25586 ( .A(n20523), .B(n20799), .Y(n19165) );
  sky130_fd_sc_hd__o21ai_1 U25588 ( .A1(n20630), .A2(n19167), .B1(n19166), .Y(
        n19168) );
  sky130_fd_sc_hd__a211o_1 U25589 ( .A1(n20856), .A2(n19170), .B1(n19169), 
        .C1(n19168), .X(n19171) );
  sky130_fd_sc_hd__nand2_1 U25590 ( .A(n19171), .B(n20505), .Y(n19172) );
  sky130_fd_sc_hd__nand2_1 U25591 ( .A(n19173), .B(n19172), .Y(n19174) );
  sky130_fd_sc_hd__nand2_1 U25592 ( .A(n19174), .B(n21629), .Y(n19229) );
  sky130_fd_sc_hd__nand2_1 U25593 ( .A(n20792), .B(n20836), .Y(n20605) );
  sky130_fd_sc_hd__nor3_1 U25594 ( .A(n20634), .B(n20605), .C(n20737), .Y(
        n20803) );
  sky130_fd_sc_hd__nand2_1 U25595 ( .A(n19206), .B(
        j202_soc_core_bootrom_00_address_w[4]), .Y(n20553) );
  sky130_fd_sc_hd__nand3_1 U25596 ( .A(n19176), .B(n20803), .C(n20553), .Y(
        n19177) );
  sky130_fd_sc_hd__nand2_1 U25597 ( .A(n19177), .B(n20833), .Y(n19198) );
  sky130_fd_sc_hd__nor2_1 U25598 ( .A(n19178), .B(n20633), .Y(n20820) );
  sky130_fd_sc_hd__nand3_1 U25599 ( .A(n20742), .B(n19179), .C(n20799), .Y(
        n20563) );
  sky130_fd_sc_hd__nor2_1 U25600 ( .A(n20516), .B(n19180), .Y(n20652) );
  sky130_fd_sc_hd__nand2_1 U25601 ( .A(n20674), .B(n20673), .Y(n19181) );
  sky130_fd_sc_hd__nand2_1 U25602 ( .A(n20687), .B(n19181), .Y(n19182) );
  sky130_fd_sc_hd__nor2_1 U25603 ( .A(n20652), .B(n19182), .Y(n20518) );
  sky130_fd_sc_hd__nor2_1 U25604 ( .A(n19185), .B(n19184), .Y(n20771) );
  sky130_fd_sc_hd__a211o_1 U25605 ( .A1(n19186), .A2(n20303), .B1(n20634), 
        .C1(n20771), .X(n19187) );
  sky130_fd_sc_hd__nor2_1 U25606 ( .A(n19187), .B(n20765), .Y(n19188) );
  sky130_fd_sc_hd__nand4_1 U25607 ( .A(n20820), .B(n20551), .C(n20518), .D(
        n19188), .Y(n19189) );
  sky130_fd_sc_hd__nand2_1 U25608 ( .A(n19189), .B(n20804), .Y(n19197) );
  sky130_fd_sc_hd__nand4_1 U25609 ( .A(n20830), .B(n20793), .C(n20528), .D(
        n20775), .Y(n19190) );
  sky130_fd_sc_hd__nand3_1 U25610 ( .A(n20742), .B(n20741), .C(n20680), .Y(
        n20554) );
  sky130_fd_sc_hd__nor2_1 U25611 ( .A(n19190), .B(n20554), .Y(n19191) );
  sky130_fd_sc_hd__nand2_1 U25612 ( .A(n20798), .B(n19191), .Y(n19192) );
  sky130_fd_sc_hd__nand2_1 U25613 ( .A(n19192), .B(n20856), .Y(n19196) );
  sky130_fd_sc_hd__nand4_1 U25614 ( .A(n20635), .B(n20775), .C(n19193), .D(
        n20774), .Y(n19194) );
  sky130_fd_sc_hd__nand2_1 U25615 ( .A(n19194), .B(n20850), .Y(n19195) );
  sky130_fd_sc_hd__nand4_1 U25616 ( .A(n19198), .B(n19197), .C(n19196), .D(
        n19195), .Y(n19199) );
  sky130_fd_sc_hd__a22oi_1 U25617 ( .A1(n21446), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[106]), .B1(n19199), .B2(
        n20784), .Y(n19228) );
  sky130_fd_sc_hd__nand2_1 U25618 ( .A(n20759), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[74]), .Y(n19223) );
  sky130_fd_sc_hd__nand2b_1 U25619 ( .A_N(n21515), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[42]), .Y(n19222) );
  sky130_fd_sc_hd__nand2_1 U25620 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[10]), .Y(n19221) );
  sky130_fd_sc_hd__nand4_1 U25621 ( .A(n19223), .B(n19222), .C(n21768), .D(
        n19221), .Y(n19200) );
  sky130_fd_sc_hd__nor2_1 U25622 ( .A(n28546), .B(n21517), .Y(n19224) );
  sky130_fd_sc_hd__nor2_1 U25623 ( .A(n19200), .B(n19224), .Y(n19215) );
  sky130_fd_sc_hd__nand3_1 U25624 ( .A(n20736), .B(n19203), .C(n20623), .Y(
        n19201) );
  sky130_fd_sc_hd__nor2_1 U25625 ( .A(n19201), .B(n20625), .Y(n20734) );
  sky130_fd_sc_hd__nand2b_1 U25626 ( .A_N(n20734), .B(n20850), .Y(n19213) );
  sky130_fd_sc_hd__nor2_1 U25627 ( .A(n19202), .B(n20765), .Y(n20637) );
  sky130_fd_sc_hd__nand2_1 U25628 ( .A(n20637), .B(n20841), .Y(n20601) );
  sky130_fd_sc_hd__nand2_1 U25629 ( .A(n20817), .B(n19203), .Y(n20612) );
  sky130_fd_sc_hd__nand3_1 U25630 ( .A(n19204), .B(n20551), .C(n20665), .Y(
        n19205) );
  sky130_fd_sc_hd__nand2_1 U25631 ( .A(n19205), .B(n20804), .Y(n19212) );
  sky130_fd_sc_hd__inv_1 U25632 ( .A(n20743), .Y(n20662) );
  sky130_fd_sc_hd__nand2_1 U25633 ( .A(n20662), .B(n20635), .Y(n20568) );
  sky130_fd_sc_hd__nand3_1 U25634 ( .A(n20551), .B(n20560), .C(n19207), .Y(
        n19208) );
  sky130_fd_sc_hd__o21ai_1 U25635 ( .A1(n20568), .A2(n19208), .B1(n20833), .Y(
        n19211) );
  sky130_fd_sc_hd__nand2_1 U25636 ( .A(n20799), .B(n20560), .Y(n19209) );
  sky130_fd_sc_hd__nand2_1 U25637 ( .A(n20762), .B(n20482), .Y(n20646) );
  sky130_fd_sc_hd__nand4_1 U25639 ( .A(n19213), .B(n19212), .C(n19211), .D(
        n19210), .Y(n19214) );
  sky130_fd_sc_hd__nand2_1 U25640 ( .A(n19214), .B(n20757), .Y(n19226) );
  sky130_fd_sc_hd__nand2_1 U25641 ( .A(j202_soc_core_memory0_ram_dout0[42]), 
        .B(n21633), .Y(n19219) );
  sky130_fd_sc_hd__nand2_1 U25642 ( .A(j202_soc_core_memory0_ram_dout0[170]), 
        .B(n21487), .Y(n19218) );
  sky130_fd_sc_hd__nand2_1 U25643 ( .A(j202_soc_core_memory0_ram_dout0[138]), 
        .B(n21489), .Y(n19217) );
  sky130_fd_sc_hd__nand2_1 U25644 ( .A(j202_soc_core_memory0_ram_dout0[74]), 
        .B(n21642), .Y(n19216) );
  sky130_fd_sc_hd__nand2_1 U25645 ( .A(j202_soc_core_memory0_ram_dout0[490]), 
        .B(n21650), .Y(n19233) );
  sky130_fd_sc_hd__nand4_1 U25646 ( .A(n19223), .B(n19222), .C(n21653), .D(
        n19221), .Y(n19225) );
  sky130_fd_sc_hd__nor2_1 U25647 ( .A(n19225), .B(n19224), .Y(n19227) );
  sky130_fd_sc_hd__nand3_1 U25648 ( .A(n19228), .B(n19227), .C(n19226), .Y(
        n19231) );
  sky130_fd_sc_hd__nor2_1 U25649 ( .A(n19231), .B(n19230), .Y(n19232) );
  sky130_fd_sc_hd__nand2_1 U25650 ( .A(n19233), .B(n19232), .Y(n20716) );
  sky130_fd_sc_hd__nand2_1 U25651 ( .A(j202_soc_core_j22_cpu_ma_M_address[0]), 
        .B(j202_soc_core_j22_cpu_ma_M_address[1]), .Y(n19234) );
  sky130_fd_sc_hd__nand2_1 U25652 ( .A(n25940), .B(n19234), .Y(n22232) );
  sky130_fd_sc_hd__nand2_1 U25653 ( .A(n19235), .B(n24069), .Y(n22230) );
  sky130_fd_sc_hd__nand2_1 U25654 ( .A(n25263), .B(n26144), .Y(n25824) );
  sky130_fd_sc_hd__nand2_1 U25655 ( .A(n19237), .B(n26929), .Y(n19260) );
  sky130_fd_sc_hd__nand2_1 U25657 ( .A(n19241), .B(n19240), .Y(n19242) );
  sky130_fd_sc_hd__xnor2_1 U25658 ( .A(n19243), .B(n19242), .Y(n22364) );
  sky130_fd_sc_hd__nand2_1 U25659 ( .A(n22364), .B(n24461), .Y(n22431) );
  sky130_fd_sc_hd__nor2_1 U25660 ( .A(n19244), .B(n24463), .Y(n22427) );
  sky130_fd_sc_hd__nand2_1 U25661 ( .A(n27115), .B(n26003), .Y(n19246) );
  sky130_fd_sc_hd__nand2_1 U25662 ( .A(n26937), .B(n26034), .Y(n19245) );
  sky130_fd_sc_hd__o211ai_1 U25663 ( .A1(n26926), .A2(n22429), .B1(n19246), 
        .C1(n19245), .Y(n19247) );
  sky130_fd_sc_hd__a21oi_1 U25664 ( .A1(n26414), .A2(n22427), .B1(n19247), .Y(
        n19248) );
  sky130_fd_sc_hd__o21ai_0 U25665 ( .A1(n27798), .A2(n26943), .B1(n19248), .Y(
        n19251) );
  sky130_fd_sc_hd__o22ai_1 U25666 ( .A1(n26284), .A2(n27795), .B1(n27800), 
        .B2(n25996), .Y(n19250) );
  sky130_fd_sc_hd__o22ai_1 U25667 ( .A1(n27816), .A2(n26936), .B1(n26272), 
        .B2(n26932), .Y(n19249) );
  sky130_fd_sc_hd__nor3_1 U25668 ( .A(n19251), .B(n19250), .C(n19249), .Y(
        n19255) );
  sky130_fd_sc_hd__xor2_1 U25669 ( .A(n26929), .B(n26937), .X(n26252) );
  sky130_fd_sc_hd__o22a_1 U25670 ( .A1(n11190), .A2(n27803), .B1(n25872), .B2(
        n26252), .X(n19253) );
  sky130_fd_sc_hd__a22oi_1 U25671 ( .A1(n27810), .A2(n22136), .B1(n27808), 
        .B2(n26377), .Y(n19252) );
  sky130_fd_sc_hd__o211a_2 U25672 ( .A1(n26937), .A2(n22251), .B1(n19253), 
        .C1(n19252), .X(n19254) );
  sky130_fd_sc_hd__o211ai_1 U25673 ( .A1(n26926), .A2(n22431), .B1(n19255), 
        .C1(n19254), .Y(n19256) );
  sky130_fd_sc_hd__a21oi_1 U25674 ( .A1(n27789), .A2(n24048), .B1(n19256), .Y(
        n19259) );
  sky130_fd_sc_hd__nand2_1 U25676 ( .A(n19264), .B(n22996), .Y(n19276) );
  sky130_fd_sc_hd__o22ai_1 U25677 ( .A1(n19266), .A2(n22983), .B1(n19265), 
        .B2(n22982), .Y(n19267) );
  sky130_fd_sc_hd__a21oi_1 U25678 ( .A1(n22986), .A2(
        j202_soc_core_j22_cpu_rf_gpr[2]), .B1(n19267), .Y(n19275) );
  sky130_fd_sc_hd__nand2_1 U25679 ( .A(n22988), .B(j202_soc_core_j22_cpu_pc[2]), .Y(n19269) );
  sky130_fd_sc_hd__nand2_1 U25680 ( .A(n22987), .B(
        j202_soc_core_j22_cpu_rf_gbr[2]), .Y(n19268) );
  sky130_fd_sc_hd__nand2_1 U25681 ( .A(n19269), .B(n19268), .Y(n19273) );
  sky130_fd_sc_hd__o22ai_1 U25682 ( .A1(n19271), .A2(n22897), .B1(n19270), 
        .B2(n22285), .Y(n19272) );
  sky130_fd_sc_hd__nor2_1 U25683 ( .A(n19273), .B(n19272), .Y(n19274) );
  sky130_fd_sc_hd__nand3_1 U25684 ( .A(n19276), .B(n19275), .C(n19274), .Y(
        n22428) );
  sky130_fd_sc_hd__nand2_1 U25685 ( .A(n22428), .B(n22950), .Y(n19277) );
  sky130_fd_sc_hd__nand2_1 U25686 ( .A(n13076), .B(n19278), .Y(n19280) );
  sky130_fd_sc_hd__inv_1 U25687 ( .A(n19279), .Y(n21284) );
  sky130_fd_sc_hd__xnor2_1 U25688 ( .A(n19280), .B(n21284), .Y(n24313) );
  sky130_fd_sc_hd__nand2_1 U25689 ( .A(n24313), .B(n24461), .Y(n26958) );
  sky130_fd_sc_hd__o22a_1 U25690 ( .A1(n19308), .A2(n26001), .B1(n19281), .B2(
        n24463), .X(n26927) );
  sky130_fd_sc_hd__o22ai_1 U25691 ( .A1(n19283), .A2(n22983), .B1(n22982), 
        .B2(n19282), .Y(n19284) );
  sky130_fd_sc_hd__a21oi_1 U25692 ( .A1(n22986), .A2(
        j202_soc_core_j22_cpu_rf_gpr[10]), .B1(n19284), .Y(n19288) );
  sky130_fd_sc_hd__a22oi_1 U25693 ( .A1(n22988), .A2(
        j202_soc_core_j22_cpu_pc[10]), .B1(n22987), .B2(
        j202_soc_core_j22_cpu_rf_gbr[10]), .Y(n19287) );
  sky130_fd_sc_hd__nand2_1 U25694 ( .A(n22989), .B(
        j202_soc_core_j22_cpu_rf_tmp[10]), .Y(n19286) );
  sky130_fd_sc_hd__nand2_1 U25695 ( .A(n22990), .B(
        j202_soc_core_j22_cpu_rf_vbr[10]), .Y(n19285) );
  sky130_fd_sc_hd__nand4_1 U25696 ( .A(n19288), .B(n19287), .C(n19286), .D(
        n19285), .Y(n19289) );
  sky130_fd_sc_hd__a21o_1 U25697 ( .A1(n19290), .A2(n22996), .B1(n19289), .X(
        n22668) );
  sky130_fd_sc_hd__nand2_1 U25698 ( .A(n22668), .B(n24450), .Y(n19291) );
  sky130_fd_sc_hd__nand3_1 U25699 ( .A(n26958), .B(n26927), .C(n19291), .Y(
        n19293) );
  sky130_fd_sc_hd__nand2_1 U25700 ( .A(n19291), .B(n24467), .Y(n19292) );
  sky130_fd_sc_hd__nand2_1 U25701 ( .A(n19293), .B(n19292), .Y(n19313) );
  sky130_fd_sc_hd__nand2_1 U25702 ( .A(n19294), .B(n21258), .Y(n19302) );
  sky130_fd_sc_hd__inv_1 U25703 ( .A(n19295), .Y(n21257) );
  sky130_fd_sc_hd__nor2_1 U25704 ( .A(n21257), .B(n22918), .Y(n19298) );
  sky130_fd_sc_hd__nand2_1 U25705 ( .A(n23030), .B(n19298), .Y(n19300) );
  sky130_fd_sc_hd__inv_1 U25706 ( .A(n19296), .Y(n21259) );
  sky130_fd_sc_hd__o21ai_1 U25707 ( .A1(n21257), .A2(n22921), .B1(n21259), .Y(
        n19297) );
  sky130_fd_sc_hd__xnor2_2 U25708 ( .A(n19302), .B(n19301), .Y(n23471) );
  sky130_fd_sc_hd__nand2_1 U25709 ( .A(n23471), .B(n24452), .Y(n19311) );
  sky130_fd_sc_hd__nand2_1 U25710 ( .A(n21275), .B(n21273), .Y(n19306) );
  sky130_fd_sc_hd__xnor2_1 U25712 ( .A(n19306), .B(n19305), .Y(n22657) );
  sky130_fd_sc_hd__o22ai_1 U25713 ( .A1(n24456), .A2(n19308), .B1(n19307), 
        .B2(n28045), .Y(n19309) );
  sky130_fd_sc_hd__a21oi_1 U25714 ( .A1(n22657), .A2(n22940), .B1(n19309), .Y(
        n19310) );
  sky130_fd_sc_hd__nand2_1 U25715 ( .A(n27773), .B(n23044), .Y(n19312) );
  sky130_fd_sc_hd__nand2_1 U25717 ( .A(j202_soc_core_qspi_wb_wdat[10]), .B(
        n29745), .Y(n29156) );
  sky130_fd_sc_hd__o21ai_0 U25718 ( .A1(n11150), .A2(n20515), .B1(n20372), .Y(
        n19315) );
  sky130_fd_sc_hd__nand2_1 U25719 ( .A(n20379), .B(n19612), .Y(n19314) );
  sky130_fd_sc_hd__nor3_1 U25720 ( .A(n19315), .B(n20296), .C(n19314), .Y(
        n19316) );
  sky130_fd_sc_hd__nand2_1 U25721 ( .A(n19562), .B(n20268), .Y(n20312) );
  sky130_fd_sc_hd__nor2_1 U25722 ( .A(n19607), .B(n19574), .Y(n20340) );
  sky130_fd_sc_hd__nand3_1 U25723 ( .A(n19316), .B(n19657), .C(n20340), .Y(
        n19318) );
  sky130_fd_sc_hd__o21ai_0 U25724 ( .A1(n19318), .A2(n19317), .B1(n20385), .Y(
        n19334) );
  sky130_fd_sc_hd__nand2_1 U25725 ( .A(n19369), .B(n20268), .Y(n19320) );
  sky130_fd_sc_hd__nor3_1 U25726 ( .A(n19320), .B(n19319), .C(n19651), .Y(
        n19323) );
  sky130_fd_sc_hd__nor2_1 U25727 ( .A(n19581), .B(n19321), .Y(n19624) );
  sky130_fd_sc_hd__nand3_1 U25728 ( .A(n19323), .B(n19624), .C(n20392), .Y(
        n19328) );
  sky130_fd_sc_hd__nor2_1 U25729 ( .A(n19561), .B(n19324), .Y(n19325) );
  sky130_fd_sc_hd__nand4_1 U25730 ( .A(n20380), .B(n19325), .C(n20306), .D(
        n19575), .Y(n19326) );
  sky130_fd_sc_hd__nand3_1 U25731 ( .A(n20344), .B(n20363), .C(n20371), .Y(
        n20278) );
  sky130_fd_sc_hd__o31a_1 U25732 ( .A1(n19326), .A2(n20278), .A3(n19579), .B1(
        n20393), .X(n19327) );
  sky130_fd_sc_hd__a21oi_1 U25733 ( .A1(n19328), .A2(n20368), .B1(n19327), .Y(
        n19333) );
  sky130_fd_sc_hd__nand4_1 U25734 ( .A(n20311), .B(n19397), .C(n20360), .D(
        n20293), .Y(n19331) );
  sky130_fd_sc_hd__and3_1 U25735 ( .A(n19622), .B(n19329), .C(n19612), .X(
        n19330) );
  sky130_fd_sc_hd__nand3_1 U25736 ( .A(n20392), .B(n19330), .C(n20363), .Y(
        n19620) );
  sky130_fd_sc_hd__nand3_1 U25738 ( .A(n19334), .B(n19333), .C(n19332), .Y(
        n19335) );
  sky130_fd_sc_hd__nand2_1 U25739 ( .A(n19335), .B(n20643), .Y(n19359) );
  sky130_fd_sc_hd__and3_1 U25740 ( .A(n29435), .B(j202_soc_core_aquc_ADR__2_), 
        .C(n25179), .X(n19596) );
  sky130_fd_sc_hd__a2bb2oi_1 U25741 ( .B1(n19596), .B2(
        j202_soc_core_bldc_core_00_adc_en), .A1_N(n29121), .A2_N(n19595), .Y(
        n19336) );
  sky130_fd_sc_hd__nand2_1 U25743 ( .A(n19338), .B(n19605), .Y(n19358) );
  sky130_fd_sc_hd__nand3_1 U25744 ( .A(n19562), .B(n20343), .C(n20326), .Y(
        n19339) );
  sky130_fd_sc_hd__o31ai_1 U25745 ( .A1(n19339), .A2(n19373), .A3(n19579), 
        .B1(n20385), .Y(n19355) );
  sky130_fd_sc_hd__nand4b_1 U25746 ( .A_N(n19574), .B(n20348), .C(n20307), .D(
        n19649), .Y(n19340) );
  sky130_fd_sc_hd__nand2_1 U25747 ( .A(n20389), .B(n20343), .Y(n19341) );
  sky130_fd_sc_hd__nor2_1 U25748 ( .A(n19341), .B(n20278), .Y(n19342) );
  sky130_fd_sc_hd__nand3_1 U25749 ( .A(n20367), .B(n19558), .C(n19342), .Y(
        n19343) );
  sky130_fd_sc_hd__nand2_1 U25750 ( .A(n19343), .B(n20374), .Y(n19354) );
  sky130_fd_sc_hd__nand4_1 U25751 ( .A(n19346), .B(n20311), .C(n20271), .D(
        n19345), .Y(n19347) );
  sky130_fd_sc_hd__nand2_1 U25752 ( .A(n19347), .B(n20393), .Y(n19353) );
  sky130_fd_sc_hd__nand2_1 U25753 ( .A(n19649), .B(n20339), .Y(n19655) );
  sky130_fd_sc_hd__nor2_1 U25754 ( .A(n19608), .B(n19655), .Y(n19572) );
  sky130_fd_sc_hd__and3_1 U25755 ( .A(n20306), .B(n20364), .C(n19348), .X(
        n19349) );
  sky130_fd_sc_hd__nand3_1 U25756 ( .A(n19350), .B(n19572), .C(n19349), .Y(
        n19351) );
  sky130_fd_sc_hd__nand2_1 U25757 ( .A(n19351), .B(n20368), .Y(n19352) );
  sky130_fd_sc_hd__nand4_1 U25758 ( .A(n19355), .B(n19354), .C(n19353), .D(
        n19352), .Y(n19356) );
  sky130_fd_sc_hd__nand2_1 U25759 ( .A(n19356), .B(n20757), .Y(n19357) );
  sky130_fd_sc_hd__nand3_1 U25760 ( .A(n19359), .B(n19358), .C(n19357), .Y(
        n19425) );
  sky130_fd_sc_hd__nand2b_1 U25761 ( .A_N(n21515), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[33]), .Y(n19416) );
  sky130_fd_sc_hd__nand2_1 U25762 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[1]), .Y(n19415) );
  sky130_fd_sc_hd__nand3_1 U25763 ( .A(n19416), .B(n21768), .C(n19415), .Y(
        n19368) );
  sky130_fd_sc_hd__o22a_1 U25764 ( .A1(n19361), .A2(n21512), .B1(n19360), .B2(
        n21519), .X(n19414) );
  sky130_fd_sc_hd__nand2_1 U25765 ( .A(n21504), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[9]), .Y(n19365) );
  sky130_fd_sc_hd__nand2_1 U25766 ( .A(n24720), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[17]), .Y(n19364) );
  sky130_fd_sc_hd__nand2_1 U25767 ( .A(n21505), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[1]), .Y(n19363) );
  sky130_fd_sc_hd__nand2_1 U25768 ( .A(n21506), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[25]), .Y(n19362) );
  sky130_fd_sc_hd__nand4_1 U25769 ( .A(n19365), .B(n19364), .C(n19363), .D(
        n19362), .Y(n19366) );
  sky130_fd_sc_hd__nand2_1 U25770 ( .A(n21513), .B(n19366), .Y(n19417) );
  sky130_fd_sc_hd__nand2_1 U25771 ( .A(n19414), .B(n19417), .Y(n19367) );
  sky130_fd_sc_hd__nor2_1 U25772 ( .A(n28307), .B(n21517), .Y(n19418) );
  sky130_fd_sc_hd__nor3_1 U25773 ( .A(n19368), .B(n19367), .C(n19418), .Y(
        n19412) );
  sky130_fd_sc_hd__nand4_1 U25774 ( .A(n19371), .B(n20292), .C(n19659), .D(
        n19404), .Y(n19372) );
  sky130_fd_sc_hd__nand2_1 U25775 ( .A(n19624), .B(n19612), .Y(n20282) );
  sky130_fd_sc_hd__o21ai_0 U25776 ( .A1(n19372), .A2(n20282), .B1(n20385), .Y(
        n19386) );
  sky130_fd_sc_hd__nand4_1 U25777 ( .A(n19564), .B(n20349), .C(n20360), .D(
        n19612), .Y(n19375) );
  sky130_fd_sc_hd__nand3_1 U25779 ( .A(n20344), .B(n20310), .C(n20348), .Y(
        n19666) );
  sky130_fd_sc_hd__nor2_1 U25780 ( .A(n20345), .B(n19666), .Y(n19376) );
  sky130_fd_sc_hd__nand2_1 U25781 ( .A(n19377), .B(n19376), .Y(n19378) );
  sky130_fd_sc_hd__nand2_1 U25782 ( .A(n19378), .B(n20393), .Y(n19384) );
  sky130_fd_sc_hd__nand3b_1 U25783 ( .A_N(n20345), .B(n20364), .C(n19575), .Y(
        n19379) );
  sky130_fd_sc_hd__nor2_1 U25784 ( .A(n19579), .B(n19379), .Y(n19618) );
  sky130_fd_sc_hd__nand4_1 U25785 ( .A(n20307), .B(n20387), .C(n19571), .D(
        n19397), .Y(n19380) );
  sky130_fd_sc_hd__nor3_1 U25786 ( .A(n19655), .B(n19380), .C(n20395), .Y(
        n19381) );
  sky130_fd_sc_hd__nand2_1 U25787 ( .A(n19618), .B(n19381), .Y(n19382) );
  sky130_fd_sc_hd__nand2_1 U25788 ( .A(n19382), .B(n20374), .Y(n19383) );
  sky130_fd_sc_hd__nand4_1 U25789 ( .A(n19386), .B(n19385), .C(n19384), .D(
        n19383), .Y(n19387) );
  sky130_fd_sc_hd__nand2_1 U25790 ( .A(n19387), .B(n20617), .Y(n19421) );
  sky130_fd_sc_hd__nand3_1 U25791 ( .A(n19610), .B(n19575), .C(n20389), .Y(
        n19388) );
  sky130_fd_sc_hd__nor2_1 U25792 ( .A(n19388), .B(n20282), .Y(n19647) );
  sky130_fd_sc_hd__nand4_1 U25793 ( .A(n20392), .B(n20390), .C(n20339), .D(
        n20387), .Y(n19389) );
  sky130_fd_sc_hd__nor2_1 U25794 ( .A(n19643), .B(n19389), .Y(n19390) );
  sky130_fd_sc_hd__nand2_1 U25795 ( .A(n19647), .B(n19390), .Y(n19391) );
  sky130_fd_sc_hd__nand2_1 U25796 ( .A(n19391), .B(n20393), .Y(n19410) );
  sky130_fd_sc_hd__nor3_1 U25797 ( .A(n19615), .B(n19392), .C(n20381), .Y(
        n19393) );
  sky130_fd_sc_hd__nand4_1 U25798 ( .A(n19618), .B(n20317), .C(n20271), .D(
        n19393), .Y(n19396) );
  sky130_fd_sc_hd__o2bb2ai_1 U25799 ( .B1(n19394), .B2(n20372), .A1_N(n19394), 
        .A2_N(n20278), .Y(n19395) );
  sky130_fd_sc_hd__a21oi_1 U25800 ( .A1(n19396), .A2(n20374), .B1(n19395), .Y(
        n19409) );
  sky130_fd_sc_hd__o211ai_1 U25801 ( .A1(n20515), .A2(n20043), .B1(n19397), 
        .C1(n20389), .Y(n19399) );
  sky130_fd_sc_hd__nor2_1 U25802 ( .A(n19399), .B(n19398), .Y(n19401) );
  sky130_fd_sc_hd__nand2_1 U25803 ( .A(n20360), .B(n20390), .Y(n19644) );
  sky130_fd_sc_hd__nor2_1 U25804 ( .A(n19644), .B(n20381), .Y(n19400) );
  sky130_fd_sc_hd__nand4_1 U25805 ( .A(n19565), .B(n19402), .C(n19401), .D(
        n19400), .Y(n19403) );
  sky130_fd_sc_hd__nand2_1 U25806 ( .A(n19403), .B(n20385), .Y(n19408) );
  sky130_fd_sc_hd__nand3_1 U25807 ( .A(n20360), .B(n19562), .C(n20292), .Y(
        n19406) );
  sky130_fd_sc_hd__nand3_1 U25808 ( .A(n19565), .B(n19660), .C(n19405), .Y(
        n19671) );
  sky130_fd_sc_hd__o21ai_1 U25809 ( .A1(n19406), .A2(n19671), .B1(n20368), .Y(
        n19407) );
  sky130_fd_sc_hd__nand4_1 U25810 ( .A(n19410), .B(n19409), .C(n19408), .D(
        n19407), .Y(n19411) );
  sky130_fd_sc_hd__nand2_1 U25811 ( .A(n19411), .B(n20784), .Y(n19423) );
  sky130_fd_sc_hd__nand2_1 U25812 ( .A(j202_soc_core_memory0_ram_dout0[481]), 
        .B(n21650), .Y(n19427) );
  sky130_fd_sc_hd__nand4_1 U25813 ( .A(n19417), .B(n19416), .C(n21653), .D(
        n19415), .Y(n19419) );
  sky130_fd_sc_hd__nor3_1 U25814 ( .A(n19420), .B(n19419), .C(n19418), .Y(
        n19422) );
  sky130_fd_sc_hd__nand3_1 U25815 ( .A(n19423), .B(n19422), .C(n19421), .Y(
        n19424) );
  sky130_fd_sc_hd__nor2_1 U25816 ( .A(n19425), .B(n19424), .Y(n19426) );
  sky130_fd_sc_hd__nand2_1 U25817 ( .A(n19427), .B(n19426), .Y(n19428) );
  sky130_fd_sc_hd__nand3_1 U25818 ( .A(n19429), .B(
        j202_soc_core_j22_cpu_ifetchl), .C(n19539), .Y(n19430) );
  sky130_fd_sc_hd__nand2_1 U25819 ( .A(j202_soc_core_memory0_ram_dout0[81]), 
        .B(n20458), .Y(n19431) );
  sky130_fd_sc_hd__nand2_1 U25820 ( .A(n19763), .B(n19432), .Y(n19433) );
  sky130_fd_sc_hd__nor2_1 U25821 ( .A(n19507), .B(n19433), .Y(n19745) );
  sky130_fd_sc_hd__nand2_1 U25822 ( .A(n19745), .B(n19694), .Y(n19438) );
  sky130_fd_sc_hd__nor2_1 U25823 ( .A(n19435), .B(n19434), .Y(n19436) );
  sky130_fd_sc_hd__nand2_1 U25824 ( .A(n19437), .B(n19436), .Y(n19805) );
  sky130_fd_sc_hd__nand2_1 U25826 ( .A(n19522), .B(n19810), .Y(n19494) );
  sky130_fd_sc_hd__nand4_1 U25827 ( .A(n19440), .B(n19439), .C(n19813), .D(
        n19764), .Y(n19443) );
  sky130_fd_sc_hd__nand3_1 U25828 ( .A(n19768), .B(n19441), .C(n19517), .Y(
        n19442) );
  sky130_fd_sc_hd__o21ai_1 U25829 ( .A1(n19443), .A2(n19442), .B1(n21103), .Y(
        n19454) );
  sky130_fd_sc_hd__nor3_1 U25830 ( .A(n19444), .B(n19507), .C(n19494), .Y(
        n19445) );
  sky130_fd_sc_hd__nand4_1 U25831 ( .A(n19513), .B(n19446), .C(n19445), .D(
        n19754), .Y(n19447) );
  sky130_fd_sc_hd__nand2_1 U25832 ( .A(n19447), .B(n17237), .Y(n19453) );
  sky130_fd_sc_hd__nor2_1 U25833 ( .A(n19448), .B(n19819), .Y(n19449) );
  sky130_fd_sc_hd__nand4_1 U25834 ( .A(n19450), .B(n19512), .C(n19720), .D(
        n19449), .Y(n19451) );
  sky130_fd_sc_hd__nand2_1 U25835 ( .A(n19451), .B(n19804), .Y(n19452) );
  sky130_fd_sc_hd__nand4_1 U25836 ( .A(n19455), .B(n19454), .C(n19453), .D(
        n19452), .Y(n19456) );
  sky130_fd_sc_hd__nand2_1 U25837 ( .A(n19456), .B(n20194), .Y(n19534) );
  sky130_fd_sc_hd__nand2_1 U25838 ( .A(n19783), .B(n19714), .Y(n19458) );
  sky130_fd_sc_hd__nand3b_1 U25839 ( .A_N(n19470), .B(n19701), .C(n19728), .Y(
        n19457) );
  sky130_fd_sc_hd__nor2_1 U25840 ( .A(n19458), .B(n19457), .Y(n19519) );
  sky130_fd_sc_hd__nand2_1 U25841 ( .A(n19813), .B(n19777), .Y(n19460) );
  sky130_fd_sc_hd__nand4_1 U25842 ( .A(n19765), .B(n19764), .C(n19781), .D(
        n19809), .Y(n19459) );
  sky130_fd_sc_hd__nor2_1 U25843 ( .A(n19460), .B(n19459), .Y(n19461) );
  sky130_fd_sc_hd__nand3_1 U25844 ( .A(n19519), .B(n19768), .C(n19461), .Y(
        n19462) );
  sky130_fd_sc_hd__nand2_1 U25845 ( .A(n19462), .B(n19804), .Y(n19479) );
  sky130_fd_sc_hd__nand2_1 U25846 ( .A(n19734), .B(n19463), .Y(n19464) );
  sky130_fd_sc_hd__nor2_1 U25847 ( .A(n19465), .B(n19464), .Y(n19466) );
  sky130_fd_sc_hd__nand4_1 U25848 ( .A(n19467), .B(n19466), .C(n19813), .D(
        n19523), .Y(n19469) );
  sky130_fd_sc_hd__a2bb2oi_1 U25849 ( .B1(n21103), .B2(n19469), .A1_N(n19468), 
        .A2_N(n19781), .Y(n19478) );
  sky130_fd_sc_hd__nor2_1 U25850 ( .A(n19470), .B(n19698), .Y(n19471) );
  sky130_fd_sc_hd__nand3_1 U25851 ( .A(n19472), .B(n19719), .C(n19471), .Y(
        n19473) );
  sky130_fd_sc_hd__nand2_1 U25852 ( .A(n19473), .B(n19816), .Y(n19477) );
  sky130_fd_sc_hd__nand3_1 U25853 ( .A(n19814), .B(n19715), .C(n19782), .Y(
        n19475) );
  sky130_fd_sc_hd__o21ai_1 U25854 ( .A1(n19475), .A2(n19474), .B1(n17237), .Y(
        n19476) );
  sky130_fd_sc_hd__nand4_1 U25855 ( .A(n19479), .B(n19478), .C(n19477), .D(
        n19476), .Y(n19503) );
  sky130_fd_sc_hd__nand2_1 U25856 ( .A(n19481), .B(n19480), .Y(n19704) );
  sky130_fd_sc_hd__o31a_1 U25858 ( .A1(n19484), .A2(n19483), .A3(n19821), .B1(
        n19816), .X(n19485) );
  sky130_fd_sc_hd__a21oi_1 U25859 ( .A1(n19487), .A2(n19486), .B1(n19485), .Y(
        n19500) );
  sky130_fd_sc_hd__nand2_1 U25860 ( .A(n19738), .B(n19523), .Y(n19488) );
  sky130_fd_sc_hd__nor2_1 U25861 ( .A(n19488), .B(n19698), .Y(n19787) );
  sky130_fd_sc_hd__nand2_1 U25862 ( .A(n19801), .B(n19810), .Y(n19489) );
  sky130_fd_sc_hd__nor2_1 U25863 ( .A(n19797), .B(n19489), .Y(n19492) );
  sky130_fd_sc_hd__nand2_1 U25864 ( .A(n19812), .B(n19490), .Y(n19491) );
  sky130_fd_sc_hd__nor2_1 U25865 ( .A(n19491), .B(n19699), .Y(n19730) );
  sky130_fd_sc_hd__nand3_1 U25866 ( .A(n19787), .B(n19492), .C(n19730), .Y(
        n19493) );
  sky130_fd_sc_hd__nand2_1 U25867 ( .A(n19493), .B(n17237), .Y(n19499) );
  sky130_fd_sc_hd__nor2_1 U25868 ( .A(n19494), .B(n19798), .Y(n19495) );
  sky130_fd_sc_hd__nand4_1 U25869 ( .A(n19496), .B(n19739), .C(n19495), .D(
        n19755), .Y(n19497) );
  sky130_fd_sc_hd__nand2_1 U25870 ( .A(n19497), .B(n21103), .Y(n19498) );
  sky130_fd_sc_hd__nand4_1 U25871 ( .A(n19501), .B(n19500), .C(n19499), .D(
        n19498), .Y(n19502) );
  sky130_fd_sc_hd__a22oi_1 U25872 ( .A1(n19503), .A2(n20235), .B1(n19502), 
        .B2(n20196), .Y(n19533) );
  sky130_fd_sc_hd__nand2_1 U25873 ( .A(n19505), .B(n19504), .Y(n19506) );
  sky130_fd_sc_hd__nand4b_1 U25874 ( .A_N(n19507), .B(n19809), .C(n19706), .D(
        n19506), .Y(n19508) );
  sky130_fd_sc_hd__nor2_1 U25875 ( .A(n19509), .B(n19508), .Y(n19510) );
  sky130_fd_sc_hd__nand4_1 U25876 ( .A(n19720), .B(n19510), .C(n19734), .D(
        n19701), .Y(n19515) );
  sky130_fd_sc_hd__nand3_1 U25877 ( .A(n19513), .B(n19512), .C(n19746), .Y(
        n19514) );
  sky130_fd_sc_hd__nor2_1 U25878 ( .A(n19515), .B(n19514), .Y(n19530) );
  sky130_fd_sc_hd__o21ai_0 U25879 ( .A1(n19516), .A2(n19696), .B1(n21103), .Y(
        n19529) );
  sky130_fd_sc_hd__nand4_1 U25880 ( .A(n19519), .B(n19518), .C(n19825), .D(
        n19517), .Y(n19527) );
  sky130_fd_sc_hd__nand2_1 U25881 ( .A(n19811), .B(n19753), .Y(n19520) );
  sky130_fd_sc_hd__nor2_1 U25882 ( .A(n19521), .B(n19520), .Y(n19829) );
  sky130_fd_sc_hd__nand4_1 U25883 ( .A(n19829), .B(n19809), .C(n19522), .D(
        n19743), .Y(n19525) );
  sky130_fd_sc_hd__nand3_1 U25884 ( .A(n19773), .B(n19714), .C(n19523), .Y(
        n19524) );
  sky130_fd_sc_hd__o31a_1 U25885 ( .A1(n19779), .A2(n19525), .A3(n19524), .B1(
        n19804), .X(n19526) );
  sky130_fd_sc_hd__a21oi_1 U25886 ( .A1(n19527), .A2(n17237), .B1(n19526), .Y(
        n19528) );
  sky130_fd_sc_hd__nand2_1 U25888 ( .A(n19531), .B(n20126), .Y(n19532) );
  sky130_fd_sc_hd__nand3_1 U25889 ( .A(n19534), .B(n19533), .C(n19532), .Y(
        n19538) );
  sky130_fd_sc_hd__a22oi_1 U25890 ( .A1(n21516), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[17]), .B1(n20540), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[49]), .Y(n19536) );
  sky130_fd_sc_hd__a22oi_1 U25891 ( .A1(n20759), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[81]), .B1(n21513), .B2(
        j202_soc_core_uart_div1[1]), .Y(n19535) );
  sky130_fd_sc_hd__o211ai_1 U25892 ( .A1(n25759), .A2(n21517), .B1(n19536), 
        .C1(n19535), .Y(n19537) );
  sky130_fd_sc_hd__a21oi_1 U25893 ( .A1(n19538), .A2(n21629), .B1(n19537), .Y(
        n21933) );
  sky130_fd_sc_hd__nand2_1 U25894 ( .A(n19539), .B(
        j202_soc_core_j22_cpu_id_opn_v_), .Y(n19857) );
  sky130_fd_sc_hd__a22oi_1 U25895 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__1_), .B1(n21916), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__1_), .Y(n19540) );
  sky130_fd_sc_hd__nand3_1 U25898 ( .A(n19544), .B(n20390), .C(n20344), .Y(
        n19545) );
  sky130_fd_sc_hd__nor2_1 U25899 ( .A(n20350), .B(n19545), .Y(n19547) );
  sky130_fd_sc_hd__nand3_1 U25900 ( .A(n19547), .B(n19546), .C(n19572), .Y(
        n19548) );
  sky130_fd_sc_hd__o21ai_0 U25901 ( .A1(n20282), .A2(n19548), .B1(n20368), .Y(
        n19570) );
  sky130_fd_sc_hd__nand2_1 U25902 ( .A(n20349), .B(n19549), .Y(n19550) );
  sky130_fd_sc_hd__nor2_1 U25903 ( .A(n19550), .B(n20278), .Y(n19551) );
  sky130_fd_sc_hd__nand3_1 U25904 ( .A(n19552), .B(n20280), .C(n19551), .Y(
        n19553) );
  sky130_fd_sc_hd__nand2_1 U25906 ( .A(n20363), .B(n19575), .Y(n20294) );
  sky130_fd_sc_hd__nor2_1 U25907 ( .A(n19555), .B(n19554), .Y(n19556) );
  sky130_fd_sc_hd__nand3_1 U25908 ( .A(n19558), .B(n19557), .C(n19556), .Y(
        n19560) );
  sky130_fd_sc_hd__a21oi_1 U25909 ( .A1(n19560), .A2(n20374), .B1(n19559), .Y(
        n19568) );
  sky130_fd_sc_hd__nand2b_1 U25910 ( .A_N(n19561), .B(n20371), .Y(n19667) );
  sky130_fd_sc_hd__nor2_1 U25911 ( .A(n19667), .B(n20270), .Y(n19563) );
  sky130_fd_sc_hd__nand4_1 U25912 ( .A(n19565), .B(n19564), .C(n19563), .D(
        n20363), .Y(n19566) );
  sky130_fd_sc_hd__nand2_1 U25913 ( .A(n19566), .B(n20385), .Y(n19567) );
  sky130_fd_sc_hd__nand4_1 U25914 ( .A(n19570), .B(n19569), .C(n19568), .D(
        n19567), .Y(n19592) );
  sky130_fd_sc_hd__nand4_1 U25915 ( .A(n19647), .B(n20311), .C(n19572), .D(
        n19571), .Y(n19573) );
  sky130_fd_sc_hd__nand2_1 U25916 ( .A(n19573), .B(n20385), .Y(n19590) );
  sky130_fd_sc_hd__nand2_1 U25917 ( .A(n19575), .B(n20333), .Y(n19577) );
  sky130_fd_sc_hd__nor2_1 U25918 ( .A(n19577), .B(n19576), .Y(n20330) );
  sky130_fd_sc_hd__nand4_1 U25919 ( .A(n20330), .B(n19657), .C(n19612), .D(
        n20348), .Y(n19578) );
  sky130_fd_sc_hd__nand2_1 U25920 ( .A(n19578), .B(n20393), .Y(n19589) );
  sky130_fd_sc_hd__nor3_1 U25921 ( .A(n19581), .B(n19580), .C(n19579), .Y(
        n19582) );
  sky130_fd_sc_hd__nand3_1 U25922 ( .A(n19617), .B(n19582), .C(n20280), .Y(
        n19583) );
  sky130_fd_sc_hd__nand2_1 U25923 ( .A(n19583), .B(n20368), .Y(n19588) );
  sky130_fd_sc_hd__nand4_1 U25924 ( .A(n19585), .B(n20343), .C(n19642), .D(
        n20338), .Y(n19586) );
  sky130_fd_sc_hd__o21ai_0 U25925 ( .A1(n19586), .A2(n20282), .B1(n20374), .Y(
        n19587) );
  sky130_fd_sc_hd__nand4_1 U25926 ( .A(n19590), .B(n19589), .C(n19588), .D(
        n19587), .Y(n19591) );
  sky130_fd_sc_hd__a22oi_1 U25927 ( .A1(n20757), .A2(n19592), .B1(n19591), 
        .B2(n20617), .Y(n19687) );
  sky130_fd_sc_hd__nand2_1 U25928 ( .A(n28203), .B(n28202), .Y(n28161) );
  sky130_fd_sc_hd__nand2_1 U25929 ( .A(n19594), .B(n19593), .Y(n19597) );
  sky130_fd_sc_hd__nor2_1 U25930 ( .A(n28161), .B(n19597), .Y(n27696) );
  sky130_fd_sc_hd__nand3_1 U25931 ( .A(n27696), .B(n29435), .C(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_), .Y(n19604) );
  sky130_fd_sc_hd__a2bb2oi_1 U25932 ( .B1(n19596), .B2(
        j202_soc_core_bldc_core_00_pwm_en), .A1_N(n29126), .A2_N(n19595), .Y(
        n19603) );
  sky130_fd_sc_hd__nand3_1 U25933 ( .A(n19599), .B(n19598), .C(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_0_), .Y(n27703) );
  sky130_fd_sc_hd__nand2_1 U25934 ( .A(n19601), .B(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[0]), .Y(n19602) );
  sky130_fd_sc_hd__nand4_1 U25935 ( .A(n19604), .B(n19603), .C(n27703), .D(
        n19602), .Y(n19606) );
  sky130_fd_sc_hd__nand2_1 U25936 ( .A(n19606), .B(n19605), .Y(n19633) );
  sky130_fd_sc_hd__nand2_1 U25937 ( .A(n21446), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[96]), .Y(n19632) );
  sky130_fd_sc_hd__nor3_1 U25938 ( .A(n19608), .B(n19615), .C(n19607), .Y(
        n19609) );
  sky130_fd_sc_hd__nand4_1 U25939 ( .A(n19610), .B(n19609), .C(n20366), .D(
        n19623), .Y(n19611) );
  sky130_fd_sc_hd__o21ai_1 U25940 ( .A1(n20282), .A2(n19611), .B1(n20393), .Y(
        n19629) );
  sky130_fd_sc_hd__nand3_1 U25941 ( .A(n20307), .B(n20339), .C(n19612), .Y(
        n19614) );
  sky130_fd_sc_hd__nor3_1 U25942 ( .A(n19615), .B(n19614), .C(n19613), .Y(
        n19616) );
  sky130_fd_sc_hd__nand3_1 U25943 ( .A(n19618), .B(n19617), .C(n19616), .Y(
        n19619) );
  sky130_fd_sc_hd__nand2_1 U25944 ( .A(n19619), .B(n20385), .Y(n19628) );
  sky130_fd_sc_hd__o21ai_1 U25945 ( .A1(n19621), .A2(n19620), .B1(n20374), .Y(
        n19627) );
  sky130_fd_sc_hd__nand3_1 U25946 ( .A(n19624), .B(n19623), .C(n19622), .Y(
        n19625) );
  sky130_fd_sc_hd__nand2_1 U25947 ( .A(n19625), .B(n20368), .Y(n19626) );
  sky130_fd_sc_hd__nand4_1 U25948 ( .A(n19629), .B(n19628), .C(n19627), .D(
        n19626), .Y(n19630) );
  sky130_fd_sc_hd__nand2_1 U25949 ( .A(n19630), .B(n20643), .Y(n19631) );
  sky130_fd_sc_hd__nand3_1 U25950 ( .A(n19633), .B(n19632), .C(n19631), .Y(
        n19689) );
  sky130_fd_sc_hd__nand2_1 U25951 ( .A(n21504), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[8]), .Y(n19637) );
  sky130_fd_sc_hd__nand2_1 U25952 ( .A(n24720), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[16]), .Y(n19636) );
  sky130_fd_sc_hd__nand2_1 U25953 ( .A(n21505), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[0]), .Y(n19635) );
  sky130_fd_sc_hd__nand2_1 U25954 ( .A(n21506), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[24]), .Y(n19634) );
  sky130_fd_sc_hd__nand4_1 U25955 ( .A(n19637), .B(n19636), .C(n19635), .D(
        n19634), .Y(n19639) );
  sky130_fd_sc_hd__a2bb2oi_1 U25956 ( .B1(n19639), .B2(n21513), .A1_N(n21515), 
        .A2_N(n19638), .Y(n19680) );
  sky130_fd_sc_hd__nand2_1 U25957 ( .A(n20759), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[64]), .Y(n19679) );
  sky130_fd_sc_hd__nand2_1 U25958 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[0]), .Y(n19678) );
  sky130_fd_sc_hd__nand4_1 U25959 ( .A(n19680), .B(n21768), .C(n19679), .D(
        n19678), .Y(n19640) );
  sky130_fd_sc_hd__nor2_1 U25960 ( .A(n28228), .B(n21517), .Y(n19683) );
  sky130_fd_sc_hd__nor2_1 U25961 ( .A(n19640), .B(n19683), .Y(n19676) );
  sky130_fd_sc_hd__nand2_1 U25962 ( .A(n19642), .B(n19641), .Y(n19645) );
  sky130_fd_sc_hd__nor3_1 U25963 ( .A(n19645), .B(n19644), .C(n19643), .Y(
        n19646) );
  sky130_fd_sc_hd__nand2_1 U25964 ( .A(n19647), .B(n19646), .Y(n19648) );
  sky130_fd_sc_hd__nand2_1 U25965 ( .A(n19648), .B(n20385), .Y(n19674) );
  sky130_fd_sc_hd__nand4_1 U25966 ( .A(n20310), .B(n19649), .C(n20292), .D(
        n20364), .Y(n19650) );
  sky130_fd_sc_hd__nor3_1 U25967 ( .A(n20312), .B(n19651), .C(n19650), .Y(
        n19653) );
  sky130_fd_sc_hd__nand2_1 U25968 ( .A(n19653), .B(n19652), .Y(n19663) );
  sky130_fd_sc_hd__nor2_1 U25969 ( .A(n19655), .B(n19654), .Y(n19658) );
  sky130_fd_sc_hd__nand4_1 U25970 ( .A(n19658), .B(n19657), .C(n19656), .D(
        n20387), .Y(n19661) );
  sky130_fd_sc_hd__nand3_1 U25971 ( .A(n19660), .B(n19659), .C(n20364), .Y(
        n20341) );
  sky130_fd_sc_hd__o31a_1 U25972 ( .A1(n19664), .A2(n19661), .A3(n20341), .B1(
        n20393), .X(n19662) );
  sky130_fd_sc_hd__a21oi_1 U25973 ( .A1(n20374), .A2(n19663), .B1(n19662), .Y(
        n19673) );
  sky130_fd_sc_hd__nor2_1 U25974 ( .A(n19665), .B(n19664), .Y(n20319) );
  sky130_fd_sc_hd__nand3_1 U25975 ( .A(n20319), .B(n19669), .C(n19668), .Y(
        n19670) );
  sky130_fd_sc_hd__nand3_1 U25977 ( .A(n19674), .B(n19673), .C(n19672), .Y(
        n19675) );
  sky130_fd_sc_hd__nand2_1 U25978 ( .A(n19675), .B(n20784), .Y(n19685) );
  sky130_fd_sc_hd__nand2_1 U25979 ( .A(j202_soc_core_memory0_ram_dout0[480]), 
        .B(n21650), .Y(n19691) );
  sky130_fd_sc_hd__nand3_1 U25980 ( .A(n19679), .B(n21653), .C(n19678), .Y(
        n19682) );
  sky130_fd_sc_hd__nor2_1 U25981 ( .A(n19682), .B(n19681), .Y(n19686) );
  sky130_fd_sc_hd__nand4_1 U25982 ( .A(n19687), .B(n19686), .C(n19685), .D(
        n19684), .Y(n19688) );
  sky130_fd_sc_hd__nor2_1 U25983 ( .A(n19689), .B(n19688), .Y(n19690) );
  sky130_fd_sc_hd__nand2_1 U25984 ( .A(n19691), .B(n19690), .Y(n19692) );
  sky130_fd_sc_hd__nand4_1 U25985 ( .A(n19695), .B(n19811), .C(n19694), .D(
        n19693), .Y(n19697) );
  sky130_fd_sc_hd__nor3_1 U25986 ( .A(n19698), .B(n19697), .C(n19696), .Y(
        n19727) );
  sky130_fd_sc_hd__nor2_1 U25987 ( .A(n19699), .B(n19821), .Y(n19703) );
  sky130_fd_sc_hd__nand4_1 U25988 ( .A(n19703), .B(n19702), .C(n19783), .D(
        n19701), .Y(n19705) );
  sky130_fd_sc_hd__o21ai_1 U25989 ( .A1(n19705), .A2(n19704), .B1(n21103), .Y(
        n19725) );
  sky130_fd_sc_hd__nand3_1 U25990 ( .A(n19734), .B(n19707), .C(n19706), .Y(
        n19709) );
  sky130_fd_sc_hd__nor3_1 U25991 ( .A(n19733), .B(n19709), .C(n19708), .Y(
        n19710) );
  sky130_fd_sc_hd__nand2_1 U25992 ( .A(n19711), .B(n19710), .Y(n19723) );
  sky130_fd_sc_hd__nand4_1 U25993 ( .A(n19715), .B(n19714), .C(n19713), .D(
        n19734), .Y(n19717) );
  sky130_fd_sc_hd__nor2_1 U25994 ( .A(n19717), .B(n19716), .Y(n19718) );
  sky130_fd_sc_hd__nand4_1 U25995 ( .A(n19721), .B(n19720), .C(n19719), .D(
        n19718), .Y(n19722) );
  sky130_fd_sc_hd__a22oi_1 U25996 ( .A1(n19723), .A2(n19804), .B1(n19722), 
        .B2(n17237), .Y(n19724) );
  sky130_fd_sc_hd__nand4_1 U25997 ( .A(n19730), .B(n19811), .C(n19729), .D(
        n19728), .Y(n19731) );
  sky130_fd_sc_hd__nand2_1 U25998 ( .A(n19731), .B(n17237), .Y(n19752) );
  sky130_fd_sc_hd__and4_1 U25999 ( .A(n19740), .B(n19783), .C(n19770), .D(
        n19734), .X(n19735) );
  sky130_fd_sc_hd__nand4_1 U26000 ( .A(n19736), .B(n19825), .C(n19823), .D(
        n19735), .Y(n19737) );
  sky130_fd_sc_hd__nand2_1 U26001 ( .A(n19737), .B(n19816), .Y(n19751) );
  sky130_fd_sc_hd__nand4_1 U26002 ( .A(n19740), .B(n19739), .C(n19781), .D(
        n19738), .Y(n19741) );
  sky130_fd_sc_hd__o21ai_1 U26003 ( .A1(n19742), .A2(n19741), .B1(n19804), .Y(
        n19750) );
  sky130_fd_sc_hd__nand4_1 U26004 ( .A(n19813), .B(n19770), .C(n19782), .D(
        n19743), .Y(n19747) );
  sky130_fd_sc_hd__nand4b_1 U26005 ( .A_N(n19747), .B(n19746), .C(n19745), .D(
        n19744), .Y(n19748) );
  sky130_fd_sc_hd__nand2_1 U26006 ( .A(n19748), .B(n21103), .Y(n19749) );
  sky130_fd_sc_hd__nand4_1 U26007 ( .A(n19752), .B(n19751), .C(n19750), .D(
        n19749), .Y(n19794) );
  sky130_fd_sc_hd__nand3_1 U26008 ( .A(n19754), .B(n19753), .C(n19782), .Y(
        n19757) );
  sky130_fd_sc_hd__nand2_1 U26009 ( .A(n19813), .B(n19755), .Y(n19756) );
  sky130_fd_sc_hd__nor2_1 U26010 ( .A(n19757), .B(n19756), .Y(n19758) );
  sky130_fd_sc_hd__nand3_1 U26011 ( .A(n19759), .B(n19768), .C(n19758), .Y(
        n19760) );
  sky130_fd_sc_hd__nand2_1 U26012 ( .A(n19760), .B(n19804), .Y(n19792) );
  sky130_fd_sc_hd__and4_1 U26013 ( .A(n19765), .B(n19764), .C(n19763), .D(
        n19762), .X(n19766) );
  sky130_fd_sc_hd__nand4_1 U26014 ( .A(n19768), .B(n19823), .C(n19767), .D(
        n19766), .Y(n19769) );
  sky130_fd_sc_hd__nand2_1 U26015 ( .A(n19769), .B(n17237), .Y(n19791) );
  sky130_fd_sc_hd__and3_1 U26016 ( .A(n19801), .B(n19771), .C(n19770), .X(
        n19772) );
  sky130_fd_sc_hd__nand4_1 U26017 ( .A(n19775), .B(n19774), .C(n19773), .D(
        n19772), .Y(n19776) );
  sky130_fd_sc_hd__nand2_1 U26018 ( .A(n19776), .B(n21103), .Y(n19790) );
  sky130_fd_sc_hd__nand2_1 U26019 ( .A(n19778), .B(n19777), .Y(n19780) );
  sky130_fd_sc_hd__nor2_1 U26020 ( .A(n19780), .B(n19779), .Y(n19786) );
  sky130_fd_sc_hd__nand2_1 U26021 ( .A(n19782), .B(n19781), .Y(n19799) );
  sky130_fd_sc_hd__nor2_1 U26022 ( .A(n19799), .B(n19784), .Y(n19785) );
  sky130_fd_sc_hd__nand4_1 U26023 ( .A(n19787), .B(n19786), .C(n19823), .D(
        n19785), .Y(n19788) );
  sky130_fd_sc_hd__nand2_1 U26024 ( .A(n19788), .B(n19816), .Y(n19789) );
  sky130_fd_sc_hd__nand4_1 U26025 ( .A(n19792), .B(n19791), .C(n19790), .D(
        n19789), .Y(n19793) );
  sky130_fd_sc_hd__a22oi_1 U26026 ( .A1(n19794), .A2(n20194), .B1(n19793), 
        .B2(n20126), .Y(n19838) );
  sky130_fd_sc_hd__nor2_1 U26027 ( .A(n19796), .B(n19795), .Y(n19803) );
  sky130_fd_sc_hd__nor2_1 U26028 ( .A(n19799), .B(n19798), .Y(n19800) );
  sky130_fd_sc_hd__nand4_1 U26029 ( .A(n19803), .B(n19802), .C(n19801), .D(
        n19800), .Y(n19806) );
  sky130_fd_sc_hd__o21ai_1 U26030 ( .A1(n19806), .A2(n19805), .B1(n19804), .Y(
        n19835) );
  sky130_fd_sc_hd__nand4_1 U26031 ( .A(n19811), .B(n19810), .C(n19809), .D(
        n19808), .Y(n19815) );
  sky130_fd_sc_hd__nand4b_1 U26032 ( .A_N(n19815), .B(n19814), .C(n19813), .D(
        n19812), .Y(n19818) );
  sky130_fd_sc_hd__nor2_1 U26034 ( .A(n19820), .B(n19819), .Y(n19824) );
  sky130_fd_sc_hd__nand4_1 U26035 ( .A(n19825), .B(n19824), .C(n19823), .D(
        n19822), .Y(n19826) );
  sky130_fd_sc_hd__nand2_1 U26036 ( .A(n19826), .B(n17237), .Y(n19833) );
  sky130_fd_sc_hd__nand3_1 U26037 ( .A(n19830), .B(n19829), .C(n19828), .Y(
        n19831) );
  sky130_fd_sc_hd__nand2_1 U26038 ( .A(n19831), .B(n21103), .Y(n19832) );
  sky130_fd_sc_hd__nand4_1 U26039 ( .A(n19835), .B(n19834), .C(n19833), .D(
        n19832), .Y(n19836) );
  sky130_fd_sc_hd__nand2_1 U26040 ( .A(n19836), .B(n20196), .Y(n19837) );
  sky130_fd_sc_hd__o211ai_1 U26041 ( .A1(n19840), .A2(n19839), .B1(n19838), 
        .C1(n19837), .Y(n19841) );
  sky130_fd_sc_hd__nand2_1 U26042 ( .A(n19841), .B(n21629), .Y(n19845) );
  sky130_fd_sc_hd__a22oi_1 U26043 ( .A1(n21516), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[16]), .B1(n20759), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[80]), .Y(n19844) );
  sky130_fd_sc_hd__a22oi_1 U26044 ( .A1(n20540), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[48]), .B1(n21513), .B2(
        j202_soc_core_uart_div1[0]), .Y(n19843) );
  sky130_fd_sc_hd__nand2_1 U26045 ( .A(n20786), .B(
        j202_soc_core_bldc_core_00_pwm_duty[4]), .Y(n19842) );
  sky130_fd_sc_hd__nand4_1 U26046 ( .A(n19845), .B(n19844), .C(n19843), .D(
        n19842), .Y(n21691) );
  sky130_fd_sc_hd__a22oi_1 U26047 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__0_), .B1(n21916), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__0_), .Y(n19846) );
  sky130_fd_sc_hd__nand2_1 U26049 ( .A(j202_soc_core_memory0_ram_dout0[80]), 
        .B(n20458), .Y(n19848) );
  sky130_fd_sc_hd__nor2_1 U26051 ( .A(n19856), .B(n19857), .Y(n20885) );
  sky130_fd_sc_hd__nor2_1 U26052 ( .A(n19858), .B(n19857), .Y(n21173) );
  sky130_fd_sc_hd__nand3_1 U26054 ( .A(n19861), .B(n19860), .C(n19859), .Y(
        n19862) );
  sky130_fd_sc_hd__nand2_1 U26055 ( .A(j202_soc_core_memory0_ram_dout0[364]), 
        .B(n21495), .Y(n20915) );
  sky130_fd_sc_hd__nand3_1 U26056 ( .A(n20187), .B(n19897), .C(n20152), .Y(
        n19871) );
  sky130_fd_sc_hd__a31oi_1 U26057 ( .A1(n19877), .A2(n19863), .A3(n20181), 
        .B1(n19910), .Y(n19870) );
  sky130_fd_sc_hd__nand3b_1 U26058 ( .A_N(n20056), .B(n20020), .C(n20181), .Y(
        n19864) );
  sky130_fd_sc_hd__nand2_1 U26059 ( .A(n19864), .B(n20179), .Y(n19869) );
  sky130_fd_sc_hd__nand2_1 U26060 ( .A(n20215), .B(n20216), .Y(n19867) );
  sky130_fd_sc_hd__nand3_1 U26061 ( .A(n19866), .B(n21359), .C(n19865), .Y(
        n20204) );
  sky130_fd_sc_hd__nand3_1 U26062 ( .A(n20181), .B(n20113), .C(n20204), .Y(
        n20198) );
  sky130_fd_sc_hd__nand2_1 U26064 ( .A(n19869), .B(n19868), .Y(n20170) );
  sky130_fd_sc_hd__a211o_1 U26065 ( .A1(n20225), .A2(n19871), .B1(n19870), 
        .C1(n20170), .X(n19872) );
  sky130_fd_sc_hd__nand2_1 U26066 ( .A(n19872), .B(n20194), .Y(n19919) );
  sky130_fd_sc_hd__nand2_1 U26067 ( .A(n20000), .B(n20139), .Y(n19955) );
  sky130_fd_sc_hd__nor2_1 U26068 ( .A(n20015), .B(n19955), .Y(n20155) );
  sky130_fd_sc_hd__nand2_1 U26069 ( .A(n20128), .B(n20033), .Y(n20140) );
  sky130_fd_sc_hd__nand4_1 U26070 ( .A(n20155), .B(n19935), .C(n20003), .D(
        n20153), .Y(n19873) );
  sky130_fd_sc_hd__nand2_1 U26071 ( .A(n19873), .B(n20179), .Y(n19886) );
  sky130_fd_sc_hd__a21oi_1 U26072 ( .A1(n20199), .A2(
        j202_soc_core_bootrom_00_address_w[2]), .B1(n19874), .Y(n19875) );
  sky130_fd_sc_hd__nand2_1 U26073 ( .A(n20130), .B(n19875), .Y(n19878) );
  sky130_fd_sc_hd__nand3_1 U26074 ( .A(n19889), .B(n19877), .C(n19876), .Y(
        n20229) );
  sky130_fd_sc_hd__a22oi_1 U26075 ( .A1(n19878), .A2(n20227), .B1(n20229), 
        .B2(n20225), .Y(n19885) );
  sky130_fd_sc_hd__nor2_1 U26076 ( .A(n19880), .B(n19879), .Y(n19883) );
  sky130_fd_sc_hd__nand3_1 U26077 ( .A(n19883), .B(n20003), .C(n19882), .Y(
        n20188) );
  sky130_fd_sc_hd__nand2_1 U26078 ( .A(n20188), .B(n20210), .Y(n19884) );
  sky130_fd_sc_hd__nand3_1 U26079 ( .A(n19886), .B(n19885), .C(n19884), .Y(
        n19887) );
  sky130_fd_sc_hd__nand2_1 U26080 ( .A(n19887), .B(n20196), .Y(n19918) );
  sky130_fd_sc_hd__and3_1 U26081 ( .A(n20215), .B(n20000), .C(n20033), .X(
        n19888) );
  sky130_fd_sc_hd__nand4_1 U26082 ( .A(n20163), .B(n20186), .C(n19889), .D(
        n19888), .Y(n19890) );
  sky130_fd_sc_hd__nand2_1 U26083 ( .A(n19890), .B(n20227), .Y(n19901) );
  sky130_fd_sc_hd__nand4_1 U26084 ( .A(n19891), .B(n20000), .C(n20183), .D(
        n20204), .Y(n19893) );
  sky130_fd_sc_hd__nand3b_1 U26085 ( .A_N(n19893), .B(n19892), .C(n20186), .Y(
        n19894) );
  sky130_fd_sc_hd__nand2_1 U26086 ( .A(n19894), .B(n20225), .Y(n19900) );
  sky130_fd_sc_hd__nor2_1 U26087 ( .A(n20013), .B(n19981), .Y(n19896) );
  sky130_fd_sc_hd__nand4_1 U26088 ( .A(n20023), .B(n19896), .C(n20139), .D(
        n19895), .Y(n19898) );
  sky130_fd_sc_hd__nand3_1 U26089 ( .A(n19965), .B(n19897), .C(n20033), .Y(
        n20219) );
  sky130_fd_sc_hd__a22oi_1 U26090 ( .A1(n19898), .A2(n20210), .B1(n20219), 
        .B2(n20179), .Y(n19899) );
  sky130_fd_sc_hd__nand3_1 U26091 ( .A(n19901), .B(n19900), .C(n19899), .Y(
        n19902) );
  sky130_fd_sc_hd__nand2_1 U26092 ( .A(n19902), .B(n20235), .Y(n19917) );
  sky130_fd_sc_hd__nor2_1 U26093 ( .A(n19957), .B(n20046), .Y(n20108) );
  sky130_fd_sc_hd__nand2_1 U26094 ( .A(n20108), .B(n20102), .Y(n19907) );
  sky130_fd_sc_hd__nor2_1 U26095 ( .A(n20060), .B(n19956), .Y(n19950) );
  sky130_fd_sc_hd__nor2_1 U26096 ( .A(n19904), .B(n19903), .Y(n19906) );
  sky130_fd_sc_hd__nand3_1 U26097 ( .A(n19950), .B(n19906), .C(n19905), .Y(
        n20228) );
  sky130_fd_sc_hd__o21a_1 U26098 ( .A1(n19907), .A2(n20228), .B1(n20225), .X(
        n20110) );
  sky130_fd_sc_hd__and3_1 U26099 ( .A(n20167), .B(n20047), .C(n20052), .X(
        n20177) );
  sky130_fd_sc_hd__and3_1 U26100 ( .A(n19965), .B(n20216), .C(n20113), .X(
        n19908) );
  sky130_fd_sc_hd__a31oi_1 U26101 ( .A1(n20177), .A2(n20003), .A3(n19908), 
        .B1(n20038), .Y(n19914) );
  sky130_fd_sc_hd__nor2_1 U26102 ( .A(n20060), .B(n20046), .Y(n19909) );
  sky130_fd_sc_hd__a31oi_1 U26103 ( .A1(n20003), .A2(n19909), .A3(n20167), 
        .B1(n20200), .Y(n19913) );
  sky130_fd_sc_hd__nor4_1 U26104 ( .A(n20100), .B(n12841), .C(n20037), .D(
        n20140), .Y(n19911) );
  sky130_fd_sc_hd__nor2_1 U26105 ( .A(n19911), .B(n19910), .Y(n19912) );
  sky130_fd_sc_hd__nor4_1 U26106 ( .A(n20110), .B(n19914), .C(n19913), .D(
        n19912), .Y(n19915) );
  sky130_fd_sc_hd__nand2b_1 U26107 ( .A_N(n19915), .B(n20126), .Y(n19916) );
  sky130_fd_sc_hd__nand4_1 U26108 ( .A(n19919), .B(n19918), .C(n19917), .D(
        n19916), .Y(n19920) );
  sky130_fd_sc_hd__nand2_1 U26109 ( .A(n19920), .B(n21629), .Y(n20925) );
  sky130_fd_sc_hd__nand2b_1 U26110 ( .A_N(n21515), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[44]), .Y(n21817) );
  sky130_fd_sc_hd__nor2_1 U26111 ( .A(n19921), .B(n21519), .Y(n19929) );
  sky130_fd_sc_hd__nand2_1 U26112 ( .A(n19927), .B(n21768), .Y(n19922) );
  sky130_fd_sc_hd__nand2b_1 U26113 ( .A_N(n21512), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[76]), .Y(n21818) );
  sky130_fd_sc_hd__nand2_1 U26114 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[12]), .Y(n21815) );
  sky130_fd_sc_hd__nand2_1 U26115 ( .A(n21818), .B(n21815), .Y(n20923) );
  sky130_fd_sc_hd__nor3_1 U26116 ( .A(n19923), .B(n19922), .C(n20923), .Y(
        n19925) );
  sky130_fd_sc_hd__nor2_1 U26117 ( .A(n25182), .B(n21517), .Y(n21821) );
  sky130_fd_sc_hd__nand3_1 U26118 ( .A(n20925), .B(n19925), .C(n19924), .Y(
        n21826) );
  sky130_fd_sc_hd__nand2_1 U26119 ( .A(j202_soc_core_memory0_ram_dout0[460]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n20911) );
  sky130_fd_sc_hd__nand2_1 U26120 ( .A(j202_soc_core_memory0_ram_dout0[428]), 
        .B(n12156), .Y(n20910) );
  sky130_fd_sc_hd__nand2_1 U26122 ( .A(j202_soc_core_memory0_ram_dout0[12]), 
        .B(n21639), .Y(n20902) );
  sky130_fd_sc_hd__nand2_1 U26123 ( .A(j202_soc_core_memory0_ram_dout0[236]), 
        .B(n21641), .Y(n20901) );
  sky130_fd_sc_hd__nand2_1 U26124 ( .A(j202_soc_core_memory0_ram_dout0[172]), 
        .B(n21487), .Y(n20912) );
  sky130_fd_sc_hd__nand2_1 U26125 ( .A(j202_soc_core_memory0_ram_dout0[204]), 
        .B(n21640), .Y(n20907) );
  sky130_fd_sc_hd__nand2_1 U26126 ( .A(j202_soc_core_memory0_ram_dout0[76]), 
        .B(n21642), .Y(n20906) );
  sky130_fd_sc_hd__nand2_1 U26127 ( .A(j202_soc_core_memory0_ram_dout0[140]), 
        .B(n21489), .Y(n20905) );
  sky130_fd_sc_hd__nand4b_1 U26128 ( .A_N(n21821), .B(n19926), .C(n21816), .D(
        n21818), .Y(n19928) );
  sky130_fd_sc_hd__nand2_1 U26129 ( .A(n20925), .B(n19927), .Y(n21819) );
  sky130_fd_sc_hd__nor2_1 U26131 ( .A(n19929), .B(n21821), .Y(n20926) );
  sky130_fd_sc_hd__nand2_1 U26132 ( .A(n21817), .B(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n19930) );
  sky130_fd_sc_hd__nor2_1 U26133 ( .A(n19930), .B(n20923), .Y(n19931) );
  sky130_fd_sc_hd__nand3_1 U26134 ( .A(n20926), .B(n20925), .C(n19931), .Y(
        n19932) );
  sky130_fd_sc_hd__nor2_1 U26135 ( .A(n19932), .B(
        j202_soc_core_memory0_ram_dout0[492]), .Y(n21822) );
  sky130_fd_sc_hd__nor2_1 U26136 ( .A(n19933), .B(n21822), .Y(n19934) );
  sky130_fd_sc_hd__nand2_1 U26137 ( .A(n20047), .B(n20183), .Y(n20016) );
  sky130_fd_sc_hd__nand4_1 U26138 ( .A(n19935), .B(n20216), .C(n20000), .D(
        n20152), .Y(n19936) );
  sky130_fd_sc_hd__nor2_1 U26139 ( .A(n20016), .B(n19936), .Y(n20203) );
  sky130_fd_sc_hd__nand3_1 U26140 ( .A(n21097), .B(n19949), .C(n19951), .Y(
        n19939) );
  sky130_fd_sc_hd__nand2_1 U26141 ( .A(n19937), .B(n20128), .Y(n19938) );
  sky130_fd_sc_hd__nor2_1 U26142 ( .A(n19939), .B(n19938), .Y(n19940) );
  sky130_fd_sc_hd__nand4_1 U26143 ( .A(n20203), .B(n19940), .C(n20153), .D(
        n20214), .Y(n19941) );
  sky130_fd_sc_hd__nand2_1 U26144 ( .A(n19941), .B(n20179), .Y(n19964) );
  sky130_fd_sc_hd__nand4_1 U26145 ( .A(n20173), .B(n20058), .C(n19942), .D(
        n20002), .Y(n19944) );
  sky130_fd_sc_hd__nor2_1 U26146 ( .A(n19944), .B(n19943), .Y(n20143) );
  sky130_fd_sc_hd__nand2_1 U26147 ( .A(n20153), .B(n19949), .Y(n19945) );
  sky130_fd_sc_hd__nor2_1 U26148 ( .A(n20175), .B(n19945), .Y(n20149) );
  sky130_fd_sc_hd__nor2_1 U26149 ( .A(n19946), .B(n20060), .Y(n19947) );
  sky130_fd_sc_hd__nand4_1 U26150 ( .A(n20143), .B(n20149), .C(n19947), .D(
        n20181), .Y(n19948) );
  sky130_fd_sc_hd__nand2_1 U26151 ( .A(n19948), .B(n20225), .Y(n19963) );
  sky130_fd_sc_hd__nand4_1 U26152 ( .A(n20148), .B(n19950), .C(n20173), .D(
        n19949), .Y(n19954) );
  sky130_fd_sc_hd__nand4_1 U26153 ( .A(n20130), .B(n20000), .C(n19951), .D(
        n20052), .Y(n19952) );
  sky130_fd_sc_hd__nor2_1 U26154 ( .A(n20037), .B(n19952), .Y(n19979) );
  sky130_fd_sc_hd__o21ai_1 U26155 ( .A1(n19954), .A2(n19953), .B1(n20210), .Y(
        n19962) );
  sky130_fd_sc_hd__nor2_1 U26156 ( .A(n19957), .B(n19956), .Y(n19958) );
  sky130_fd_sc_hd__nand3_1 U26157 ( .A(n20021), .B(n19959), .C(n19958), .Y(
        n20136) );
  sky130_fd_sc_hd__nand4_1 U26158 ( .A(n20162), .B(n20119), .C(n19965), .D(
        n20058), .Y(n19960) );
  sky130_fd_sc_hd__o21ai_1 U26159 ( .A1(n20136), .A2(n19960), .B1(n20227), .Y(
        n19961) );
  sky130_fd_sc_hd__nand4_1 U26160 ( .A(n19964), .B(n19963), .C(n19962), .D(
        n19961), .Y(n19992) );
  sky130_fd_sc_hd__nand3_1 U26161 ( .A(n19996), .B(n19965), .C(n20003), .Y(
        n20164) );
  sky130_fd_sc_hd__nor2_1 U26162 ( .A(n19967), .B(n20060), .Y(n19968) );
  sky130_fd_sc_hd__nand4_1 U26163 ( .A(n20203), .B(n19968), .C(n20167), .D(
        n20139), .Y(n19969) );
  sky130_fd_sc_hd__nand3_1 U26165 ( .A(n20214), .B(n20216), .C(n20181), .Y(
        n19973) );
  sky130_fd_sc_hd__nand2_1 U26166 ( .A(n20108), .B(n19971), .Y(n19972) );
  sky130_fd_sc_hd__nor2_1 U26167 ( .A(n19973), .B(n19972), .Y(n19974) );
  sky130_fd_sc_hd__nand3_1 U26168 ( .A(n19996), .B(n20120), .C(n19974), .Y(
        n19975) );
  sky130_fd_sc_hd__nand2_1 U26169 ( .A(n19975), .B(n20179), .Y(n19989) );
  sky130_fd_sc_hd__nand2_1 U26170 ( .A(n20152), .B(n20128), .Y(n19977) );
  sky130_fd_sc_hd__nor2_1 U26171 ( .A(n19977), .B(n19976), .Y(n19978) );
  sky130_fd_sc_hd__nand4_1 U26172 ( .A(n19979), .B(n19978), .C(n20153), .D(
        n20181), .Y(n19980) );
  sky130_fd_sc_hd__nand2_1 U26173 ( .A(n19980), .B(n20227), .Y(n19988) );
  sky130_fd_sc_hd__nand3_1 U26174 ( .A(n20023), .B(n19982), .C(n19999), .Y(
        n20230) );
  sky130_fd_sc_hd__nand2_1 U26175 ( .A(n20000), .B(n20181), .Y(n20031) );
  sky130_fd_sc_hd__nand3_1 U26176 ( .A(n19985), .B(n19984), .C(n19983), .Y(
        n19986) );
  sky130_fd_sc_hd__nand3_1 U26177 ( .A(n20186), .B(n20173), .C(n20052), .Y(
        n20019) );
  sky130_fd_sc_hd__o21ai_1 U26178 ( .A1(n19986), .A2(n20019), .B1(n20210), .Y(
        n19987) );
  sky130_fd_sc_hd__nand4_1 U26179 ( .A(n19990), .B(n19989), .C(n19988), .D(
        n19987), .Y(n19991) );
  sky130_fd_sc_hd__a22o_1 U26180 ( .A1(n20235), .A2(n19992), .B1(n19991), .B2(
        n20194), .X(n20070) );
  sky130_fd_sc_hd__nand3_1 U26181 ( .A(n20128), .B(n20103), .C(n20129), .Y(
        n19994) );
  sky130_fd_sc_hd__nor2_1 U26182 ( .A(n19994), .B(n19993), .Y(n19995) );
  sky130_fd_sc_hd__nand3_1 U26183 ( .A(n19997), .B(n19996), .C(n19995), .Y(
        n19998) );
  sky130_fd_sc_hd__nand2_1 U26184 ( .A(n19998), .B(n20227), .Y(n20012) );
  sky130_fd_sc_hd__nand3_1 U26185 ( .A(n20000), .B(n19999), .C(n20052), .Y(
        n20221) );
  sky130_fd_sc_hd__nand4_1 U26186 ( .A(n20119), .B(n20185), .C(n20002), .D(
        n20001), .Y(n20004) );
  sky130_fd_sc_hd__nand3_1 U26187 ( .A(n20003), .B(n20118), .C(n20214), .Y(
        n20022) );
  sky130_fd_sc_hd__o21ai_1 U26188 ( .A1(n20004), .A2(n20022), .B1(n20210), .Y(
        n20011) );
  sky130_fd_sc_hd__nand3_1 U26189 ( .A(n20173), .B(n20033), .C(n20138), .Y(
        n20005) );
  sky130_fd_sc_hd__nor2_1 U26190 ( .A(n20005), .B(n20221), .Y(n20007) );
  sky130_fd_sc_hd__nand4_1 U26191 ( .A(n20008), .B(n20007), .C(n20006), .D(
        n20023), .Y(n20009) );
  sky130_fd_sc_hd__nand2_1 U26192 ( .A(n20009), .B(n20179), .Y(n20010) );
  sky130_fd_sc_hd__nand3_1 U26193 ( .A(n20012), .B(n20011), .C(n20010), .Y(
        n20018) );
  sky130_fd_sc_hd__nor2_1 U26194 ( .A(n20013), .B(n20136), .Y(n20050) );
  sky130_fd_sc_hd__nand2_1 U26195 ( .A(n20050), .B(n20014), .Y(n20105) );
  sky130_fd_sc_hd__o31a_1 U26196 ( .A1(n20016), .A2(n20015), .A3(n20105), .B1(
        n20225), .X(n20017) );
  sky130_fd_sc_hd__o21ai_1 U26197 ( .A1(n20018), .A2(n20017), .B1(n20196), .Y(
        n20068) );
  sky130_fd_sc_hd__nand3_1 U26198 ( .A(n20021), .B(n20020), .C(n20047), .Y(
        n20053) );
  sky130_fd_sc_hd__nand3_1 U26199 ( .A(n20023), .B(n20153), .C(n20102), .Y(
        n20025) );
  sky130_fd_sc_hd__nor2_1 U26200 ( .A(n20025), .B(n20024), .Y(n20026) );
  sky130_fd_sc_hd__nand4_1 U26201 ( .A(n20028), .B(n20209), .C(n20027), .D(
        n20026), .Y(n20042) );
  sky130_fd_sc_hd__nand3_1 U26202 ( .A(n20173), .B(n20030), .C(n20112), .Y(
        n20032) );
  sky130_fd_sc_hd__nor2_1 U26203 ( .A(n20032), .B(n20031), .Y(n20040) );
  sky130_fd_sc_hd__nor2_1 U26204 ( .A(n20036), .B(n20035), .Y(n20178) );
  sky130_fd_sc_hd__a31oi_1 U26205 ( .A1(n20040), .A2(n20178), .A3(n20039), 
        .B1(n20038), .Y(n20041) );
  sky130_fd_sc_hd__a21oi_1 U26206 ( .A1(n20042), .A2(n20225), .B1(n20041), .Y(
        n20065) );
  sky130_fd_sc_hd__and3_1 U26207 ( .A(n20215), .B(n20103), .C(n20058), .X(
        n20049) );
  sky130_fd_sc_hd__nor2_1 U26209 ( .A(n20046), .B(n20045), .Y(n20048) );
  sky130_fd_sc_hd__nand4_1 U26210 ( .A(n20050), .B(n20049), .C(n20048), .D(
        n20047), .Y(n20051) );
  sky130_fd_sc_hd__nand2_1 U26211 ( .A(n20051), .B(n20210), .Y(n20064) );
  sky130_fd_sc_hd__nand2_1 U26212 ( .A(n20172), .B(n20052), .Y(n20054) );
  sky130_fd_sc_hd__nor2_1 U26213 ( .A(n20054), .B(n20053), .Y(n20109) );
  sky130_fd_sc_hd__nand2_1 U26214 ( .A(n20145), .B(n20138), .Y(n20057) );
  sky130_fd_sc_hd__nor2_1 U26215 ( .A(n20057), .B(n20056), .Y(n20134) );
  sky130_fd_sc_hd__nand2_1 U26216 ( .A(n20058), .B(n20204), .Y(n20059) );
  sky130_fd_sc_hd__nor2_1 U26217 ( .A(n20060), .B(n20059), .Y(n20061) );
  sky130_fd_sc_hd__nand4_1 U26218 ( .A(n20109), .B(n20134), .C(n20061), .D(
        n20153), .Y(n20062) );
  sky130_fd_sc_hd__nand2_1 U26219 ( .A(n20062), .B(n20179), .Y(n20063) );
  sky130_fd_sc_hd__nand3_1 U26220 ( .A(n20065), .B(n20064), .C(n20063), .Y(
        n20066) );
  sky130_fd_sc_hd__nand2_1 U26221 ( .A(n20066), .B(n20126), .Y(n20067) );
  sky130_fd_sc_hd__nand2_1 U26222 ( .A(n20068), .B(n20067), .Y(n20069) );
  sky130_fd_sc_hd__o21a_1 U26223 ( .A1(n20070), .A2(n20069), .B1(n21629), .X(
        n20088) );
  sky130_fd_sc_hd__nand2b_1 U26224 ( .A_N(n21512), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[77]), .Y(n20953) );
  sky130_fd_sc_hd__nor2_1 U26225 ( .A(n20071), .B(n21515), .Y(n20077) );
  sky130_fd_sc_hd__nand2_1 U26226 ( .A(n20953), .B(n20072), .Y(n20074) );
  sky130_fd_sc_hd__nand2_1 U26227 ( .A(n21446), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[109]), .Y(n20082) );
  sky130_fd_sc_hd__nand2_1 U26228 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[13]), .Y(n20076) );
  sky130_fd_sc_hd__nand3_1 U26229 ( .A(n20082), .B(n21768), .C(n20076), .Y(
        n20073) );
  sky130_fd_sc_hd__nor2_1 U26230 ( .A(n20074), .B(n20073), .Y(n20075) );
  sky130_fd_sc_hd__nand2b_1 U26231 ( .A_N(n21517), .B(
        j202_soc_core_bldc_core_00_pwm_duty[1]), .Y(n20083) );
  sky130_fd_sc_hd__nand3_1 U26232 ( .A(n20957), .B(n20075), .C(n20083), .Y(
        n22225) );
  sky130_fd_sc_hd__nand3_1 U26233 ( .A(n20082), .B(n20953), .C(n21816), .Y(
        n20080) );
  sky130_fd_sc_hd__nor2_1 U26234 ( .A(n20078), .B(n20077), .Y(n20954) );
  sky130_fd_sc_hd__nor2_1 U26235 ( .A(n20080), .B(n20079), .Y(n20081) );
  sky130_fd_sc_hd__nand2_1 U26236 ( .A(n20083), .B(n20081), .Y(n20087) );
  sky130_fd_sc_hd__nand3_1 U26237 ( .A(n20954), .B(
        j202_soc_core_memory0_ram_dout0_sel[15]), .C(n20953), .Y(n20084) );
  sky130_fd_sc_hd__nand2_1 U26238 ( .A(n20083), .B(n20082), .Y(n20955) );
  sky130_fd_sc_hd__nor2_1 U26239 ( .A(n20084), .B(n20955), .Y(n20085) );
  sky130_fd_sc_hd__nand2_1 U26240 ( .A(n20957), .B(n20085), .Y(n20086) );
  sky130_fd_sc_hd__o22ai_1 U26241 ( .A1(n20088), .A2(n20087), .B1(n20086), 
        .B2(j202_soc_core_memory0_ram_dout0[493]), .Y(n22222) );
  sky130_fd_sc_hd__nand2_1 U26242 ( .A(j202_soc_core_j22_cpu_id_op2_v_), .B(
        j202_soc_core_j22_cpu_id_op2_inst__14_), .Y(n20092) );
  sky130_fd_sc_hd__nand2_1 U26243 ( .A(n11203), .B(n20092), .Y(n20093) );
  sky130_fd_sc_hd__nand2_1 U26244 ( .A(j202_soc_core_memory0_ram_dout0[174]), 
        .B(n21487), .Y(n20094) );
  sky130_fd_sc_hd__nand2_1 U26245 ( .A(j202_soc_core_memory0_ram_dout0[302]), 
        .B(n21503), .Y(n20096) );
  sky130_fd_sc_hd__nand2_1 U26246 ( .A(j202_soc_core_memory0_ram_dout0[46]), 
        .B(n21633), .Y(n20095) );
  sky130_fd_sc_hd__nand2_1 U26247 ( .A(j202_soc_core_memory0_ram_dout0[78]), 
        .B(n21642), .Y(n20097) );
  sky130_fd_sc_hd__o2bb2ai_1 U26248 ( .B1(n20098), .B2(n21515), .A1_N(
        j202_soc_core_ahblite_interconnect_s_hrdata[110]), .A2_N(n21446), .Y(
        n20242) );
  sky130_fd_sc_hd__nand2_1 U26249 ( .A(n20759), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[78]), .Y(n20244) );
  sky130_fd_sc_hd__nand2_1 U26250 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[14]), .Y(n20243) );
  sky130_fd_sc_hd__nand3_1 U26251 ( .A(n20244), .B(n21768), .C(n20243), .Y(
        n20099) );
  sky130_fd_sc_hd__nor2_1 U26252 ( .A(n20242), .B(n20099), .Y(n20241) );
  sky130_fd_sc_hd__nor2_1 U26253 ( .A(n20101), .B(n20100), .Y(n20104) );
  sky130_fd_sc_hd__nand4_1 U26254 ( .A(n20104), .B(n20103), .C(n20181), .D(
        n20102), .Y(n20106) );
  sky130_fd_sc_hd__o21ai_1 U26255 ( .A1(n20106), .A2(n20105), .B1(n20210), .Y(
        n20125) );
  sky130_fd_sc_hd__nand2_1 U26256 ( .A(n20181), .B(n20204), .Y(n20220) );
  sky130_fd_sc_hd__nand3_1 U26257 ( .A(n20109), .B(n20108), .C(n20107), .Y(
        n20111) );
  sky130_fd_sc_hd__a21oi_1 U26258 ( .A1(n20111), .A2(n20179), .B1(n20110), .Y(
        n20124) );
  sky130_fd_sc_hd__nand3_1 U26259 ( .A(n20215), .B(n20113), .C(n20112), .Y(
        n20114) );
  sky130_fd_sc_hd__nand2_1 U26260 ( .A(n20153), .B(n20138), .Y(n20169) );
  sky130_fd_sc_hd__nor3_1 U26261 ( .A(n20114), .B(n20140), .C(n20169), .Y(
        n20116) );
  sky130_fd_sc_hd__nand3_1 U26262 ( .A(n20116), .B(n20209), .C(n20115), .Y(
        n20117) );
  sky130_fd_sc_hd__nand2_1 U26263 ( .A(n20117), .B(n20227), .Y(n20123) );
  sky130_fd_sc_hd__nand4_1 U26264 ( .A(n20120), .B(n20155), .C(n20119), .D(
        n20118), .Y(n20121) );
  sky130_fd_sc_hd__nand2_1 U26265 ( .A(n20121), .B(n20225), .Y(n20122) );
  sky130_fd_sc_hd__nand4_1 U26266 ( .A(n20125), .B(n20124), .C(n20123), .D(
        n20122), .Y(n20127) );
  sky130_fd_sc_hd__nand2_1 U26267 ( .A(n20127), .B(n20126), .Y(n20239) );
  sky130_fd_sc_hd__nand3_1 U26268 ( .A(n20130), .B(n20129), .C(n20128), .Y(
        n20131) );
  sky130_fd_sc_hd__nor2_1 U26269 ( .A(n20132), .B(n20131), .Y(n20133) );
  sky130_fd_sc_hd__nand2_1 U26270 ( .A(n20134), .B(n20133), .Y(n20135) );
  sky130_fd_sc_hd__nand4_1 U26272 ( .A(n20139), .B(n20138), .C(n20137), .D(
        n20204), .Y(n20141) );
  sky130_fd_sc_hd__nor2_1 U26273 ( .A(n20141), .B(n20140), .Y(n20142) );
  sky130_fd_sc_hd__nand2_1 U26274 ( .A(n20143), .B(n20142), .Y(n20144) );
  sky130_fd_sc_hd__nand2_1 U26275 ( .A(n20144), .B(n20210), .Y(n20160) );
  sky130_fd_sc_hd__nand2_1 U26276 ( .A(n20183), .B(n20145), .Y(n20147) );
  sky130_fd_sc_hd__nor2_1 U26277 ( .A(n20147), .B(n20146), .Y(n20150) );
  sky130_fd_sc_hd__nand4_1 U26278 ( .A(n20150), .B(n20149), .C(n20148), .D(
        n20178), .Y(n20151) );
  sky130_fd_sc_hd__nand2_1 U26279 ( .A(n20151), .B(n20179), .Y(n20159) );
  sky130_fd_sc_hd__nand3_1 U26280 ( .A(n20153), .B(n20183), .C(n20152), .Y(
        n20154) );
  sky130_fd_sc_hd__nor2_1 U26281 ( .A(n20154), .B(n20219), .Y(n20156) );
  sky130_fd_sc_hd__nand3_1 U26282 ( .A(n20156), .B(n20155), .C(n20163), .Y(
        n20157) );
  sky130_fd_sc_hd__nand2_1 U26283 ( .A(n20157), .B(n20225), .Y(n20158) );
  sky130_fd_sc_hd__nand4_1 U26284 ( .A(n20161), .B(n20160), .C(n20159), .D(
        n20158), .Y(n20197) );
  sky130_fd_sc_hd__nand2_1 U26285 ( .A(n20163), .B(n20162), .Y(n20165) );
  sky130_fd_sc_hd__o21ai_1 U26286 ( .A1(n20165), .A2(n20164), .B1(n20225), .Y(
        n20193) );
  sky130_fd_sc_hd__nand2_1 U26287 ( .A(n20167), .B(n20166), .Y(n20168) );
  sky130_fd_sc_hd__o31a_1 U26288 ( .A1(n20169), .A2(n20221), .A3(n20168), .B1(
        n20227), .X(n20171) );
  sky130_fd_sc_hd__nor2_1 U26289 ( .A(n20171), .B(n20170), .Y(n20192) );
  sky130_fd_sc_hd__nand2_1 U26290 ( .A(n20173), .B(n20172), .Y(n20174) );
  sky130_fd_sc_hd__nor2_1 U26291 ( .A(n20175), .B(n20174), .Y(n20176) );
  sky130_fd_sc_hd__nand3_1 U26292 ( .A(n20178), .B(n20177), .C(n20176), .Y(
        n20180) );
  sky130_fd_sc_hd__nand2_1 U26293 ( .A(n20180), .B(n20179), .Y(n20191) );
  sky130_fd_sc_hd__and4_1 U26294 ( .A(n20214), .B(n20183), .C(n20182), .D(
        n20181), .X(n20184) );
  sky130_fd_sc_hd__nand4_1 U26295 ( .A(n20187), .B(n20186), .C(n20185), .D(
        n20184), .Y(n20189) );
  sky130_fd_sc_hd__o21ai_1 U26296 ( .A1(n20189), .A2(n20188), .B1(n20210), .Y(
        n20190) );
  sky130_fd_sc_hd__nand4_1 U26297 ( .A(n20193), .B(n20192), .C(n20191), .D(
        n20190), .Y(n20195) );
  sky130_fd_sc_hd__a22oi_1 U26298 ( .A1(n20197), .A2(n20196), .B1(n20195), 
        .B2(n20194), .Y(n20238) );
  sky130_fd_sc_hd__a21oi_1 U26299 ( .A1(n19148), .A2(n20199), .B1(n20198), .Y(
        n20201) );
  sky130_fd_sc_hd__a31oi_1 U26300 ( .A1(n20203), .A2(n20202), .A3(n20201), 
        .B1(n20200), .Y(n20234) );
  sky130_fd_sc_hd__nand3_1 U26301 ( .A(n20205), .B(n20215), .C(n20204), .Y(
        n20207) );
  sky130_fd_sc_hd__nor2_1 U26302 ( .A(n20207), .B(n20206), .Y(n20208) );
  sky130_fd_sc_hd__nand2_1 U26303 ( .A(n20209), .B(n20208), .Y(n20211) );
  sky130_fd_sc_hd__nand4_1 U26305 ( .A(n20217), .B(n20216), .C(n20215), .D(
        n20214), .Y(n20218) );
  sky130_fd_sc_hd__nor2_1 U26306 ( .A(n20219), .B(n20218), .Y(n20224) );
  sky130_fd_sc_hd__nor2_1 U26307 ( .A(n20221), .B(n20220), .Y(n20222) );
  sky130_fd_sc_hd__nand3_1 U26308 ( .A(n20224), .B(n20223), .C(n20222), .Y(
        n20226) );
  sky130_fd_sc_hd__nand2_1 U26309 ( .A(n20226), .B(n20225), .Y(n20232) );
  sky130_fd_sc_hd__o31ai_1 U26310 ( .A1(n20230), .A2(n20229), .A3(n20228), 
        .B1(n20227), .Y(n20231) );
  sky130_fd_sc_hd__nand4b_1 U26311 ( .A_N(n20234), .B(n20233), .C(n20232), .D(
        n20231), .Y(n20236) );
  sky130_fd_sc_hd__nand2_1 U26312 ( .A(n20236), .B(n20235), .Y(n20237) );
  sky130_fd_sc_hd__nand3_1 U26313 ( .A(n20239), .B(n20238), .C(n20237), .Y(
        n20240) );
  sky130_fd_sc_hd__nand2_1 U26314 ( .A(n20240), .B(n21629), .Y(n20249) );
  sky130_fd_sc_hd__nand2_1 U26315 ( .A(n20786), .B(
        j202_soc_core_bldc_core_00_pwm_duty[2]), .Y(n20246) );
  sky130_fd_sc_hd__nand2_1 U26316 ( .A(j202_soc_core_memory0_ram_dout0[494]), 
        .B(n21650), .Y(n20251) );
  sky130_fd_sc_hd__nand4_1 U26317 ( .A(n20245), .B(n21653), .C(n20244), .D(
        n20243), .Y(n20248) );
  sky130_fd_sc_hd__nor2_1 U26318 ( .A(n20248), .B(n20247), .Y(n20250) );
  sky130_fd_sc_hd__nand3_1 U26319 ( .A(n20251), .B(n20250), .C(n20249), .Y(
        n21001) );
  sky130_fd_sc_hd__nand2_1 U26320 ( .A(n21916), .B(
        j202_soc_core_j22_cpu_id_opn_inst__14_), .Y(n20252) );
  sky130_fd_sc_hd__a22oi_1 U26321 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__2_), .B1(n21916), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__2_), .Y(n20256) );
  sky130_fd_sc_hd__o21a_1 U26322 ( .A1(n11203), .A2(n20257), .B1(n20256), .X(
        n20258) );
  sky130_fd_sc_hd__nand2_1 U26323 ( .A(j202_soc_core_memory0_ram_dout0[131]), 
        .B(n21489), .Y(n20262) );
  sky130_fd_sc_hd__nand2_1 U26324 ( .A(j202_soc_core_memory0_ram_dout0[67]), 
        .B(n21642), .Y(n20261) );
  sky130_fd_sc_hd__nand2_1 U26325 ( .A(j202_soc_core_memory0_ram_dout0[163]), 
        .B(n21487), .Y(n20260) );
  sky130_fd_sc_hd__nand2_1 U26326 ( .A(j202_soc_core_memory0_ram_dout0[323]), 
        .B(n21490), .Y(n20259) );
  sky130_fd_sc_hd__nand2_1 U26327 ( .A(j202_soc_core_memory0_ram_dout0[451]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n20266) );
  sky130_fd_sc_hd__nand2_1 U26328 ( .A(j202_soc_core_memory0_ram_dout0[419]), 
        .B(n12156), .Y(n20265) );
  sky130_fd_sc_hd__nand2_1 U26329 ( .A(j202_soc_core_memory0_ram_dout0[355]), 
        .B(n21495), .Y(n20264) );
  sky130_fd_sc_hd__nand2_1 U26330 ( .A(j202_soc_core_memory0_ram_dout0[387]), 
        .B(n21496), .Y(n20263) );
  sky130_fd_sc_hd__nand2_1 U26331 ( .A(j202_soc_core_memory0_ram_dout0[3]), 
        .B(n21639), .Y(n20414) );
  sky130_fd_sc_hd__nand2_1 U26332 ( .A(j202_soc_core_memory0_ram_dout0[195]), 
        .B(n21640), .Y(n20413) );
  sky130_fd_sc_hd__a22oi_1 U26333 ( .A1(n21516), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[3]), .B1(n20759), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[67]), .Y(n20267) );
  sky130_fd_sc_hd__o21a_1 U26334 ( .A1(n27680), .A2(n21517), .B1(n20267), .X(
        n20419) );
  sky130_fd_sc_hd__nand2b_1 U26335 ( .A_N(n21515), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[35]), .Y(n20418) );
  sky130_fd_sc_hd__nand3_1 U26336 ( .A(n20419), .B(n21768), .C(n20418), .Y(
        n20411) );
  sky130_fd_sc_hd__nand4_1 U26337 ( .A(n20367), .B(n20317), .C(n20268), .D(
        n20293), .Y(n20269) );
  sky130_fd_sc_hd__o21ai_0 U26338 ( .A1(n20282), .A2(n20269), .B1(n20368), .Y(
        n20287) );
  sky130_fd_sc_hd__nor2_1 U26339 ( .A(n20291), .B(n20270), .Y(n20384) );
  sky130_fd_sc_hd__nand4_1 U26340 ( .A(n20384), .B(n20271), .C(n20348), .D(
        n20339), .Y(n20273) );
  sky130_fd_sc_hd__o21ai_0 U26341 ( .A1(n20273), .A2(n20272), .B1(n20385), .Y(
        n20286) );
  sky130_fd_sc_hd__nand3_1 U26342 ( .A(n20379), .B(n20364), .C(n20289), .Y(
        n20274) );
  sky130_fd_sc_hd__nor2_1 U26343 ( .A(n20274), .B(n20297), .Y(n20275) );
  sky130_fd_sc_hd__nand3_1 U26344 ( .A(n20275), .B(n20334), .C(n20392), .Y(
        n20276) );
  sky130_fd_sc_hd__nand2_1 U26345 ( .A(n20276), .B(n20374), .Y(n20285) );
  sky130_fd_sc_hd__nand4_1 U26346 ( .A(n20277), .B(n20360), .C(n20339), .D(
        n20377), .Y(n20281) );
  sky130_fd_sc_hd__nand4b_1 U26347 ( .A_N(n20281), .B(n20280), .C(n20317), .D(
        n20279), .Y(n20283) );
  sky130_fd_sc_hd__nand4_1 U26349 ( .A(n20287), .B(n20286), .C(n20285), .D(
        n20284), .Y(n20288) );
  sky130_fd_sc_hd__nand2_1 U26350 ( .A(n20288), .B(n20643), .Y(n20410) );
  sky130_fd_sc_hd__nand2_1 U26351 ( .A(n20380), .B(n20289), .Y(n20290) );
  sky130_fd_sc_hd__nor2_1 U26352 ( .A(n20291), .B(n20290), .Y(n20332) );
  sky130_fd_sc_hd__nand3_1 U26353 ( .A(n20332), .B(n20292), .C(n20390), .Y(
        n20308) );
  sky130_fd_sc_hd__nor3_1 U26354 ( .A(n20296), .B(n20295), .C(n20294), .Y(
        n20298) );
  sky130_fd_sc_hd__nand4_1 U26355 ( .A(n20299), .B(n20317), .C(n20298), .D(
        n20353), .Y(n20300) );
  sky130_fd_sc_hd__nand2_1 U26356 ( .A(n20300), .B(n20385), .Y(n20324) );
  sky130_fd_sc_hd__nand3_1 U26358 ( .A(n20307), .B(n20306), .C(n20305), .Y(
        n20309) );
  sky130_fd_sc_hd__o21ai_1 U26359 ( .A1(n20309), .A2(n20308), .B1(n20374), .Y(
        n20323) );
  sky130_fd_sc_hd__nand4b_1 U26360 ( .A_N(n20312), .B(n20311), .C(n20310), .D(
        n20349), .Y(n20313) );
  sky130_fd_sc_hd__o21ai_1 U26361 ( .A1(n20313), .A2(n20395), .B1(n20393), .Y(
        n20322) );
  sky130_fd_sc_hd__nor2_1 U26362 ( .A(n20315), .B(n20314), .Y(n20318) );
  sky130_fd_sc_hd__nand4_1 U26363 ( .A(n20319), .B(n20318), .C(n20317), .D(
        n20316), .Y(n20320) );
  sky130_fd_sc_hd__nand2_1 U26364 ( .A(n20320), .B(n20368), .Y(n20321) );
  sky130_fd_sc_hd__nand4_1 U26365 ( .A(n20324), .B(n20323), .C(n20322), .D(
        n20321), .Y(n20325) );
  sky130_fd_sc_hd__nand2_1 U26366 ( .A(n20325), .B(n20784), .Y(n20409) );
  sky130_fd_sc_hd__nor2_1 U26367 ( .A(n20328), .B(n20327), .Y(n20329) );
  sky130_fd_sc_hd__nand2_1 U26368 ( .A(n20330), .B(n20329), .Y(n20331) );
  sky130_fd_sc_hd__nand2_1 U26369 ( .A(n20331), .B(n20393), .Y(n20358) );
  sky130_fd_sc_hd__nand4_1 U26370 ( .A(n20335), .B(n20334), .C(n20379), .D(
        n20333), .Y(n20336) );
  sky130_fd_sc_hd__o21ai_0 U26371 ( .A1(n20337), .A2(n20336), .B1(n20385), .Y(
        n20357) );
  sky130_fd_sc_hd__nand4_1 U26372 ( .A(n20340), .B(n20339), .C(n20338), .D(
        n20379), .Y(n20342) );
  sky130_fd_sc_hd__o21ai_0 U26373 ( .A1(n20342), .A2(n20341), .B1(n20368), .Y(
        n20356) );
  sky130_fd_sc_hd__nand2_1 U26374 ( .A(n20344), .B(n20343), .Y(n20346) );
  sky130_fd_sc_hd__nor2_1 U26375 ( .A(n20346), .B(n20345), .Y(n20352) );
  sky130_fd_sc_hd__nand3_1 U26376 ( .A(n20349), .B(n20348), .C(n20347), .Y(
        n20351) );
  sky130_fd_sc_hd__nor2_1 U26377 ( .A(n20351), .B(n20350), .Y(n20373) );
  sky130_fd_sc_hd__nand4_1 U26378 ( .A(n20367), .B(n20353), .C(n20352), .D(
        n20373), .Y(n20354) );
  sky130_fd_sc_hd__nand2_1 U26379 ( .A(n20354), .B(n20374), .Y(n20355) );
  sky130_fd_sc_hd__nand4_1 U26380 ( .A(n20358), .B(n20357), .C(n20356), .D(
        n20355), .Y(n20359) );
  sky130_fd_sc_hd__nand2_1 U26381 ( .A(n20359), .B(n20617), .Y(n20408) );
  sky130_fd_sc_hd__nor2_1 U26382 ( .A(n20362), .B(n20361), .Y(n20365) );
  sky130_fd_sc_hd__nand4_1 U26383 ( .A(n20366), .B(n20365), .C(n20364), .D(
        n20363), .Y(n20370) );
  sky130_fd_sc_hd__o21ai_1 U26384 ( .A1(n20370), .A2(n20369), .B1(n20368), .Y(
        n20399) );
  sky130_fd_sc_hd__nand4_1 U26385 ( .A(n20373), .B(n20384), .C(n20372), .D(
        n20371), .Y(n20375) );
  sky130_fd_sc_hd__nand2_1 U26386 ( .A(n20375), .B(n20374), .Y(n20398) );
  sky130_fd_sc_hd__nand4_1 U26387 ( .A(n20380), .B(n20379), .C(n20378), .D(
        n20377), .Y(n20382) );
  sky130_fd_sc_hd__nor2_1 U26388 ( .A(n20382), .B(n20381), .Y(n20383) );
  sky130_fd_sc_hd__nand2_1 U26389 ( .A(n20384), .B(n20383), .Y(n20386) );
  sky130_fd_sc_hd__nand2_1 U26390 ( .A(n20386), .B(n20385), .Y(n20397) );
  sky130_fd_sc_hd__o21a_1 U26391 ( .A1(n20388), .A2(n21595), .B1(n20387), .X(
        n20391) );
  sky130_fd_sc_hd__nand4_1 U26392 ( .A(n20392), .B(n20391), .C(n20390), .D(
        n20389), .Y(n20394) );
  sky130_fd_sc_hd__nand4_1 U26394 ( .A(n20399), .B(n20398), .C(n20397), .D(
        n20396), .Y(n20406) );
  sky130_fd_sc_hd__nand2_1 U26395 ( .A(n21504), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[11]), .Y(n20403) );
  sky130_fd_sc_hd__nand2_1 U26396 ( .A(n24720), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[19]), .Y(n20402) );
  sky130_fd_sc_hd__nand2_1 U26397 ( .A(n21505), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[3]), .Y(n20401) );
  sky130_fd_sc_hd__nand2_1 U26398 ( .A(n21506), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[27]), .Y(n20400) );
  sky130_fd_sc_hd__nand4_1 U26399 ( .A(n20403), .B(n20402), .C(n20401), .D(
        n20400), .Y(n20404) );
  sky130_fd_sc_hd__a22oi_1 U26400 ( .A1(n21446), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[99]), .B1(n21513), .B2(
        n20404), .Y(n20405) );
  sky130_fd_sc_hd__nand4_1 U26401 ( .A(n20410), .B(n20409), .C(n20408), .D(
        n20407), .Y(n20420) );
  sky130_fd_sc_hd__nor2_1 U26402 ( .A(n20411), .B(n20420), .Y(n20412) );
  sky130_fd_sc_hd__nand2_1 U26403 ( .A(j202_soc_core_memory0_ram_dout0[483]), 
        .B(n21650), .Y(n20423) );
  sky130_fd_sc_hd__nand3_1 U26404 ( .A(n20419), .B(n21653), .C(n20418), .Y(
        n20421) );
  sky130_fd_sc_hd__nor2_1 U26405 ( .A(n20421), .B(n20420), .Y(n20422) );
  sky130_fd_sc_hd__nand2_1 U26406 ( .A(n20423), .B(n20422), .Y(n20440) );
  sky130_fd_sc_hd__a22oi_1 U26407 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__3_), .B1(n21916), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__3_), .Y(n20424) );
  sky130_fd_sc_hd__nand2b_1 U26408 ( .A_N(n12399), .B(n28417), .Y(n20430) );
  sky130_fd_sc_hd__nand3_1 U26409 ( .A(n28360), .B(n20429), .C(n20428), .Y(
        n28155) );
  sky130_fd_sc_hd__nand2_1 U26410 ( .A(n24602), .B(n28402), .Y(n24570) );
  sky130_fd_sc_hd__nand2_1 U26411 ( .A(n20430), .B(n24570), .Y(n29540) );
  sky130_fd_sc_hd__nand2_1 U26412 ( .A(n11102), .B(n22739), .Y(n20439) );
  sky130_fd_sc_hd__nand2_1 U26413 ( .A(n20433), .B(n20432), .Y(n20434) );
  sky130_fd_sc_hd__xor2_1 U26414 ( .A(n20435), .B(n20434), .X(n24052) );
  sky130_fd_sc_hd__o22ai_1 U26415 ( .A1(n26284), .A2(n11186), .B1(
        j202_soc_core_j22_cpu_pc[1]), .B2(n22705), .Y(n20436) );
  sky130_fd_sc_hd__a21oi_1 U26416 ( .A1(n24052), .A2(n17225), .B1(n20436), .Y(
        n20438) );
  sky130_fd_sc_hd__nand2_1 U26417 ( .A(n21924), .B(n12354), .Y(n20437) );
  sky130_fd_sc_hd__nand3_2 U26418 ( .A(n20439), .B(n20438), .C(n20437), .Y(
        n29581) );
  sky130_fd_sc_hd__nand2_1 U26419 ( .A(n20441), .B(n20440), .Y(n24027) );
  sky130_fd_sc_hd__nand2b_1 U26420 ( .A_N(n24027), .B(n22739), .Y(n20452) );
  sky130_fd_sc_hd__nand2_1 U26421 ( .A(n21787), .B(n21785), .Y(n20444) );
  sky130_fd_sc_hd__xnor2_1 U26422 ( .A(n20444), .B(n21788), .Y(n24082) );
  sky130_fd_sc_hd__xnor2_1 U26423 ( .A(n20446), .B(n21781), .Y(n24773) );
  sky130_fd_sc_hd__nor2_1 U26424 ( .A(n20447), .B(n22705), .Y(n20449) );
  sky130_fd_sc_hd__o22ai_1 U26425 ( .A1(n20447), .A2(n13365), .B1(n11190), 
        .B2(n11186), .Y(n20448) );
  sky130_fd_sc_hd__a211oi_1 U26426 ( .A1(n24082), .A2(n17225), .B1(n20449), 
        .C1(n20448), .Y(n20451) );
  sky130_fd_sc_hd__nand2_1 U26427 ( .A(n21924), .B(n28515), .Y(n20450) );
  sky130_fd_sc_hd__nand3_1 U26428 ( .A(n20452), .B(n20451), .C(n20450), .Y(
        n29553) );
  sky130_fd_sc_hd__a22oi_1 U26430 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__7_), .B1(n21916), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__7_), .Y(n20453) );
  sky130_fd_sc_hd__nand2_1 U26431 ( .A(j202_soc_core_memory0_ram_dout0[72]), 
        .B(n20458), .Y(n20461) );
  sky130_fd_sc_hd__nand2b_1 U26432 ( .A_N(n20656), .B(n13199), .Y(n20842) );
  sky130_fd_sc_hd__nand2_1 U26433 ( .A(n20775), .B(n20842), .Y(n20663) );
  sky130_fd_sc_hd__nor2_1 U26434 ( .A(n20463), .B(n20663), .Y(n20566) );
  sky130_fd_sc_hd__nand2_1 U26435 ( .A(n20490), .B(n20464), .Y(n20840) );
  sky130_fd_sc_hd__nand2_1 U26436 ( .A(n20840), .B(n20623), .Y(n20769) );
  sky130_fd_sc_hd__nand2_1 U26437 ( .A(n20566), .B(n20519), .Y(n20465) );
  sky130_fd_sc_hd__o21ai_1 U26438 ( .A1(n20625), .A2(n20465), .B1(n20833), .Y(
        n20481) );
  sky130_fd_sc_hd__nand3_1 U26439 ( .A(n20467), .B(n20466), .C(n20528), .Y(
        n20469) );
  sky130_fd_sc_hd__nor2_1 U26440 ( .A(n20468), .B(n20605), .Y(n20847) );
  sky130_fd_sc_hd__nand2_1 U26441 ( .A(n20847), .B(n20774), .Y(n20569) );
  sky130_fd_sc_hd__o21ai_1 U26442 ( .A1(n20469), .A2(n20569), .B1(n20804), .Y(
        n20480) );
  sky130_fd_sc_hd__and3_1 U26443 ( .A(n20830), .B(n20603), .C(n20623), .X(
        n20470) );
  sky130_fd_sc_hd__nand3_1 U26444 ( .A(n20635), .B(n20471), .C(n20470), .Y(
        n20473) );
  sky130_fd_sc_hd__nand2_1 U26445 ( .A(n20472), .B(n20528), .Y(n20789) );
  sky130_fd_sc_hd__nand4b_1 U26446 ( .A_N(n20633), .B(n20790), .C(n20842), .D(
        n20661), .Y(n20807) );
  sky130_fd_sc_hd__o21ai_1 U26447 ( .A1(n20473), .A2(n20807), .B1(n20856), .Y(
        n20479) );
  sky130_fd_sc_hd__nand3_1 U26448 ( .A(n20842), .B(n20560), .C(n20836), .Y(
        n20475) );
  sky130_fd_sc_hd__nor2_1 U26449 ( .A(n20475), .B(n20474), .Y(n20476) );
  sky130_fd_sc_hd__nand4_1 U26450 ( .A(n20662), .B(n20551), .C(n20664), .D(
        n20476), .Y(n20477) );
  sky130_fd_sc_hd__nand2_1 U26451 ( .A(n20477), .B(n20850), .Y(n20478) );
  sky130_fd_sc_hd__nand4_1 U26452 ( .A(n20481), .B(n20480), .C(n20479), .D(
        n20478), .Y(n20507) );
  sky130_fd_sc_hd__nand2_1 U26453 ( .A(n20820), .B(n20482), .Y(n20659) );
  sky130_fd_sc_hd__nor2_1 U26454 ( .A(n20483), .B(n20659), .Y(n20513) );
  sky130_fd_sc_hd__nand3_1 U26455 ( .A(n20837), .B(n20675), .C(n20775), .Y(
        n20484) );
  sky130_fd_sc_hd__nand2_1 U26456 ( .A(n20486), .B(n20485), .Y(n20599) );
  sky130_fd_sc_hd__nand4_1 U26457 ( .A(n20513), .B(n20610), .C(n20817), .D(
        n20599), .Y(n20488) );
  sky130_fd_sc_hd__nor3_1 U26458 ( .A(n20488), .B(n20487), .C(n20815), .Y(
        n20489) );
  sky130_fd_sc_hd__nand2_1 U26459 ( .A(n20838), .B(n20489), .Y(n20492) );
  sky130_fd_sc_hd__nand3_1 U26460 ( .A(n20798), .B(n20767), .C(n20491), .Y(
        n20686) );
  sky130_fd_sc_hd__o21ai_1 U26461 ( .A1(n20492), .A2(n20686), .B1(n20804), .Y(
        n20504) );
  sky130_fd_sc_hd__nand3_1 U26462 ( .A(n20635), .B(n20814), .C(n20599), .Y(
        n20645) );
  sky130_fd_sc_hd__nand2_1 U26463 ( .A(n20637), .B(n20519), .Y(n20493) );
  sky130_fd_sc_hd__nor2_1 U26464 ( .A(n20645), .B(n20493), .Y(n20839) );
  sky130_fd_sc_hd__nand2_1 U26465 ( .A(n20839), .B(n20494), .Y(n20495) );
  sky130_fd_sc_hd__nand2_1 U26466 ( .A(n20495), .B(n20850), .Y(n20503) );
  sky130_fd_sc_hd__nand2_1 U26467 ( .A(n20742), .B(n20840), .Y(n20732) );
  sky130_fd_sc_hd__nand2_1 U26468 ( .A(n20610), .B(n20799), .Y(n20788) );
  sky130_fd_sc_hd__nand2_1 U26469 ( .A(n20496), .B(n20746), .Y(n20593) );
  sky130_fd_sc_hd__nor4_1 U26470 ( .A(n20807), .B(n20732), .C(n20788), .D(
        n20593), .Y(n20497) );
  sky130_fd_sc_hd__nand2b_1 U26471 ( .A_N(n20497), .B(n20856), .Y(n20502) );
  sky130_fd_sc_hd__nor3_1 U26472 ( .A(n20821), .B(n20626), .C(n20844), .Y(
        n20498) );
  sky130_fd_sc_hd__nand2_1 U26473 ( .A(n20799), .B(n20498), .Y(n20500) );
  sky130_fd_sc_hd__nand4_1 U26475 ( .A(n20504), .B(n20503), .C(n20502), .D(
        n20501), .Y(n20506) );
  sky130_fd_sc_hd__a22oi_1 U26476 ( .A1(n20508), .A2(n20507), .B1(n20506), 
        .B2(n20505), .Y(n20579) );
  sky130_fd_sc_hd__nor2_1 U26477 ( .A(n20509), .B(n20765), .Y(n20510) );
  sky130_fd_sc_hd__nand4_1 U26478 ( .A(n20510), .B(n20852), .C(n20793), .D(
        n20837), .Y(n20511) );
  sky130_fd_sc_hd__nor2_1 U26479 ( .A(n20511), .B(n20612), .Y(n20512) );
  sky130_fd_sc_hd__nand2_1 U26480 ( .A(n20513), .B(n20512), .Y(n20514) );
  sky130_fd_sc_hd__nand2_1 U26481 ( .A(n20514), .B(n20850), .Y(n20539) );
  sky130_fd_sc_hd__o21a_1 U26482 ( .A1(n20516), .A2(n20515), .B1(n20560), .X(
        n20517) );
  sky130_fd_sc_hd__nand4_1 U26483 ( .A(n20551), .B(n20519), .C(n20518), .D(
        n20517), .Y(n20527) );
  sky130_fd_sc_hd__nor2_1 U26484 ( .A(n20663), .B(n20737), .Y(n20524) );
  sky130_fd_sc_hd__nand2b_1 U26485 ( .A_N(n20520), .B(n21088), .Y(n20794) );
  sky130_fd_sc_hd__and4_1 U26486 ( .A(n20794), .B(n20521), .C(n20623), .D(
        n20680), .X(n20522) );
  sky130_fd_sc_hd__nand4_1 U26487 ( .A(n20525), .B(n20524), .C(n20523), .D(
        n20522), .Y(n20526) );
  sky130_fd_sc_hd__a22oi_1 U26488 ( .A1(n20527), .A2(n20804), .B1(n20526), 
        .B2(n20856), .Y(n20538) );
  sky130_fd_sc_hd__nand2_1 U26489 ( .A(n20842), .B(n20528), .Y(n20777) );
  sky130_fd_sc_hd__nand3_1 U26490 ( .A(n20530), .B(n20820), .C(n20529), .Y(
        n20596) );
  sky130_fd_sc_hd__nand2_1 U26491 ( .A(n20532), .B(n20531), .Y(n20533) );
  sky130_fd_sc_hd__nand3_1 U26492 ( .A(n20664), .B(n20534), .C(n20635), .Y(
        n20763) );
  sky130_fd_sc_hd__nand3_1 U26493 ( .A(n20535), .B(n20740), .C(n20831), .Y(
        n20536) );
  sky130_fd_sc_hd__nand3_1 U26495 ( .A(n20539), .B(n20538), .C(n20537), .Y(
        n20548) );
  sky130_fd_sc_hd__nand2_1 U26496 ( .A(n20786), .B(
        j202_soc_core_bldc_core_00_pwm_period[8]), .Y(n20546) );
  sky130_fd_sc_hd__a22oi_1 U26497 ( .A1(n20759), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[72]), .B1(n20540), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[40]), .Y(n20545) );
  sky130_fd_sc_hd__a22oi_1 U26498 ( .A1(n21516), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[8]), .B1(n21446), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[104]), .Y(n20544) );
  sky130_fd_sc_hd__xnor2_1 U26499 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[1]), 
        .B(j202_soc_core_uart_TOP_rx_fifo_wp[1]), .Y(n27960) );
  sky130_fd_sc_hd__xnor2_1 U26500 ( .A(j202_soc_core_uart_TOP_rx_fifo_wp[0]), 
        .B(j202_soc_core_uart_TOP_rx_fifo_rp[0]), .Y(n20541) );
  sky130_fd_sc_hd__nand2_1 U26501 ( .A(n27960), .B(n20541), .Y(n23895) );
  sky130_fd_sc_hd__nor2_1 U26502 ( .A(j202_soc_core_uart_TOP_rx_fifo_gb), .B(
        n23895), .Y(n20542) );
  sky130_fd_sc_hd__nand2_1 U26503 ( .A(n21513), .B(n20542), .Y(n20543) );
  sky130_fd_sc_hd__nand4_1 U26504 ( .A(n20546), .B(n20545), .C(n20544), .D(
        n20543), .Y(n20547) );
  sky130_fd_sc_hd__a21oi_1 U26505 ( .A1(n20548), .A2(n20784), .B1(n20547), .Y(
        n20578) );
  sky130_fd_sc_hd__nor2_1 U26506 ( .A(n20612), .B(n20821), .Y(n20557) );
  sky130_fd_sc_hd__nand2_1 U26507 ( .A(n20836), .B(n20687), .Y(n20653) );
  sky130_fd_sc_hd__nor3_1 U26508 ( .A(n20653), .B(n20549), .C(n20595), .Y(
        n20550) );
  sky130_fd_sc_hd__nand3_1 U26509 ( .A(n20557), .B(n20551), .C(n20550), .Y(
        n20552) );
  sky130_fd_sc_hd__nand2_1 U26510 ( .A(n20552), .B(n20804), .Y(n20575) );
  sky130_fd_sc_hd__nand3_1 U26511 ( .A(n20553), .B(n20675), .C(n20559), .Y(
        n20555) );
  sky130_fd_sc_hd__nor3_1 U26512 ( .A(n20555), .B(n20777), .C(n20554), .Y(
        n20556) );
  sky130_fd_sc_hd__nand2_1 U26513 ( .A(n20557), .B(n20556), .Y(n20558) );
  sky130_fd_sc_hd__nand2_1 U26514 ( .A(n20558), .B(n20850), .Y(n20574) );
  sky130_fd_sc_hd__and3_1 U26515 ( .A(n20817), .B(n20793), .C(n20766), .X(
        n20649) );
  sky130_fd_sc_hd__nand3_1 U26516 ( .A(n20741), .B(n20560), .C(n20559), .Y(
        n20562) );
  sky130_fd_sc_hd__nor2_1 U26517 ( .A(n20562), .B(n20561), .Y(n20565) );
  sky130_fd_sc_hd__nor2_1 U26518 ( .A(n20563), .B(n20743), .Y(n20564) );
  sky130_fd_sc_hd__nand4_1 U26519 ( .A(n20649), .B(n20566), .C(n20565), .D(
        n20564), .Y(n20572) );
  sky130_fd_sc_hd__nand2_1 U26520 ( .A(n20610), .B(n20687), .Y(n20567) );
  sky130_fd_sc_hd__nor2_1 U26521 ( .A(n20568), .B(n20567), .Y(n20854) );
  sky130_fd_sc_hd__nor2_1 U26522 ( .A(n20598), .B(n20569), .Y(n20570) );
  sky130_fd_sc_hd__nand2_1 U26523 ( .A(n20854), .B(n20570), .Y(n20571) );
  sky130_fd_sc_hd__a22oi_1 U26524 ( .A1(n20856), .A2(n20572), .B1(n20571), 
        .B2(n20833), .Y(n20573) );
  sky130_fd_sc_hd__nand3_1 U26525 ( .A(n20575), .B(n20574), .C(n20573), .Y(
        n20576) );
  sky130_fd_sc_hd__nand2_1 U26526 ( .A(n20576), .B(n20757), .Y(n20577) );
  sky130_fd_sc_hd__o211ai_1 U26527 ( .A1(n20580), .A2(n20579), .B1(n20578), 
        .C1(n20577), .Y(n20581) );
  sky130_fd_sc_hd__a21oi_1 U26528 ( .A1(j202_soc_core_memory0_ram_dout0[488]), 
        .A2(n11207), .B1(n20581), .Y(n20582) );
  sky130_fd_sc_hd__nand2_1 U26529 ( .A(n21693), .B(n21919), .Y(n20584) );
  sky130_fd_sc_hd__a22oi_1 U26530 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__8_), .B1(n21916), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__8_), .Y(n20583) );
  sky130_fd_sc_hd__a22oi_1 U26531 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__9_), .B1(n21916), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__9_), .Y(n20587) );
  sky130_fd_sc_hd__nand2_1 U26532 ( .A(j202_soc_core_memory0_ram_dout0[137]), 
        .B(n21489), .Y(n20592) );
  sky130_fd_sc_hd__nand2_1 U26533 ( .A(j202_soc_core_memory0_ram_dout0[73]), 
        .B(n21642), .Y(n20591) );
  sky130_fd_sc_hd__nand2_1 U26534 ( .A(j202_soc_core_memory0_ram_dout0[201]), 
        .B(n21640), .Y(n20590) );
  sky130_fd_sc_hd__nand2_1 U26535 ( .A(j202_soc_core_memory0_ram_dout0[105]), 
        .B(n21488), .Y(n20589) );
  sky130_fd_sc_hd__nand2b_1 U26536 ( .A_N(n20595), .B(n20594), .Y(n20597) );
  sky130_fd_sc_hd__o21ai_1 U26537 ( .A1(n20597), .A2(n20596), .B1(n20856), .Y(
        n20616) );
  sky130_fd_sc_hd__nand4_1 U26538 ( .A(n20794), .B(n20793), .C(n20741), .D(
        n20799), .Y(n20600) );
  sky130_fd_sc_hd__nor2_1 U26539 ( .A(n20598), .B(n20737), .Y(n20747) );
  sky130_fd_sc_hd__nand3_1 U26540 ( .A(n20739), .B(n20687), .C(n20599), .Y(
        n20628) );
  sky130_fd_sc_hd__nand2_1 U26541 ( .A(n20602), .B(n20850), .Y(n20615) );
  sky130_fd_sc_hd__nand3_1 U26542 ( .A(n20852), .B(n20793), .C(n20623), .Y(
        n20683) );
  sky130_fd_sc_hd__nor2_1 U26543 ( .A(n20605), .B(n20604), .Y(n20606) );
  sky130_fd_sc_hd__nand4_1 U26544 ( .A(n20608), .B(n20607), .C(n20606), .D(
        n20746), .Y(n20609) );
  sky130_fd_sc_hd__nand2_1 U26545 ( .A(n20609), .B(n20804), .Y(n20614) );
  sky130_fd_sc_hd__nand4_1 U26546 ( .A(n20610), .B(n20840), .C(n20767), .D(
        n20766), .Y(n20611) );
  sky130_fd_sc_hd__o21ai_1 U26547 ( .A1(n20612), .A2(n20611), .B1(n20833), .Y(
        n20613) );
  sky130_fd_sc_hd__nand4_1 U26548 ( .A(n20616), .B(n20615), .C(n20614), .D(
        n20613), .Y(n20618) );
  sky130_fd_sc_hd__nand2_1 U26549 ( .A(n20618), .B(n20617), .Y(n20710) );
  sky130_fd_sc_hd__o2bb2ai_1 U26550 ( .B1(n20619), .B2(n21515), .A1_N(
        j202_soc_core_ahblite_interconnect_s_hrdata[105]), .A2_N(n21446), .Y(
        n20703) );
  sky130_fd_sc_hd__nor2_1 U26551 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[0]), 
        .B(n29278), .Y(n20620) );
  sky130_fd_sc_hd__xor2_1 U26552 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[1]), 
        .B(j202_soc_core_uart_TOP_tx_fifo_wp[1]), .X(n27925) );
  sky130_fd_sc_hd__nor2_1 U26553 ( .A(n20620), .B(n27925), .Y(n28586) );
  sky130_fd_sc_hd__nand2_1 U26554 ( .A(n29278), .B(
        j202_soc_core_uart_TOP_tx_fifo_wp[0]), .Y(n28584) );
  sky130_fd_sc_hd__nand4_1 U26555 ( .A(n21513), .B(n28586), .C(
        j202_soc_core_uart_TOP_tx_fifo_gb), .D(n28584), .Y(n20704) );
  sky130_fd_sc_hd__nand2b_1 U26556 ( .A_N(n21512), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[73]), .Y(n20702) );
  sky130_fd_sc_hd__nand2_1 U26557 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[9]), .Y(n20701) );
  sky130_fd_sc_hd__nand4_1 U26558 ( .A(n20704), .B(n21768), .C(n20702), .D(
        n20701), .Y(n20621) );
  sky130_fd_sc_hd__nor2_1 U26559 ( .A(n20703), .B(n20621), .Y(n20622) );
  sky130_fd_sc_hd__nand2_1 U26560 ( .A(n20786), .B(
        j202_soc_core_bldc_core_00_pwm_period[9]), .Y(n20709) );
  sky130_fd_sc_hd__nand3_1 U26561 ( .A(n20710), .B(n20622), .C(n20709), .Y(
        n20696) );
  sky130_fd_sc_hd__nand2_1 U26562 ( .A(n20817), .B(n20741), .Y(n20651) );
  sky130_fd_sc_hd__nand3_1 U26563 ( .A(n20664), .B(n20623), .C(n20675), .Y(
        n20808) );
  sky130_fd_sc_hd__nor2_1 U26564 ( .A(n20626), .B(n20625), .Y(n20631) );
  sky130_fd_sc_hd__nand4_1 U26565 ( .A(n20637), .B(n20814), .C(n20774), .D(
        n20680), .Y(n20627) );
  sky130_fd_sc_hd__nor2_1 U26566 ( .A(n20628), .B(n20627), .Y(n20629) );
  sky130_fd_sc_hd__o22a_1 U26567 ( .A1(n20632), .A2(n20631), .B1(n20630), .B2(
        n20629), .X(n20641) );
  sky130_fd_sc_hd__nor3_1 U26568 ( .A(n20634), .B(n20633), .C(n20663), .Y(
        n20636) );
  sky130_fd_sc_hd__nand4_1 U26569 ( .A(n20638), .B(n20637), .C(n20636), .D(
        n20635), .Y(n20639) );
  sky130_fd_sc_hd__nand2_1 U26570 ( .A(n20639), .B(n20856), .Y(n20640) );
  sky130_fd_sc_hd__nand3_1 U26571 ( .A(n20642), .B(n20641), .C(n20640), .Y(
        n20644) );
  sky130_fd_sc_hd__nand2_1 U26572 ( .A(n20644), .B(n20643), .Y(n20695) );
  sky130_fd_sc_hd__nand2_1 U26573 ( .A(n20775), .B(n20799), .Y(n20647) );
  sky130_fd_sc_hd__nor2_1 U26574 ( .A(n20647), .B(n20646), .Y(n20648) );
  sky130_fd_sc_hd__nand3_1 U26575 ( .A(n20649), .B(n20802), .C(n20648), .Y(
        n20650) );
  sky130_fd_sc_hd__nor2_1 U26577 ( .A(n20652), .B(n20651), .Y(n20752) );
  sky130_fd_sc_hd__nand4_1 U26578 ( .A(n20752), .B(n20654), .C(n20775), .D(
        n20794), .Y(n20655) );
  sky130_fd_sc_hd__nand2_1 U26579 ( .A(n20655), .B(n20850), .Y(n20670) );
  sky130_fd_sc_hd__nand2_1 U26580 ( .A(n20767), .B(n20656), .Y(n20657) );
  sky130_fd_sc_hd__nor2_1 U26581 ( .A(n20657), .B(n20765), .Y(n20658) );
  sky130_fd_sc_hd__nand3_1 U26582 ( .A(n20740), .B(n20658), .C(n20794), .Y(
        n20660) );
  sky130_fd_sc_hd__o21ai_0 U26583 ( .A1(n20660), .A2(n20659), .B1(n20856), .Y(
        n20669) );
  sky130_fd_sc_hd__nand4_1 U26584 ( .A(n20662), .B(n20847), .C(n20661), .D(
        n20736), .Y(n20666) );
  sky130_fd_sc_hd__nand4b_1 U26585 ( .A_N(n20666), .B(n20665), .C(n20664), .D(
        n20819), .Y(n20667) );
  sky130_fd_sc_hd__nand2_1 U26586 ( .A(n20667), .B(n20804), .Y(n20668) );
  sky130_fd_sc_hd__nand4_1 U26587 ( .A(n20671), .B(n20670), .C(n20669), .D(
        n20668), .Y(n20672) );
  sky130_fd_sc_hd__nand2_1 U26588 ( .A(n20672), .B(n20757), .Y(n20694) );
  sky130_fd_sc_hd__nand3_1 U26589 ( .A(n20674), .B(
        j202_soc_core_bootrom_00_address_w[4]), .C(n20673), .Y(n20676) );
  sky130_fd_sc_hd__nand2_1 U26590 ( .A(n20676), .B(n20675), .Y(n20770) );
  sky130_fd_sc_hd__nor2_1 U26591 ( .A(n20677), .B(n20770), .Y(n20678) );
  sky130_fd_sc_hd__nand4_1 U26592 ( .A(n20679), .B(n20678), .C(n20840), .D(
        n20794), .Y(n20685) );
  sky130_fd_sc_hd__nand2_1 U26593 ( .A(n20680), .B(n20799), .Y(n20681) );
  sky130_fd_sc_hd__nand4b_1 U26594 ( .A_N(n20681), .B(n20742), .C(n20830), .D(
        n20829), .Y(n20682) );
  sky130_fd_sc_hd__nor2_1 U26595 ( .A(n20683), .B(n20682), .Y(n20779) );
  sky130_fd_sc_hd__a2bb2oi_1 U26596 ( .B1(n20804), .B2(n20685), .A1_N(n20684), 
        .A2_N(n20779), .Y(n20691) );
  sky130_fd_sc_hd__nand2_1 U26597 ( .A(n20686), .B(n20850), .Y(n20690) );
  sky130_fd_sc_hd__nand3_1 U26598 ( .A(n20774), .B(n20687), .C(n20767), .Y(
        n20688) );
  sky130_fd_sc_hd__o21ai_1 U26599 ( .A1(n20688), .A2(n20763), .B1(n20833), .Y(
        n20689) );
  sky130_fd_sc_hd__nand3_1 U26600 ( .A(n20691), .B(n20690), .C(n20689), .Y(
        n20692) );
  sky130_fd_sc_hd__nand2_1 U26601 ( .A(n20692), .B(n20784), .Y(n20693) );
  sky130_fd_sc_hd__nand3_1 U26602 ( .A(n20695), .B(n20694), .C(n20693), .Y(
        n20700) );
  sky130_fd_sc_hd__nor2_1 U26603 ( .A(n20696), .B(n20700), .Y(n20697) );
  sky130_fd_sc_hd__nand2_1 U26604 ( .A(j202_soc_core_memory0_ram_dout0[329]), 
        .B(n21490), .Y(n20699) );
  sky130_fd_sc_hd__nand2_1 U26605 ( .A(j202_soc_core_memory0_ram_dout0[265]), 
        .B(n21634), .Y(n20698) );
  sky130_fd_sc_hd__nand2_1 U26606 ( .A(j202_soc_core_memory0_ram_dout0[489]), 
        .B(n21650), .Y(n20715) );
  sky130_fd_sc_hd__nand3_1 U26607 ( .A(n20702), .B(n21653), .C(n20701), .Y(
        n20707) );
  sky130_fd_sc_hd__nand2_1 U26608 ( .A(n20705), .B(n20704), .Y(n20706) );
  sky130_fd_sc_hd__nor2_1 U26609 ( .A(n20707), .B(n20706), .Y(n20708) );
  sky130_fd_sc_hd__nand2_1 U26610 ( .A(n20709), .B(n20708), .Y(n20712) );
  sky130_fd_sc_hd__nor2_1 U26611 ( .A(n20712), .B(n20711), .Y(n20713) );
  sky130_fd_sc_hd__nand3_1 U26612 ( .A(n20715), .B(n20714), .C(n20713), .Y(
        n21335) );
  sky130_fd_sc_hd__a22oi_1 U26613 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__10_), .B1(n21916), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__10_), .Y(n20718) );
  sky130_fd_sc_hd__nand2_1 U26614 ( .A(j202_soc_core_memory0_ram_dout0[459]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n20724) );
  sky130_fd_sc_hd__nand2_1 U26615 ( .A(j202_soc_core_memory0_ram_dout0[235]), 
        .B(n21641), .Y(n20723) );
  sky130_fd_sc_hd__nand2_1 U26616 ( .A(j202_soc_core_memory0_ram_dout0[11]), 
        .B(n21639), .Y(n20722) );
  sky130_fd_sc_hd__nand2_1 U26617 ( .A(j202_soc_core_memory0_ram_dout0[299]), 
        .B(n21503), .Y(n20721) );
  sky130_fd_sc_hd__nand2_1 U26619 ( .A(j202_soc_core_memory0_ram_dout0[43]), 
        .B(n21633), .Y(n20728) );
  sky130_fd_sc_hd__nand2_1 U26620 ( .A(j202_soc_core_memory0_ram_dout0[331]), 
        .B(n21490), .Y(n20727) );
  sky130_fd_sc_hd__nand2_1 U26621 ( .A(j202_soc_core_memory0_ram_dout0[267]), 
        .B(n21634), .Y(n20726) );
  sky130_fd_sc_hd__nand2_1 U26622 ( .A(j202_soc_core_memory0_ram_dout0[395]), 
        .B(n21496), .Y(n20725) );
  sky130_fd_sc_hd__nand2_1 U26624 ( .A(j202_soc_core_memory0_ram_dout0[171]), 
        .B(n21487), .Y(n20867) );
  sky130_fd_sc_hd__nand2_1 U26625 ( .A(j202_soc_core_memory0_ram_dout0[139]), 
        .B(n21489), .Y(n20866) );
  sky130_fd_sc_hd__nor2_1 U26626 ( .A(n20732), .B(n20731), .Y(n20733) );
  sky130_fd_sc_hd__nand4b_1 U26627 ( .A_N(n20821), .B(n20847), .C(n20734), .D(
        n20733), .Y(n20735) );
  sky130_fd_sc_hd__nand2_1 U26628 ( .A(n20735), .B(n20804), .Y(n20756) );
  sky130_fd_sc_hd__nand2_1 U26629 ( .A(n20794), .B(n20736), .Y(n20738) );
  sky130_fd_sc_hd__nor2_1 U26630 ( .A(n20738), .B(n20737), .Y(n20751) );
  sky130_fd_sc_hd__nand4_1 U26631 ( .A(n20751), .B(n20740), .C(n20739), .D(
        n20799), .Y(n20750) );
  sky130_fd_sc_hd__nand3_1 U26632 ( .A(n20794), .B(n20742), .C(n20741), .Y(
        n20748) );
  sky130_fd_sc_hd__nor2_1 U26633 ( .A(n20744), .B(n20743), .Y(n20745) );
  sky130_fd_sc_hd__nand4b_1 U26634 ( .A_N(n20748), .B(n20747), .C(n20746), .D(
        n20745), .Y(n20749) );
  sky130_fd_sc_hd__a22oi_1 U26635 ( .A1(n20750), .A2(n20856), .B1(n20749), 
        .B2(n20833), .Y(n20755) );
  sky130_fd_sc_hd__nand4_1 U26636 ( .A(n20752), .B(n20751), .C(n20852), .D(
        n20837), .Y(n20753) );
  sky130_fd_sc_hd__nand2_1 U26637 ( .A(n20753), .B(n20850), .Y(n20754) );
  sky130_fd_sc_hd__nand3_1 U26638 ( .A(n20756), .B(n20755), .C(n20754), .Y(
        n20758) );
  sky130_fd_sc_hd__nand2_1 U26639 ( .A(n20758), .B(n20757), .Y(n20879) );
  sky130_fd_sc_hd__nand2b_1 U26640 ( .A_N(n21515), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[43]), .Y(n20873) );
  sky130_fd_sc_hd__nand2_1 U26641 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[11]), .Y(n20872) );
  sky130_fd_sc_hd__nand3_1 U26642 ( .A(n20873), .B(n21768), .C(n20872), .Y(
        n20761) );
  sky130_fd_sc_hd__o2bb2ai_1 U26643 ( .B1(n20760), .B2(n21519), .A1_N(
        j202_soc_core_ahblite_interconnect_s_hrdata[75]), .A2_N(n20759), .Y(
        n20874) );
  sky130_fd_sc_hd__nor2_1 U26644 ( .A(n20761), .B(n20874), .Y(n20787) );
  sky130_fd_sc_hd__nand2_1 U26645 ( .A(n20838), .B(n20762), .Y(n20764) );
  sky130_fd_sc_hd__nand4b_1 U26647 ( .A_N(n20844), .B(n20768), .C(n20767), .D(
        n20766), .Y(n20773) );
  sky130_fd_sc_hd__nor3_1 U26648 ( .A(n20771), .B(n20770), .C(n20769), .Y(
        n20772) );
  sky130_fd_sc_hd__a2bb2oi_1 U26649 ( .B1(n20850), .B2(n20773), .A1_N(n20772), 
        .A2_N(n20846), .Y(n20782) );
  sky130_fd_sc_hd__nand4_1 U26650 ( .A(n20775), .B(n20831), .C(n20774), .D(
        n20840), .Y(n20776) );
  sky130_fd_sc_hd__nor2_1 U26651 ( .A(n20777), .B(n20776), .Y(n20778) );
  sky130_fd_sc_hd__nand2_1 U26652 ( .A(n20779), .B(n20778), .Y(n20780) );
  sky130_fd_sc_hd__nand2_1 U26653 ( .A(n20780), .B(n20856), .Y(n20781) );
  sky130_fd_sc_hd__nand3_1 U26654 ( .A(n20783), .B(n20782), .C(n20781), .Y(
        n20785) );
  sky130_fd_sc_hd__nand2_1 U26655 ( .A(n20785), .B(n20784), .Y(n20877) );
  sky130_fd_sc_hd__nand2_1 U26656 ( .A(n20786), .B(
        j202_soc_core_bldc_core_00_pwm_period[11]), .Y(n20876) );
  sky130_fd_sc_hd__nand4_1 U26657 ( .A(n20879), .B(n20787), .C(n20877), .D(
        n20876), .Y(n20864) );
  sky130_fd_sc_hd__nor2_1 U26658 ( .A(n20789), .B(n20788), .Y(n20791) );
  sky130_fd_sc_hd__nand4_1 U26659 ( .A(n20840), .B(n20792), .C(n20791), .D(
        n20790), .Y(n20796) );
  sky130_fd_sc_hd__nand2_1 U26660 ( .A(n20794), .B(n20793), .Y(n20795) );
  sky130_fd_sc_hd__nor2_1 U26661 ( .A(n20796), .B(n20795), .Y(n20797) );
  sky130_fd_sc_hd__nand3_1 U26662 ( .A(n20798), .B(n20820), .C(n20797), .Y(
        n20806) );
  sky130_fd_sc_hd__nor2_1 U26663 ( .A(n20800), .B(n20815), .Y(n20801) );
  sky130_fd_sc_hd__nand4_1 U26664 ( .A(n20803), .B(n20802), .C(n20838), .D(
        n20801), .Y(n20805) );
  sky130_fd_sc_hd__a22oi_1 U26665 ( .A1(n20806), .A2(n20850), .B1(n20805), 
        .B2(n20804), .Y(n20826) );
  sky130_fd_sc_hd__nand3_1 U26666 ( .A(n20810), .B(n20809), .C(n13182), .Y(
        n20811) );
  sky130_fd_sc_hd__nand3_1 U26667 ( .A(n20853), .B(n20812), .C(n20811), .Y(
        n20813) );
  sky130_fd_sc_hd__nand2_1 U26668 ( .A(n20813), .B(n20856), .Y(n20825) );
  sky130_fd_sc_hd__nor2_1 U26669 ( .A(n20816), .B(n20815), .Y(n20818) );
  sky130_fd_sc_hd__nand4_1 U26670 ( .A(n20820), .B(n20819), .C(n20818), .D(
        n20817), .Y(n20822) );
  sky130_fd_sc_hd__o21ai_1 U26671 ( .A1(n20822), .A2(n20821), .B1(n20833), .Y(
        n20824) );
  sky130_fd_sc_hd__a31oi_1 U26672 ( .A1(n20826), .A2(n20825), .A3(n20824), 
        .B1(n20823), .Y(n20863) );
  sky130_fd_sc_hd__nor2_1 U26673 ( .A(n20828), .B(n20827), .Y(n20832) );
  sky130_fd_sc_hd__nand4_1 U26674 ( .A(n20832), .B(n20831), .C(n20830), .D(
        n20829), .Y(n20835) );
  sky130_fd_sc_hd__nand4_1 U26676 ( .A(n20839), .B(n20838), .C(n20837), .D(
        n20836), .Y(n20851) );
  sky130_fd_sc_hd__nand4_1 U26677 ( .A(n20843), .B(n20842), .C(n20841), .D(
        n20840), .Y(n20845) );
  sky130_fd_sc_hd__nor2_1 U26678 ( .A(n20845), .B(n20844), .Y(n20848) );
  sky130_fd_sc_hd__a21oi_1 U26679 ( .A1(n20848), .A2(n20847), .B1(n20846), .Y(
        n20849) );
  sky130_fd_sc_hd__a21oi_1 U26680 ( .A1(n20851), .A2(n20850), .B1(n20849), .Y(
        n20860) );
  sky130_fd_sc_hd__nand3_1 U26681 ( .A(n20854), .B(n20853), .C(n20852), .Y(
        n20857) );
  sky130_fd_sc_hd__a21oi_1 U26682 ( .A1(n20857), .A2(n20856), .B1(n20855), .Y(
        n20859) );
  sky130_fd_sc_hd__a31oi_1 U26683 ( .A1(n20861), .A2(n20860), .A3(n20859), 
        .B1(n20858), .Y(n20862) );
  sky130_fd_sc_hd__nor2_1 U26684 ( .A(n20864), .B(n20880), .Y(n20865) );
  sky130_fd_sc_hd__nand2_1 U26685 ( .A(j202_soc_core_memory0_ram_dout0[203]), 
        .B(n21640), .Y(n20871) );
  sky130_fd_sc_hd__nand2_1 U26686 ( .A(j202_soc_core_memory0_ram_dout0[107]), 
        .B(n21488), .Y(n20870) );
  sky130_fd_sc_hd__nand2_1 U26687 ( .A(j202_soc_core_memory0_ram_dout0[427]), 
        .B(n12156), .Y(n20869) );
  sky130_fd_sc_hd__nand2_1 U26688 ( .A(j202_soc_core_memory0_ram_dout0[363]), 
        .B(n21495), .Y(n20868) );
  sky130_fd_sc_hd__nand2_1 U26689 ( .A(j202_soc_core_memory0_ram_dout0[491]), 
        .B(n21650), .Y(n20883) );
  sky130_fd_sc_hd__nand3_1 U26690 ( .A(n20873), .B(n21653), .C(n20872), .Y(
        n20875) );
  sky130_fd_sc_hd__nor2_1 U26691 ( .A(n20875), .B(n20874), .Y(n20878) );
  sky130_fd_sc_hd__nand4_1 U26692 ( .A(n20879), .B(n20878), .C(n20877), .D(
        n20876), .Y(n20881) );
  sky130_fd_sc_hd__nor2_1 U26693 ( .A(n20881), .B(n20880), .Y(n20882) );
  sky130_fd_sc_hd__nand2_1 U26694 ( .A(n20883), .B(n20882), .Y(n21175) );
  sky130_fd_sc_hd__a22oi_1 U26695 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__11_), .B1(n21916), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__11_), .Y(n20884) );
  sky130_fd_sc_hd__a21oi_1 U26696 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__12_), .B1(n20885), .Y(n20887) );
  sky130_fd_sc_hd__nor2_1 U26697 ( .A(n21042), .B(n24143), .Y(n20891) );
  sky130_fd_sc_hd__xnor2_1 U26698 ( .A(n20889), .B(n12421), .Y(n20890) );
  sky130_fd_sc_hd__nand3_1 U26699 ( .A(n20895), .B(n11208), .C(n20894), .Y(
        n20896) );
  sky130_fd_sc_hd__nand3_1 U26701 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[2]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_sck), .C(n29828), .Y(n25202) );
  sky130_fd_sc_hd__nor2_1 U26702 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .B(n25202), .Y(n23852) );
  sky130_fd_sc_hd__nand2_1 U26703 ( .A(n23852), .B(n24030), .Y(n28692) );
  sky130_fd_sc_hd__nand2b_1 U26704 ( .A_N(n29603), .B(n28692), .Y(n29267) );
  sky130_fd_sc_hd__nand2_1 U26705 ( .A(n26623), .B(
        j202_soc_core_wbqspiflash_00_spi_wr), .Y(n26600) );
  sky130_fd_sc_hd__nand2_1 U26706 ( .A(n29267), .B(n26600), .Y(n26665) );
  sky130_fd_sc_hd__nor2_1 U26707 ( .A(n24030), .B(n25202), .Y(n24029) );
  sky130_fd_sc_hd__nand2_1 U26708 ( .A(n26665), .B(n26664), .Y(n29563) );
  sky130_fd_sc_hd__nand4_1 U26709 ( .A(n20904), .B(n20901), .C(n20903), .D(
        n20902), .Y(n20909) );
  sky130_fd_sc_hd__nor2_1 U26710 ( .A(n20909), .B(n20908), .Y(n20920) );
  sky130_fd_sc_hd__nand3_1 U26711 ( .A(n20912), .B(n20911), .C(n20910), .Y(
        n20918) );
  sky130_fd_sc_hd__nand4_1 U26712 ( .A(n20916), .B(n20915), .C(n20913), .D(
        n20914), .Y(n20917) );
  sky130_fd_sc_hd__nor2_1 U26713 ( .A(n20918), .B(n20917), .Y(n20919) );
  sky130_fd_sc_hd__nand2_1 U26714 ( .A(n20920), .B(n20919), .Y(n21825) );
  sky130_fd_sc_hd__nor2_1 U26715 ( .A(n21768), .B(
        j202_soc_core_memory0_ram_dout0[492]), .Y(n20921) );
  sky130_fd_sc_hd__nor2_1 U26716 ( .A(n21816), .B(n20921), .Y(n20922) );
  sky130_fd_sc_hd__and4_1 U26718 ( .A(n20926), .B(n20925), .C(n20924), .D(
        n21817), .X(n20927) );
  sky130_fd_sc_hd__nand2_1 U26719 ( .A(n20928), .B(n20927), .Y(n29487) );
  sky130_fd_sc_hd__nand2_1 U26720 ( .A(n29487), .B(n22739), .Y(n20947) );
  sky130_fd_sc_hd__nand2_1 U26721 ( .A(n22698), .B(n20931), .Y(n21177) );
  sky130_fd_sc_hd__nor2_1 U26722 ( .A(n14009), .B(n21177), .Y(n20932) );
  sky130_fd_sc_hd__xnor2_1 U26723 ( .A(n20933), .B(n20932), .Y(n26026) );
  sky130_fd_sc_hd__nand2_1 U26724 ( .A(n22747), .B(n26026), .Y(n20935) );
  sky130_fd_sc_hd__nand2_1 U26725 ( .A(n21924), .B(n28460), .Y(n20934) );
  sky130_fd_sc_hd__o211a_2 U26726 ( .A1(n26318), .A2(n11186), .B1(n20935), 
        .C1(n20934), .X(n20946) );
  sky130_fd_sc_hd__o21ai_1 U26727 ( .A1(n20937), .A2(n22752), .B1(n20936), .Y(
        n20965) );
  sky130_fd_sc_hd__a21oi_1 U26728 ( .A1(n20965), .A2(n21181), .B1(n20939), .Y(
        n20944) );
  sky130_fd_sc_hd__nand2_1 U26729 ( .A(n20942), .B(n20941), .Y(n20943) );
  sky130_fd_sc_hd__xor2_1 U26730 ( .A(n20944), .B(n20943), .X(n26016) );
  sky130_fd_sc_hd__nand2_1 U26731 ( .A(n26016), .B(n17225), .Y(n20945) );
  sky130_fd_sc_hd__nor2_1 U26732 ( .A(n20948), .B(n11378), .Y(n20949) );
  sky130_fd_sc_hd__nor2_1 U26733 ( .A(n21768), .B(
        j202_soc_core_memory0_ram_dout0[493]), .Y(n20951) );
  sky130_fd_sc_hd__nor2_1 U26734 ( .A(n21816), .B(n20951), .Y(n20952) );
  sky130_fd_sc_hd__o21ai_1 U26735 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .A2(n22224), .B1(n20952), 
        .Y(n20959) );
  sky130_fd_sc_hd__nand2_1 U26736 ( .A(n20954), .B(n20953), .Y(n20956) );
  sky130_fd_sc_hd__nor2_1 U26737 ( .A(n20956), .B(n20955), .Y(n20958) );
  sky130_fd_sc_hd__nand3_1 U26738 ( .A(n20959), .B(n20958), .C(n20957), .Y(
        n29564) );
  sky130_fd_sc_hd__nand2_1 U26739 ( .A(n29564), .B(n22739), .Y(n20972) );
  sky130_fd_sc_hd__nand2_1 U26740 ( .A(n22698), .B(n20960), .Y(n21003) );
  sky130_fd_sc_hd__xnor2_1 U26741 ( .A(n14175), .B(n20978), .Y(n25423) );
  sky130_fd_sc_hd__o21ai_1 U26742 ( .A1(n25428), .A2(n22705), .B1(n20961), .Y(
        n20962) );
  sky130_fd_sc_hd__a21oi_1 U26743 ( .A1(n21924), .A2(n28454), .B1(n20962), .Y(
        n20971) );
  sky130_fd_sc_hd__nand2_1 U26744 ( .A(n21009), .B(n21007), .Y(n20969) );
  sky130_fd_sc_hd__o21ai_1 U26745 ( .A1(n20968), .A2(n21183), .B1(n20967), .Y(
        n21010) );
  sky130_fd_sc_hd__xnor2_1 U26746 ( .A(n20969), .B(n21010), .Y(n25430) );
  sky130_fd_sc_hd__nand2_1 U26747 ( .A(n25430), .B(n17225), .Y(n20970) );
  sky130_fd_sc_hd__nand3_1 U26748 ( .A(n20972), .B(n20971), .C(n20970), .Y(
        n29474) );
  sky130_fd_sc_hd__nand2_1 U26749 ( .A(n20973), .B(n21020), .Y(n20974) );
  sky130_fd_sc_hd__a21oi_1 U26750 ( .A1(n21689), .A2(n21690), .B1(n21691), .Y(
        n26181) );
  sky130_fd_sc_hd__nand2b_1 U26751 ( .A_N(n26181), .B(n22739), .Y(n20991) );
  sky130_fd_sc_hd__nand2_1 U26752 ( .A(n20978), .B(n20977), .Y(n20992) );
  sky130_fd_sc_hd__nor2_1 U26753 ( .A(n14563), .B(n20992), .Y(n20979) );
  sky130_fd_sc_hd__xnor2_1 U26754 ( .A(n22769), .B(n20979), .Y(n24862) );
  sky130_fd_sc_hd__o21ai_0 U26755 ( .A1(n28532), .A2(n22745), .B1(n20980), .Y(
        n20981) );
  sky130_fd_sc_hd__a21oi_1 U26756 ( .A1(n24862), .A2(n22747), .B1(n20981), .Y(
        n20990) );
  sky130_fd_sc_hd__a21oi_1 U26757 ( .A1(n17040), .A2(n20996), .B1(n20983), .Y(
        n20988) );
  sky130_fd_sc_hd__nand2_1 U26758 ( .A(n20986), .B(n20985), .Y(n20987) );
  sky130_fd_sc_hd__xor2_1 U26759 ( .A(n20988), .B(n20987), .X(n24865) );
  sky130_fd_sc_hd__nand2_1 U26760 ( .A(n24865), .B(n17225), .Y(n20989) );
  sky130_fd_sc_hd__nand3_1 U26761 ( .A(n20991), .B(n20990), .C(n20989), .Y(
        n29482) );
  sky130_fd_sc_hd__nand2b_1 U26762 ( .A_N(n26169), .B(n22739), .Y(n21000) );
  sky130_fd_sc_hd__xor2_1 U26763 ( .A(n20992), .B(n14563), .X(n26074) );
  sky130_fd_sc_hd__nand2_1 U26764 ( .A(n22747), .B(n26074), .Y(n20994) );
  sky130_fd_sc_hd__nand2_1 U26765 ( .A(n21924), .B(n28443), .Y(n20993) );
  sky130_fd_sc_hd__o211a_2 U26766 ( .A1(n26430), .A2(n11186), .B1(n20994), 
        .C1(n20993), .X(n20999) );
  sky130_fd_sc_hd__nand2_1 U26767 ( .A(n20996), .B(n20995), .Y(n20997) );
  sky130_fd_sc_hd__xnor2_1 U26768 ( .A(n20997), .B(n17040), .Y(n26069) );
  sky130_fd_sc_hd__nand2_1 U26769 ( .A(n26069), .B(n17225), .Y(n20998) );
  sky130_fd_sc_hd__nand3_1 U26770 ( .A(n21000), .B(n20999), .C(n20998), .Y(
        n29550) );
  sky130_fd_sc_hd__nand2_1 U26771 ( .A(n21002), .B(n21001), .Y(n25939) );
  sky130_fd_sc_hd__nand2b_1 U26772 ( .A_N(n25939), .B(n22739), .Y(n21018) );
  sky130_fd_sc_hd__nor2_1 U26773 ( .A(n14175), .B(n21003), .Y(n21004) );
  sky130_fd_sc_hd__xnor2_1 U26774 ( .A(n14143), .B(n21004), .Y(n25971) );
  sky130_fd_sc_hd__nand2_1 U26775 ( .A(n22747), .B(n25971), .Y(n21006) );
  sky130_fd_sc_hd__nand2_1 U26776 ( .A(n21924), .B(n28449), .Y(n21005) );
  sky130_fd_sc_hd__o211a_2 U26777 ( .A1(n26319), .A2(n11186), .B1(n21006), 
        .C1(n21005), .X(n21017) );
  sky130_fd_sc_hd__a21oi_1 U26778 ( .A1(n21010), .A2(n21009), .B1(n21008), .Y(
        n21015) );
  sky130_fd_sc_hd__nand2_1 U26779 ( .A(n21013), .B(n21012), .Y(n21014) );
  sky130_fd_sc_hd__xor2_1 U26780 ( .A(n21015), .B(n21014), .X(n25975) );
  sky130_fd_sc_hd__nand2_1 U26781 ( .A(n25975), .B(n17225), .Y(n21016) );
  sky130_fd_sc_hd__nand2_1 U26782 ( .A(n21021), .B(n21020), .Y(n21023) );
  sky130_fd_sc_hd__nand2_1 U26783 ( .A(n21932), .B(n21933), .Y(n26177) );
  sky130_fd_sc_hd__nand2_1 U26784 ( .A(n26177), .B(n22739), .Y(n21039) );
  sky130_fd_sc_hd__xor2_1 U26785 ( .A(n21026), .B(n22849), .X(n25725) );
  sky130_fd_sc_hd__nand2_1 U26786 ( .A(n22747), .B(n25725), .Y(n21028) );
  sky130_fd_sc_hd__nand2_1 U26787 ( .A(n21924), .B(n28526), .Y(n21027) );
  sky130_fd_sc_hd__a21oi_1 U26788 ( .A1(n17040), .A2(n21030), .B1(n21029), .Y(
        n21036) );
  sky130_fd_sc_hd__nand2_1 U26789 ( .A(n21034), .B(n21033), .Y(n21035) );
  sky130_fd_sc_hd__xor2_1 U26790 ( .A(n21036), .B(n21035), .X(n25728) );
  sky130_fd_sc_hd__nand2_1 U26791 ( .A(n25728), .B(n17225), .Y(n21037) );
  sky130_fd_sc_hd__nand3_1 U26792 ( .A(n21039), .B(n21038), .C(n21037), .Y(
        n29441) );
  sky130_fd_sc_hd__nor2_1 U26793 ( .A(n29473), .B(n29474), .Y(n25029) );
  sky130_fd_sc_hd__nand3_1 U26794 ( .A(n25029), .B(n21040), .C(n23623), .Y(
        n21048) );
  sky130_fd_sc_hd__nor2_1 U26795 ( .A(n29088), .B(n29547), .Y(n21047) );
  sky130_fd_sc_hd__nor2_2 U26796 ( .A(n21046), .B(n21045), .Y(n21316) );
  sky130_fd_sc_hd__nand3_1 U26797 ( .A(n24725), .B(n21049), .C(
        j202_soc_core_ahb2apb_00_state[1]), .Y(n24726) );
  sky130_fd_sc_hd__nand2_1 U26798 ( .A(n21050), .B(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[0]), .Y(n24728) );
  sky130_fd_sc_hd__nor2_1 U26799 ( .A(n24726), .B(n24728), .Y(n29485) );
  sky130_fd_sc_hd__nand2_1 U26800 ( .A(
        j202_soc_core_intc_core_00_in_intreq[16]), .B(
        j202_soc_core_intc_core_00_rg_itgt[16]), .Y(n23286) );
  sky130_fd_sc_hd__nand2_1 U26801 ( .A(
        j202_soc_core_intc_core_00_in_intreq[17]), .B(
        j202_soc_core_intc_core_00_rg_itgt[17]), .Y(n23285) );
  sky130_fd_sc_hd__nand2_1 U26802 ( .A(n23286), .B(n23285), .Y(n23313) );
  sky130_fd_sc_hd__nand2_1 U26803 ( .A(
        j202_soc_core_intc_core_00_in_intreq[19]), .B(
        j202_soc_core_intc_core_00_rg_itgt[19]), .Y(n23295) );
  sky130_fd_sc_hd__nand2_1 U26804 ( .A(
        j202_soc_core_intc_core_00_in_intreq[18]), .B(
        j202_soc_core_intc_core_00_rg_itgt[18]), .Y(n23294) );
  sky130_fd_sc_hd__nand2_1 U26805 ( .A(n23295), .B(n23294), .Y(n23307) );
  sky130_fd_sc_hd__nor2_1 U26806 ( .A(n23313), .B(n23307), .Y(n23344) );
  sky130_fd_sc_hd__nand2_1 U26807 ( .A(
        j202_soc_core_intc_core_00_in_intreq[20]), .B(
        j202_soc_core_intc_core_00_rg_itgt[20]), .Y(n23341) );
  sky130_fd_sc_hd__nand2_1 U26808 ( .A(n23344), .B(n23341), .Y(n23372) );
  sky130_fd_sc_hd__nand2_1 U26809 ( .A(j202_soc_core_intc_core_00_in_intreq[0]), .B(j202_soc_core_intc_core_00_rg_itgt[0]), .Y(n23169) );
  sky130_fd_sc_hd__nand2_1 U26810 ( .A(j202_soc_core_intc_core_00_in_intreq[1]), .B(j202_soc_core_intc_core_00_rg_itgt[1]), .Y(n23166) );
  sky130_fd_sc_hd__nand2_1 U26811 ( .A(n23169), .B(n23166), .Y(n23180) );
  sky130_fd_sc_hd__nand2_1 U26812 ( .A(j202_soc_core_intc_core_00_in_intreq[3]), .B(j202_soc_core_intc_core_00_rg_itgt[3]), .Y(n23157) );
  sky130_fd_sc_hd__nand2_1 U26813 ( .A(j202_soc_core_intc_core_00_in_intreq[2]), .B(j202_soc_core_intc_core_00_rg_itgt[2]), .Y(n23158) );
  sky130_fd_sc_hd__nand2_1 U26814 ( .A(n23157), .B(n23158), .Y(n23173) );
  sky130_fd_sc_hd__nor2_1 U26815 ( .A(n23180), .B(n23173), .Y(n23248) );
  sky130_fd_sc_hd__nand2_1 U26816 ( .A(j202_soc_core_intc_core_00_in_intreq[4]), .B(j202_soc_core_intc_core_00_rg_itgt[4]), .Y(n23189) );
  sky130_fd_sc_hd__nand2_1 U26817 ( .A(j202_soc_core_intc_core_00_in_intreq[5]), .B(j202_soc_core_intc_core_00_rg_itgt[5]), .Y(n23192) );
  sky130_fd_sc_hd__nand2_1 U26818 ( .A(n23189), .B(n23192), .Y(n23217) );
  sky130_fd_sc_hd__nand2_1 U26819 ( .A(j202_soc_core_intc_core_00_in_intreq[6]), .B(j202_soc_core_intc_core_00_rg_itgt[6]), .Y(n23199) );
  sky130_fd_sc_hd__nand2_1 U26820 ( .A(j202_soc_core_intc_core_00_in_intreq[7]), .B(j202_soc_core_intc_core_00_rg_itgt[7]), .Y(n23200) );
  sky130_fd_sc_hd__nand2_1 U26821 ( .A(n23199), .B(n23200), .Y(n23215) );
  sky130_fd_sc_hd__nor2_1 U26822 ( .A(n23217), .B(n23215), .Y(n23241) );
  sky130_fd_sc_hd__nand2_1 U26823 ( .A(n23248), .B(n23241), .Y(n23278) );
  sky130_fd_sc_hd__nand2_1 U26824 ( .A(
        j202_soc_core_intc_core_00_in_intreq[12]), .B(
        j202_soc_core_intc_core_00_rg_itgt[12]), .Y(n23062) );
  sky130_fd_sc_hd__nand2_1 U26825 ( .A(
        j202_soc_core_intc_core_00_in_intreq[13]), .B(
        j202_soc_core_intc_core_00_rg_itgt[13]), .Y(n23065) );
  sky130_fd_sc_hd__nand2_1 U26826 ( .A(n23062), .B(n23065), .Y(n23141) );
  sky130_fd_sc_hd__nand2_1 U26827 ( .A(j202_soc_core_intc_core_00_rg_itgt[8]), 
        .B(j202_soc_core_intc_core_00_in_intreq[8]), .Y(n23090) );
  sky130_fd_sc_hd__nand2_1 U26828 ( .A(j202_soc_core_intc_core_00_rg_itgt[9]), 
        .B(j202_soc_core_intc_core_00_in_intreq[9]), .Y(n23093) );
  sky130_fd_sc_hd__nand2_1 U26829 ( .A(n23090), .B(n23093), .Y(n23119) );
  sky130_fd_sc_hd__nand2_1 U26830 ( .A(
        j202_soc_core_intc_core_00_in_intreq[10]), .B(
        j202_soc_core_intc_core_00_rg_itgt[10]), .Y(n23100) );
  sky130_fd_sc_hd__nand2_1 U26831 ( .A(j202_soc_core_intc_core_00_rg_itgt[11]), 
        .B(j202_soc_core_intc_core_00_in_intreq[11]), .Y(n23101) );
  sky130_fd_sc_hd__nand2_1 U26832 ( .A(n23100), .B(n23101), .Y(n23117) );
  sky130_fd_sc_hd__nand2_1 U26833 ( .A(n21052), .B(n21051), .Y(n23146) );
  sky130_fd_sc_hd__nor2_1 U26834 ( .A(n23141), .B(n23146), .Y(n23272) );
  sky130_fd_sc_hd__nand2_1 U26835 ( .A(j202_soc_core_intc_core_00_rg_itgt[14]), 
        .B(j202_soc_core_intc_core_00_in_intreq[14]), .Y(n23072) );
  sky130_fd_sc_hd__nand2_1 U26836 ( .A(
        j202_soc_core_intc_core_00_in_intreq[15]), .B(
        j202_soc_core_intc_core_00_rg_itgt[15]), .Y(n23073) );
  sky130_fd_sc_hd__nand2_1 U26837 ( .A(n23072), .B(n23073), .Y(n23275) );
  sky130_fd_sc_hd__nand3_1 U26838 ( .A(n21054), .B(n23272), .C(n21053), .Y(
        n23376) );
  sky130_fd_sc_hd__nor2_1 U26839 ( .A(n23372), .B(n23376), .Y(n28377) );
  sky130_fd_sc_hd__nand2_1 U26840 ( .A(n28377), .B(n12069), .Y(n27711) );
  sky130_fd_sc_hd__nor2_1 U26841 ( .A(n29088), .B(n28377), .Y(n29480) );
  sky130_fd_sc_hd__nor3_1 U26843 ( .A(n28275), .B(n24302), .C(n21055), .Y(
        n21056) );
  sky130_fd_sc_hd__nand2_1 U26844 ( .A(j202_soc_core_memory0_ram_dout0[38]), 
        .B(n21633), .Y(n21059) );
  sky130_fd_sc_hd__nand2_1 U26845 ( .A(j202_soc_core_memory0_ram_dout0[230]), 
        .B(n21641), .Y(n21058) );
  sky130_fd_sc_hd__nand2_1 U26846 ( .A(j202_soc_core_memory0_ram_dout0[6]), 
        .B(n21639), .Y(n21057) );
  sky130_fd_sc_hd__nand2_1 U26847 ( .A(j202_soc_core_memory0_ram_dout0[134]), 
        .B(n21489), .Y(n21063) );
  sky130_fd_sc_hd__nand2_1 U26848 ( .A(j202_soc_core_memory0_ram_dout0[70]), 
        .B(n21642), .Y(n21062) );
  sky130_fd_sc_hd__nand2_1 U26849 ( .A(j202_soc_core_memory0_ram_dout0[198]), 
        .B(n21640), .Y(n21061) );
  sky130_fd_sc_hd__nand2_1 U26850 ( .A(j202_soc_core_memory0_ram_dout0[102]), 
        .B(n21488), .Y(n21060) );
  sky130_fd_sc_hd__nand2b_1 U26851 ( .A_N(n21515), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[38]), .Y(n21164) );
  sky130_fd_sc_hd__nand2_1 U26852 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[6]), .Y(n21163) );
  sky130_fd_sc_hd__nand3_1 U26853 ( .A(n21164), .B(n21768), .C(n21163), .Y(
        n21073) );
  sky130_fd_sc_hd__o22a_1 U26854 ( .A1(n21066), .A2(n21512), .B1(n21065), .B2(
        n21519), .X(n21162) );
  sky130_fd_sc_hd__nand2_1 U26855 ( .A(n21504), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[14]), .Y(n21070) );
  sky130_fd_sc_hd__nand2_1 U26856 ( .A(n24720), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[22]), .Y(n21069) );
  sky130_fd_sc_hd__nand2_1 U26857 ( .A(n21505), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[6]), .Y(n21068) );
  sky130_fd_sc_hd__nand2_1 U26858 ( .A(n21506), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[30]), .Y(n21067) );
  sky130_fd_sc_hd__nand4_1 U26859 ( .A(n21070), .B(n21069), .C(n21068), .D(
        n21067), .Y(n21071) );
  sky130_fd_sc_hd__nand2_1 U26860 ( .A(n21513), .B(n21071), .Y(n21165) );
  sky130_fd_sc_hd__nand2_1 U26861 ( .A(n21162), .B(n21165), .Y(n21072) );
  sky130_fd_sc_hd__nor2_1 U26862 ( .A(n27445), .B(n21517), .Y(n21166) );
  sky130_fd_sc_hd__nor3_1 U26863 ( .A(n21073), .B(n21072), .C(n21166), .Y(
        n21161) );
  sky130_fd_sc_hd__nand3_1 U26864 ( .A(n21360), .B(n21075), .C(n21074), .Y(
        n21394) );
  sky130_fd_sc_hd__nand4_1 U26865 ( .A(n21572), .B(n21607), .C(n21399), .D(
        n21365), .Y(n21618) );
  sky130_fd_sc_hd__o21ai_1 U26866 ( .A1(n21526), .A2(n21618), .B1(n21617), .Y(
        n21080) );
  sky130_fd_sc_hd__nand3_1 U26867 ( .A(n21380), .B(n21607), .C(n21593), .Y(
        n21078) );
  sky130_fd_sc_hd__nand2_1 U26868 ( .A(n21412), .B(n21395), .Y(n21087) );
  sky130_fd_sc_hd__o2bb2ai_1 U26869 ( .B1(n21395), .B2(n21550), .A1_N(n21087), 
        .A2_N(n21076), .Y(n21077) );
  sky130_fd_sc_hd__a21oi_1 U26870 ( .A1(n21078), .A2(n21610), .B1(n21077), .Y(
        n21079) );
  sky130_fd_sc_hd__nand2_1 U26871 ( .A(n21080), .B(n21079), .Y(n21540) );
  sky130_fd_sc_hd__nand4_1 U26872 ( .A(n21125), .B(n21575), .C(n21527), .D(
        n21568), .Y(n21081) );
  sky130_fd_sc_hd__nor2_1 U26873 ( .A(n21599), .B(n21081), .Y(n21539) );
  sky130_fd_sc_hd__nor2_1 U26874 ( .A(n21083), .B(n21082), .Y(n21084) );
  sky130_fd_sc_hd__nand4_1 U26875 ( .A(n21539), .B(n21085), .C(n21084), .D(
        n21521), .Y(n21086) );
  sky130_fd_sc_hd__nand2_1 U26876 ( .A(n21086), .B(n21598), .Y(n21094) );
  sky130_fd_sc_hd__a2bb2oi_1 U26877 ( .B1(n21087), .B2(n21426), .A1_N(n21412), 
        .A2_N(n21375), .Y(n21093) );
  sky130_fd_sc_hd__nand2b_1 U26878 ( .A_N(n21097), .B(n21088), .Y(n21576) );
  sky130_fd_sc_hd__nand2_1 U26879 ( .A(n21576), .B(n21567), .Y(n21089) );
  sky130_fd_sc_hd__nand2_1 U26880 ( .A(n21089), .B(n21603), .Y(n21092) );
  sky130_fd_sc_hd__nand4_1 U26882 ( .A(n21094), .B(n21093), .C(n21092), .D(
        n21091), .Y(n21095) );
  sky130_fd_sc_hd__nor2_1 U26883 ( .A(n21540), .B(n21095), .Y(n21159) );
  sky130_fd_sc_hd__nand2_1 U26884 ( .A(n21096), .B(n21388), .Y(n21366) );
  sky130_fd_sc_hd__nand4_1 U26885 ( .A(n21098), .B(n21408), .C(n21097), .D(
        n21573), .Y(n21100) );
  sky130_fd_sc_hd__o21ai_1 U26886 ( .A1(n21100), .A2(n21099), .B1(n21603), .Y(
        n21119) );
  sky130_fd_sc_hd__nand2_1 U26887 ( .A(n21102), .B(n21101), .Y(n21582) );
  sky130_fd_sc_hd__nand3_1 U26888 ( .A(n21365), .B(n21582), .C(n21606), .Y(
        n21108) );
  sky130_fd_sc_hd__nand3_1 U26889 ( .A(n21104), .B(n11150), .C(n21103), .Y(
        n21105) );
  sky130_fd_sc_hd__nand4_1 U26890 ( .A(n21380), .B(n21574), .C(n21394), .D(
        n21105), .Y(n21106) );
  sky130_fd_sc_hd__nor3_1 U26891 ( .A(n21108), .B(n21107), .C(n21106), .Y(
        n21113) );
  sky130_fd_sc_hd__nor2_1 U26892 ( .A(n21109), .B(n21142), .Y(n21111) );
  sky130_fd_sc_hd__nand4_1 U26893 ( .A(n21111), .B(n21110), .C(n21521), .D(
        n21606), .Y(n21414) );
  sky130_fd_sc_hd__nor3_1 U26894 ( .A(n21526), .B(n21137), .C(n21414), .Y(
        n21112) );
  sky130_fd_sc_hd__o22a_1 U26895 ( .A1(n21412), .A2(n21113), .B1(n21580), .B2(
        n21112), .X(n21118) );
  sky130_fd_sc_hd__nand2_1 U26896 ( .A(n21574), .B(n21415), .Y(n21601) );
  sky130_fd_sc_hd__nor2_1 U26897 ( .A(n21114), .B(n21601), .Y(n21115) );
  sky130_fd_sc_hd__nand4_1 U26898 ( .A(n21428), .B(n21413), .C(n21423), .D(
        n21115), .Y(n21116) );
  sky130_fd_sc_hd__nand2_1 U26899 ( .A(n21116), .B(n21598), .Y(n21117) );
  sky130_fd_sc_hd__nand3_1 U26900 ( .A(n21119), .B(n21118), .C(n21117), .Y(
        n21120) );
  sky130_fd_sc_hd__nand2_1 U26901 ( .A(n21120), .B(n21589), .Y(n21158) );
  sky130_fd_sc_hd__o31a_1 U26902 ( .A1(n21122), .A2(n21389), .A3(n21126), .B1(
        n21610), .X(n21123) );
  sky130_fd_sc_hd__nor2_1 U26903 ( .A(n21124), .B(n21123), .Y(n21136) );
  sky130_fd_sc_hd__and3_1 U26904 ( .A(n21576), .B(n21125), .C(n21607), .X(
        n21373) );
  sky130_fd_sc_hd__nand4_1 U26905 ( .A(n21373), .B(n21121), .C(n21593), .D(
        n21379), .Y(n21128) );
  sky130_fd_sc_hd__nand2_1 U26906 ( .A(n21128), .B(n21598), .Y(n21135) );
  sky130_fd_sc_hd__nor2_1 U26907 ( .A(n21129), .B(n21525), .Y(n21416) );
  sky130_fd_sc_hd__nand2b_1 U26908 ( .A_N(n21349), .B(n21416), .Y(n21130) );
  sky130_fd_sc_hd__nand2_1 U26909 ( .A(n21130), .B(n21617), .Y(n21370) );
  sky130_fd_sc_hd__nand2_1 U26910 ( .A(n21360), .B(n13179), .Y(n21594) );
  sky130_fd_sc_hd__o211ai_1 U26911 ( .A1(n21132), .A2(n21594), .B1(n21573), 
        .C1(n21593), .Y(n21133) );
  sky130_fd_sc_hd__nand2b_1 U26912 ( .A_N(n21605), .B(n21616), .Y(n21523) );
  sky130_fd_sc_hd__nand4_1 U26914 ( .A(n21136), .B(n21135), .C(n21370), .D(
        n21134), .Y(n21156) );
  sky130_fd_sc_hd__nor2_1 U26915 ( .A(n21138), .B(n21137), .Y(n21396) );
  sky130_fd_sc_hd__nor2_1 U26916 ( .A(n21146), .B(n21139), .Y(n21140) );
  sky130_fd_sc_hd__nand2_1 U26917 ( .A(n21396), .B(n21140), .Y(n21154) );
  sky130_fd_sc_hd__nor2_1 U26918 ( .A(n21556), .B(n21141), .Y(n21563) );
  sky130_fd_sc_hd__a31oi_1 U26919 ( .A1(n21563), .A2(n21394), .A3(n21399), 
        .B1(n21580), .Y(n21153) );
  sky130_fd_sc_hd__nand2_1 U26920 ( .A(n21616), .B(n21554), .Y(n21144) );
  sky130_fd_sc_hd__nand4_1 U26921 ( .A(n21555), .B(n21147), .C(n21364), .D(
        n21536), .Y(n21143) );
  sky130_fd_sc_hd__nor2_1 U26922 ( .A(n21144), .B(n21143), .Y(n21151) );
  sky130_fd_sc_hd__nand2_1 U26923 ( .A(n21146), .B(n21145), .Y(n21351) );
  sky130_fd_sc_hd__nand3_1 U26924 ( .A(n21351), .B(n21394), .C(n21147), .Y(
        n21609) );
  sky130_fd_sc_hd__nand3_1 U26925 ( .A(n21380), .B(n21415), .C(n21616), .Y(
        n21562) );
  sky130_fd_sc_hd__nor3_1 U26926 ( .A(n21609), .B(n21148), .C(n21562), .Y(
        n21149) );
  sky130_fd_sc_hd__o22ai_1 U26927 ( .A1(n21151), .A2(n21395), .B1(n21150), 
        .B2(n21149), .Y(n21152) );
  sky130_fd_sc_hd__a211o_1 U26928 ( .A1(n21617), .A2(n21154), .B1(n21153), 
        .C1(n21152), .X(n21155) );
  sky130_fd_sc_hd__a22oi_1 U26929 ( .A1(n21624), .A2(n21156), .B1(n21155), 
        .B2(n21591), .Y(n21157) );
  sky130_fd_sc_hd__o211ai_1 U26930 ( .A1(n21405), .A2(n21159), .B1(n21158), 
        .C1(n21157), .Y(n21160) );
  sky130_fd_sc_hd__nand2_1 U26931 ( .A(n21160), .B(n21629), .Y(n21169) );
  sky130_fd_sc_hd__nand2_1 U26932 ( .A(j202_soc_core_memory0_ram_dout0[486]), 
        .B(n21650), .Y(n21171) );
  sky130_fd_sc_hd__nand4_1 U26933 ( .A(n21165), .B(n21164), .C(n21653), .D(
        n21163), .Y(n21167) );
  sky130_fd_sc_hd__nor3_1 U26934 ( .A(n21168), .B(n21167), .C(n21166), .Y(
        n21170) );
  sky130_fd_sc_hd__nand3_1 U26935 ( .A(n21171), .B(n21170), .C(n21169), .Y(
        n21318) );
  sky130_fd_sc_hd__a22oi_1 U26936 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__6_), .B1(n21916), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__6_), .Y(n21172) );
  sky130_fd_sc_hd__nand2_1 U26938 ( .A(n21176), .B(n21175), .Y(n24068) );
  sky130_fd_sc_hd__nand2b_1 U26939 ( .A_N(n12409), .B(n22739), .Y(n21186) );
  sky130_fd_sc_hd__xor2_1 U26940 ( .A(n21177), .B(n14009), .X(n24070) );
  sky130_fd_sc_hd__a21oi_1 U26942 ( .A1(n21924), .A2(n28467), .B1(n21179), .Y(
        n21185) );
  sky130_fd_sc_hd__nand2_1 U26943 ( .A(n21181), .B(n21180), .Y(n21182) );
  sky130_fd_sc_hd__xor2_1 U26944 ( .A(n21183), .B(n21182), .X(n25926) );
  sky130_fd_sc_hd__nand2_1 U26945 ( .A(n25926), .B(n17225), .Y(n21184) );
  sky130_fd_sc_hd__nand2_1 U26946 ( .A(n24589), .B(n24912), .Y(n25025) );
  sky130_fd_sc_hd__nand3_1 U26947 ( .A(n11854), .B(n21188), .C(n25025), .Y(
        n25022) );
  sky130_fd_sc_hd__inv_1 U26948 ( .A(n25022), .Y(n23049) );
  sky130_fd_sc_hd__nand3_1 U26949 ( .A(n23049), .B(n23048), .C(n25052), .Y(
        n23051) );
  sky130_fd_sc_hd__nor2_1 U26950 ( .A(n23053), .B(n23051), .Y(n29532) );
  sky130_fd_sc_hd__nand2_1 U26951 ( .A(n21191), .B(n21190), .Y(n21199) );
  sky130_fd_sc_hd__nand2_1 U26952 ( .A(n22195), .B(n21195), .Y(n21197) );
  sky130_fd_sc_hd__a21oi_1 U26953 ( .A1(n22202), .A2(n21195), .B1(n21194), .Y(
        n21196) );
  sky130_fd_sc_hd__o21ai_2 U26954 ( .A1(n21197), .A2(n11866), .B1(n21196), .Y(
        n21198) );
  sky130_fd_sc_hd__xnor2_2 U26955 ( .A(n21199), .B(n21198), .Y(n23485) );
  sky130_fd_sc_hd__nand2_1 U26956 ( .A(n25263), .B(n21200), .Y(n21696) );
  sky130_fd_sc_hd__nand2_1 U26957 ( .A(n11190), .B(n26135), .Y(n26248) );
  sky130_fd_sc_hd__nand2_1 U26958 ( .A(n26334), .B(n28515), .Y(n26307) );
  sky130_fd_sc_hd__nand3_1 U26959 ( .A(n26248), .B(n25827), .C(n26307), .Y(
        n21202) );
  sky130_fd_sc_hd__o2bb2ai_1 U26961 ( .B1(n25818), .B2(n28515), .A1_N(n23532), 
        .A2_N(n25697), .Y(n21203) );
  sky130_fd_sc_hd__a21oi_1 U26962 ( .A1(n26334), .A2(n25824), .B1(n21203), .Y(
        n21205) );
  sky130_fd_sc_hd__nand2_1 U26963 ( .A(n23533), .B(n25692), .Y(n21204) );
  sky130_fd_sc_hd__o211ai_1 U26964 ( .A1(n26307), .A2(n21206), .B1(n21205), 
        .C1(n21204), .Y(n21207) );
  sky130_fd_sc_hd__nor2_1 U26965 ( .A(n21208), .B(n21207), .Y(n21209) );
  sky130_fd_sc_hd__o21a_1 U26966 ( .A1(n26135), .A2(n21210), .B1(n21209), .X(
        n21211) );
  sky130_fd_sc_hd__nand2_1 U26967 ( .A(n21212), .B(n21211), .Y(n21213) );
  sky130_fd_sc_hd__nand2_1 U26968 ( .A(n21213), .B(n26426), .Y(n21229) );
  sky130_fd_sc_hd__nand2_1 U26969 ( .A(n21216), .B(n21215), .Y(n21218) );
  sky130_fd_sc_hd__xor2_1 U26970 ( .A(n21218), .B(n21217), .X(n24329) );
  sky130_fd_sc_hd__nand2_1 U26971 ( .A(n24329), .B(n24461), .Y(n22442) );
  sky130_fd_sc_hd__nand2_1 U26972 ( .A(n23004), .B(n21219), .Y(n21220) );
  sky130_fd_sc_hd__o21a_1 U26973 ( .A1(n21221), .A2(n24463), .B1(n21220), .X(
        n22441) );
  sky130_fd_sc_hd__o22ai_1 U26974 ( .A1(n22441), .A2(n26926), .B1(n27025), 
        .B2(n26943), .Y(n21222) );
  sky130_fd_sc_hd__a21oi_1 U26975 ( .A1(n27808), .A2(n26375), .B1(n21222), .Y(
        n21226) );
  sky130_fd_sc_hd__o22ai_1 U26976 ( .A1(n27147), .A2(n27795), .B1(n27365), 
        .B2(n27803), .Y(n21224) );
  sky130_fd_sc_hd__o2bb2ai_1 U26977 ( .B1(n27027), .B2(n25996), .A1_N(n22260), 
        .A2_N(n27810), .Y(n21223) );
  sky130_fd_sc_hd__nor2_1 U26978 ( .A(n21224), .B(n21223), .Y(n21225) );
  sky130_fd_sc_hd__o211ai_1 U26979 ( .A1(n26926), .A2(n22442), .B1(n21226), 
        .C1(n21225), .Y(n21227) );
  sky130_fd_sc_hd__a21oi_1 U26980 ( .A1(n27789), .A2(n24082), .B1(n21227), .Y(
        n21228) );
  sky130_fd_sc_hd__nand2_1 U26981 ( .A(n21229), .B(n21228), .Y(n21231) );
  sky130_fd_sc_hd__a21oi_1 U26982 ( .A1(n22213), .A2(n21234), .B1(n21233), .Y(
        n21239) );
  sky130_fd_sc_hd__nand2_1 U26983 ( .A(n21237), .B(n21236), .Y(n21238) );
  sky130_fd_sc_hd__xor2_1 U26984 ( .A(n21239), .B(n21238), .X(n22817) );
  sky130_fd_sc_hd__a22oi_1 U26985 ( .A1(j202_soc_core_j22_cpu_ml_mach[3]), 
        .A2(n23041), .B1(n22817), .B2(n25679), .Y(n22438) );
  sky130_fd_sc_hd__nand3_1 U26986 ( .A(n24769), .B(n22439), .C(n22438), .Y(
        n21241) );
  sky130_fd_sc_hd__nand2_1 U26987 ( .A(n24769), .B(n27355), .Y(n21240) );
  sky130_fd_sc_hd__nand2_1 U26988 ( .A(n21242), .B(n22996), .Y(n21254) );
  sky130_fd_sc_hd__o22ai_1 U26989 ( .A1(n21244), .A2(n22983), .B1(n21243), 
        .B2(n22982), .Y(n21245) );
  sky130_fd_sc_hd__a21oi_1 U26990 ( .A1(n22986), .A2(
        j202_soc_core_j22_cpu_rf_gpr[3]), .B1(n21245), .Y(n21253) );
  sky130_fd_sc_hd__nand2_1 U26991 ( .A(n22988), .B(j202_soc_core_j22_cpu_pc[3]), .Y(n21247) );
  sky130_fd_sc_hd__nand2_1 U26992 ( .A(n22987), .B(
        j202_soc_core_j22_cpu_rf_gbr[3]), .Y(n21246) );
  sky130_fd_sc_hd__nand2_1 U26993 ( .A(n21247), .B(n21246), .Y(n21251) );
  sky130_fd_sc_hd__o22ai_1 U26994 ( .A1(n21249), .A2(n22897), .B1(n21248), 
        .B2(n22285), .Y(n21250) );
  sky130_fd_sc_hd__nor2_1 U26995 ( .A(n21251), .B(n21250), .Y(n21252) );
  sky130_fd_sc_hd__nand3_1 U26996 ( .A(n21254), .B(n21253), .C(n21252), .Y(
        n22440) );
  sky130_fd_sc_hd__nand2_1 U26997 ( .A(n22440), .B(n22862), .Y(n22825) );
  sky130_fd_sc_hd__nand2b_1 U26998 ( .A_N(n22825), .B(n24587), .Y(n21255) );
  sky130_fd_sc_hd__nand2_1 U26999 ( .A(n21256), .B(n21905), .Y(n21267) );
  sky130_fd_sc_hd__nor2_1 U27000 ( .A(n21260), .B(n21257), .Y(n21262) );
  sky130_fd_sc_hd__nand2_1 U27001 ( .A(n21762), .B(n21262), .Y(n21904) );
  sky130_fd_sc_hd__nand2_1 U27002 ( .A(n23030), .B(n21263), .Y(n21265) );
  sky130_fd_sc_hd__o21ai_1 U27003 ( .A1(n21260), .A2(n21259), .B1(n21258), .Y(
        n21261) );
  sky130_fd_sc_hd__a21oi_1 U27004 ( .A1(n21761), .A2(n21262), .B1(n21261), .Y(
        n21906) );
  sky130_fd_sc_hd__o21ai_2 U27005 ( .A1(n21265), .A2(n11866), .B1(n21264), .Y(
        n21266) );
  sky130_fd_sc_hd__xnor2_2 U27006 ( .A(n21267), .B(n21266), .Y(n23476) );
  sky130_fd_sc_hd__nand2_1 U27008 ( .A(n21270), .B(n21269), .Y(n21279) );
  sky130_fd_sc_hd__nand2_1 U27009 ( .A(n22958), .B(n21275), .Y(n21277) );
  sky130_fd_sc_hd__a21oi_1 U27010 ( .A1(n22965), .A2(n21275), .B1(n21274), .Y(
        n21276) );
  sky130_fd_sc_hd__o21ai_1 U27011 ( .A1(n21277), .A2(n22967), .B1(n21276), .Y(
        n21278) );
  sky130_fd_sc_hd__xnor2_1 U27012 ( .A(n21279), .B(n21278), .Y(n22525) );
  sky130_fd_sc_hd__nand2_1 U27013 ( .A(n22525), .B(n22940), .Y(n25907) );
  sky130_fd_sc_hd__nand2b_1 U27014 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[11]), .Y(n25906) );
  sky130_fd_sc_hd__nand2_1 U27015 ( .A(n23004), .B(n21280), .Y(n25910) );
  sky130_fd_sc_hd__nand4_1 U27016 ( .A(n25908), .B(n25907), .C(n25906), .D(
        n25910), .Y(n21282) );
  sky130_fd_sc_hd__nand2_1 U27017 ( .A(n25910), .B(n27052), .Y(n21281) );
  sky130_fd_sc_hd__nand2_1 U27018 ( .A(n21282), .B(n21281), .Y(n21289) );
  sky130_fd_sc_hd__a21oi_1 U27019 ( .A1(n21284), .A2(n13076), .B1(n21283), .Y(
        n21288) );
  sky130_fd_sc_hd__nand2_1 U27020 ( .A(n21286), .B(n21285), .Y(n21287) );
  sky130_fd_sc_hd__xor2_1 U27021 ( .A(n21288), .B(n21287), .X(n24341) );
  sky130_fd_sc_hd__nand2_1 U27022 ( .A(n24341), .B(n24461), .Y(n25928) );
  sky130_fd_sc_hd__nand2b_1 U27023 ( .A_N(n24463), .B(
        j202_soc_core_j22_cpu_ml_macl[11]), .Y(n25911) );
  sky130_fd_sc_hd__nand3_1 U27024 ( .A(n21289), .B(n25928), .C(n25911), .Y(
        n21290) );
  sky130_fd_sc_hd__nand2_1 U27025 ( .A(n21291), .B(n22996), .Y(n21303) );
  sky130_fd_sc_hd__o22ai_1 U27026 ( .A1(n21293), .A2(n22983), .B1(n21292), 
        .B2(n22982), .Y(n21294) );
  sky130_fd_sc_hd__a21oi_1 U27027 ( .A1(n22986), .A2(
        j202_soc_core_j22_cpu_rf_gpr[11]), .B1(n21294), .Y(n21302) );
  sky130_fd_sc_hd__nand2_1 U27028 ( .A(n22988), .B(
        j202_soc_core_j22_cpu_pc[11]), .Y(n21296) );
  sky130_fd_sc_hd__nand2_1 U27029 ( .A(n22987), .B(
        j202_soc_core_j22_cpu_rf_gbr[11]), .Y(n21295) );
  sky130_fd_sc_hd__nand2_1 U27030 ( .A(n21296), .B(n21295), .Y(n21300) );
  sky130_fd_sc_hd__o22ai_1 U27031 ( .A1(n21298), .A2(n22897), .B1(n21297), 
        .B2(n22285), .Y(n21299) );
  sky130_fd_sc_hd__nor2_1 U27032 ( .A(n21300), .B(n21299), .Y(n21301) );
  sky130_fd_sc_hd__nand3_1 U27033 ( .A(n21303), .B(n21302), .C(n21301), .Y(
        n22538) );
  sky130_fd_sc_hd__nand2_1 U27034 ( .A(n22538), .B(n24450), .Y(n21304) );
  sky130_fd_sc_hd__nand2_1 U27035 ( .A(j202_soc_core_qspi_wb_wdat[11]), .B(
        n29827), .Y(n29155) );
  sky130_fd_sc_hd__nor4_1 U27036 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[10]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[11]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[13]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[14]), .Y(n21308) );
  sky130_fd_sc_hd__nor4_1 U27037 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[15]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[17]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[19]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[18]), .Y(n21307) );
  sky130_fd_sc_hd__nor4_1 U27038 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[0]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[4]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[8]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[12]), .Y(n21306) );
  sky130_fd_sc_hd__nor4_1 U27039 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[16]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[20]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[24]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[28]), .Y(n21305) );
  sky130_fd_sc_hd__nand4_1 U27040 ( .A(n21308), .B(n21307), .C(n21306), .D(
        n21305), .Y(n21315) );
  sky130_fd_sc_hd__nor4_1 U27041 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[30]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[31]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[22]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[23]), .Y(n21311) );
  sky130_fd_sc_hd__nor4_1 U27042 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[1]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[21]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[25]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[29]), .Y(n21310) );
  sky130_fd_sc_hd__nand4_1 U27043 ( .A(n21311), .B(n21310), .C(n21309), .D(
        n26813), .Y(n21314) );
  sky130_fd_sc_hd__nor4_1 U27044 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[5]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[6]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[7]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[9]), .Y(n21312) );
  sky130_fd_sc_hd__or3b_2 U27045 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[3]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[2]), .C_N(n21312), .X(
        n21313) );
  sky130_fd_sc_hd__o31a_1 U27046 ( .A1(n21315), .A2(n21314), .A3(n21313), .B1(
        n29827), .X(n29580) );
  sky130_fd_sc_hd__nand2_1 U27047 ( .A(n21316), .B(n29482), .Y(n21317) );
  sky130_fd_sc_hd__nor2_1 U27049 ( .A(n13640), .B(n21660), .Y(n21319) );
  sky130_fd_sc_hd__xnor2_1 U27050 ( .A(n13576), .B(n21319), .Y(n25152) );
  sky130_fd_sc_hd__o22ai_1 U27051 ( .A1(n21320), .A2(n13365), .B1(n11191), 
        .B2(n11186), .Y(n21321) );
  sky130_fd_sc_hd__a21oi_1 U27052 ( .A1(n22701), .A2(n28495), .B1(n21321), .Y(
        n21324) );
  sky130_fd_sc_hd__nand2_1 U27053 ( .A(n21322), .B(n25152), .Y(n21323) );
  sky130_fd_sc_hd__o211a_2 U27054 ( .A1(n25944), .A2(n22745), .B1(n21324), 
        .C1(n21323), .X(n21333) );
  sky130_fd_sc_hd__nand2_1 U27055 ( .A(n21327), .B(n21326), .Y(n21331) );
  sky130_fd_sc_hd__a21oi_1 U27056 ( .A1(n21788), .A2(n21329), .B1(n21328), .Y(
        n21667) );
  sky130_fd_sc_hd__o21ai_0 U27057 ( .A1(n21663), .A2(n21667), .B1(n21664), .Y(
        n21330) );
  sky130_fd_sc_hd__xnor2_1 U27058 ( .A(n21331), .B(n21330), .Y(n24056) );
  sky130_fd_sc_hd__nand2_1 U27059 ( .A(n24056), .B(n17225), .Y(n21332) );
  sky130_fd_sc_hd__nand3_1 U27060 ( .A(n21334), .B(n21333), .C(n21332), .Y(
        n29555) );
  sky130_fd_sc_hd__nand2b_1 U27061 ( .A_N(n24074), .B(n22739), .Y(n21348) );
  sky130_fd_sc_hd__xnor2_1 U27062 ( .A(n14375), .B(n22698), .Y(n24075) );
  sky130_fd_sc_hd__o22ai_1 U27063 ( .A1(n24905), .A2(n13365), .B1(n26944), 
        .B2(n11186), .Y(n21337) );
  sky130_fd_sc_hd__a21oi_1 U27064 ( .A1(n22701), .A2(n28478), .B1(n21337), .Y(
        n21339) );
  sky130_fd_sc_hd__nand2_1 U27065 ( .A(n22702), .B(n28478), .Y(n21338) );
  sky130_fd_sc_hd__o211a_2 U27066 ( .A1(n24905), .A2(n22705), .B1(n21339), 
        .C1(n21338), .X(n21347) );
  sky130_fd_sc_hd__nand2_1 U27067 ( .A(n22691), .B(n22689), .Y(n21345) );
  sky130_fd_sc_hd__xnor2_1 U27069 ( .A(n21345), .B(n22692), .Y(n24873) );
  sky130_fd_sc_hd__nand2_1 U27070 ( .A(n24873), .B(n17225), .Y(n21346) );
  sky130_fd_sc_hd__nand3_1 U27071 ( .A(n21348), .B(n21347), .C(n21346), .Y(
        n29546) );
  sky130_fd_sc_hd__nand3_1 U27072 ( .A(n21423), .B(n21380), .C(n21536), .Y(
        n21611) );
  sky130_fd_sc_hd__nand2_1 U27073 ( .A(n21355), .B(n21521), .Y(n21350) );
  sky130_fd_sc_hd__nor2_1 U27074 ( .A(n21350), .B(n21349), .Y(n21392) );
  sky130_fd_sc_hd__nand4_1 U27075 ( .A(n21352), .B(n21392), .C(n21430), .D(
        n21607), .Y(n21357) );
  sky130_fd_sc_hd__nand2_1 U27076 ( .A(n21364), .B(n21415), .Y(n21531) );
  sky130_fd_sc_hd__nor2_1 U27077 ( .A(n21531), .B(n21353), .Y(n21537) );
  sky130_fd_sc_hd__and3_1 U27078 ( .A(n21362), .B(n21573), .C(n21354), .X(
        n21529) );
  sky130_fd_sc_hd__a31oi_1 U27079 ( .A1(n21537), .A2(n21355), .A3(n21529), 
        .B1(n21412), .Y(n21356) );
  sky130_fd_sc_hd__a21oi_1 U27080 ( .A1(n21357), .A2(n21603), .B1(n21356), .Y(
        n21371) );
  sky130_fd_sc_hd__nand3_1 U27081 ( .A(n21360), .B(n21359), .C(n21358), .Y(
        n21361) );
  sky130_fd_sc_hd__nand3_1 U27082 ( .A(n21584), .B(n21362), .C(n21361), .Y(
        n21363) );
  sky130_fd_sc_hd__nand2_1 U27083 ( .A(n21363), .B(n21610), .Y(n21369) );
  sky130_fd_sc_hd__nand4_1 U27084 ( .A(n21365), .B(n21384), .C(n21394), .D(
        n21364), .Y(n21367) );
  sky130_fd_sc_hd__o21ai_1 U27085 ( .A1(n21367), .A2(n21366), .B1(n21598), .Y(
        n21368) );
  sky130_fd_sc_hd__nand4_1 U27086 ( .A(n21371), .B(n21370), .C(n21369), .D(
        n21368), .Y(n21372) );
  sky130_fd_sc_hd__nand2_1 U27087 ( .A(n21372), .B(n21591), .Y(n21439) );
  sky130_fd_sc_hd__nand2_1 U27088 ( .A(n21373), .B(n21575), .Y(n21374) );
  sky130_fd_sc_hd__nand2_1 U27089 ( .A(n21374), .B(n21598), .Y(n21621) );
  sky130_fd_sc_hd__a21oi_1 U27090 ( .A1(n21392), .A2(n21385), .B1(n21412), .Y(
        n21378) );
  sky130_fd_sc_hd__a21oi_1 U27091 ( .A1(n21376), .A2(n21375), .B1(n21395), .Y(
        n21377) );
  sky130_fd_sc_hd__nor2_1 U27092 ( .A(n21378), .B(n21377), .Y(n21383) );
  sky130_fd_sc_hd__nand4_1 U27093 ( .A(n21380), .B(n21554), .C(n21606), .D(
        n21379), .Y(n21381) );
  sky130_fd_sc_hd__nand2_1 U27094 ( .A(n21381), .B(n21610), .Y(n21382) );
  sky130_fd_sc_hd__nand3_1 U27095 ( .A(n21621), .B(n21383), .C(n21382), .Y(
        n21407) );
  sky130_fd_sc_hd__nand4_1 U27096 ( .A(n21584), .B(n21386), .C(n21385), .D(
        n21384), .Y(n21387) );
  sky130_fd_sc_hd__nand2_1 U27097 ( .A(n21387), .B(n21617), .Y(n21404) );
  sky130_fd_sc_hd__nand3_1 U27098 ( .A(n21388), .B(n21583), .C(n21606), .Y(
        n21390) );
  sky130_fd_sc_hd__nor3_1 U27099 ( .A(n21556), .B(n21390), .C(n21389), .Y(
        n21391) );
  sky130_fd_sc_hd__a21oi_1 U27100 ( .A1(n21393), .A2(n13044), .B1(n21580), .Y(
        n21398) );
  sky130_fd_sc_hd__a31oi_1 U27101 ( .A1(n21551), .A2(n21529), .A3(n21396), 
        .B1(n21395), .Y(n21397) );
  sky130_fd_sc_hd__nor2_1 U27102 ( .A(n21398), .B(n21397), .Y(n21403) );
  sky130_fd_sc_hd__nand4_1 U27103 ( .A(n21399), .B(n21551), .C(n21567), .D(
        n21606), .Y(n21400) );
  sky130_fd_sc_hd__o21ai_1 U27104 ( .A1(n21401), .A2(n21400), .B1(n21598), .Y(
        n21402) );
  sky130_fd_sc_hd__nand3_1 U27105 ( .A(n21404), .B(n21403), .C(n21402), .Y(
        n21406) );
  sky130_fd_sc_hd__a22oi_1 U27106 ( .A1(n21407), .A2(n21624), .B1(n21406), 
        .B2(n21545), .Y(n21438) );
  sky130_fd_sc_hd__nand4_1 U27107 ( .A(n21410), .B(n21409), .C(n21584), .D(
        n21408), .Y(n21411) );
  sky130_fd_sc_hd__nand2_1 U27108 ( .A(n21411), .B(n21603), .Y(n21435) );
  sky130_fd_sc_hd__a21oi_1 U27109 ( .A1(n21416), .A2(n21413), .B1(n21412), .Y(
        n21549) );
  sky130_fd_sc_hd__and4_1 U27110 ( .A(n21416), .B(n21576), .C(n21415), .D(
        n21421), .X(n21417) );
  sky130_fd_sc_hd__a31oi_1 U27111 ( .A1(n21419), .A2(n21418), .A3(n21417), 
        .B1(n21580), .Y(n21420) );
  sky130_fd_sc_hd__nor2_1 U27112 ( .A(n21549), .B(n21420), .Y(n21434) );
  sky130_fd_sc_hd__nand2_1 U27113 ( .A(n21574), .B(n21421), .Y(n21422) );
  sky130_fd_sc_hd__nor2_1 U27114 ( .A(n21422), .B(n21609), .Y(n21424) );
  sky130_fd_sc_hd__nand3_1 U27115 ( .A(n21537), .B(n21424), .C(n21423), .Y(
        n21425) );
  sky130_fd_sc_hd__nand2_1 U27116 ( .A(n21425), .B(n21598), .Y(n21433) );
  sky130_fd_sc_hd__nor2_1 U27117 ( .A(n21427), .B(n21426), .Y(n21429) );
  sky130_fd_sc_hd__nand4_1 U27118 ( .A(n21430), .B(n21429), .C(n21428), .D(
        n21606), .Y(n21431) );
  sky130_fd_sc_hd__nand2_1 U27119 ( .A(n21617), .B(n21431), .Y(n21432) );
  sky130_fd_sc_hd__nand4_1 U27120 ( .A(n21435), .B(n21434), .C(n21433), .D(
        n21432), .Y(n21436) );
  sky130_fd_sc_hd__nand2_1 U27121 ( .A(n21436), .B(n21589), .Y(n21437) );
  sky130_fd_sc_hd__nand2b_1 U27122 ( .A_N(n21517), .B(
        j202_soc_core_bldc_core_00_pwm_period[4]), .Y(n21775) );
  sky130_fd_sc_hd__nand2_1 U27123 ( .A(n21504), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[12]), .Y(n21444) );
  sky130_fd_sc_hd__nand2_1 U27124 ( .A(n24720), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[20]), .Y(n21443) );
  sky130_fd_sc_hd__nand2_1 U27125 ( .A(n21505), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[4]), .Y(n21442) );
  sky130_fd_sc_hd__nand2_1 U27126 ( .A(n21506), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[28]), .Y(n21441) );
  sky130_fd_sc_hd__nand4_1 U27127 ( .A(n21444), .B(n21443), .C(n21442), .D(
        n21441), .Y(n21445) );
  sky130_fd_sc_hd__nand2_1 U27128 ( .A(n21513), .B(n21445), .Y(n21776) );
  sky130_fd_sc_hd__nand2_1 U27129 ( .A(n21446), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[100]), .Y(n21773) );
  sky130_fd_sc_hd__nand2_1 U27130 ( .A(n21776), .B(n21773), .Y(n21454) );
  sky130_fd_sc_hd__nand2_1 U27131 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[4]), .Y(n21453) );
  sky130_fd_sc_hd__nor2_1 U27132 ( .A(n21447), .B(n21512), .Y(n21452) );
  sky130_fd_sc_hd__nor2_1 U27133 ( .A(n21448), .B(n21452), .Y(n21829) );
  sky130_fd_sc_hd__nand2b_1 U27134 ( .A_N(n21515), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[36]), .Y(n21457) );
  sky130_fd_sc_hd__nor2_1 U27135 ( .A(n21650), .B(n21449), .Y(n21828) );
  sky130_fd_sc_hd__and4_1 U27136 ( .A(n21775), .B(n21450), .C(n21829), .D(
        n21828), .X(n21451) );
  sky130_fd_sc_hd__nand2_1 U27137 ( .A(n21772), .B(n21768), .Y(n21455) );
  sky130_fd_sc_hd__nand2_1 U27138 ( .A(n21457), .B(n21453), .Y(n21771) );
  sky130_fd_sc_hd__nor3_1 U27139 ( .A(n21455), .B(n21771), .C(n21454), .Y(
        n21456) );
  sky130_fd_sc_hd__nand3_1 U27140 ( .A(n21777), .B(n21456), .C(n21775), .Y(
        n21837) );
  sky130_fd_sc_hd__nand2_1 U27141 ( .A(n21484), .B(n21837), .Y(n21462) );
  sky130_fd_sc_hd__nand4_1 U27142 ( .A(n21829), .B(
        j202_soc_core_memory0_ram_dout0_sel[15]), .C(n21776), .D(n21457), .Y(
        n21458) );
  sky130_fd_sc_hd__nand2_1 U27143 ( .A(n21775), .B(n21773), .Y(n21827) );
  sky130_fd_sc_hd__nor2_1 U27144 ( .A(n21458), .B(n21827), .Y(n21459) );
  sky130_fd_sc_hd__nand2_1 U27145 ( .A(n21777), .B(n21459), .Y(n21460) );
  sky130_fd_sc_hd__a22oi_1 U27146 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__4_), .B1(n21916), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__4_), .Y(n21461) );
  sky130_fd_sc_hd__nand2_1 U27147 ( .A(j202_soc_core_memory0_ram_dout0[68]), 
        .B(n21642), .Y(n21465) );
  sky130_fd_sc_hd__nand2_1 U27148 ( .A(j202_soc_core_memory0_ram_dout0[452]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n21464) );
  sky130_fd_sc_hd__nand2_1 U27149 ( .A(j202_soc_core_memory0_ram_dout0[356]), 
        .B(n21495), .Y(n21463) );
  sky130_fd_sc_hd__nand3_1 U27150 ( .A(n21465), .B(n21464), .C(n21463), .Y(
        n21471) );
  sky130_fd_sc_hd__nand2_1 U27151 ( .A(j202_soc_core_memory0_ram_dout0[420]), 
        .B(n12156), .Y(n21469) );
  sky130_fd_sc_hd__nand2_1 U27152 ( .A(j202_soc_core_memory0_ram_dout0[324]), 
        .B(n21490), .Y(n21468) );
  sky130_fd_sc_hd__nand2_1 U27153 ( .A(j202_soc_core_memory0_ram_dout0[388]), 
        .B(n21496), .Y(n21467) );
  sky130_fd_sc_hd__nand2_1 U27154 ( .A(j202_soc_core_memory0_ram_dout0[292]), 
        .B(n21503), .Y(n21466) );
  sky130_fd_sc_hd__nand4_1 U27155 ( .A(n21469), .B(n21468), .C(n21467), .D(
        n21466), .Y(n21470) );
  sky130_fd_sc_hd__nor2_1 U27156 ( .A(n21471), .B(n21470), .Y(n21482) );
  sky130_fd_sc_hd__nand2_1 U27157 ( .A(j202_soc_core_memory0_ram_dout0[260]), 
        .B(n21634), .Y(n21475) );
  sky130_fd_sc_hd__nand2_1 U27158 ( .A(j202_soc_core_memory0_ram_dout0[228]), 
        .B(n21641), .Y(n21474) );
  sky130_fd_sc_hd__nand2_1 U27159 ( .A(j202_soc_core_memory0_ram_dout0[36]), 
        .B(n21633), .Y(n21473) );
  sky130_fd_sc_hd__nand2_1 U27160 ( .A(j202_soc_core_memory0_ram_dout0[196]), 
        .B(n21640), .Y(n21472) );
  sky130_fd_sc_hd__and4_1 U27161 ( .A(n21475), .B(n21474), .C(n21473), .D(
        n21472), .X(n21481) );
  sky130_fd_sc_hd__nand2_1 U27162 ( .A(j202_soc_core_memory0_ram_dout0[4]), 
        .B(n21639), .Y(n21479) );
  sky130_fd_sc_hd__nand2_1 U27163 ( .A(j202_soc_core_memory0_ram_dout0[132]), 
        .B(n21489), .Y(n21478) );
  sky130_fd_sc_hd__nand2_1 U27164 ( .A(j202_soc_core_memory0_ram_dout0[100]), 
        .B(n21488), .Y(n21477) );
  sky130_fd_sc_hd__nand2_1 U27165 ( .A(j202_soc_core_memory0_ram_dout0[164]), 
        .B(n21487), .Y(n21476) );
  sky130_fd_sc_hd__and4_1 U27166 ( .A(n21479), .B(n21478), .C(n21477), .D(
        n21476), .X(n21480) );
  sky130_fd_sc_hd__nand3_1 U27167 ( .A(n21836), .B(n21484), .C(n21483), .Y(
        n21485) );
  sky130_fd_sc_hd__nand2_1 U27168 ( .A(j202_soc_core_memory0_ram_dout0[165]), 
        .B(n21487), .Y(n21494) );
  sky130_fd_sc_hd__nand2_1 U27169 ( .A(j202_soc_core_memory0_ram_dout0[101]), 
        .B(n21488), .Y(n21493) );
  sky130_fd_sc_hd__nand2_1 U27170 ( .A(j202_soc_core_memory0_ram_dout0[133]), 
        .B(n21489), .Y(n21492) );
  sky130_fd_sc_hd__nand2_1 U27171 ( .A(j202_soc_core_memory0_ram_dout0[325]), 
        .B(n21490), .Y(n21491) );
  sky130_fd_sc_hd__nand4_1 U27172 ( .A(n21494), .B(n21493), .C(n21492), .D(
        n21491), .Y(n21502) );
  sky130_fd_sc_hd__nand2_1 U27173 ( .A(j202_soc_core_memory0_ram_dout0[357]), 
        .B(n21495), .Y(n21500) );
  sky130_fd_sc_hd__nand2_1 U27174 ( .A(j202_soc_core_memory0_ram_dout0[389]), 
        .B(n21496), .Y(n21499) );
  sky130_fd_sc_hd__nand2_1 U27175 ( .A(j202_soc_core_memory0_ram_dout0[453]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n21498) );
  sky130_fd_sc_hd__nand2_1 U27176 ( .A(j202_soc_core_memory0_ram_dout0[421]), 
        .B(n12156), .Y(n21497) );
  sky130_fd_sc_hd__nand4_1 U27177 ( .A(n21500), .B(n21499), .C(n21498), .D(
        n21497), .Y(n21501) );
  sky130_fd_sc_hd__nor2_1 U27178 ( .A(n21502), .B(n21501), .Y(n21649) );
  sky130_fd_sc_hd__nand2_1 U27179 ( .A(j202_soc_core_memory0_ram_dout0[293]), 
        .B(n21503), .Y(n21632) );
  sky130_fd_sc_hd__nand2_1 U27180 ( .A(n21504), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[13]), .Y(n21510) );
  sky130_fd_sc_hd__nand2_1 U27181 ( .A(n24720), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[21]), .Y(n21509) );
  sky130_fd_sc_hd__nand2_1 U27182 ( .A(n21505), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[5]), .Y(n21508) );
  sky130_fd_sc_hd__nand2_1 U27183 ( .A(n21506), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[29]), .Y(n21507) );
  sky130_fd_sc_hd__nand4_1 U27184 ( .A(n21510), .B(n21509), .C(n21508), .D(
        n21507), .Y(n21514) );
  sky130_fd_sc_hd__a2bb2oi_1 U27185 ( .B1(n21514), .B2(n21513), .A1_N(n21512), 
        .A2_N(n21511), .Y(n21654) );
  sky130_fd_sc_hd__nand2b_1 U27186 ( .A_N(n21515), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[37]), .Y(n21652) );
  sky130_fd_sc_hd__nand2_1 U27187 ( .A(n21516), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[5]), .Y(n21651) );
  sky130_fd_sc_hd__nand4_1 U27188 ( .A(n21654), .B(n21768), .C(n21652), .D(
        n21651), .Y(n21520) );
  sky130_fd_sc_hd__o22ai_1 U27189 ( .A1(n21519), .A2(n21518), .B1(n27409), 
        .B2(n21517), .Y(n21655) );
  sky130_fd_sc_hd__nor2_1 U27190 ( .A(n21520), .B(n21655), .Y(n21631) );
  sky130_fd_sc_hd__nor3_1 U27191 ( .A(n21524), .B(n21523), .C(n21522), .Y(
        n21544) );
  sky130_fd_sc_hd__nor2_1 U27192 ( .A(n21526), .B(n21525), .Y(n21528) );
  sky130_fd_sc_hd__nand4_1 U27193 ( .A(n21529), .B(n21528), .C(n21527), .D(
        n21593), .Y(n21535) );
  sky130_fd_sc_hd__nor3_1 U27194 ( .A(n21532), .B(n21531), .C(n21530), .Y(
        n21533) );
  sky130_fd_sc_hd__nand2_1 U27195 ( .A(n21584), .B(n21533), .Y(n21534) );
  sky130_fd_sc_hd__a22oi_1 U27196 ( .A1(n21603), .A2(n21535), .B1(n21534), 
        .B2(n21617), .Y(n21543) );
  sky130_fd_sc_hd__nand4_1 U27197 ( .A(n21539), .B(n21538), .C(n21537), .D(
        n21536), .Y(n21541) );
  sky130_fd_sc_hd__a21oi_1 U27198 ( .A1(n21598), .A2(n21541), .B1(n21540), .Y(
        n21542) );
  sky130_fd_sc_hd__o211ai_1 U27199 ( .A1(n21580), .A2(n21544), .B1(n21543), 
        .C1(n21542), .Y(n21546) );
  sky130_fd_sc_hd__nand2_1 U27200 ( .A(n21546), .B(n21545), .Y(n21628) );
  sky130_fd_sc_hd__nand2_1 U27201 ( .A(n21547), .B(n21576), .Y(n21548) );
  sky130_fd_sc_hd__nand2_1 U27202 ( .A(n21548), .B(n21598), .Y(n21561) );
  sky130_fd_sc_hd__nand3_1 U27203 ( .A(n21551), .B(n21550), .C(n21615), .Y(
        n21553) );
  sky130_fd_sc_hd__o21ai_1 U27204 ( .A1(n21553), .A2(n21552), .B1(n21610), .Y(
        n21559) );
  sky130_fd_sc_hd__nand4b_1 U27205 ( .A_N(n21556), .B(n21555), .C(n21575), .D(
        n21554), .Y(n21557) );
  sky130_fd_sc_hd__nand4_1 U27207 ( .A(n21561), .B(n21560), .C(n21559), .D(
        n21558), .Y(n21592) );
  sky130_fd_sc_hd__nand3b_1 U27208 ( .A_N(n21565), .B(n21564), .C(n21563), .Y(
        n21566) );
  sky130_fd_sc_hd__nand2_1 U27209 ( .A(n21566), .B(n21603), .Y(n21588) );
  sky130_fd_sc_hd__nand4_1 U27210 ( .A(n21569), .B(n21615), .C(n21568), .D(
        n21567), .Y(n21581) );
  sky130_fd_sc_hd__nand3_1 U27211 ( .A(n21572), .B(n21571), .C(n21570), .Y(
        n21578) );
  sky130_fd_sc_hd__nand4_1 U27212 ( .A(n21576), .B(n21575), .C(n21574), .D(
        n21573), .Y(n21577) );
  sky130_fd_sc_hd__nor2_1 U27213 ( .A(n21578), .B(n21577), .Y(n21579) );
  sky130_fd_sc_hd__a2bb2oi_1 U27214 ( .B1(n21598), .B2(n21581), .A1_N(n21580), 
        .A2_N(n21579), .Y(n21587) );
  sky130_fd_sc_hd__nand3_1 U27215 ( .A(n21584), .B(n21583), .C(n21582), .Y(
        n21585) );
  sky130_fd_sc_hd__nand2_1 U27216 ( .A(n21585), .B(n21617), .Y(n21586) );
  sky130_fd_sc_hd__nand3_1 U27217 ( .A(n21588), .B(n21587), .C(n21586), .Y(
        n21590) );
  sky130_fd_sc_hd__a22oi_1 U27218 ( .A1(n21592), .A2(n21591), .B1(n21590), 
        .B2(n21589), .Y(n21627) );
  sky130_fd_sc_hd__o21a_1 U27219 ( .A1(n21595), .A2(n21594), .B1(n21593), .X(
        n21596) );
  sky130_fd_sc_hd__nand3_1 U27220 ( .A(n21597), .B(n21596), .C(n21606), .Y(
        n21604) );
  sky130_fd_sc_hd__o31a_1 U27221 ( .A1(n21601), .A2(n21600), .A3(n21599), .B1(
        n21598), .X(n21602) );
  sky130_fd_sc_hd__a21oi_1 U27222 ( .A1(n21604), .A2(n21603), .B1(n21602), .Y(
        n21623) );
  sky130_fd_sc_hd__nand4b_1 U27223 ( .A_N(n21609), .B(n21608), .C(n21607), .D(
        n21606), .Y(n21612) );
  sky130_fd_sc_hd__o21ai_1 U27224 ( .A1(n21612), .A2(n21611), .B1(n21610), .Y(
        n21622) );
  sky130_fd_sc_hd__nand3_1 U27225 ( .A(n21616), .B(n21615), .C(n21614), .Y(
        n21619) );
  sky130_fd_sc_hd__nand4_1 U27227 ( .A(n21623), .B(n21622), .C(n21621), .D(
        n21620), .Y(n21625) );
  sky130_fd_sc_hd__nand2_1 U27228 ( .A(n21625), .B(n21624), .Y(n21626) );
  sky130_fd_sc_hd__nand3_1 U27229 ( .A(n21628), .B(n21627), .C(n21626), .Y(
        n21630) );
  sky130_fd_sc_hd__nand2_1 U27230 ( .A(n21630), .B(n21629), .Y(n21657) );
  sky130_fd_sc_hd__nand3_1 U27231 ( .A(n21632), .B(n21631), .C(n21657), .Y(
        n21638) );
  sky130_fd_sc_hd__nand2_1 U27232 ( .A(j202_soc_core_memory0_ram_dout0[37]), 
        .B(n21633), .Y(n21636) );
  sky130_fd_sc_hd__nand2_1 U27233 ( .A(j202_soc_core_memory0_ram_dout0[261]), 
        .B(n21634), .Y(n21635) );
  sky130_fd_sc_hd__nand2_1 U27234 ( .A(n21636), .B(n21635), .Y(n21637) );
  sky130_fd_sc_hd__nor2_1 U27235 ( .A(n21638), .B(n21637), .Y(n21648) );
  sky130_fd_sc_hd__nand2_1 U27236 ( .A(j202_soc_core_memory0_ram_dout0[5]), 
        .B(n21639), .Y(n21646) );
  sky130_fd_sc_hd__nand2_1 U27237 ( .A(j202_soc_core_memory0_ram_dout0[197]), 
        .B(n21640), .Y(n21645) );
  sky130_fd_sc_hd__nand2_1 U27238 ( .A(j202_soc_core_memory0_ram_dout0[229]), 
        .B(n21641), .Y(n21644) );
  sky130_fd_sc_hd__nand2_1 U27239 ( .A(j202_soc_core_memory0_ram_dout0[69]), 
        .B(n21642), .Y(n21643) );
  sky130_fd_sc_hd__nand2_1 U27240 ( .A(j202_soc_core_memory0_ram_dout0[485]), 
        .B(n21650), .Y(n21659) );
  sky130_fd_sc_hd__nand4_1 U27241 ( .A(n21654), .B(n21653), .C(n21652), .D(
        n21651), .Y(n21656) );
  sky130_fd_sc_hd__nor2_1 U27242 ( .A(n21656), .B(n21655), .Y(n21658) );
  sky130_fd_sc_hd__nand3_1 U27243 ( .A(n21659), .B(n21658), .C(n21657), .Y(
        n21918) );
  sky130_fd_sc_hd__nand2_1 U27244 ( .A(n21920), .B(n21918), .Y(n22233) );
  sky130_fd_sc_hd__nand2b_1 U27245 ( .A_N(n22233), .B(n22739), .Y(n21670) );
  sky130_fd_sc_hd__xor2_1 U27246 ( .A(n21660), .B(n13640), .X(n24803) );
  sky130_fd_sc_hd__o22a_1 U27247 ( .A1(n26421), .A2(n22743), .B1(n11189), .B2(
        n11186), .X(n21661) );
  sky130_fd_sc_hd__o21ai_0 U27248 ( .A1(n26421), .A2(n22745), .B1(n21661), .Y(
        n21662) );
  sky130_fd_sc_hd__a21oi_1 U27249 ( .A1(n24803), .A2(n22747), .B1(n21662), .Y(
        n21669) );
  sky130_fd_sc_hd__nand2_1 U27250 ( .A(n21665), .B(n21664), .Y(n21666) );
  sky130_fd_sc_hd__xor2_1 U27251 ( .A(n21667), .B(n21666), .X(n24044) );
  sky130_fd_sc_hd__nand2_1 U27252 ( .A(n24044), .B(n17225), .Y(n21668) );
  sky130_fd_sc_hd__nand3_1 U27253 ( .A(n21670), .B(n21669), .C(n21668), .Y(
        n29554) );
  sky130_fd_sc_hd__o22ai_1 U27254 ( .A1(n21672), .A2(n22983), .B1(n21671), 
        .B2(n22982), .Y(n21673) );
  sky130_fd_sc_hd__a21oi_1 U27255 ( .A1(n22990), .A2(
        j202_soc_core_j22_cpu_rf_vbr[0]), .B1(n21673), .Y(n21678) );
  sky130_fd_sc_hd__a22oi_1 U27256 ( .A1(n22988), .A2(
        j202_soc_core_j22_cpu_pc[0]), .B1(j202_soc_core_j22_cpu_rf_gbr[0]), 
        .B2(n22987), .Y(n21677) );
  sky130_fd_sc_hd__o22a_1 U27257 ( .A1(n21674), .A2(n22897), .B1(n21717), .B2(
        n22894), .X(n21676) );
  sky130_fd_sc_hd__nand2_1 U27258 ( .A(n22986), .B(
        j202_soc_core_j22_cpu_rf_gpr[0]), .Y(n21675) );
  sky130_fd_sc_hd__nand4_1 U27259 ( .A(n21678), .B(n21677), .C(n21676), .D(
        n21675), .Y(n21679) );
  sky130_fd_sc_hd__a21oi_1 U27260 ( .A1(n21680), .A2(n22996), .B1(n21679), .Y(
        n22780) );
  sky130_fd_sc_hd__nand2_1 U27261 ( .A(n21685), .B(n21972), .Y(n21686) );
  sky130_fd_sc_hd__xor2_1 U27262 ( .A(n21973), .B(n21686), .X(n22766) );
  sky130_fd_sc_hd__o22ai_1 U27263 ( .A1(n24456), .A2(n18188), .B1(n21687), 
        .B2(n28045), .Y(n21688) );
  sky130_fd_sc_hd__a21oi_1 U27264 ( .A1(n22766), .A2(n25679), .B1(n21688), .Y(
        n22416) );
  sky130_fd_sc_hd__nand2_1 U27265 ( .A(n21691), .B(n22230), .Y(n21692) );
  sky130_fd_sc_hd__nand2_1 U27266 ( .A(n21693), .B(n22114), .Y(n21695) );
  sky130_fd_sc_hd__nand2b_1 U27267 ( .A_N(n26048), .B(n21696), .Y(n26922) );
  sky130_fd_sc_hd__o21ai_1 U27268 ( .A1(n11123), .A2(n26377), .B1(n26922), .Y(
        n21697) );
  sky130_fd_sc_hd__nand2_1 U27269 ( .A(n12284), .B(n21697), .Y(n21728) );
  sky130_fd_sc_hd__nand2_1 U27270 ( .A(n21700), .B(n21699), .Y(n21701) );
  sky130_fd_sc_hd__xnor2_1 U27271 ( .A(n21702), .B(n21701), .Y(n24078) );
  sky130_fd_sc_hd__nand2_1 U27272 ( .A(n24353), .B(n24461), .Y(n22421) );
  sky130_fd_sc_hd__nand2_1 U27273 ( .A(n25996), .B(n21707), .Y(n26935) );
  sky130_fd_sc_hd__nand2_1 U27274 ( .A(n28541), .B(n26377), .Y(n26293) );
  sky130_fd_sc_hd__nor2_1 U27275 ( .A(n21708), .B(n24463), .Y(n22420) );
  sky130_fd_sc_hd__nand4_1 U27276 ( .A(n21709), .B(n26270), .C(
        j202_soc_core_j22_cpu_exuop_EXU_[5]), .D(
        j202_soc_core_j22_cpu_rfuo_sr__t_), .Y(n21710) );
  sky130_fd_sc_hd__nand2b_1 U27277 ( .A_N(n26001), .B(
        j202_soc_core_j22_cpu_ml_bufa[0]), .Y(n22418) );
  sky130_fd_sc_hd__o22ai_1 U27278 ( .A1(n26048), .A2(n21710), .B1(n26926), 
        .B2(n22418), .Y(n21711) );
  sky130_fd_sc_hd__a21oi_1 U27279 ( .A1(n22420), .A2(n26414), .B1(n21711), .Y(
        n21713) );
  sky130_fd_sc_hd__nand2_1 U27280 ( .A(n25685), .B(n26945), .Y(n21712) );
  sky130_fd_sc_hd__o211ai_1 U27281 ( .A1(n26293), .A2(n26939), .B1(n21713), 
        .C1(n21712), .Y(n21714) );
  sky130_fd_sc_hd__a21oi_1 U27282 ( .A1(n27111), .A2(n26935), .B1(n21714), .Y(
        n21722) );
  sky130_fd_sc_hd__nand2_1 U27283 ( .A(n11188), .B(n26265), .Y(n26242) );
  sky130_fd_sc_hd__nand3_1 U27284 ( .A(n26242), .B(n27806), .C(n26293), .Y(
        n21715) );
  sky130_fd_sc_hd__o21ai_0 U27285 ( .A1(n26284), .A2(n27803), .B1(n21715), .Y(
        n21716) );
  sky130_fd_sc_hd__a21oi_1 U27286 ( .A1(n27810), .A2(n26929), .B1(n21716), .Y(
        n21720) );
  sky130_fd_sc_hd__mux2i_1 U27287 ( .A0(n21717), .A1(n28429), .S(n26421), .Y(
        n21718) );
  sky130_fd_sc_hd__nand3_1 U27288 ( .A(n21718), .B(n25999), .C(n28521), .Y(
        n21719) );
  sky130_fd_sc_hd__nand4_1 U27289 ( .A(n21722), .B(n21721), .C(n21720), .D(
        n21719), .Y(n21724) );
  sky130_fd_sc_hd__mux2i_1 U27290 ( .A0(n22251), .A1(n27793), .S(n26265), .Y(
        n21723) );
  sky130_fd_sc_hd__nor2_1 U27291 ( .A(n21724), .B(n21723), .Y(n21725) );
  sky130_fd_sc_hd__a21oi_1 U27293 ( .A1(n27789), .A2(n24078), .B1(n21726), .Y(
        n21727) );
  sky130_fd_sc_hd__nand2_1 U27294 ( .A(n21731), .B(n22883), .Y(n21732) );
  sky130_fd_sc_hd__xor2_1 U27295 ( .A(n22884), .B(n21732), .X(n26966) );
  sky130_fd_sc_hd__nand2_1 U27296 ( .A(n26966), .B(n24461), .Y(n24950) );
  sky130_fd_sc_hd__nor2_1 U27297 ( .A(n21733), .B(n24463), .Y(n24933) );
  sky130_fd_sc_hd__o22ai_1 U27298 ( .A1(n21735), .A2(n22983), .B1(n22982), 
        .B2(n21734), .Y(n21736) );
  sky130_fd_sc_hd__a21oi_1 U27299 ( .A1(n22990), .A2(
        j202_soc_core_j22_cpu_rf_vbr[8]), .B1(n21736), .Y(n21742) );
  sky130_fd_sc_hd__a22oi_1 U27300 ( .A1(n22988), .A2(
        j202_soc_core_j22_cpu_pc[8]), .B1(n22987), .B2(
        j202_soc_core_j22_cpu_rf_gbr[8]), .Y(n21741) );
  sky130_fd_sc_hd__o22a_1 U27301 ( .A1(n22897), .A2(n21738), .B1(n21737), .B2(
        n22894), .X(n21740) );
  sky130_fd_sc_hd__nand2_1 U27302 ( .A(n22986), .B(
        j202_soc_core_j22_cpu_rf_gpr[8]), .Y(n21739) );
  sky130_fd_sc_hd__nand4_1 U27303 ( .A(n21742), .B(n21741), .C(n21740), .D(
        n21739), .Y(n21743) );
  sky130_fd_sc_hd__a21oi_1 U27304 ( .A1(n21744), .A2(n22996), .B1(n21743), .Y(
        n22735) );
  sky130_fd_sc_hd__nor2_1 U27305 ( .A(n21745), .B(n28045), .Y(n24921) );
  sky130_fd_sc_hd__nand2_1 U27306 ( .A(n27717), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .Y(n21746) );
  sky130_fd_sc_hd__a2bb2oi_1 U27307 ( .B1(n23044), .B2(n24921), .A1_N(n21747), 
        .A2_N(n21746), .Y(n21748) );
  sky130_fd_sc_hd__a21oi_1 U27309 ( .A1(n27717), .A2(n24933), .B1(n21750), .Y(
        n21751) );
  sky130_fd_sc_hd__o21ai_1 U27310 ( .A1(n24467), .A2(n24950), .B1(n21751), .Y(
        n21759) );
  sky130_fd_sc_hd__nand2_1 U27311 ( .A(n22875), .B(n22873), .Y(n21757) );
  sky130_fd_sc_hd__o21ai_1 U27312 ( .A1(n21755), .A2(n22967), .B1(n21754), .Y(
        n21756) );
  sky130_fd_sc_hd__xnor2_1 U27313 ( .A(n21757), .B(n21756), .Y(n22731) );
  sky130_fd_sc_hd__nand2_1 U27314 ( .A(n22731), .B(n22940), .Y(n24922) );
  sky130_fd_sc_hd__nor2_1 U27315 ( .A(n22309), .B(n24922), .Y(n21758) );
  sky130_fd_sc_hd__nor2_1 U27316 ( .A(n21759), .B(n21758), .Y(n21767) );
  sky130_fd_sc_hd__nand2_1 U27317 ( .A(n23030), .B(n21762), .Y(n21764) );
  sky130_fd_sc_hd__nand2_1 U27319 ( .A(n24153), .B(n24452), .Y(n24924) );
  sky130_fd_sc_hd__nand2_1 U27320 ( .A(n21765), .B(n23044), .Y(n21766) );
  sky130_fd_sc_hd__nor2_1 U27321 ( .A(n21768), .B(
        j202_soc_core_memory0_ram_dout0[484]), .Y(n21769) );
  sky130_fd_sc_hd__nor2_1 U27322 ( .A(n21816), .B(n21769), .Y(n21770) );
  sky130_fd_sc_hd__nand4_1 U27324 ( .A(n21775), .B(n21774), .C(n21773), .D(
        n21772), .Y(n21778) );
  sky130_fd_sc_hd__nand2_1 U27325 ( .A(n21777), .B(n21776), .Y(n21831) );
  sky130_fd_sc_hd__nor2_1 U27326 ( .A(n21778), .B(n21831), .Y(n21779) );
  sky130_fd_sc_hd__nand2_1 U27327 ( .A(n21780), .B(n21779), .Y(n29443) );
  sky130_fd_sc_hd__nand2_1 U27328 ( .A(n29443), .B(n22739), .Y(n21796) );
  sky130_fd_sc_hd__nand2_1 U27329 ( .A(n21781), .B(j202_soc_core_j22_cpu_pc[3]), .Y(n21782) );
  sky130_fd_sc_hd__xor2_1 U27330 ( .A(n21782), .B(n13750), .X(n27507) );
  sky130_fd_sc_hd__o22a_1 U27331 ( .A1(n26240), .A2(n22743), .B1(n27365), .B2(
        n11186), .X(n21783) );
  sky130_fd_sc_hd__o21ai_1 U27332 ( .A1(n26240), .A2(n22745), .B1(n21783), .Y(
        n21784) );
  sky130_fd_sc_hd__a21oi_1 U27333 ( .A1(n27507), .A2(n22747), .B1(n21784), .Y(
        n21795) );
  sky130_fd_sc_hd__a21oi_1 U27334 ( .A1(n21788), .A2(n21787), .B1(n21786), .Y(
        n21793) );
  sky130_fd_sc_hd__nand2_1 U27335 ( .A(n21791), .B(n21790), .Y(n21792) );
  sky130_fd_sc_hd__xor2_1 U27336 ( .A(n21793), .B(n21792), .X(n24035) );
  sky130_fd_sc_hd__nand2_1 U27337 ( .A(n24035), .B(n17225), .Y(n21794) );
  sky130_fd_sc_hd__nand3_1 U27338 ( .A(n21796), .B(n21795), .C(n21794), .Y(
        n29545) );
  sky130_fd_sc_hd__nand2_1 U27339 ( .A(n21797), .B(n22996), .Y(n21809) );
  sky130_fd_sc_hd__a22oi_1 U27340 ( .A1(n22988), .A2(
        j202_soc_core_j22_cpu_pc[4]), .B1(j202_soc_core_j22_cpu_rf_gbr[4]), 
        .B2(n22987), .Y(n21808) );
  sky130_fd_sc_hd__nand2_1 U27341 ( .A(n22986), .B(
        j202_soc_core_j22_cpu_rf_gpr[4]), .Y(n21807) );
  sky130_fd_sc_hd__o22ai_1 U27342 ( .A1(n21799), .A2(n22983), .B1(n21798), 
        .B2(n22982), .Y(n21805) );
  sky130_fd_sc_hd__nor2_1 U27343 ( .A(n21800), .B(n22285), .Y(n21804) );
  sky130_fd_sc_hd__o22ai_1 U27344 ( .A1(n21802), .A2(n22897), .B1(n21801), 
        .B2(n22894), .Y(n21803) );
  sky130_fd_sc_hd__nor3_1 U27345 ( .A(n21805), .B(n21804), .C(n21803), .Y(
        n21806) );
  sky130_fd_sc_hd__nand4_1 U27346 ( .A(n21809), .B(n21808), .C(n21807), .D(
        n21806), .Y(n22453) );
  sky130_fd_sc_hd__nand2_1 U27347 ( .A(n22453), .B(n22862), .Y(n22330) );
  sky130_fd_sc_hd__nand2_1 U27349 ( .A(n21810), .B(n22197), .Y(n21814) );
  sky130_fd_sc_hd__nand2_1 U27350 ( .A(n22195), .B(n22193), .Y(n21812) );
  sky130_fd_sc_hd__a21oi_1 U27351 ( .A1(n22202), .A2(n22193), .B1(n22196), .Y(
        n21811) );
  sky130_fd_sc_hd__o21ai_2 U27352 ( .A1(n21812), .A2(n11866), .B1(n21811), .Y(
        n21813) );
  sky130_fd_sc_hd__xnor2_2 U27353 ( .A(n21814), .B(n21813), .Y(n27362) );
  sky130_fd_sc_hd__nand2_1 U27354 ( .A(n27362), .B(n24452), .Y(n22450) );
  sky130_fd_sc_hd__nand4_1 U27355 ( .A(n21818), .B(n21817), .C(n21816), .D(
        n21815), .Y(n21820) );
  sky130_fd_sc_hd__nor3_1 U27356 ( .A(n21821), .B(n21820), .C(n21819), .Y(
        n21823) );
  sky130_fd_sc_hd__nor3_1 U27357 ( .A(n21823), .B(n11149), .C(n21822), .Y(
        n21824) );
  sky130_fd_sc_hd__o21ai_1 U27358 ( .A1(n21826), .A2(n21825), .B1(n21824), .Y(
        n21840) );
  sky130_fd_sc_hd__nand3_1 U27359 ( .A(n21830), .B(n21829), .C(n21828), .Y(
        n21832) );
  sky130_fd_sc_hd__nor2_1 U27361 ( .A(n21834), .B(n21833), .Y(n21835) );
  sky130_fd_sc_hd__o21ai_1 U27362 ( .A1(n21837), .A2(n21836), .B1(n21835), .Y(
        n21839) );
  sky130_fd_sc_hd__nand2b_1 U27363 ( .A_N(n26240), .B(n22136), .Y(n26299) );
  sky130_fd_sc_hd__nand2_1 U27364 ( .A(n26299), .B(n27806), .Y(n21847) );
  sky130_fd_sc_hd__and2_0 U27365 ( .A(n21847), .B(n26919), .X(n21842) );
  sky130_fd_sc_hd__o21ai_1 U27366 ( .A1(n26411), .A2(n22136), .B1(n27787), .Y(
        n21863) );
  sky130_fd_sc_hd__nand2_1 U27367 ( .A(n21844), .B(n21843), .Y(n21845) );
  sky130_fd_sc_hd__xnor2_1 U27368 ( .A(n21846), .B(n21845), .Y(n22317) );
  sky130_fd_sc_hd__nand2_1 U27369 ( .A(n22317), .B(n24461), .Y(n22456) );
  sky130_fd_sc_hd__nand2_1 U27370 ( .A(n22251), .B(n21847), .Y(n21848) );
  sky130_fd_sc_hd__mux2i_1 U27371 ( .A0(n21848), .A1(n26034), .S(n26240), .Y(
        n21859) );
  sky130_fd_sc_hd__nor2_1 U27372 ( .A(n21849), .B(n24463), .Y(n22451) );
  sky130_fd_sc_hd__nand2_1 U27373 ( .A(n23004), .B(
        j202_soc_core_j22_cpu_ml_bufa[4]), .Y(n22454) );
  sky130_fd_sc_hd__o2bb2ai_1 U27374 ( .B1(n22454), .B2(n26926), .A1_N(n26003), 
        .A2_N(n26331), .Y(n21850) );
  sky130_fd_sc_hd__a21oi_1 U27375 ( .A1(n22451), .A2(n26414), .B1(n21850), .Y(
        n21851) );
  sky130_fd_sc_hd__o21ai_0 U27376 ( .A1(n26939), .A2(n26299), .B1(n21851), .Y(
        n21852) );
  sky130_fd_sc_hd__a21oi_1 U27377 ( .A1(n27810), .A2(n26378), .B1(n21852), .Y(
        n21853) );
  sky130_fd_sc_hd__o21a_1 U27378 ( .A1(n28506), .A2(n26932), .B1(n21853), .X(
        n21858) );
  sky130_fd_sc_hd__o22ai_1 U27379 ( .A1(n11189), .A2(n27803), .B1(n26318), 
        .B2(n26943), .Y(n21854) );
  sky130_fd_sc_hd__a21oi_1 U27380 ( .A1(n27808), .A2(n26929), .B1(n21854), .Y(
        n21857) );
  sky130_fd_sc_hd__o22ai_1 U27381 ( .A1(n11190), .A2(n27795), .B1(n27383), 
        .B2(n25996), .Y(n21855) );
  sky130_fd_sc_hd__a21oi_1 U27382 ( .A1(n21949), .A2(n28460), .B1(n21855), .Y(
        n21856) );
  sky130_fd_sc_hd__nand4_1 U27383 ( .A(n21859), .B(n21858), .C(n21857), .D(
        n21856), .Y(n21860) );
  sky130_fd_sc_hd__a21oi_1 U27384 ( .A1(n24035), .A2(n27789), .B1(n21860), .Y(
        n21861) );
  sky130_fd_sc_hd__inv_1 U27386 ( .A(n21866), .Y(n22210) );
  sky130_fd_sc_hd__a21oi_1 U27387 ( .A1(n22213), .A2(n22207), .B1(n21867), .Y(
        n21870) );
  sky130_fd_sc_hd__nand2_1 U27388 ( .A(n21868), .B(n22209), .Y(n21869) );
  sky130_fd_sc_hd__xor2_1 U27389 ( .A(n21870), .B(n21869), .X(n22320) );
  sky130_fd_sc_hd__nand2_1 U27390 ( .A(n22320), .B(n25679), .Y(n27357) );
  sky130_fd_sc_hd__nand2b_1 U27391 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[4]), .Y(n27356) );
  sky130_fd_sc_hd__nand2_1 U27392 ( .A(n27357), .B(n27356), .Y(n22448) );
  sky130_fd_sc_hd__nor2_1 U27393 ( .A(n22448), .B(n27359), .Y(n21871) );
  sky130_fd_sc_hd__nand3_2 U27394 ( .A(n21874), .B(n21873), .C(n22266), .Y(
        n22316) );
  sky130_fd_sc_hd__nand2_1 U27395 ( .A(n21875), .B(n22960), .Y(n21879) );
  sky130_fd_sc_hd__nand2_1 U27396 ( .A(n22958), .B(n12331), .Y(n21877) );
  sky130_fd_sc_hd__a21oi_1 U27397 ( .A1(n22965), .A2(n12331), .B1(n11426), .Y(
        n21876) );
  sky130_fd_sc_hd__o21ai_1 U27398 ( .A1(n21877), .A2(n22967), .B1(n21876), .Y(
        n21878) );
  sky130_fd_sc_hd__xnor2_1 U27399 ( .A(n21879), .B(n21878), .Y(n24765) );
  sky130_fd_sc_hd__nand2_1 U27400 ( .A(n24765), .B(n25679), .Y(n25991) );
  sky130_fd_sc_hd__inv_1 U27401 ( .A(n21880), .Y(n22975) );
  sky130_fd_sc_hd__nand2_1 U27402 ( .A(n21881), .B(n22974), .Y(n21882) );
  sky130_fd_sc_hd__xor2_1 U27403 ( .A(n22975), .B(n21882), .X(n24349) );
  sky130_fd_sc_hd__nand2_1 U27404 ( .A(n24349), .B(n24461), .Y(n26018) );
  sky130_fd_sc_hd__nor2_1 U27405 ( .A(n21883), .B(n24463), .Y(n26004) );
  sky130_fd_sc_hd__o22ai_1 U27406 ( .A1(n21885), .A2(n22983), .B1(n22982), 
        .B2(n21884), .Y(n21886) );
  sky130_fd_sc_hd__a21oi_1 U27407 ( .A1(n22986), .A2(
        j202_soc_core_j22_cpu_rf_gpr[12]), .B1(n21886), .Y(n21890) );
  sky130_fd_sc_hd__a22oi_1 U27408 ( .A1(n22988), .A2(
        j202_soc_core_j22_cpu_pc[12]), .B1(n22987), .B2(
        j202_soc_core_j22_cpu_rf_gbr[12]), .Y(n21889) );
  sky130_fd_sc_hd__nand2_1 U27409 ( .A(n22989), .B(
        j202_soc_core_j22_cpu_rf_tmp[12]), .Y(n21888) );
  sky130_fd_sc_hd__nand2_1 U27410 ( .A(n22990), .B(n12042), .Y(n21887) );
  sky130_fd_sc_hd__nand4_1 U27411 ( .A(n21890), .B(n21889), .C(n21888), .D(
        n21887), .Y(n21891) );
  sky130_fd_sc_hd__a21o_1 U27412 ( .A1(n21892), .A2(n22996), .B1(n21891), .X(
        n22650) );
  sky130_fd_sc_hd__nand2_1 U27413 ( .A(n22650), .B(n24450), .Y(n21896) );
  sky130_fd_sc_hd__nand3_1 U27414 ( .A(n23004), .B(n27717), .C(
        j202_soc_core_j22_cpu_ml_bufa[12]), .Y(n21895) );
  sky130_fd_sc_hd__nor2_1 U27415 ( .A(n21893), .B(n28045), .Y(n25990) );
  sky130_fd_sc_hd__nand2_1 U27416 ( .A(n25990), .B(n23044), .Y(n21894) );
  sky130_fd_sc_hd__nand3_1 U27417 ( .A(n21896), .B(n21895), .C(n21894), .Y(
        n21897) );
  sky130_fd_sc_hd__a21oi_1 U27418 ( .A1(n26004), .A2(n27717), .B1(n21897), .Y(
        n21898) );
  sky130_fd_sc_hd__o21ai_0 U27419 ( .A1(n24467), .A2(n26018), .B1(n21898), .Y(
        n21899) );
  sky130_fd_sc_hd__nand2_1 U27420 ( .A(n21903), .B(n21902), .Y(n21913) );
  sky130_fd_sc_hd__nor2_1 U27421 ( .A(n21907), .B(n21904), .Y(n21909) );
  sky130_fd_sc_hd__nand2_1 U27422 ( .A(n23030), .B(n21909), .Y(n21911) );
  sky130_fd_sc_hd__o21a_1 U27423 ( .A1(n21907), .A2(n21906), .B1(n21905), .X(
        n21908) );
  sky130_fd_sc_hd__xnor2_1 U27424 ( .A(n21913), .B(n21912), .Y(n23470) );
  sky130_fd_sc_hd__nor2_1 U27425 ( .A(n22309), .B(n25993), .Y(n21914) );
  sky130_fd_sc_hd__nor2_1 U27426 ( .A(n21901), .B(n21914), .Y(n21915) );
  sky130_fd_sc_hd__inv_1 U27427 ( .A(n22233), .Y(n29445) );
  sky130_fd_sc_hd__a22oi_1 U27428 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__5_), .B1(n21916), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__5_), .Y(n21923) );
  sky130_fd_sc_hd__nand2_1 U27429 ( .A(n12292), .B(n21917), .Y(n21922) );
  sky130_fd_sc_hd__nand2_1 U27432 ( .A(n29444), .B(n22739), .Y(n21931) );
  sky130_fd_sc_hd__nand2_1 U27433 ( .A(n24078), .B(n17225), .Y(n21928) );
  sky130_fd_sc_hd__nand2_1 U27434 ( .A(n21924), .B(n28541), .Y(n21927) );
  sky130_fd_sc_hd__nand2_1 U27435 ( .A(n21925), .B(n26377), .Y(n21926) );
  sky130_fd_sc_hd__and3_1 U27436 ( .A(n21928), .B(n21927), .C(n21926), .X(
        n21930) );
  sky130_fd_sc_hd__nand2_1 U27437 ( .A(n22747), .B(j202_soc_core_j22_cpu_pc[0]), .Y(n21929) );
  sky130_fd_sc_hd__nand3_1 U27438 ( .A(n21931), .B(n21930), .C(n21929), .Y(
        n29565) );
  sky130_fd_sc_hd__a21oi_1 U27439 ( .A1(n12354), .A2(n27791), .B1(n27790), .Y(
        n21935) );
  sky130_fd_sc_hd__o21ai_1 U27440 ( .A1(n26411), .A2(n26375), .B1(n27787), .Y(
        n21937) );
  sky130_fd_sc_hd__nand2_1 U27441 ( .A(n28528), .B(n21937), .Y(n21956) );
  sky130_fd_sc_hd__nand2_1 U27442 ( .A(n21939), .B(n21938), .Y(n21940) );
  sky130_fd_sc_hd__xnor2_1 U27443 ( .A(n11143), .B(n21940), .Y(n24320) );
  sky130_fd_sc_hd__nand2_1 U27444 ( .A(n24320), .B(n24461), .Y(n21996) );
  sky130_fd_sc_hd__xnor2_1 U27445 ( .A(n12354), .B(n26375), .Y(n26250) );
  sky130_fd_sc_hd__o22a_1 U27446 ( .A1(n26944), .A2(n26943), .B1(n25872), .B2(
        n26250), .X(n21941) );
  sky130_fd_sc_hd__nor2_1 U27448 ( .A(n21942), .B(n24463), .Y(n21983) );
  sky130_fd_sc_hd__nand2b_1 U27449 ( .A_N(n26001), .B(n21943), .Y(n21994) );
  sky130_fd_sc_hd__o2bb2ai_1 U27450 ( .B1(n26926), .B2(n21994), .A1_N(n26003), 
        .A2_N(n26051), .Y(n21944) );
  sky130_fd_sc_hd__a21oi_1 U27451 ( .A1(n21983), .A2(n26414), .B1(n21944), .Y(
        n21946) );
  sky130_fd_sc_hd__nand2_1 U27452 ( .A(n27810), .B(n26334), .Y(n21945) );
  sky130_fd_sc_hd__o211ai_1 U27453 ( .A1(n26320), .A2(n25996), .B1(n21946), 
        .C1(n21945), .Y(n21948) );
  sky130_fd_sc_hd__o22ai_1 U27454 ( .A1(n11188), .A2(n27795), .B1(n27147), 
        .B2(n27803), .Y(n21947) );
  sky130_fd_sc_hd__a211o_1 U27455 ( .A1(n21949), .A2(n28478), .B1(n21948), 
        .C1(n21947), .X(n21951) );
  sky130_fd_sc_hd__mux2i_1 U27456 ( .A0(n22251), .A1(n27793), .S(n11144), .Y(
        n21950) );
  sky130_fd_sc_hd__nor3_1 U27457 ( .A(n21952), .B(n21951), .C(n21950), .Y(
        n21953) );
  sky130_fd_sc_hd__o21ai_1 U27458 ( .A1(n26926), .A2(n21996), .B1(n21953), .Y(
        n21954) );
  sky130_fd_sc_hd__a21oi_1 U27459 ( .A1(n27789), .A2(n24052), .B1(n21954), .Y(
        n21955) );
  sky130_fd_sc_hd__nand2_1 U27460 ( .A(n21959), .B(n21958), .Y(n21968) );
  sky130_fd_sc_hd__nand2_1 U27461 ( .A(n10972), .B(n21963), .Y(n21966) );
  sky130_fd_sc_hd__a21oi_1 U27462 ( .A1(n21963), .A2(n11349), .B1(n21962), .Y(
        n21965) );
  sky130_fd_sc_hd__o21ai_2 U27463 ( .A1(n21966), .A2(n12349), .B1(n21965), .Y(
        n21967) );
  sky130_fd_sc_hd__xnor2_2 U27464 ( .A(n21968), .B(n21967), .Y(n23479) );
  sky130_fd_sc_hd__nand2_2 U27465 ( .A(n23479), .B(n24452), .Y(n21982) );
  sky130_fd_sc_hd__nand2_1 U27466 ( .A(n21971), .B(n21970), .Y(n21976) );
  sky130_fd_sc_hd__o21ai_1 U27467 ( .A1(n21974), .A2(n21973), .B1(n21972), .Y(
        n21975) );
  sky130_fd_sc_hd__xnor2_1 U27468 ( .A(n21976), .B(n21975), .Y(n22848) );
  sky130_fd_sc_hd__nand2_1 U27469 ( .A(n22848), .B(n25679), .Y(n21979) );
  sky130_fd_sc_hd__nand2b_1 U27470 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[1]), .Y(n21978) );
  sky130_fd_sc_hd__nand2_1 U27471 ( .A(n28056), .B(n21943), .Y(n21977) );
  sky130_fd_sc_hd__and3_1 U27472 ( .A(n21979), .B(n21978), .C(n21977), .X(
        n21981) );
  sky130_fd_sc_hd__nand2_1 U27473 ( .A(n21982), .B(n21981), .Y(n24794) );
  sky130_fd_sc_hd__nand2_1 U27474 ( .A(n24794), .B(n23044), .Y(n22001) );
  sky130_fd_sc_hd__o22ai_1 U27475 ( .A1(n21985), .A2(n22983), .B1(n21984), 
        .B2(n22982), .Y(n21986) );
  sky130_fd_sc_hd__a21oi_1 U27476 ( .A1(n22990), .A2(
        j202_soc_core_j22_cpu_rf_vbr[1]), .B1(n21986), .Y(n21991) );
  sky130_fd_sc_hd__a22oi_1 U27477 ( .A1(n22988), .A2(
        j202_soc_core_j22_cpu_pc[1]), .B1(n22987), .B2(
        j202_soc_core_j22_cpu_rf_gbr[1]), .Y(n21990) );
  sky130_fd_sc_hd__o22a_1 U27478 ( .A1(n21987), .A2(n22897), .B1(n24668), .B2(
        n22894), .X(n21989) );
  sky130_fd_sc_hd__nand2_1 U27479 ( .A(n22986), .B(
        j202_soc_core_j22_cpu_rf_gpr[1]), .Y(n21988) );
  sky130_fd_sc_hd__nand4_1 U27480 ( .A(n21991), .B(n21990), .C(n21989), .D(
        n21988), .Y(n21992) );
  sky130_fd_sc_hd__nand2_1 U27481 ( .A(n22866), .B(n22452), .Y(n21997) );
  sky130_fd_sc_hd__nand4_1 U27482 ( .A(n21996), .B(n21995), .C(n21994), .D(
        n21997), .Y(n21999) );
  sky130_fd_sc_hd__nand2_1 U27483 ( .A(n21997), .B(n24467), .Y(n21998) );
  sky130_fd_sc_hd__nand2_1 U27484 ( .A(n21999), .B(n21998), .Y(n22000) );
  sky130_fd_sc_hd__nand3_1 U27485 ( .A(n22868), .B(n22001), .C(n22000), .Y(
        n29507) );
  sky130_fd_sc_hd__inv_2 U27486 ( .A(n22002), .Y(n25148) );
  sky130_fd_sc_hd__nand2_1 U27488 ( .A(n24127), .B(n11140), .Y(n27898) );
  sky130_fd_sc_hd__nand2_1 U27489 ( .A(n23391), .B(n28417), .Y(n22012) );
  sky130_fd_sc_hd__nor2_1 U27490 ( .A(j202_soc_core_j22_cpu_opst[2]), .B(
        j202_soc_core_j22_cpu_opst[1]), .Y(n23414) );
  sky130_fd_sc_hd__nand2_1 U27491 ( .A(n22011), .B(n23414), .Y(n24702) );
  sky130_fd_sc_hd__nand2_1 U27492 ( .A(n22012), .B(n28394), .Y(n29597) );
  sky130_fd_sc_hd__nor2_1 U27493 ( .A(n22013), .B(n24613), .Y(n29542) );
  sky130_fd_sc_hd__nor2_1 U27494 ( .A(n22014), .B(n11145), .Y(n22020) );
  sky130_fd_sc_hd__nor2_1 U27495 ( .A(n22015), .B(n11145), .Y(n22486) );
  sky130_fd_sc_hd__nor2_1 U27496 ( .A(n22020), .B(n22016), .Y(n22714) );
  sky130_fd_sc_hd__nand2_1 U27497 ( .A(n22016), .B(n22020), .Y(n22712) );
  sky130_fd_sc_hd__nand2_1 U27498 ( .A(n22483), .B(n22712), .Y(n22077) );
  sky130_fd_sc_hd__nor2_1 U27499 ( .A(n22018), .B(n11145), .Y(n22062) );
  sky130_fd_sc_hd__nor2_1 U27500 ( .A(n22019), .B(n11145), .Y(n22064) );
  sky130_fd_sc_hd__nor2_1 U27501 ( .A(n22062), .B(n22063), .Y(n22178) );
  sky130_fd_sc_hd__nand2_1 U27502 ( .A(n11187), .B(n22173), .Y(n22069) );
  sky130_fd_sc_hd__nor2_1 U27503 ( .A(n22021), .B(n11145), .Y(n22056) );
  sky130_fd_sc_hd__nor2_1 U27504 ( .A(n22022), .B(n11145), .Y(n22058) );
  sky130_fd_sc_hd__nor2_1 U27505 ( .A(n22056), .B(n22057), .Y(n22338) );
  sky130_fd_sc_hd__nand2_1 U27506 ( .A(n22801), .B(n22333), .Y(n22175) );
  sky130_fd_sc_hd__xnor2_1 U27507 ( .A(n22024), .B(n22023), .Y(n22025) );
  sky130_fd_sc_hd__o21ai_1 U27508 ( .A1(n22027), .A2(n11145), .B1(n22026), .Y(
        n22036) );
  sky130_fd_sc_hd__fa_1 U27509 ( .A(n22033), .B(n22032), .CIN(n22031), .COUT(
        n22041), .SUM(n18918) );
  sky130_fd_sc_hd__nor2_1 U27510 ( .A(n22040), .B(n22041), .Y(n22833) );
  sky130_fd_sc_hd__nor2_1 U27511 ( .A(n22034), .B(n11145), .Y(n22037) );
  sky130_fd_sc_hd__fa_1 U27512 ( .A(n22038), .B(n22036), .CIN(n22035), .COUT(
        n22043), .SUM(n22040) );
  sky130_fd_sc_hd__nand2_1 U27513 ( .A(n22782), .B(n22829), .Y(n22047) );
  sky130_fd_sc_hd__nand2_1 U27514 ( .A(n12098), .B(n22050), .Y(n22052) );
  sky130_fd_sc_hd__nor2_1 U27515 ( .A(n22052), .B(n22593), .Y(n22352) );
  sky130_fd_sc_hd__fa_1 U27516 ( .A(n22039), .B(n22038), .CIN(n22037), .COUT(
        n22054), .SUM(n22042) );
  sky130_fd_sc_hd__nand2_1 U27517 ( .A(n22352), .B(n22351), .Y(n22334) );
  sky130_fd_sc_hd__nor2_1 U27518 ( .A(n22071), .B(n22334), .Y(n22542) );
  sky130_fd_sc_hd__nand2_1 U27519 ( .A(n22017), .B(n22542), .Y(n22711) );
  sky130_fd_sc_hd__nand2_1 U27520 ( .A(n23030), .B(n22073), .Y(n22075) );
  sky130_fd_sc_hd__nand2_1 U27521 ( .A(n22041), .B(n22040), .Y(n22831) );
  sky130_fd_sc_hd__nand2_1 U27522 ( .A(n22043), .B(n22042), .Y(n22828) );
  sky130_fd_sc_hd__a21oi_1 U27523 ( .A1(n22045), .A2(n22829), .B1(n22044), .Y(
        n22046) );
  sky130_fd_sc_hd__a21oi_1 U27525 ( .A1(n22050), .A2(n22049), .B1(n22048), .Y(
        n22051) );
  sky130_fd_sc_hd__o21ai_1 U27526 ( .A1(n23019), .A2(n22052), .B1(n22051), .Y(
        n22353) );
  sky130_fd_sc_hd__nand2_1 U27527 ( .A(n22054), .B(n22053), .Y(n22350) );
  sky130_fd_sc_hd__a21oi_2 U27528 ( .A1(n22353), .A2(n22351), .B1(n22055), .Y(
        n22335) );
  sky130_fd_sc_hd__nand2_1 U27529 ( .A(n22057), .B(n22056), .Y(n22800) );
  sky130_fd_sc_hd__nand2_1 U27530 ( .A(n22059), .B(n22058), .Y(n22332) );
  sky130_fd_sc_hd__a21oi_1 U27531 ( .A1(n22333), .A2(n22061), .B1(n22060), .Y(
        n22174) );
  sky130_fd_sc_hd__nand2_1 U27532 ( .A(n22063), .B(n22062), .Y(n22268) );
  sky130_fd_sc_hd__nand2_1 U27533 ( .A(n22065), .B(n22064), .Y(n22172) );
  sky130_fd_sc_hd__a21oi_1 U27534 ( .A1(n22173), .A2(n22067), .B1(n22066), .Y(
        n22068) );
  sky130_fd_sc_hd__o21a_1 U27535 ( .A1(n22069), .A2(n22174), .B1(n22068), .X(
        n22070) );
  sky130_fd_sc_hd__a21oi_1 U27536 ( .A1(n22789), .A2(n22542), .B1(n22543), .Y(
        n22713) );
  sky130_fd_sc_hd__a21oi_1 U27537 ( .A1(n23036), .A2(n22073), .B1(n22072), .Y(
        n22074) );
  sky130_fd_sc_hd__xnor2_1 U27538 ( .A(n22077), .B(n22076), .Y(n22078) );
  sky130_fd_sc_hd__nand2_1 U27539 ( .A(n22078), .B(n24452), .Y(n25220) );
  sky130_fd_sc_hd__nand2_1 U27540 ( .A(n27717), .B(n27052), .Y(n23018) );
  sky130_fd_sc_hd__nand2_1 U27541 ( .A(n27768), .B(n22087), .Y(n22080) );
  sky130_fd_sc_hd__nand2_1 U27542 ( .A(n24324), .B(n22979), .Y(n22079) );
  sky130_fd_sc_hd__o211ai_1 U27543 ( .A1(n22980), .A2(n22081), .B1(n22080), 
        .C1(n22079), .Y(n22082) );
  sky130_fd_sc_hd__a21oi_1 U27544 ( .A1(n22083), .A2(n24764), .B1(n22082), .Y(
        n25224) );
  sky130_fd_sc_hd__nand2b_1 U27545 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[23]), .Y(n25219) );
  sky130_fd_sc_hd__nand2_1 U27546 ( .A(n22988), .B(n22089), .Y(n23000) );
  sky130_fd_sc_hd__nor2_1 U27547 ( .A(n24304), .B(n22983), .Y(n23006) );
  sky130_fd_sc_hd__nand2_1 U27548 ( .A(n23006), .B(
        j202_soc_core_j22_cpu_rf_pr[23]), .Y(n22086) );
  sky130_fd_sc_hd__nor2_1 U27549 ( .A(n24304), .B(n22084), .Y(n23003) );
  sky130_fd_sc_hd__nand2_1 U27550 ( .A(n23003), .B(
        j202_soc_core_j22_cpu_rf_gpr[23]), .Y(n22085) );
  sky130_fd_sc_hd__o211a_2 U27551 ( .A1(n23000), .A2(n15260), .B1(n22086), 
        .C1(n22085), .X(n22097) );
  sky130_fd_sc_hd__nor2_1 U27552 ( .A(j202_soc_core_j22_cpu_regop_Rs__1_), .B(
        n24304), .Y(n23010) );
  sky130_fd_sc_hd__nor2_1 U27553 ( .A(n24304), .B(n22982), .Y(n23005) );
  sky130_fd_sc_hd__nand2_1 U27554 ( .A(n28056), .B(n22087), .Y(n25218) );
  sky130_fd_sc_hd__nor2_1 U27555 ( .A(n27052), .B(n25218), .Y(n22088) );
  sky130_fd_sc_hd__a22oi_1 U27556 ( .A1(n23005), .A2(
        j202_soc_core_j22_cpu_rf_gpr[502]), .B1(n22088), .B2(n27717), .Y(
        n22093) );
  sky130_fd_sc_hd__nor2_1 U27557 ( .A(n24304), .B(n22285), .Y(n23008) );
  sky130_fd_sc_hd__nand2_1 U27558 ( .A(n23008), .B(
        j202_soc_core_j22_cpu_rf_vbr[23]), .Y(n22092) );
  sky130_fd_sc_hd__nand2_1 U27559 ( .A(n22987), .B(n22089), .Y(n22998) );
  sky130_fd_sc_hd__nand2_1 U27560 ( .A(n22722), .B(
        j202_soc_core_j22_cpu_rf_gbr[23]), .Y(n22091) );
  sky130_fd_sc_hd__nor2_1 U27561 ( .A(n24304), .B(n22897), .Y(n23009) );
  sky130_fd_sc_hd__nand2_1 U27562 ( .A(n23009), .B(
        j202_soc_core_j22_cpu_rf_tmp[23]), .Y(n22090) );
  sky130_fd_sc_hd__nand4_1 U27563 ( .A(n22093), .B(n22092), .C(n22091), .D(
        n22090), .Y(n22094) );
  sky130_fd_sc_hd__a21oi_1 U27564 ( .A1(n23010), .A2(n22095), .B1(n22094), .Y(
        n22096) );
  sky130_fd_sc_hd__o211ai_1 U27565 ( .A1(n22309), .A2(n25219), .B1(n22097), 
        .C1(n22096), .Y(n22098) );
  sky130_fd_sc_hd__a21oi_1 U27566 ( .A1(n22862), .A2(n22384), .B1(n22098), .Y(
        n22099) );
  sky130_fd_sc_hd__a21oi_1 U27568 ( .A1(n22101), .A2(n23044), .B1(n22100), .Y(
        n22104) );
  sky130_fd_sc_hd__nand2_1 U27569 ( .A(n23478), .B(n25679), .Y(n25222) );
  sky130_fd_sc_hd__nand2_1 U27570 ( .A(n22102), .B(n23044), .Y(n22103) );
  sky130_fd_sc_hd__nand3_1 U27571 ( .A(n12206), .B(n22104), .C(n22103), .Y(
        n29511) );
  sky130_fd_sc_hd__inv_2 U27572 ( .A(n23036), .Y(n22106) );
  sky130_fd_sc_hd__nand2_1 U27573 ( .A(n22110), .B(n22109), .Y(n22111) );
  sky130_fd_sc_hd__xor2_1 U27574 ( .A(n22967), .B(n22111), .X(n22150) );
  sky130_fd_sc_hd__o22ai_1 U27575 ( .A1(n24456), .A2(n17449), .B1(n22112), 
        .B2(n28045), .Y(n22113) );
  sky130_fd_sc_hd__a21oi_1 U27576 ( .A1(n22150), .A2(n22940), .B1(n22113), .Y(
        n22393) );
  sky130_fd_sc_hd__nand2_1 U27578 ( .A(n11191), .B(n22117), .Y(n22118) );
  sky130_fd_sc_hd__nand2_1 U27579 ( .A(n25642), .B(n23532), .Y(n22120) );
  sky130_fd_sc_hd__nand2_1 U27580 ( .A(n26378), .B(n27785), .Y(n22122) );
  sky130_fd_sc_hd__nand2_1 U27581 ( .A(n22122), .B(n27787), .Y(n22123) );
  sky130_fd_sc_hd__nand2_1 U27582 ( .A(n12039), .B(n22123), .Y(n22145) );
  sky130_fd_sc_hd__nand2_1 U27583 ( .A(n22126), .B(n22125), .Y(n22127) );
  sky130_fd_sc_hd__xnor2_1 U27584 ( .A(n22124), .B(n22127), .Y(n24308) );
  sky130_fd_sc_hd__nand2_1 U27585 ( .A(n24308), .B(n24461), .Y(n22398) );
  sky130_fd_sc_hd__nand2_1 U27586 ( .A(n24056), .B(n27789), .Y(n22141) );
  sky130_fd_sc_hd__o22ai_1 U27587 ( .A1(n11189), .A2(n27795), .B1(n26319), 
        .B2(n26943), .Y(n22130) );
  sky130_fd_sc_hd__o22ai_1 U27588 ( .A1(n27616), .A2(n27803), .B1(n26324), 
        .B2(n25996), .Y(n22129) );
  sky130_fd_sc_hd__o22ai_1 U27589 ( .A1(n25973), .A2(n26936), .B1(n26277), 
        .B2(n26932), .Y(n22128) );
  sky130_fd_sc_hd__nor3_1 U27590 ( .A(n22130), .B(n22129), .C(n22128), .Y(
        n22140) );
  sky130_fd_sc_hd__nand2_1 U27591 ( .A(n26378), .B(n28495), .Y(n26306) );
  sky130_fd_sc_hd__nor2_1 U27592 ( .A(n22131), .B(n24463), .Y(n22395) );
  sky130_fd_sc_hd__nand2_1 U27593 ( .A(n22395), .B(n26414), .Y(n22134) );
  sky130_fd_sc_hd__nand2b_1 U27594 ( .A_N(n26001), .B(
        j202_soc_core_j22_cpu_ml_bufa[6]), .Y(n22397) );
  sky130_fd_sc_hd__o22ai_1 U27595 ( .A1(n26926), .A2(n22397), .B1(n27793), 
        .B2(n28495), .Y(n22132) );
  sky130_fd_sc_hd__a21oi_1 U27596 ( .A1(n25109), .A2(n26378), .B1(n22132), .Y(
        n22133) );
  sky130_fd_sc_hd__o211ai_1 U27597 ( .A1(n26306), .A2(n26939), .B1(n22134), 
        .C1(n22133), .Y(n22135) );
  sky130_fd_sc_hd__a21oi_1 U27598 ( .A1(n26247), .A2(n27806), .B1(n22135), .Y(
        n22138) );
  sky130_fd_sc_hd__a22oi_1 U27599 ( .A1(n27810), .A2(n26945), .B1(n27808), 
        .B2(n22136), .Y(n22137) );
  sky130_fd_sc_hd__o211a_2 U27600 ( .A1(n25944), .A2(n22251), .B1(n22138), 
        .C1(n22137), .X(n22139) );
  sky130_fd_sc_hd__nand3_1 U27601 ( .A(n22141), .B(n22140), .C(n22139), .Y(
        n22142) );
  sky130_fd_sc_hd__a21oi_1 U27602 ( .A1(n22143), .A2(n26414), .B1(n22142), .Y(
        n22144) );
  sky130_fd_sc_hd__nand2_1 U27603 ( .A(n22145), .B(n22144), .Y(n22146) );
  sky130_fd_sc_hd__o2bb2ai_1 U27604 ( .B1(n22980), .B2(n22148), .A1_N(n24308), 
        .A2_N(n22979), .Y(n22149) );
  sky130_fd_sc_hd__a21oi_1 U27605 ( .A1(n22150), .A2(n24764), .B1(n22149), .Y(
        n25371) );
  sky130_fd_sc_hd__o22ai_1 U27606 ( .A1(n22152), .A2(n22983), .B1(n22982), 
        .B2(n22151), .Y(n22153) );
  sky130_fd_sc_hd__a21oi_1 U27607 ( .A1(n22990), .A2(
        j202_soc_core_j22_cpu_rf_vbr[6]), .B1(n22153), .Y(n22159) );
  sky130_fd_sc_hd__a22oi_1 U27608 ( .A1(n22988), .A2(
        j202_soc_core_j22_cpu_pc[6]), .B1(n22987), .B2(
        j202_soc_core_j22_cpu_rf_gbr[6]), .Y(n22158) );
  sky130_fd_sc_hd__o22a_1 U27609 ( .A1(n22897), .A2(n22155), .B1(n22154), .B2(
        n22894), .X(n22157) );
  sky130_fd_sc_hd__nand2_1 U27610 ( .A(n22986), .B(
        j202_soc_core_j22_cpu_rf_gpr[6]), .Y(n22156) );
  sky130_fd_sc_hd__nand4_1 U27611 ( .A(n22159), .B(n22158), .C(n22157), .D(
        n22156), .Y(n22160) );
  sky130_fd_sc_hd__a21o_1 U27612 ( .A1(n22161), .A2(n22996), .B1(n22160), .X(
        n22558) );
  sky130_fd_sc_hd__nand2_1 U27613 ( .A(n23003), .B(
        j202_soc_core_j22_cpu_rf_gpr[22]), .Y(n22163) );
  sky130_fd_sc_hd__nand2_1 U27614 ( .A(n22722), .B(
        j202_soc_core_j22_cpu_rf_gbr[22]), .Y(n22162) );
  sky130_fd_sc_hd__o211ai_1 U27615 ( .A1(n22164), .A2(n23000), .B1(n22163), 
        .C1(n22162), .Y(n22168) );
  sky130_fd_sc_hd__nand2_1 U27616 ( .A(n23004), .B(n25627), .Y(n25358) );
  sky130_fd_sc_hd__a22oi_1 U27617 ( .A1(n23006), .A2(
        j202_soc_core_j22_cpu_rf_pr[22]), .B1(n23005), .B2(
        j202_soc_core_j22_cpu_rf_gpr[501]), .Y(n22166) );
  sky130_fd_sc_hd__a22oi_1 U27618 ( .A1(n23009), .A2(
        j202_soc_core_j22_cpu_rf_tmp[22]), .B1(n23008), .B2(
        j202_soc_core_j22_cpu_rf_vbr[22]), .Y(n22165) );
  sky130_fd_sc_hd__o211ai_1 U27619 ( .A1(n24467), .A2(n25358), .B1(n22166), 
        .C1(n22165), .Y(n22167) );
  sky130_fd_sc_hd__a211o_1 U27620 ( .A1(n22169), .A2(n23010), .B1(n22168), 
        .C1(n22167), .X(n22170) );
  sky130_fd_sc_hd__a21oi_1 U27621 ( .A1(n22558), .A2(n22862), .B1(n22170), .Y(
        n22171) );
  sky130_fd_sc_hd__o21a_1 U27622 ( .A1(n23018), .A2(n25371), .B1(n22171), .X(
        n22189) );
  sky130_fd_sc_hd__nand2_1 U27623 ( .A(n23477), .B(n25679), .Y(n22187) );
  sky130_fd_sc_hd__nand2_1 U27624 ( .A(n22173), .B(n22172), .Y(n22184) );
  sky130_fd_sc_hd__nor2_1 U27625 ( .A(n22175), .B(n22334), .Y(n22177) );
  sky130_fd_sc_hd__nand2_1 U27626 ( .A(n22017), .B(n22177), .Y(n22269) );
  sky130_fd_sc_hd__nor2_1 U27627 ( .A(n22178), .B(n22269), .Y(n22180) );
  sky130_fd_sc_hd__nand2_1 U27628 ( .A(n23030), .B(n22180), .Y(n22182) );
  sky130_fd_sc_hd__a21oi_1 U27629 ( .A1(n23036), .A2(n22180), .B1(n22179), .Y(
        n22181) );
  sky130_fd_sc_hd__xnor2_1 U27630 ( .A(n22184), .B(n22183), .Y(n22185) );
  sky130_fd_sc_hd__nand2_1 U27631 ( .A(n25626), .B(n23044), .Y(n22188) );
  sky130_fd_sc_hd__nand3_1 U27632 ( .A(n22560), .B(n22189), .C(n22188), .Y(
        n29510) );
  sky130_fd_sc_hd__nand2_1 U27633 ( .A(n22192), .B(n22191), .Y(n22206) );
  sky130_fd_sc_hd__nor2_1 U27634 ( .A(n22199), .B(n22194), .Y(n22201) );
  sky130_fd_sc_hd__nand2_1 U27635 ( .A(n22201), .B(n22195), .Y(n22204) );
  sky130_fd_sc_hd__a21oi_1 U27637 ( .A1(n22202), .A2(n22201), .B1(n22200), .Y(
        n22203) );
  sky130_fd_sc_hd__o21ai_2 U27638 ( .A1(n22204), .A2(n11866), .B1(n22203), .Y(
        n22205) );
  sky130_fd_sc_hd__xnor2_2 U27639 ( .A(n22206), .B(n22205), .Y(n23469) );
  sky130_fd_sc_hd__nor2_1 U27640 ( .A(n12435), .B(n22208), .Y(n22214) );
  sky130_fd_sc_hd__nand2_1 U27643 ( .A(n22217), .B(n22216), .Y(n22218) );
  sky130_fd_sc_hd__xor2_1 U27644 ( .A(n22219), .B(n22218), .X(n22281) );
  sky130_fd_sc_hd__a22oi_1 U27645 ( .A1(j202_soc_core_j22_cpu_ml_mach[5]), 
        .A2(n23041), .B1(n22281), .B2(n25679), .Y(n22404) );
  sky130_fd_sc_hd__nand3_1 U27646 ( .A(n29445), .B(n22232), .C(n22260), .Y(
        n22220) );
  sky130_fd_sc_hd__nor2_1 U27647 ( .A(n11149), .B(n22222), .Y(n22223) );
  sky130_fd_sc_hd__buf_2 U27649 ( .A(n12292), .X(n23516) );
  sky130_fd_sc_hd__nand2_1 U27650 ( .A(n23516), .B(n22227), .Y(n22228) );
  sky130_fd_sc_hd__nand2_1 U27651 ( .A(n22259), .B(n26922), .Y(n22237) );
  sky130_fd_sc_hd__nand2b_1 U27652 ( .A_N(n22233), .B(n22232), .Y(n22234) );
  sky130_fd_sc_hd__nand2_1 U27653 ( .A(n22237), .B(n28501), .Y(n22263) );
  sky130_fd_sc_hd__nand2_1 U27654 ( .A(n22240), .B(n22239), .Y(n22242) );
  sky130_fd_sc_hd__xor2_1 U27655 ( .A(n22242), .B(n22241), .X(n24364) );
  sky130_fd_sc_hd__nand2_1 U27656 ( .A(n24364), .B(n24461), .Y(n22407) );
  sky130_fd_sc_hd__o22ai_1 U27657 ( .A1(n27365), .A2(n27795), .B1(n26321), 
        .B2(n26943), .Y(n22243) );
  sky130_fd_sc_hd__a21oi_1 U27658 ( .A1(n26329), .A2(n26935), .B1(n22243), .Y(
        n22250) );
  sky130_fd_sc_hd__o22a_1 U27659 ( .A1(n25451), .A2(n26936), .B1(n26281), .B2(
        n26932), .X(n22249) );
  sky130_fd_sc_hd__xnor2_1 U27660 ( .A(n22260), .B(n26421), .Y(n26245) );
  sky130_fd_sc_hd__a22oi_1 U27661 ( .A1(n27808), .A2(n26334), .B1(n26245), 
        .B2(n27806), .Y(n22248) );
  sky130_fd_sc_hd__nand2_1 U27662 ( .A(n23004), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .Y(n22244) );
  sky130_fd_sc_hd__o21a_1 U27663 ( .A1(n22245), .A2(n24463), .B1(n22244), .X(
        n22406) );
  sky130_fd_sc_hd__o22ai_1 U27664 ( .A1(n22406), .A2(n26926), .B1(n11191), 
        .B2(n27803), .Y(n22246) );
  sky130_fd_sc_hd__a21oi_1 U27665 ( .A1(n27810), .A2(n24879), .B1(n22246), .Y(
        n22247) );
  sky130_fd_sc_hd__nand4_1 U27666 ( .A(n22250), .B(n22249), .C(n22248), .D(
        n22247), .Y(n22253) );
  sky130_fd_sc_hd__mux2i_1 U27667 ( .A0(n22251), .A1(n27793), .S(n26421), .Y(
        n22252) );
  sky130_fd_sc_hd__nor2_1 U27668 ( .A(n22253), .B(n22252), .Y(n22254) );
  sky130_fd_sc_hd__a21oi_1 U27670 ( .A1(n22257), .A2(n27785), .B1(n22256), .Y(
        n22262) );
  sky130_fd_sc_hd__o21a_1 U27671 ( .A1(n26421), .A2(n26939), .B1(n26919), .X(
        n22258) );
  sky130_fd_sc_hd__nand2_1 U27672 ( .A(n11187), .B(n22268), .Y(n22275) );
  sky130_fd_sc_hd__nand2_1 U27673 ( .A(n23030), .B(n22271), .Y(n22273) );
  sky130_fd_sc_hd__a21oi_1 U27674 ( .A1(n23036), .A2(n22271), .B1(n22270), .Y(
        n22272) );
  sky130_fd_sc_hd__xnor2_1 U27675 ( .A(n22275), .B(n22274), .Y(n22276) );
  sky130_fd_sc_hd__nand2_1 U27676 ( .A(n22276), .B(n24452), .Y(n25378) );
  sky130_fd_sc_hd__nand2_1 U27677 ( .A(n27768), .B(n22299), .Y(n22278) );
  sky130_fd_sc_hd__nand2_1 U27678 ( .A(n24364), .B(n22979), .Y(n22277) );
  sky130_fd_sc_hd__o211ai_1 U27679 ( .A1(n22980), .A2(n22279), .B1(n22278), 
        .C1(n22277), .Y(n22280) );
  sky130_fd_sc_hd__nand2_1 U27680 ( .A(n22282), .B(n22996), .Y(n22295) );
  sky130_fd_sc_hd__a22oi_1 U27681 ( .A1(n22988), .A2(
        j202_soc_core_j22_cpu_pc[5]), .B1(j202_soc_core_j22_cpu_rf_gbr[5]), 
        .B2(n22987), .Y(n22294) );
  sky130_fd_sc_hd__nand2_1 U27682 ( .A(n22986), .B(
        j202_soc_core_j22_cpu_rf_gpr[5]), .Y(n22293) );
  sky130_fd_sc_hd__o22ai_1 U27683 ( .A1(n22284), .A2(n22983), .B1(n22283), 
        .B2(n22982), .Y(n22291) );
  sky130_fd_sc_hd__nor2_1 U27684 ( .A(n22286), .B(n22285), .Y(n22290) );
  sky130_fd_sc_hd__o22ai_1 U27685 ( .A1(n22288), .A2(n22897), .B1(n22287), 
        .B2(n22894), .Y(n22289) );
  sky130_fd_sc_hd__nor3_1 U27686 ( .A(n22291), .B(n22290), .C(n22289), .Y(
        n22292) );
  sky130_fd_sc_hd__nand4_1 U27687 ( .A(n22295), .B(n22294), .C(n22293), .D(
        n22292), .Y(n22951) );
  sky130_fd_sc_hd__nand2b_1 U27688 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[21]), .Y(n25377) );
  sky130_fd_sc_hd__nand2_1 U27689 ( .A(n23005), .B(
        j202_soc_core_j22_cpu_rf_gpr[500]), .Y(n22297) );
  sky130_fd_sc_hd__nand2_1 U27690 ( .A(n23003), .B(
        j202_soc_core_j22_cpu_rf_gpr[21]), .Y(n22296) );
  sky130_fd_sc_hd__o211a_2 U27691 ( .A1(n23000), .A2(n22298), .B1(n22297), 
        .C1(n22296), .X(n22308) );
  sky130_fd_sc_hd__nand2_1 U27692 ( .A(n28056), .B(n22299), .Y(n25376) );
  sky130_fd_sc_hd__nor2_1 U27693 ( .A(n27052), .B(n25376), .Y(n22300) );
  sky130_fd_sc_hd__a22oi_1 U27694 ( .A1(n23006), .A2(
        j202_soc_core_j22_cpu_rf_pr[21]), .B1(n22300), .B2(n27717), .Y(n22304)
         );
  sky130_fd_sc_hd__nand2_1 U27695 ( .A(n23008), .B(
        j202_soc_core_j22_cpu_rf_vbr[21]), .Y(n22303) );
  sky130_fd_sc_hd__nand2_1 U27696 ( .A(n23009), .B(
        j202_soc_core_j22_cpu_rf_tmp[21]), .Y(n22302) );
  sky130_fd_sc_hd__nand2_1 U27697 ( .A(n22722), .B(
        j202_soc_core_j22_cpu_rf_gbr[21]), .Y(n22301) );
  sky130_fd_sc_hd__nand4_1 U27698 ( .A(n22304), .B(n22303), .C(n22302), .D(
        n22301), .Y(n22305) );
  sky130_fd_sc_hd__a21oi_1 U27699 ( .A1(n22306), .A2(n23010), .B1(n22305), .Y(
        n22307) );
  sky130_fd_sc_hd__o211ai_1 U27700 ( .A1(n22309), .A2(n25377), .B1(n22308), 
        .C1(n22307), .Y(n22310) );
  sky130_fd_sc_hd__a21oi_1 U27701 ( .A1(n22862), .A2(n22951), .B1(n22310), .Y(
        n22311) );
  sky130_fd_sc_hd__o21ai_0 U27702 ( .A1(n23018), .A2(n25375), .B1(n22311), .Y(
        n22312) );
  sky130_fd_sc_hd__a21oi_1 U27703 ( .A1(n23544), .A2(n23044), .B1(n22312), .Y(
        n22315) );
  sky130_fd_sc_hd__nand2_1 U27704 ( .A(n23469), .B(n25679), .Y(n25379) );
  sky130_fd_sc_hd__nand2_1 U27705 ( .A(n22313), .B(n23044), .Y(n22314) );
  sky130_fd_sc_hd__nand3_1 U27706 ( .A(n12241), .B(n22315), .C(n22314), .Y(
        n29509) );
  sky130_fd_sc_hd__o22ai_1 U27707 ( .A1(n22980), .A2(n22318), .B1(n22365), 
        .B2(n23589), .Y(n22319) );
  sky130_fd_sc_hd__a21oi_1 U27708 ( .A1(n22320), .A2(n24764), .B1(n22319), .Y(
        n25664) );
  sky130_fd_sc_hd__o22ai_1 U27709 ( .A1(n22322), .A2(n23000), .B1(n22321), 
        .B2(n22998), .Y(n22323) );
  sky130_fd_sc_hd__a21oi_1 U27710 ( .A1(j202_soc_core_j22_cpu_rf_gpr[20]), 
        .A2(n23003), .B1(n22323), .Y(n22329) );
  sky130_fd_sc_hd__nand2_1 U27711 ( .A(n23004), .B(n11474), .Y(n25640) );
  sky130_fd_sc_hd__a22oi_1 U27712 ( .A1(n23006), .A2(
        j202_soc_core_j22_cpu_rf_pr[20]), .B1(n23005), .B2(
        j202_soc_core_j22_cpu_rf_gpr[499]), .Y(n22325) );
  sky130_fd_sc_hd__a22oi_1 U27713 ( .A1(n23009), .A2(
        j202_soc_core_j22_cpu_rf_tmp[20]), .B1(n23008), .B2(
        j202_soc_core_j22_cpu_rf_vbr[20]), .Y(n22324) );
  sky130_fd_sc_hd__o211a_2 U27714 ( .A1(n24467), .A2(n25640), .B1(n22325), 
        .C1(n22324), .X(n22328) );
  sky130_fd_sc_hd__nand2_1 U27715 ( .A(n22326), .B(n23010), .Y(n22327) );
  sky130_fd_sc_hd__nand4_1 U27716 ( .A(n22330), .B(n22329), .C(n22328), .D(
        n22327), .Y(n22331) );
  sky130_fd_sc_hd__o21ba_2 U27717 ( .A1(n23018), .A2(n25664), .B1_N(n22331), 
        .X(n22349) );
  sky130_fd_sc_hd__nand2_1 U27718 ( .A(n27362), .B(n25679), .Y(n22347) );
  sky130_fd_sc_hd__nand2_1 U27719 ( .A(n22333), .B(n22332), .Y(n22344) );
  sky130_fd_sc_hd__inv_1 U27720 ( .A(n22334), .Y(n22337) );
  sky130_fd_sc_hd__nand2_1 U27721 ( .A(n22017), .B(n22337), .Y(n22802) );
  sky130_fd_sc_hd__nor2_1 U27722 ( .A(n22338), .B(n22802), .Y(n22340) );
  sky130_fd_sc_hd__nand2_1 U27723 ( .A(n23030), .B(n22340), .Y(n22342) );
  sky130_fd_sc_hd__a21oi_1 U27724 ( .A1(n22789), .A2(n22337), .B1(n22336), .Y(
        n22803) );
  sky130_fd_sc_hd__o21ai_1 U27725 ( .A1(n22338), .A2(n22803), .B1(n22800), .Y(
        n22339) );
  sky130_fd_sc_hd__a21oi_1 U27726 ( .A1(n23036), .A2(n22340), .B1(n22339), .Y(
        n22341) );
  sky130_fd_sc_hd__xnor2_1 U27727 ( .A(n22344), .B(n22343), .Y(n22345) );
  sky130_fd_sc_hd__nand2_1 U27728 ( .A(n25665), .B(n23044), .Y(n22348) );
  sky130_fd_sc_hd__nand3_1 U27729 ( .A(n22316), .B(n22349), .C(n22348), .Y(
        n29508) );
  sky130_fd_sc_hd__nand2_1 U27730 ( .A(n22351), .B(n22350), .Y(n22361) );
  sky130_fd_sc_hd__inv_1 U27731 ( .A(n22352), .Y(n22355) );
  sky130_fd_sc_hd__nor2_1 U27732 ( .A(n22355), .B(n22602), .Y(n22357) );
  sky130_fd_sc_hd__nand2_1 U27733 ( .A(n23030), .B(n22357), .Y(n22359) );
  sky130_fd_sc_hd__o21ai_1 U27734 ( .A1(n22355), .A2(n22604), .B1(n22354), .Y(
        n22356) );
  sky130_fd_sc_hd__a21oi_1 U27735 ( .A1(n23036), .A2(n22357), .B1(n22356), .Y(
        n22358) );
  sky130_fd_sc_hd__o21ai_1 U27736 ( .A1(n22359), .A2(n12349), .B1(n22358), .Y(
        n22360) );
  sky130_fd_sc_hd__xnor2_1 U27737 ( .A(n22361), .B(n22360), .Y(n22362) );
  sky130_fd_sc_hd__a22oi_1 U27738 ( .A1(j202_soc_core_j22_cpu_ml_mach[18]), 
        .A2(n23041), .B1(n22362), .B2(n24452), .Y(n25866) );
  sky130_fd_sc_hd__nand2_1 U27739 ( .A(n25890), .B(n25679), .Y(n22363) );
  sky130_fd_sc_hd__nand2_1 U27740 ( .A(n25866), .B(n22363), .Y(n27117) );
  sky130_fd_sc_hd__nand2_1 U27741 ( .A(n27117), .B(n23044), .Y(n22379) );
  sky130_fd_sc_hd__o22ai_1 U27742 ( .A1(n22980), .A2(n22366), .B1(n22365), 
        .B2(n23593), .Y(n22367) );
  sky130_fd_sc_hd__a21oi_1 U27743 ( .A1(n22368), .A2(n24764), .B1(n22367), .Y(
        n25869) );
  sky130_fd_sc_hd__nand2_1 U27744 ( .A(n23003), .B(
        j202_soc_core_j22_cpu_rf_gpr[18]), .Y(n22370) );
  sky130_fd_sc_hd__nand2_1 U27745 ( .A(n22722), .B(
        j202_soc_core_j22_cpu_rf_gbr[18]), .Y(n22369) );
  sky130_fd_sc_hd__o211ai_1 U27746 ( .A1(n13377), .A2(n23000), .B1(n22370), 
        .C1(n22369), .Y(n22374) );
  sky130_fd_sc_hd__nand2_1 U27747 ( .A(n23004), .B(n11392), .Y(n25873) );
  sky130_fd_sc_hd__a22oi_1 U27748 ( .A1(n23006), .A2(
        j202_soc_core_j22_cpu_rf_pr[18]), .B1(n23005), .B2(
        j202_soc_core_j22_cpu_rf_gpr[497]), .Y(n22372) );
  sky130_fd_sc_hd__a22oi_1 U27749 ( .A1(n23009), .A2(
        j202_soc_core_j22_cpu_rf_tmp[18]), .B1(n23008), .B2(
        j202_soc_core_j22_cpu_rf_vbr[18]), .Y(n22371) );
  sky130_fd_sc_hd__o211ai_1 U27750 ( .A1(n24467), .A2(n25873), .B1(n22372), 
        .C1(n22371), .Y(n22373) );
  sky130_fd_sc_hd__a211o_1 U27751 ( .A1(n23010), .A2(n22375), .B1(n22374), 
        .C1(n22373), .X(n22376) );
  sky130_fd_sc_hd__a21oi_1 U27752 ( .A1(n22862), .A2(n22428), .B1(n22376), .Y(
        n22377) );
  sky130_fd_sc_hd__o21a_1 U27753 ( .A1(n23018), .A2(n25869), .B1(n22377), .X(
        n22378) );
  sky130_fd_sc_hd__nand3_1 U27754 ( .A(n22379), .B(n22437), .C(n22378), .Y(
        n29505) );
  sky130_fd_sc_hd__nand2_1 U27755 ( .A(n27617), .B(n23044), .Y(n22392) );
  sky130_fd_sc_hd__nand2_1 U27756 ( .A(n22384), .B(n22452), .Y(n22388) );
  sky130_fd_sc_hd__nand4_1 U27757 ( .A(n22387), .B(n22386), .C(n22385), .D(
        n22388), .Y(n22390) );
  sky130_fd_sc_hd__nand2_1 U27758 ( .A(n22388), .B(n24467), .Y(n22389) );
  sky130_fd_sc_hd__nand2_1 U27759 ( .A(n22390), .B(n22389), .Y(n22391) );
  sky130_fd_sc_hd__nand3_1 U27760 ( .A(n22392), .B(n12206), .C(n22391), .Y(
        n29525) );
  sky130_fd_sc_hd__nand2_1 U27761 ( .A(n27462), .B(n23044), .Y(n22403) );
  sky130_fd_sc_hd__nand2_1 U27762 ( .A(n22558), .B(n22452), .Y(n22399) );
  sky130_fd_sc_hd__nand4_1 U27763 ( .A(n22398), .B(n22397), .C(n22396), .D(
        n22399), .Y(n22401) );
  sky130_fd_sc_hd__nand2_1 U27764 ( .A(n22399), .B(n24467), .Y(n22400) );
  sky130_fd_sc_hd__nand2_1 U27765 ( .A(n22401), .B(n22400), .Y(n22402) );
  sky130_fd_sc_hd__nand3_1 U27766 ( .A(n22560), .B(n22403), .C(n22402), .Y(
        n29524) );
  sky130_fd_sc_hd__nand2_1 U27767 ( .A(n27153), .B(n23044), .Y(n22412) );
  sky130_fd_sc_hd__nand2_1 U27768 ( .A(n22951), .B(n22452), .Y(n22408) );
  sky130_fd_sc_hd__nand3_1 U27769 ( .A(n22407), .B(n22406), .C(n22408), .Y(
        n22410) );
  sky130_fd_sc_hd__nand2_1 U27770 ( .A(n22408), .B(n24467), .Y(n22409) );
  sky130_fd_sc_hd__nand2_1 U27771 ( .A(n22410), .B(n22409), .Y(n22411) );
  sky130_fd_sc_hd__nand3_1 U27772 ( .A(n12241), .B(n22412), .C(n22411), .Y(
        n29523) );
  sky130_fd_sc_hd__nor3_1 U27773 ( .A(j202_soc_core_aquc_WE_), .B(n22413), .C(
        n22414), .Y(n29541) );
  sky130_fd_sc_hd__nand2_1 U27774 ( .A(j202_soc_core_aquc_WE_), .B(
        j202_soc_core_aquc_CE__1_), .Y(n25316) );
  sky130_fd_sc_hd__nor2_1 U27775 ( .A(n22414), .B(n25316), .Y(n29483) );
  sky130_fd_sc_hd__nand2_1 U27776 ( .A(n27645), .B(n23044), .Y(n22425) );
  sky130_fd_sc_hd__nor2_1 U27777 ( .A(n22417), .B(n22780), .Y(n22423) );
  sky130_fd_sc_hd__nor3_1 U27778 ( .A(n22420), .B(n22419), .C(n22423), .Y(
        n22422) );
  sky130_fd_sc_hd__o2bb2ai_1 U27779 ( .B1(n27717), .B2(n22423), .A1_N(n22422), 
        .A2_N(n22421), .Y(n22424) );
  sky130_fd_sc_hd__nand2_1 U27780 ( .A(n11460), .B(n30015), .Y(n27144) );
  sky130_fd_sc_hd__nand2_1 U27781 ( .A(n27144), .B(n23044), .Y(n22436) );
  sky130_fd_sc_hd__nand2_1 U27782 ( .A(n22428), .B(n22452), .Y(n22432) );
  sky130_fd_sc_hd__nand4_1 U27783 ( .A(n22431), .B(n22430), .C(n22429), .D(
        n22432), .Y(n22434) );
  sky130_fd_sc_hd__nand2_1 U27784 ( .A(n22432), .B(n24467), .Y(n22433) );
  sky130_fd_sc_hd__nand2_1 U27785 ( .A(n22434), .B(n22433), .Y(n22435) );
  sky130_fd_sc_hd__nand3_1 U27786 ( .A(n22437), .B(n22436), .C(n22435), .Y(
        n29518) );
  sky130_fd_sc_hd__nand2_1 U27787 ( .A(n24772), .B(n23044), .Y(n22447) );
  sky130_fd_sc_hd__nand2_1 U27788 ( .A(n22440), .B(n22452), .Y(n22443) );
  sky130_fd_sc_hd__nand3_1 U27789 ( .A(n22442), .B(n22441), .C(n22443), .Y(
        n22445) );
  sky130_fd_sc_hd__nand2_1 U27790 ( .A(n22443), .B(n24467), .Y(n22444) );
  sky130_fd_sc_hd__nand2_1 U27791 ( .A(n22445), .B(n22444), .Y(n22446) );
  sky130_fd_sc_hd__nand3_1 U27792 ( .A(n22826), .B(n22447), .C(n22446), .Y(
        n29521) );
  sky130_fd_sc_hd__nand2_1 U27793 ( .A(n22450), .B(n22449), .Y(n28054) );
  sky130_fd_sc_hd__nand2_1 U27794 ( .A(n28054), .B(n23044), .Y(n22461) );
  sky130_fd_sc_hd__nand2_1 U27795 ( .A(n22453), .B(n22452), .Y(n22457) );
  sky130_fd_sc_hd__nand4_1 U27796 ( .A(n22456), .B(n22455), .C(n22454), .D(
        n22457), .Y(n22459) );
  sky130_fd_sc_hd__nand2_1 U27797 ( .A(n22457), .B(n24467), .Y(n22458) );
  sky130_fd_sc_hd__nand2_1 U27798 ( .A(n22459), .B(n22458), .Y(n22460) );
  sky130_fd_sc_hd__nand2_1 U27799 ( .A(n26032), .B(n24764), .Y(n26405) );
  sky130_fd_sc_hd__nand2b_1 U27800 ( .A_N(n22980), .B(
        j202_soc_core_j22_cpu_ml_macl[31]), .Y(n26401) );
  sky130_fd_sc_hd__nand2_1 U27801 ( .A(n24337), .B(n22979), .Y(n26403) );
  sky130_fd_sc_hd__nand3_1 U27802 ( .A(n26405), .B(n26401), .C(n26403), .Y(
        n25768) );
  sky130_fd_sc_hd__o22ai_1 U27803 ( .A1(n22463), .A2(n23000), .B1(n22462), 
        .B2(n22998), .Y(n22464) );
  sky130_fd_sc_hd__a21oi_1 U27804 ( .A1(j202_soc_core_j22_cpu_rf_gpr[31]), 
        .A2(n23003), .B1(n22464), .Y(n22470) );
  sky130_fd_sc_hd__nand2_1 U27805 ( .A(n23004), .B(n25777), .Y(n26400) );
  sky130_fd_sc_hd__a22oi_1 U27806 ( .A1(n23006), .A2(
        j202_soc_core_j22_cpu_rf_pr[31]), .B1(n23005), .B2(
        j202_soc_core_j22_cpu_rf_gpr[510]), .Y(n22465) );
  sky130_fd_sc_hd__o21a_1 U27807 ( .A1(n24467), .A2(n26400), .B1(n22465), .X(
        n22469) );
  sky130_fd_sc_hd__a22oi_1 U27808 ( .A1(n23009), .A2(
        j202_soc_core_j22_cpu_rf_tmp[31]), .B1(n23008), .B2(
        j202_soc_core_j22_cpu_rf_vbr[31]), .Y(n22468) );
  sky130_fd_sc_hd__nand2_1 U27809 ( .A(n22466), .B(n23010), .Y(n22467) );
  sky130_fd_sc_hd__nand4_1 U27810 ( .A(n22470), .B(n22469), .C(n22468), .D(
        n22467), .Y(n22471) );
  sky130_fd_sc_hd__a21oi_1 U27811 ( .A1(n23973), .A2(n22472), .B1(n22471), .Y(
        n22473) );
  sky130_fd_sc_hd__nand2b_1 U27812 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[31]), .Y(n26398) );
  sky130_fd_sc_hd__nor2_1 U27813 ( .A(n22474), .B(n11145), .Y(n22476) );
  sky130_fd_sc_hd__nand2_1 U27814 ( .A(n13046), .B(n22476), .Y(n22477) );
  sky130_fd_sc_hd__nand2_1 U27815 ( .A(n22478), .B(n22477), .Y(n22518) );
  sky130_fd_sc_hd__nor2_1 U27816 ( .A(n22479), .B(n11145), .Y(n22510) );
  sky130_fd_sc_hd__nor2_1 U27817 ( .A(n22510), .B(n13046), .Y(n22599) );
  sky130_fd_sc_hd__nor2_1 U27818 ( .A(n22480), .B(n11145), .Y(n22490) );
  sky130_fd_sc_hd__nor2_1 U27819 ( .A(n22481), .B(n11145), .Y(n22492) );
  sky130_fd_sc_hd__nor2_1 U27820 ( .A(n22490), .B(n22491), .Y(n22678) );
  sky130_fd_sc_hd__nor2_1 U27821 ( .A(n22482), .B(n11145), .Y(n22498) );
  sky130_fd_sc_hd__nand2_1 U27822 ( .A(n22929), .B(n22671), .Y(n22497) );
  sky130_fd_sc_hd__nand2_1 U27823 ( .A(n22483), .B(n22710), .Y(n22675) );
  sky130_fd_sc_hd__nor2_1 U27824 ( .A(n22497), .B(n22675), .Y(n22541) );
  sky130_fd_sc_hd__nor2_1 U27825 ( .A(n22484), .B(n11145), .Y(n22504) );
  sky130_fd_sc_hd__nor2_1 U27826 ( .A(n22504), .B(n22505), .Y(n23026) );
  sky130_fd_sc_hd__nor2_1 U27827 ( .A(n22485), .B(n11145), .Y(n22500) );
  sky130_fd_sc_hd__nor2_1 U27828 ( .A(n22498), .B(n22499), .Y(n22621) );
  sky130_fd_sc_hd__nand2_1 U27829 ( .A(n22540), .B(n22619), .Y(n23033) );
  sky130_fd_sc_hd__nor2_1 U27830 ( .A(n23026), .B(n23033), .Y(n22507) );
  sky130_fd_sc_hd__nand2_1 U27831 ( .A(n22542), .B(n22509), .Y(n22605) );
  sky130_fd_sc_hd__nor2_1 U27832 ( .A(n22599), .B(n22605), .Y(n22512) );
  sky130_fd_sc_hd__nand2_1 U27833 ( .A(n23030), .B(n22514), .Y(n22516) );
  sky130_fd_sc_hd__nand2_1 U27834 ( .A(n22487), .B(n22486), .Y(n22709) );
  sky130_fd_sc_hd__a21oi_1 U27835 ( .A1(n22710), .A2(n22489), .B1(n22488), .Y(
        n22673) );
  sky130_fd_sc_hd__nand2_1 U27836 ( .A(n22491), .B(n22490), .Y(n22928) );
  sky130_fd_sc_hd__nand2_1 U27837 ( .A(n22493), .B(n22492), .Y(n22670) );
  sky130_fd_sc_hd__a21oi_1 U27838 ( .A1(n22671), .A2(n22495), .B1(n22494), .Y(
        n22496) );
  sky130_fd_sc_hd__o21ai_1 U27839 ( .A1(n22497), .A2(n22673), .B1(n22496), .Y(
        n22544) );
  sky130_fd_sc_hd__nand2_1 U27840 ( .A(n22499), .B(n22498), .Y(n22620) );
  sky130_fd_sc_hd__nand2_1 U27841 ( .A(n22501), .B(n22500), .Y(n22618) );
  sky130_fd_sc_hd__a21oi_1 U27842 ( .A1(n22619), .A2(n22503), .B1(n22502), .Y(
        n23031) );
  sky130_fd_sc_hd__nand2_1 U27843 ( .A(n22505), .B(n22504), .Y(n23027) );
  sky130_fd_sc_hd__a21o_1 U27845 ( .A1(n22544), .A2(n22507), .B1(n22506), .X(
        n22508) );
  sky130_fd_sc_hd__a21oi_1 U27846 ( .A1(n22543), .A2(n22509), .B1(n22508), .Y(
        n22603) );
  sky130_fd_sc_hd__nand2_1 U27847 ( .A(n13046), .B(n22510), .Y(n22600) );
  sky130_fd_sc_hd__a21o_1 U27849 ( .A1(n23021), .A2(n22512), .B1(n22511), .X(
        n22513) );
  sky130_fd_sc_hd__a21oi_1 U27850 ( .A1(n23036), .A2(n22514), .B1(n22513), .Y(
        n22515) );
  sky130_fd_sc_hd__xnor2_1 U27851 ( .A(n22518), .B(n22517), .Y(n22519) );
  sky130_fd_sc_hd__nand2_1 U27852 ( .A(n22519), .B(n24452), .Y(n26399) );
  sky130_fd_sc_hd__nand3_1 U27853 ( .A(n26448), .B(n26398), .C(n26399), .Y(
        n25775) );
  sky130_fd_sc_hd__nor2b_1 U27854 ( .B_N(j202_soc_core_qspi_int), .A(n29088), 
        .Y(n29582) );
  sky130_fd_sc_hd__o22ai_1 U27855 ( .A1(n22526), .A2(n22845), .B1(n22522), 
        .B2(n22980), .Y(n22523) );
  sky130_fd_sc_hd__a21oi_1 U27856 ( .A1(n24341), .A2(n22979), .B1(n22523), .Y(
        n22524) );
  sky130_fd_sc_hd__nor2_1 U27857 ( .A(n22526), .B(n22850), .Y(n27051) );
  sky130_fd_sc_hd__a22oi_1 U27858 ( .A1(j202_soc_core_j22_cpu_rf_pr[27]), .A2(
        n23006), .B1(n27051), .B2(n27717), .Y(n22530) );
  sky130_fd_sc_hd__nand2_1 U27859 ( .A(n23008), .B(n30074), .Y(n22529) );
  sky130_fd_sc_hd__nand2_1 U27860 ( .A(n22722), .B(
        j202_soc_core_j22_cpu_rf_gbr[27]), .Y(n22528) );
  sky130_fd_sc_hd__nand2_1 U27861 ( .A(n23009), .B(
        j202_soc_core_j22_cpu_rf_tmp[27]), .Y(n22527) );
  sky130_fd_sc_hd__nand4_1 U27862 ( .A(n22530), .B(n22529), .C(n22528), .D(
        n22527), .Y(n22536) );
  sky130_fd_sc_hd__a2bb2oi_1 U27863 ( .B1(j202_soc_core_j22_cpu_rf_gpr[506]), 
        .B2(n23005), .A1_N(n22531), .A2_N(n23000), .Y(n22535) );
  sky130_fd_sc_hd__nand2_1 U27864 ( .A(n22532), .B(n23010), .Y(n22534) );
  sky130_fd_sc_hd__nand2_1 U27865 ( .A(n23003), .B(
        j202_soc_core_j22_cpu_rf_gpr[27]), .Y(n22533) );
  sky130_fd_sc_hd__nand4b_1 U27866 ( .A_N(n22536), .B(n22535), .C(n22534), .D(
        n22533), .Y(n22537) );
  sky130_fd_sc_hd__a21oi_1 U27867 ( .A1(n23973), .A2(n22538), .B1(n22537), .Y(
        n22539) );
  sky130_fd_sc_hd__o21a_1 U27868 ( .A1(n23018), .A2(n27021), .B1(n22539), .X(
        n22557) );
  sky130_fd_sc_hd__nand2_1 U27869 ( .A(n23476), .B(n22940), .Y(n27020) );
  sky130_fd_sc_hd__nand2b_1 U27870 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[27]), .Y(n27053) );
  sky130_fd_sc_hd__nand2_1 U27871 ( .A(n22540), .B(n22620), .Y(n22554) );
  sky130_fd_sc_hd__inv_1 U27872 ( .A(n22542), .Y(n22672) );
  sky130_fd_sc_hd__nor2_1 U27873 ( .A(n22546), .B(n22672), .Y(n22548) );
  sky130_fd_sc_hd__nand2_1 U27874 ( .A(n22017), .B(n22548), .Y(n23029) );
  sky130_fd_sc_hd__nand2_1 U27875 ( .A(n23030), .B(n22550), .Y(n22552) );
  sky130_fd_sc_hd__o21ai_1 U27876 ( .A1(n22546), .A2(n22674), .B1(n22545), .Y(
        n22547) );
  sky130_fd_sc_hd__a21oi_1 U27877 ( .A1(n22789), .A2(n22548), .B1(n22547), .Y(
        n23032) );
  sky130_fd_sc_hd__inv_1 U27878 ( .A(n23032), .Y(n22549) );
  sky130_fd_sc_hd__a21oi_1 U27879 ( .A1(n23036), .A2(n22550), .B1(n22549), .Y(
        n22551) );
  sky130_fd_sc_hd__xnor2_1 U27881 ( .A(n22554), .B(n22553), .Y(n22555) );
  sky130_fd_sc_hd__nand2_1 U27882 ( .A(n22555), .B(n24452), .Y(n27055) );
  sky130_fd_sc_hd__nand3_1 U27883 ( .A(n27020), .B(n27053), .C(n27055), .Y(
        n23570) );
  sky130_fd_sc_hd__nand2_1 U27884 ( .A(n23570), .B(n23044), .Y(n22556) );
  sky130_fd_sc_hd__nand2_1 U27885 ( .A(n22558), .B(n22950), .Y(n22559) );
  sky130_fd_sc_hd__nor2_1 U27886 ( .A(n22561), .B(n22980), .Y(n25112) );
  sky130_fd_sc_hd__nand2_1 U27887 ( .A(n22564), .B(n22563), .Y(n22565) );
  sky130_fd_sc_hd__nand2_1 U27888 ( .A(n24458), .B(n24764), .Y(n22571) );
  sky130_fd_sc_hd__nand2_1 U27889 ( .A(n22567), .B(n22566), .Y(n22569) );
  sky130_fd_sc_hd__xnor2_1 U27890 ( .A(n22569), .B(n22568), .Y(n24462) );
  sky130_fd_sc_hd__nand2_1 U27891 ( .A(n24462), .B(n22979), .Y(n22570) );
  sky130_fd_sc_hd__nand2_1 U27892 ( .A(n22571), .B(n22570), .Y(n25129) );
  sky130_fd_sc_hd__nor2_1 U27893 ( .A(n25112), .B(n25129), .Y(n25144) );
  sky130_fd_sc_hd__o22ai_1 U27894 ( .A1(n22573), .A2(n22983), .B1(n22982), 
        .B2(n22572), .Y(n22574) );
  sky130_fd_sc_hd__a21oi_1 U27895 ( .A1(n22986), .A2(
        j202_soc_core_j22_cpu_rf_gpr[14]), .B1(n22574), .Y(n22578) );
  sky130_fd_sc_hd__a22oi_1 U27896 ( .A1(n22988), .A2(
        j202_soc_core_j22_cpu_pc[14]), .B1(n22987), .B2(
        j202_soc_core_j22_cpu_rf_gbr[14]), .Y(n22577) );
  sky130_fd_sc_hd__nand2_1 U27897 ( .A(n22989), .B(
        j202_soc_core_j22_cpu_rf_tmp[14]), .Y(n22576) );
  sky130_fd_sc_hd__nand2_1 U27898 ( .A(n22990), .B(
        j202_soc_core_j22_cpu_rf_vbr[14]), .Y(n22575) );
  sky130_fd_sc_hd__nand4_1 U27899 ( .A(n22578), .B(n22577), .C(n22576), .D(
        n22575), .Y(n22579) );
  sky130_fd_sc_hd__a21o_1 U27900 ( .A1(n22580), .A2(n22996), .B1(n22579), .X(
        n24451) );
  sky130_fd_sc_hd__o22ai_1 U27901 ( .A1(n22582), .A2(n23000), .B1(n22581), 
        .B2(n22998), .Y(n22583) );
  sky130_fd_sc_hd__a21oi_1 U27902 ( .A1(j202_soc_core_j22_cpu_rf_gpr[30]), 
        .A2(n23003), .B1(n22583), .Y(n22589) );
  sky130_fd_sc_hd__nand2_1 U27903 ( .A(n23004), .B(n12425), .Y(n25111) );
  sky130_fd_sc_hd__a22oi_1 U27904 ( .A1(n23006), .A2(
        j202_soc_core_j22_cpu_rf_pr[30]), .B1(n23005), .B2(
        j202_soc_core_j22_cpu_rf_gpr[509]), .Y(n22584) );
  sky130_fd_sc_hd__o21a_1 U27905 ( .A1(n24467), .A2(n25111), .B1(n22584), .X(
        n22588) );
  sky130_fd_sc_hd__a22oi_1 U27906 ( .A1(n23009), .A2(
        j202_soc_core_j22_cpu_rf_tmp[30]), .B1(n23008), .B2(
        j202_soc_core_j22_cpu_rf_vbr[30]), .Y(n22587) );
  sky130_fd_sc_hd__nand2_1 U27907 ( .A(n22585), .B(n23010), .Y(n22586) );
  sky130_fd_sc_hd__nand4_1 U27908 ( .A(n22589), .B(n22588), .C(n22587), .D(
        n22586), .Y(n22590) );
  sky130_fd_sc_hd__a21oi_1 U27909 ( .A1(n24451), .A2(n23973), .B1(n22590), .Y(
        n22591) );
  sky130_fd_sc_hd__nand2_1 U27910 ( .A(n12098), .B(n22592), .Y(n22598) );
  sky130_fd_sc_hd__nand2_1 U27912 ( .A(n23030), .B(n22595), .Y(n22597) );
  sky130_fd_sc_hd__o21ai_1 U27913 ( .A1(n22593), .A2(n22604), .B1(n23019), .Y(
        n22594) );
  sky130_fd_sc_hd__nand2_1 U27914 ( .A(n24453), .B(n25679), .Y(n22615) );
  sky130_fd_sc_hd__nand2_1 U27915 ( .A(n22601), .B(n22600), .Y(n22611) );
  sky130_fd_sc_hd__nor2_1 U27916 ( .A(n22605), .B(n22602), .Y(n22607) );
  sky130_fd_sc_hd__nand2_1 U27917 ( .A(n23030), .B(n22607), .Y(n22609) );
  sky130_fd_sc_hd__o21ai_1 U27918 ( .A1(n22605), .A2(n22604), .B1(n22603), .Y(
        n22606) );
  sky130_fd_sc_hd__a21oi_1 U27919 ( .A1(n23036), .A2(n22607), .B1(n22606), .Y(
        n22608) );
  sky130_fd_sc_hd__xnor2_1 U27920 ( .A(n22611), .B(n22610), .Y(n22612) );
  sky130_fd_sc_hd__nand2_1 U27921 ( .A(n22612), .B(n24452), .Y(n22614) );
  sky130_fd_sc_hd__nand2_1 U27922 ( .A(n23041), .B(
        j202_soc_core_j22_cpu_ml_mach[30]), .Y(n22613) );
  sky130_fd_sc_hd__nand3_1 U27923 ( .A(n22615), .B(n22614), .C(n22613), .Y(
        n25128) );
  sky130_fd_sc_hd__nand2_1 U27924 ( .A(n25128), .B(n23044), .Y(n22616) );
  sky130_fd_sc_hd__nand2_1 U27925 ( .A(n22619), .B(n22618), .Y(n22627) );
  sky130_fd_sc_hd__nor2_1 U27926 ( .A(n22621), .B(n23029), .Y(n22623) );
  sky130_fd_sc_hd__nand2_1 U27927 ( .A(n23030), .B(n22623), .Y(n22625) );
  sky130_fd_sc_hd__o21ai_1 U27928 ( .A1(n22621), .A2(n23032), .B1(n22620), .Y(
        n22622) );
  sky130_fd_sc_hd__a21oi_1 U27929 ( .A1(n23036), .A2(n22623), .B1(n22622), .Y(
        n22624) );
  sky130_fd_sc_hd__xnor2_1 U27930 ( .A(n22627), .B(n22626), .Y(n22628) );
  sky130_fd_sc_hd__nand2_1 U27931 ( .A(n22628), .B(n24452), .Y(n23579) );
  sky130_fd_sc_hd__nand2_1 U27932 ( .A(n24349), .B(n22979), .Y(n22632) );
  sky130_fd_sc_hd__nand2_1 U27933 ( .A(n27768), .B(n23582), .Y(n22629) );
  sky130_fd_sc_hd__o21a_1 U27934 ( .A1(n22630), .A2(n22980), .B1(n22629), .X(
        n22631) );
  sky130_fd_sc_hd__nand2_1 U27935 ( .A(n22632), .B(n22631), .Y(n24763) );
  sky130_fd_sc_hd__a31oi_1 U27936 ( .A1(n22632), .A2(n25439), .A3(n22631), 
        .B1(n27828), .Y(n22633) );
  sky130_fd_sc_hd__nand2b_1 U27938 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[28]), .Y(n23578) );
  sky130_fd_sc_hd__o22ai_1 U27939 ( .A1(n22634), .A2(n22850), .B1(n27052), 
        .B2(n23578), .Y(n22635) );
  sky130_fd_sc_hd__nor2b_1 U27940 ( .B_N(n22636), .A(n22635), .Y(n22638) );
  sky130_fd_sc_hd__nor2_1 U27941 ( .A(n27052), .B(n24854), .Y(n26031) );
  sky130_fd_sc_hd__nand2_1 U27942 ( .A(n23577), .B(n26031), .Y(n22637) );
  sky130_fd_sc_hd__nand2_1 U27944 ( .A(n25817), .B(n27717), .Y(n22653) );
  sky130_fd_sc_hd__nand2_1 U27945 ( .A(n22639), .B(
        j202_soc_core_j22_cpu_pc[28]), .Y(n22643) );
  sky130_fd_sc_hd__nand2_1 U27946 ( .A(n22722), .B(
        j202_soc_core_j22_cpu_rf_gbr[28]), .Y(n22642) );
  sky130_fd_sc_hd__nand2_1 U27947 ( .A(n23009), .B(
        j202_soc_core_j22_cpu_rf_tmp[28]), .Y(n22641) );
  sky130_fd_sc_hd__nand2_1 U27948 ( .A(n23008), .B(
        j202_soc_core_j22_cpu_rf_vbr[28]), .Y(n22640) );
  sky130_fd_sc_hd__nand4_1 U27949 ( .A(n22643), .B(n22642), .C(n22641), .D(
        n22640), .Y(n22648) );
  sky130_fd_sc_hd__nand2_1 U27950 ( .A(n22644), .B(n23010), .Y(n22647) );
  sky130_fd_sc_hd__a22oi_1 U27951 ( .A1(n23006), .A2(
        j202_soc_core_j22_cpu_rf_pr[28]), .B1(n23005), .B2(
        j202_soc_core_j22_cpu_rf_gpr[507]), .Y(n22646) );
  sky130_fd_sc_hd__nand2_1 U27952 ( .A(n23003), .B(
        j202_soc_core_j22_cpu_rf_gpr[28]), .Y(n22645) );
  sky130_fd_sc_hd__nand4b_1 U27953 ( .A_N(n22648), .B(n22647), .C(n22646), .D(
        n22645), .Y(n22649) );
  sky130_fd_sc_hd__a21oi_1 U27954 ( .A1(n22650), .A2(n23973), .B1(n22649), .Y(
        n22651) );
  sky130_fd_sc_hd__nand2_1 U27955 ( .A(n24313), .B(n22979), .Y(n22654) );
  sky130_fd_sc_hd__a21oi_1 U27957 ( .A1(n22657), .A2(n24764), .B1(n22656), .Y(
        n27783) );
  sky130_fd_sc_hd__o22ai_1 U27958 ( .A1(n22659), .A2(n23000), .B1(n22658), 
        .B2(n22998), .Y(n22660) );
  sky130_fd_sc_hd__a21oi_1 U27959 ( .A1(j202_soc_core_j22_cpu_rf_gpr[26]), 
        .A2(n23003), .B1(n22660), .Y(n22666) );
  sky130_fd_sc_hd__nand2_1 U27960 ( .A(n23004), .B(n27767), .Y(n27826) );
  sky130_fd_sc_hd__a22oi_1 U27961 ( .A1(n23006), .A2(
        j202_soc_core_j22_cpu_rf_pr[26]), .B1(n23005), .B2(
        j202_soc_core_j22_cpu_rf_gpr[505]), .Y(n22661) );
  sky130_fd_sc_hd__o21a_1 U27962 ( .A1(n24467), .A2(n27826), .B1(n22661), .X(
        n22665) );
  sky130_fd_sc_hd__a22oi_1 U27963 ( .A1(n23009), .A2(
        j202_soc_core_j22_cpu_rf_tmp[26]), .B1(n23008), .B2(
        j202_soc_core_j22_cpu_rf_vbr[26]), .Y(n22664) );
  sky130_fd_sc_hd__nand2_1 U27964 ( .A(n22662), .B(n23010), .Y(n22663) );
  sky130_fd_sc_hd__nand4_1 U27965 ( .A(n22666), .B(n22665), .C(n22664), .D(
        n22663), .Y(n22667) );
  sky130_fd_sc_hd__a21oi_1 U27966 ( .A1(n22668), .A2(n23973), .B1(n22667), .Y(
        n22669) );
  sky130_fd_sc_hd__o21a_1 U27967 ( .A1(n23018), .A2(n27783), .B1(n22669), .X(
        n22687) );
  sky130_fd_sc_hd__nand2_1 U27968 ( .A(n23471), .B(n25679), .Y(n27781) );
  sky130_fd_sc_hd__nand2b_1 U27969 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[26]), .Y(n27827) );
  sky130_fd_sc_hd__nand2_1 U27970 ( .A(n22671), .B(n22670), .Y(n22684) );
  sky130_fd_sc_hd__nor2_1 U27971 ( .A(n22675), .B(n22672), .Y(n22677) );
  sky130_fd_sc_hd__nand2_1 U27972 ( .A(n22017), .B(n22677), .Y(n22930) );
  sky130_fd_sc_hd__nor2_1 U27973 ( .A(n22678), .B(n22930), .Y(n22680) );
  sky130_fd_sc_hd__nand2_1 U27974 ( .A(n23030), .B(n22680), .Y(n22682) );
  sky130_fd_sc_hd__o21ai_1 U27975 ( .A1(n22675), .A2(n22674), .B1(n22673), .Y(
        n22676) );
  sky130_fd_sc_hd__a21oi_1 U27976 ( .A1(n23036), .A2(n22680), .B1(n22679), .Y(
        n22681) );
  sky130_fd_sc_hd__o21ai_1 U27977 ( .A1(n22682), .A2(n12349), .B1(n22681), .Y(
        n22683) );
  sky130_fd_sc_hd__xnor2_1 U27978 ( .A(n22684), .B(n22683), .Y(n22685) );
  sky130_fd_sc_hd__nand2_1 U27979 ( .A(n22685), .B(n24452), .Y(n27829) );
  sky130_fd_sc_hd__nand3_1 U27980 ( .A(n27781), .B(n27827), .C(n27829), .Y(
        n23562) );
  sky130_fd_sc_hd__nand2_1 U27981 ( .A(n23562), .B(n23044), .Y(n22686) );
  sky130_fd_sc_hd__nand2b_1 U27982 ( .A_N(n24090), .B(n22739), .Y(n22708) );
  sky130_fd_sc_hd__a21oi_1 U27983 ( .A1(n22692), .A2(n22691), .B1(n22690), .Y(
        n22697) );
  sky130_fd_sc_hd__nand2_1 U27984 ( .A(n22695), .B(n22694), .Y(n22696) );
  sky130_fd_sc_hd__xor2_1 U27985 ( .A(n22697), .B(n22696), .X(n26956) );
  sky130_fd_sc_hd__nand2_1 U27986 ( .A(n22698), .B(j202_soc_core_j22_cpu_pc[9]), .Y(n22699) );
  sky130_fd_sc_hd__xor2_1 U27987 ( .A(n22699), .B(n14345), .X(n24092) );
  sky130_fd_sc_hd__o22ai_1 U27988 ( .A1(n27776), .A2(n13365), .B1(n27798), 
        .B2(n11186), .Y(n22700) );
  sky130_fd_sc_hd__a21oi_1 U27989 ( .A1(n22701), .A2(n28473), .B1(n22700), .Y(
        n22704) );
  sky130_fd_sc_hd__nand2_1 U27990 ( .A(n22702), .B(n28473), .Y(n22703) );
  sky130_fd_sc_hd__o211ai_1 U27991 ( .A1(n27776), .A2(n22705), .B1(n22704), 
        .C1(n22703), .Y(n22706) );
  sky130_fd_sc_hd__a21oi_1 U27992 ( .A1(n26956), .A2(n17225), .B1(n22706), .Y(
        n22707) );
  sky130_fd_sc_hd__nand2_1 U27993 ( .A(n22708), .B(n22707), .Y(n29548) );
  sky130_fd_sc_hd__nand2b_1 U27994 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[24]), .Y(n24155) );
  sky130_fd_sc_hd__nand2_1 U27995 ( .A(n22710), .B(n22709), .Y(n22720) );
  sky130_fd_sc_hd__nor2_1 U27996 ( .A(n22714), .B(n22711), .Y(n22716) );
  sky130_fd_sc_hd__nand2_1 U27997 ( .A(n23030), .B(n22716), .Y(n22718) );
  sky130_fd_sc_hd__o21ai_1 U27998 ( .A1(n22714), .A2(n22713), .B1(n22712), .Y(
        n22715) );
  sky130_fd_sc_hd__a21oi_1 U27999 ( .A1(n23036), .A2(n22716), .B1(n22715), .Y(
        n22717) );
  sky130_fd_sc_hd__o21ai_1 U28000 ( .A1(n22718), .A2(n12349), .B1(n22717), .Y(
        n22719) );
  sky130_fd_sc_hd__xnor2_1 U28001 ( .A(n22720), .B(n22719), .Y(n22721) );
  sky130_fd_sc_hd__nand2_1 U28002 ( .A(n22721), .B(n24452), .Y(n24147) );
  sky130_fd_sc_hd__nand2_1 U28003 ( .A(n23003), .B(
        j202_soc_core_j22_cpu_rf_gpr[24]), .Y(n22724) );
  sky130_fd_sc_hd__nand2_1 U28004 ( .A(n22722), .B(
        j202_soc_core_j22_cpu_rf_gbr[24]), .Y(n22723) );
  sky130_fd_sc_hd__o211ai_1 U28005 ( .A1(n22725), .A2(n23000), .B1(n22724), 
        .C1(n22723), .Y(n22729) );
  sky130_fd_sc_hd__nand2_1 U28006 ( .A(n23004), .B(
        j202_soc_core_j22_cpu_ml_bufa[24]), .Y(n24154) );
  sky130_fd_sc_hd__a22oi_1 U28007 ( .A1(n23006), .A2(
        j202_soc_core_j22_cpu_rf_pr[24]), .B1(n23005), .B2(
        j202_soc_core_j22_cpu_rf_gpr[503]), .Y(n22727) );
  sky130_fd_sc_hd__a22oi_1 U28008 ( .A1(n23009), .A2(
        j202_soc_core_j22_cpu_rf_tmp[24]), .B1(n23008), .B2(
        j202_soc_core_j22_cpu_rf_vbr[24]), .Y(n22726) );
  sky130_fd_sc_hd__o211ai_1 U28009 ( .A1(n24467), .A2(n24154), .B1(n22727), 
        .C1(n22726), .Y(n22728) );
  sky130_fd_sc_hd__a211oi_1 U28010 ( .A1(n23010), .A2(n22730), .B1(n22729), 
        .C1(n22728), .Y(n22734) );
  sky130_fd_sc_hd__nand2_1 U28011 ( .A(n22731), .B(n24764), .Y(n24151) );
  sky130_fd_sc_hd__nand2_1 U28012 ( .A(n26966), .B(n22979), .Y(n24149) );
  sky130_fd_sc_hd__nand2b_1 U28013 ( .A_N(n22980), .B(
        j202_soc_core_j22_cpu_ml_macl[24]), .Y(n24148) );
  sky130_fd_sc_hd__nand3_1 U28014 ( .A(n24151), .B(n24149), .C(n24148), .Y(
        n25211) );
  sky130_fd_sc_hd__nand2_1 U28015 ( .A(n25211), .B(n22732), .Y(n22733) );
  sky130_fd_sc_hd__o211ai_1 U28016 ( .A1(n22735), .A2(n24299), .B1(n22734), 
        .C1(n22733), .Y(n22736) );
  sky130_fd_sc_hd__a21oi_1 U28017 ( .A1(n23574), .A2(n23044), .B1(n22736), .Y(
        n22738) );
  sky130_fd_sc_hd__nor2b_1 U28018 ( .B_N(
        j202_soc_core_intc_core_00_rg_sint[15]), .A(n29088), .Y(n29567) );
  sky130_fd_sc_hd__nor2b_1 U28019 ( .B_N(
        j202_soc_core_intc_core_00_rg_sint[14]), .A(n29088), .Y(n29576) );
  sky130_fd_sc_hd__nor2b_1 U28020 ( .B_N(
        j202_soc_core_intc_core_00_rg_sint[13]), .A(j202_soc_core_rst), .Y(
        n29566) );
  sky130_fd_sc_hd__nor2b_1 U28021 ( .B_N(
        j202_soc_core_intc_core_00_rg_sint[12]), .A(n29088), .Y(n29562) );
  sky130_fd_sc_hd__nor2b_1 U28022 ( .B_N(
        j202_soc_core_intc_core_00_rg_sint[11]), .A(n29088), .Y(n29590) );
  sky130_fd_sc_hd__nor2b_1 U28023 ( .B_N(
        j202_soc_core_intc_core_00_rg_sint[10]), .A(n29088), .Y(n29558) );
  sky130_fd_sc_hd__nor2b_1 U28024 ( .B_N(j202_soc_core_intc_core_00_rg_sint[9]), .A(n29088), .Y(n29574) );
  sky130_fd_sc_hd__nor2b_1 U28025 ( .B_N(j202_soc_core_intc_core_00_rg_sint[8]), .A(n29088), .Y(n29575) );
  sky130_fd_sc_hd__nor2b_1 U28026 ( .B_N(j202_soc_core_intc_core_00_rg_sint[7]), .A(n29088), .Y(n29572) );
  sky130_fd_sc_hd__nor2b_1 U28027 ( .B_N(j202_soc_core_intc_core_00_rg_sint[6]), .A(n29088), .Y(n29573) );
  sky130_fd_sc_hd__nor2b_1 U28028 ( .B_N(j202_soc_core_intc_core_00_rg_sint[5]), .A(j202_soc_core_rst), .Y(n29570) );
  sky130_fd_sc_hd__nor2b_1 U28029 ( .B_N(j202_soc_core_intc_core_00_rg_sint[4]), .A(n29088), .Y(n29571) );
  sky130_fd_sc_hd__nor2b_1 U28030 ( .B_N(j202_soc_core_intc_core_00_rg_sint[3]), .A(n29088), .Y(n29584) );
  sky130_fd_sc_hd__nor2b_1 U28031 ( .B_N(j202_soc_core_intc_core_00_rg_sint[2]), .A(n29088), .Y(n29561) );
  sky130_fd_sc_hd__nor2b_1 U28032 ( .B_N(j202_soc_core_intc_core_00_rg_sint[1]), .A(n29088), .Y(n29544) );
  sky130_fd_sc_hd__nor2b_1 U28033 ( .B_N(j202_soc_core_intc_core_00_rg_sint[0]), .A(n29088), .Y(n29543) );
  sky130_fd_sc_hd__nand2_1 U28034 ( .A(n29486), .B(n22739), .Y(n22758) );
  sky130_fd_sc_hd__nand2_1 U28035 ( .A(n22740), .B(j202_soc_core_j22_cpu_pc[7]), .Y(n22742) );
  sky130_fd_sc_hd__xor2_1 U28036 ( .A(n22742), .B(n22741), .X(n26974) );
  sky130_fd_sc_hd__o22a_1 U28037 ( .A1(n26317), .A2(n11186), .B1(n24931), .B2(
        n22743), .X(n22744) );
  sky130_fd_sc_hd__a21oi_1 U28039 ( .A1(n26974), .A2(n22747), .B1(n22746), .Y(
        n22757) );
  sky130_fd_sc_hd__nand2_1 U28040 ( .A(n22750), .B(n22749), .Y(n22755) );
  sky130_fd_sc_hd__xnor2_1 U28042 ( .A(n22755), .B(n22754), .Y(n24947) );
  sky130_fd_sc_hd__nand2_1 U28043 ( .A(n24947), .B(n17225), .Y(n22756) );
  sky130_fd_sc_hd__nand3_1 U28044 ( .A(n22758), .B(n22757), .C(n22756), .Y(
        n29552) );
  sky130_fd_sc_hd__nor2_1 U28045 ( .A(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[0]), .B(n22759), .Y(
        n28201) );
  sky130_fd_sc_hd__nand2_1 U28046 ( .A(n28201), .B(n22760), .Y(n28162) );
  sky130_fd_sc_hd__nor4_1 U28047 ( .A(n28162), .B(n22761), .C(n28203), .D(
        n28164), .Y(n29585) );
  sky130_fd_sc_hd__nor2b_1 U28048 ( .B_N(j202_soc_core_bldc_int), .A(n29088), 
        .Y(n29586) );
  sky130_fd_sc_hd__buf_2 U28049 ( .A(j202_soc_core_j22_cpu_ml_bufa[16]), .X(
        n24829) );
  sky130_fd_sc_hd__nand2_1 U28050 ( .A(n27768), .B(n24829), .Y(n22763) );
  sky130_fd_sc_hd__nand2_1 U28051 ( .A(n24353), .B(n22979), .Y(n22762) );
  sky130_fd_sc_hd__o211ai_1 U28052 ( .A1(n22980), .A2(n22764), .B1(n22763), 
        .C1(n22762), .Y(n22765) );
  sky130_fd_sc_hd__a21oi_1 U28053 ( .A1(n22766), .A2(n24764), .B1(n22765), .Y(
        n24851) );
  sky130_fd_sc_hd__nand2_1 U28054 ( .A(n23003), .B(
        j202_soc_core_j22_cpu_rf_gpr[16]), .Y(n22768) );
  sky130_fd_sc_hd__nand2_1 U28055 ( .A(n23006), .B(
        j202_soc_core_j22_cpu_rf_pr[16]), .Y(n22767) );
  sky130_fd_sc_hd__o211ai_1 U28056 ( .A1(n22769), .A2(n23000), .B1(n22768), 
        .C1(n22767), .Y(n22775) );
  sky130_fd_sc_hd__nor2_1 U28057 ( .A(n22770), .B(n22850), .Y(n24835) );
  sky130_fd_sc_hd__a22oi_1 U28058 ( .A1(n23005), .A2(
        j202_soc_core_j22_cpu_rf_gpr[495]), .B1(n24835), .B2(n27717), .Y(
        n22774) );
  sky130_fd_sc_hd__a2bb2oi_1 U28059 ( .B1(j202_soc_core_j22_cpu_rf_tmp[16]), 
        .B2(n23009), .A1_N(n22771), .A2_N(n22998), .Y(n22773) );
  sky130_fd_sc_hd__nand2_1 U28060 ( .A(n23008), .B(
        j202_soc_core_j22_cpu_rf_vbr[16]), .Y(n22772) );
  sky130_fd_sc_hd__nand4b_1 U28061 ( .A_N(n22775), .B(n22774), .C(n22773), .D(
        n22772), .Y(n22776) );
  sky130_fd_sc_hd__a21oi_1 U28062 ( .A1(n23010), .A2(n22777), .B1(n22776), .Y(
        n22778) );
  sky130_fd_sc_hd__o21a_1 U28063 ( .A1(n22780), .A2(n22779), .B1(n22778), .X(
        n22781) );
  sky130_fd_sc_hd__o21a_1 U28064 ( .A1(n23018), .A2(n24851), .B1(n22781), .X(
        n22798) );
  sky130_fd_sc_hd__nand2_1 U28065 ( .A(n22782), .B(n22831), .Y(n22794) );
  sky130_fd_sc_hd__nor2_1 U28066 ( .A(n22786), .B(n22783), .Y(n22788) );
  sky130_fd_sc_hd__nand2_1 U28067 ( .A(n22017), .B(n22788), .Y(n22830) );
  sky130_fd_sc_hd__nand2_1 U28068 ( .A(n23030), .B(n22790), .Y(n22792) );
  sky130_fd_sc_hd__o21ai_1 U28069 ( .A1(n22786), .A2(n22785), .B1(n22784), .Y(
        n22787) );
  sky130_fd_sc_hd__a21oi_1 U28070 ( .A1(n22789), .A2(n22788), .B1(n22787), .Y(
        n22832) );
  sky130_fd_sc_hd__a21boi_1 U28071 ( .A1(n23036), .A2(n22790), .B1_N(n22832), 
        .Y(n22791) );
  sky130_fd_sc_hd__o21ai_1 U28072 ( .A1(n22792), .A2(n12349), .B1(n22791), .Y(
        n22793) );
  sky130_fd_sc_hd__xnor2_1 U28073 ( .A(n22794), .B(n22793), .Y(n23463) );
  sky130_fd_sc_hd__nand2_1 U28074 ( .A(n24853), .B(n24452), .Y(n22796) );
  sky130_fd_sc_hd__nand2_1 U28075 ( .A(n24855), .B(n22940), .Y(n22795) );
  sky130_fd_sc_hd__nand2b_1 U28076 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[16]), .Y(n24836) );
  sky130_fd_sc_hd__nand3_1 U28077 ( .A(n22796), .B(n22795), .C(n24836), .Y(
        n24828) );
  sky130_fd_sc_hd__nand2_1 U28078 ( .A(n24828), .B(n23044), .Y(n22797) );
  sky130_fd_sc_hd__nand3_1 U28079 ( .A(n11443), .B(n22798), .C(n22797), .Y(
        n29503) );
  sky130_fd_sc_hd__nand2_1 U28080 ( .A(n22801), .B(n22800), .Y(n22809) );
  sky130_fd_sc_hd__nand2_1 U28081 ( .A(n23030), .B(n22805), .Y(n22807) );
  sky130_fd_sc_hd__inv_1 U28082 ( .A(n22803), .Y(n22804) );
  sky130_fd_sc_hd__a21oi_1 U28083 ( .A1(n23036), .A2(n22805), .B1(n22804), .Y(
        n22806) );
  sky130_fd_sc_hd__xnor2_1 U28084 ( .A(n22809), .B(n22808), .Y(n22810) );
  sky130_fd_sc_hd__nand2_1 U28085 ( .A(n22810), .B(n24452), .Y(n25676) );
  sky130_fd_sc_hd__nand2_1 U28086 ( .A(n28056), .B(n22811), .Y(n25680) );
  sky130_fd_sc_hd__nand2b_1 U28087 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[19]), .Y(n25681) );
  sky130_fd_sc_hd__a21oi_1 U28088 ( .A1(n23485), .A2(n22940), .B1(n22812), .Y(
        n25718) );
  sky130_fd_sc_hd__nand2_1 U28089 ( .A(n27768), .B(n22811), .Y(n22814) );
  sky130_fd_sc_hd__nand2_1 U28090 ( .A(n24329), .B(n22979), .Y(n22813) );
  sky130_fd_sc_hd__o211ai_1 U28091 ( .A1(n22980), .A2(n22815), .B1(n22814), 
        .C1(n22813), .Y(n22816) );
  sky130_fd_sc_hd__a21oi_1 U28092 ( .A1(n22817), .A2(n24764), .B1(n22816), .Y(
        n25677) );
  sky130_fd_sc_hd__a22oi_1 U28093 ( .A1(n23009), .A2(
        j202_soc_core_j22_cpu_rf_tmp[19]), .B1(n23008), .B2(
        j202_soc_core_j22_cpu_rf_vbr[19]), .Y(n22822) );
  sky130_fd_sc_hd__a22oi_1 U28094 ( .A1(n23006), .A2(
        j202_soc_core_j22_cpu_rf_pr[19]), .B1(n23005), .B2(
        j202_soc_core_j22_cpu_rf_gpr[498]), .Y(n22821) );
  sky130_fd_sc_hd__o22a_1 U28095 ( .A1(n15484), .A2(n23000), .B1(n22818), .B2(
        n22998), .X(n22820) );
  sky130_fd_sc_hd__nand2_1 U28096 ( .A(n23003), .B(
        j202_soc_core_j22_cpu_rf_gpr[19]), .Y(n22819) );
  sky130_fd_sc_hd__nand4_1 U28097 ( .A(n22822), .B(n22821), .C(n22820), .D(
        n22819), .Y(n22823) );
  sky130_fd_sc_hd__a21oi_1 U28098 ( .A1(n23010), .A2(n22824), .B1(n22823), .Y(
        n22827) );
  sky130_fd_sc_hd__nand2_1 U28099 ( .A(n22829), .B(n22828), .Y(n22839) );
  sky130_fd_sc_hd__nor2_1 U28100 ( .A(n22833), .B(n22830), .Y(n22835) );
  sky130_fd_sc_hd__nand2_1 U28101 ( .A(n23030), .B(n22835), .Y(n22837) );
  sky130_fd_sc_hd__o21ai_1 U28102 ( .A1(n22833), .A2(n22832), .B1(n22831), .Y(
        n22834) );
  sky130_fd_sc_hd__a21oi_1 U28103 ( .A1(n23036), .A2(n22835), .B1(n22834), .Y(
        n22836) );
  sky130_fd_sc_hd__xnor2_1 U28104 ( .A(n22839), .B(n22838), .Y(n22840) );
  sky130_fd_sc_hd__nand2_1 U28105 ( .A(n22840), .B(n24452), .Y(n22842) );
  sky130_fd_sc_hd__nand2_1 U28106 ( .A(n23041), .B(
        j202_soc_core_j22_cpu_ml_mach[17]), .Y(n22841) );
  sky130_fd_sc_hd__nand2_1 U28107 ( .A(n22842), .B(n22841), .Y(n22843) );
  sky130_fd_sc_hd__a21oi_2 U28108 ( .A1(n23479), .A2(n25679), .B1(n22843), .Y(
        n25763) );
  sky130_fd_sc_hd__o22ai_1 U28109 ( .A1(n17785), .A2(n22845), .B1(n22844), 
        .B2(n22980), .Y(n22846) );
  sky130_fd_sc_hd__a21oi_1 U28110 ( .A1(n24320), .A2(n22979), .B1(n22846), .Y(
        n22847) );
  sky130_fd_sc_hd__a2bb2oi_1 U28111 ( .B1(j202_soc_core_j22_cpu_rf_tmp[17]), 
        .B2(n23009), .A1_N(n22849), .A2_N(n23000), .Y(n22854) );
  sky130_fd_sc_hd__nand2_1 U28112 ( .A(n23006), .B(
        j202_soc_core_j22_cpu_rf_pr[17]), .Y(n22853) );
  sky130_fd_sc_hd__nand2_1 U28113 ( .A(n23008), .B(
        j202_soc_core_j22_cpu_rf_vbr[17]), .Y(n22852) );
  sky130_fd_sc_hd__nor2_1 U28114 ( .A(n17785), .B(n22850), .Y(n25294) );
  sky130_fd_sc_hd__nand2_1 U28115 ( .A(n25294), .B(n27717), .Y(n22851) );
  sky130_fd_sc_hd__nand4_1 U28116 ( .A(n22854), .B(n22853), .C(n22852), .D(
        n22851), .Y(n22860) );
  sky130_fd_sc_hd__nand2_1 U28117 ( .A(n22855), .B(n23010), .Y(n22859) );
  sky130_fd_sc_hd__a2bb2oi_1 U28118 ( .B1(n23005), .B2(
        j202_soc_core_j22_cpu_rf_gpr[496]), .A1_N(n22856), .A2_N(n22998), .Y(
        n22858) );
  sky130_fd_sc_hd__nand2_1 U28119 ( .A(n23003), .B(
        j202_soc_core_j22_cpu_rf_gpr[17]), .Y(n22857) );
  sky130_fd_sc_hd__nand4b_1 U28120 ( .A_N(n22860), .B(n22859), .C(n22858), .D(
        n22857), .Y(n22861) );
  sky130_fd_sc_hd__a21oi_1 U28121 ( .A1(n22866), .A2(n22862), .B1(n22861), .Y(
        n22863) );
  sky130_fd_sc_hd__o21a_1 U28122 ( .A1(n23018), .A2(n25307), .B1(n22863), .X(
        n22864) );
  sky130_fd_sc_hd__nand2_1 U28123 ( .A(n22866), .B(n22950), .Y(n22867) );
  sky130_fd_sc_hd__nand2_1 U28124 ( .A(n22871), .B(n22870), .Y(n22879) );
  sky130_fd_sc_hd__nand2_1 U28125 ( .A(n11403), .B(n22875), .Y(n22877) );
  sky130_fd_sc_hd__a21oi_1 U28126 ( .A1(n22875), .A2(n21753), .B1(n22874), .Y(
        n22876) );
  sky130_fd_sc_hd__o21ai_1 U28127 ( .A1(n22877), .A2(n22967), .B1(n22876), .Y(
        n22878) );
  sky130_fd_sc_hd__xnor2_1 U28128 ( .A(n22879), .B(n22878), .Y(n22941) );
  sky130_fd_sc_hd__nand2_1 U28129 ( .A(n22882), .B(n22881), .Y(n22887) );
  sky130_fd_sc_hd__o21ai_1 U28130 ( .A1(n22885), .A2(n22884), .B1(n22883), .Y(
        n22886) );
  sky130_fd_sc_hd__xnor2_1 U28131 ( .A(n22887), .B(n22886), .Y(n24333) );
  sky130_fd_sc_hd__nand2_1 U28132 ( .A(n24333), .B(n22979), .Y(n22888) );
  sky130_fd_sc_hd__o21ai_0 U28133 ( .A1(n22980), .A2(n22889), .B1(n22888), .Y(
        n22890) );
  sky130_fd_sc_hd__a21oi_1 U28134 ( .A1(n22941), .A2(n24764), .B1(n22890), .Y(
        n25262) );
  sky130_fd_sc_hd__o22ai_1 U28135 ( .A1(n22892), .A2(n22983), .B1(n22982), 
        .B2(n22891), .Y(n22893) );
  sky130_fd_sc_hd__a21oi_1 U28136 ( .A1(n22990), .A2(
        j202_soc_core_j22_cpu_rf_vbr[9]), .B1(n22893), .Y(n22901) );
  sky130_fd_sc_hd__a22oi_1 U28137 ( .A1(n22988), .A2(
        j202_soc_core_j22_cpu_pc[9]), .B1(n22987), .B2(
        j202_soc_core_j22_cpu_rf_gbr[9]), .Y(n22900) );
  sky130_fd_sc_hd__o22a_1 U28138 ( .A1(n22897), .A2(n22896), .B1(n22895), .B2(
        n22894), .X(n22899) );
  sky130_fd_sc_hd__nand2_1 U28139 ( .A(n22986), .B(
        j202_soc_core_j22_cpu_rf_gpr[9]), .Y(n22898) );
  sky130_fd_sc_hd__nand4_1 U28140 ( .A(n22901), .B(n22900), .C(n22899), .D(
        n22898), .Y(n22902) );
  sky130_fd_sc_hd__a21o_1 U28141 ( .A1(n22903), .A2(n22996), .B1(n22902), .X(
        n22946) );
  sky130_fd_sc_hd__o22ai_1 U28142 ( .A1(n22905), .A2(n23000), .B1(n22904), 
        .B2(n22998), .Y(n22906) );
  sky130_fd_sc_hd__a21oi_1 U28143 ( .A1(j202_soc_core_j22_cpu_rf_gpr[25]), 
        .A2(n23003), .B1(n22906), .Y(n22912) );
  sky130_fd_sc_hd__nand2_1 U28144 ( .A(n23004), .B(n23567), .Y(n25261) );
  sky130_fd_sc_hd__a22oi_1 U28145 ( .A1(n23006), .A2(
        j202_soc_core_j22_cpu_rf_pr[25]), .B1(n23005), .B2(
        j202_soc_core_j22_cpu_rf_gpr[504]), .Y(n22907) );
  sky130_fd_sc_hd__o21a_1 U28146 ( .A1(n24467), .A2(n25261), .B1(n22907), .X(
        n22911) );
  sky130_fd_sc_hd__a22oi_1 U28147 ( .A1(n23009), .A2(
        j202_soc_core_j22_cpu_rf_tmp[25]), .B1(n23008), .B2(
        j202_soc_core_j22_cpu_rf_vbr[25]), .Y(n22910) );
  sky130_fd_sc_hd__nand2_1 U28148 ( .A(n22908), .B(n23010), .Y(n22909) );
  sky130_fd_sc_hd__nand4_1 U28149 ( .A(n22912), .B(n22911), .C(n22910), .D(
        n22909), .Y(n22913) );
  sky130_fd_sc_hd__a21oi_1 U28150 ( .A1(n22946), .A2(n23973), .B1(n22913), .Y(
        n22914) );
  sky130_fd_sc_hd__o21a_1 U28151 ( .A1(n23018), .A2(n25262), .B1(n22914), .X(
        n22939) );
  sky130_fd_sc_hd__nand2_1 U28153 ( .A(n22917), .B(n22916), .Y(n22927) );
  sky130_fd_sc_hd__nor2_1 U28154 ( .A(n22920), .B(n22918), .Y(n22923) );
  sky130_fd_sc_hd__o21ai_2 U28156 ( .A1(n22925), .A2(n11866), .B1(n22924), .Y(
        n22926) );
  sky130_fd_sc_hd__xnor2_2 U28157 ( .A(n22927), .B(n22926), .Y(n23483) );
  sky130_fd_sc_hd__nand2_1 U28158 ( .A(n22929), .B(n22928), .Y(n22936) );
  sky130_fd_sc_hd__inv_1 U28159 ( .A(n22930), .Y(n22932) );
  sky130_fd_sc_hd__nand2_1 U28160 ( .A(n23030), .B(n22932), .Y(n22934) );
  sky130_fd_sc_hd__a21oi_1 U28161 ( .A1(n23036), .A2(n22932), .B1(n22931), .Y(
        n22933) );
  sky130_fd_sc_hd__xnor2_1 U28162 ( .A(n22936), .B(n22935), .Y(n22937) );
  sky130_fd_sc_hd__nand2b_1 U28163 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[25]), .Y(n25255) );
  sky130_fd_sc_hd__nand3_1 U28164 ( .A(n25260), .B(n25259), .C(n25255), .Y(
        n23566) );
  sky130_fd_sc_hd__nand2_1 U28165 ( .A(n23566), .B(n23044), .Y(n22938) );
  sky130_fd_sc_hd__nand3_2 U28166 ( .A(n22949), .B(n22939), .C(n22938), .Y(
        n29513) );
  sky130_fd_sc_hd__nand2_1 U28167 ( .A(n22941), .B(n22940), .Y(n24797) );
  sky130_fd_sc_hd__nand2b_1 U28168 ( .A_N(n28045), .B(
        j202_soc_core_j22_cpu_ml_mach[9]), .Y(n24796) );
  sky130_fd_sc_hd__nand2_1 U28169 ( .A(n23004), .B(n12050), .Y(n24874) );
  sky130_fd_sc_hd__nand4_1 U28170 ( .A(n24798), .B(n24797), .C(n24796), .D(
        n24874), .Y(n22943) );
  sky130_fd_sc_hd__nand2_1 U28171 ( .A(n24874), .B(n27052), .Y(n22942) );
  sky130_fd_sc_hd__nand2_1 U28172 ( .A(n22943), .B(n22942), .Y(n22944) );
  sky130_fd_sc_hd__nand2_1 U28173 ( .A(n24333), .B(n24461), .Y(n24898) );
  sky130_fd_sc_hd__nand2b_1 U28174 ( .A_N(n24463), .B(
        j202_soc_core_j22_cpu_ml_macl[9]), .Y(n24876) );
  sky130_fd_sc_hd__nand3_1 U28175 ( .A(n22944), .B(n24898), .C(n24876), .Y(
        n22945) );
  sky130_fd_sc_hd__nand2_1 U28176 ( .A(n22945), .B(n27717), .Y(n22948) );
  sky130_fd_sc_hd__nand2_1 U28177 ( .A(n22946), .B(n24450), .Y(n22947) );
  sky130_fd_sc_hd__nand3_2 U28178 ( .A(n22949), .B(n22948), .C(n22947), .Y(
        n29527) );
  sky130_fd_sc_hd__nand2_1 U28179 ( .A(n22951), .B(n22950), .Y(n22952) );
  sky130_fd_sc_hd__nand2_1 U28182 ( .A(n22955), .B(n22954), .Y(n22970) );
  sky130_fd_sc_hd__nor2_1 U28183 ( .A(n11471), .B(n22957), .Y(n22964) );
  sky130_fd_sc_hd__nand2_1 U28184 ( .A(n22964), .B(n22958), .Y(n22968) );
  sky130_fd_sc_hd__a21oi_1 U28186 ( .A1(n22965), .A2(n22964), .B1(n22963), .Y(
        n22966) );
  sky130_fd_sc_hd__xnor2_1 U28188 ( .A(n22970), .B(n22969), .Y(n25442) );
  sky130_fd_sc_hd__inv_1 U28189 ( .A(n22971), .Y(n22973) );
  sky130_fd_sc_hd__nand2_1 U28190 ( .A(n22973), .B(n22972), .Y(n22978) );
  sky130_fd_sc_hd__o21ai_1 U28191 ( .A1(n22976), .A2(n22975), .B1(n22974), .Y(
        n22977) );
  sky130_fd_sc_hd__xnor2_1 U28192 ( .A(n22978), .B(n22977), .Y(n24444) );
  sky130_fd_sc_hd__nand2_1 U28193 ( .A(n24444), .B(n22979), .Y(n25440) );
  sky130_fd_sc_hd__nand2b_1 U28194 ( .A_N(n22980), .B(
        j202_soc_core_j22_cpu_ml_macl[29]), .Y(n25438) );
  sky130_fd_sc_hd__nand2_1 U28195 ( .A(n25440), .B(n25438), .Y(n25443) );
  sky130_fd_sc_hd__a21oi_1 U28196 ( .A1(n25442), .A2(n24764), .B1(n25443), .Y(
        n25391) );
  sky130_fd_sc_hd__o22ai_1 U28197 ( .A1(n22984), .A2(n22983), .B1(n22982), 
        .B2(n22981), .Y(n22985) );
  sky130_fd_sc_hd__a21oi_1 U28198 ( .A1(n22986), .A2(
        j202_soc_core_j22_cpu_rf_gpr[13]), .B1(n22985), .Y(n22994) );
  sky130_fd_sc_hd__a22oi_1 U28199 ( .A1(n22988), .A2(
        j202_soc_core_j22_cpu_pc[13]), .B1(n22987), .B2(
        j202_soc_core_j22_cpu_rf_gbr[13]), .Y(n22993) );
  sky130_fd_sc_hd__nand2_1 U28200 ( .A(n22989), .B(
        j202_soc_core_j22_cpu_rf_tmp[13]), .Y(n22992) );
  sky130_fd_sc_hd__nand2_1 U28201 ( .A(n22990), .B(
        j202_soc_core_j22_cpu_rf_vbr[13]), .Y(n22991) );
  sky130_fd_sc_hd__nand4_1 U28202 ( .A(n22994), .B(n22993), .C(n22992), .D(
        n22991), .Y(n22995) );
  sky130_fd_sc_hd__a21o_1 U28203 ( .A1(n22997), .A2(n22996), .B1(n22995), .X(
        n24438) );
  sky130_fd_sc_hd__o22ai_1 U28204 ( .A1(n23001), .A2(n23000), .B1(n22999), 
        .B2(n22998), .Y(n23002) );
  sky130_fd_sc_hd__a21oi_1 U28205 ( .A1(j202_soc_core_j22_cpu_rf_gpr[29]), 
        .A2(n23003), .B1(n23002), .Y(n23015) );
  sky130_fd_sc_hd__nand2_1 U28206 ( .A(n23004), .B(n25389), .Y(n25444) );
  sky130_fd_sc_hd__a22oi_1 U28207 ( .A1(n23006), .A2(
        j202_soc_core_j22_cpu_rf_pr[29]), .B1(n23005), .B2(
        j202_soc_core_j22_cpu_rf_gpr[508]), .Y(n23007) );
  sky130_fd_sc_hd__o21a_1 U28208 ( .A1(n24467), .A2(n25444), .B1(n23007), .X(
        n23014) );
  sky130_fd_sc_hd__a22oi_1 U28209 ( .A1(n23009), .A2(
        j202_soc_core_j22_cpu_rf_tmp[29]), .B1(n23008), .B2(
        j202_soc_core_j22_cpu_rf_vbr[29]), .Y(n23013) );
  sky130_fd_sc_hd__nand2_1 U28210 ( .A(n23011), .B(n23010), .Y(n23012) );
  sky130_fd_sc_hd__nand4_1 U28211 ( .A(n23015), .B(n23014), .C(n23013), .D(
        n23012), .Y(n23016) );
  sky130_fd_sc_hd__a21oi_1 U28212 ( .A1(n24438), .A2(n23973), .B1(n23016), .Y(
        n23017) );
  sky130_fd_sc_hd__nand2_1 U28213 ( .A(n23020), .B(n23019), .Y(n23025) );
  sky130_fd_sc_hd__nand2_1 U28214 ( .A(n23030), .B(n22017), .Y(n23023) );
  sky130_fd_sc_hd__nand2_1 U28215 ( .A(n24439), .B(n25679), .Y(n23043) );
  sky130_fd_sc_hd__nand2_1 U28216 ( .A(n23028), .B(n23027), .Y(n23039) );
  sky130_fd_sc_hd__nor2_1 U28217 ( .A(n23033), .B(n23029), .Y(n23035) );
  sky130_fd_sc_hd__o21ai_1 U28218 ( .A1(n23033), .A2(n23032), .B1(n23031), .Y(
        n23034) );
  sky130_fd_sc_hd__a21oi_1 U28219 ( .A1(n23036), .A2(n23035), .B1(n23034), .Y(
        n23037) );
  sky130_fd_sc_hd__xnor2_1 U28220 ( .A(n23039), .B(n23038), .Y(n23040) );
  sky130_fd_sc_hd__nand2_1 U28221 ( .A(n25464), .B(n23044), .Y(n23045) );
  sky130_fd_sc_hd__nor2_1 U28222 ( .A(j202_soc_core_uart_BRG_sio_ce_x4_r), .B(
        n28624), .Y(n29601) );
  sky130_fd_sc_hd__nand2_1 U28223 ( .A(j202_soc_core_uart_TOP_dpll_state[0]), 
        .B(n23047), .Y(n29096) );
  sky130_fd_sc_hd__nand2_1 U28224 ( .A(n29601), .B(n29827), .Y(n28598) );
  sky130_fd_sc_hd__nor2_1 U28225 ( .A(j202_soc_core_uart_BRG_cnt[0]), .B(
        n28598), .Y(n29602) );
  sky130_fd_sc_hd__nor2_1 U28226 ( .A(j202_soc_core_uart_BRG_cnt[1]), .B(
        j202_soc_core_uart_BRG_cnt[0]), .Y(n29609) );
  sky130_fd_sc_hd__nand2_1 U28227 ( .A(j202_soc_core_uart_sio_ce), .B(
        j202_soc_core_uart_TOP_shift_en), .Y(n24518) );
  sky130_fd_sc_hd__nor2_1 U28228 ( .A(n29088), .B(n24518), .Y(n29494) );
  sky130_fd_sc_hd__nand2_1 U28229 ( .A(n29474), .B(n29473), .Y(n23057) );
  sky130_fd_sc_hd__nor2_1 U28230 ( .A(n23057), .B(n23051), .Y(n29529) );
  sky130_fd_sc_hd__nand2b_1 U28231 ( .A_N(n29473), .B(n29474), .Y(n23621) );
  sky130_fd_sc_hd__nand3_1 U28232 ( .A(n23049), .B(n29547), .C(n29549), .Y(
        n23054) );
  sky130_fd_sc_hd__nor2_1 U28233 ( .A(n23621), .B(n23054), .Y(n29536) );
  sky130_fd_sc_hd__nand3_1 U28234 ( .A(n23049), .B(n25052), .C(n29547), .Y(
        n23055) );
  sky130_fd_sc_hd__nor2_1 U28235 ( .A(n23621), .B(n23055), .Y(n29535) );
  sky130_fd_sc_hd__nand3_1 U28236 ( .A(n23049), .B(n23048), .C(n29549), .Y(
        n23056) );
  sky130_fd_sc_hd__nor2_1 U28237 ( .A(n23621), .B(n23056), .Y(n29596) );
  sky130_fd_sc_hd__nor2_1 U28238 ( .A(n23621), .B(n23051), .Y(n29528) );
  sky130_fd_sc_hd__nand2_1 U28239 ( .A(j202_soc_core_qspi_wb_wdat[31]), .B(
        n29745), .Y(n27601) );
  sky130_fd_sc_hd__nand2_1 U28240 ( .A(j202_soc_core_qspi_wb_wdat[30]), .B(
        n29745), .Y(n28002) );
  sky130_fd_sc_hd__nand2_1 U28241 ( .A(j202_soc_core_qspi_wb_wdat[29]), .B(
        n12069), .Y(n25494) );
  sky130_fd_sc_hd__nand2_1 U28242 ( .A(j202_soc_core_qspi_wb_wdat[28]), .B(
        n12069), .Y(n27395) );
  sky130_fd_sc_hd__nand2_1 U28243 ( .A(j202_soc_core_qspi_wb_wdat[27]), .B(
        n29830), .Y(n27078) );
  sky130_fd_sc_hd__nand2_1 U28244 ( .A(j202_soc_core_qspi_wb_wdat[26]), .B(
        n29828), .Y(n27875) );
  sky130_fd_sc_hd__nand2_1 U28245 ( .A(j202_soc_core_qspi_wb_wdat[25]), .B(
        n12069), .Y(n27172) );
  sky130_fd_sc_hd__nand2_1 U28246 ( .A(j202_soc_core_qspi_wb_wdat[24]), .B(
        n29745), .Y(n27655) );
  sky130_fd_sc_hd__nand2_1 U28247 ( .A(j202_soc_core_qspi_wb_wdat[23]), .B(
        n29745), .Y(n27633) );
  sky130_fd_sc_hd__nand2_1 U28248 ( .A(j202_soc_core_qspi_wb_wdat[22]), .B(
        n12069), .Y(n25614) );
  sky130_fd_sc_hd__nand2_1 U28249 ( .A(j202_soc_core_qspi_wb_wdat[21]), .B(
        n12069), .Y(n25582) );
  sky130_fd_sc_hd__nand2_1 U28250 ( .A(j202_soc_core_qspi_wb_wdat[20]), .B(
        n29745), .Y(n29152) );
  sky130_fd_sc_hd__nand2_1 U28251 ( .A(j202_soc_core_qspi_wb_wdat[19]), .B(
        n29827), .Y(n29150) );
  sky130_fd_sc_hd__nand2_1 U28252 ( .A(j202_soc_core_qspi_wb_wdat[18]), .B(
        n29745), .Y(n29153) );
  sky130_fd_sc_hd__nand2_1 U28253 ( .A(j202_soc_core_qspi_wb_wdat[17]), .B(
        n29745), .Y(n29149) );
  sky130_fd_sc_hd__nand2_1 U28254 ( .A(j202_soc_core_qspi_wb_wdat[16]), .B(
        n29745), .Y(n29151) );
  sky130_fd_sc_hd__nand2_1 U28255 ( .A(j202_soc_core_qspi_wb_wdat[9]), .B(
        n29745), .Y(n29148) );
  sky130_fd_sc_hd__nand2_1 U28256 ( .A(j202_soc_core_qspi_wb_wdat[8]), .B(
        n29745), .Y(n29146) );
  sky130_fd_sc_hd__nand2_1 U28257 ( .A(j202_soc_core_qspi_wb_wdat[7]), .B(
        n12069), .Y(n29157) );
  sky130_fd_sc_hd__nand2_1 U28258 ( .A(j202_soc_core_qspi_wb_wdat[6]), .B(
        n29745), .Y(n29158) );
  sky130_fd_sc_hd__nand2_1 U28259 ( .A(j202_soc_core_qspi_wb_wdat[5]), .B(
        n12069), .Y(n29159) );
  sky130_fd_sc_hd__nand2_1 U28260 ( .A(j202_soc_core_qspi_wb_wdat[4]), .B(
        n29745), .Y(n29160) );
  sky130_fd_sc_hd__nand2_1 U28261 ( .A(j202_soc_core_qspi_wb_wdat[3]), .B(
        n29827), .Y(n29161) );
  sky130_fd_sc_hd__nand2_1 U28262 ( .A(j202_soc_core_qspi_wb_wdat[2]), .B(
        n29828), .Y(n29162) );
  sky130_fd_sc_hd__nand2_1 U28263 ( .A(j202_soc_core_qspi_wb_wdat[1]), .B(
        n29827), .Y(n29163) );
  sky130_fd_sc_hd__nand2_1 U28264 ( .A(j202_soc_core_qspi_wb_wdat[0]), .B(
        n29745), .Y(n29165) );
  sky130_fd_sc_hd__nor2_1 U28265 ( .A(n29474), .B(n23050), .Y(n23560) );
  sky130_fd_sc_hd__nor2_1 U28266 ( .A(n23052), .B(n23054), .Y(n29538) );
  sky130_fd_sc_hd__nor2_1 U28267 ( .A(n23052), .B(n23055), .Y(n29591) );
  sky130_fd_sc_hd__nor2_1 U28268 ( .A(n23052), .B(n23056), .Y(n29531) );
  sky130_fd_sc_hd__nor2_1 U28269 ( .A(n23052), .B(n23051), .Y(n29592) );
  sky130_fd_sc_hd__nor2_1 U28270 ( .A(n23053), .B(n23054), .Y(n29600) );
  sky130_fd_sc_hd__nor2_1 U28271 ( .A(n23053), .B(n23055), .Y(n29539) );
  sky130_fd_sc_hd__nor2_1 U28272 ( .A(n23053), .B(n23056), .Y(n29533) );
  sky130_fd_sc_hd__nand2_1 U28273 ( .A(j202_soc_core_qspi_wb_wdat[12]), .B(
        n12069), .Y(n29147) );
  sky130_fd_sc_hd__nand2_1 U28274 ( .A(j202_soc_core_qspi_wb_wdat[13]), .B(
        n29827), .Y(n29145) );
  sky130_fd_sc_hd__nand2_1 U28275 ( .A(j202_soc_core_qspi_wb_wdat[14]), .B(
        n29827), .Y(n29144) );
  sky130_fd_sc_hd__nor2_1 U28276 ( .A(n23057), .B(n23054), .Y(n29534) );
  sky130_fd_sc_hd__nor2_1 U28277 ( .A(n23057), .B(n23055), .Y(n29537) );
  sky130_fd_sc_hd__nor2_1 U28278 ( .A(n23057), .B(n23056), .Y(n29530) );
  sky130_fd_sc_hd__nor3_1 U28279 ( .A(j202_soc_core_bldc_core_00_comm[2]), .B(
        n29117), .C(n29121), .Y(n29608) );
  sky130_fd_sc_hd__nand2_1 U28280 ( .A(n26736), .B(
        j202_soc_core_intc_core_00_rg_ipr[54]), .Y(n23059) );
  sky130_fd_sc_hd__o2bb2ai_1 U28281 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[52]), .B2(n26739), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[49]), .A2_N(n25576), .Y(n23058) );
  sky130_fd_sc_hd__o211ai_1 U28282 ( .A1(j202_soc_core_intc_core_00_rg_ipr[49]), .A2(n25576), .B1(n23059), .C1(n23058), .Y(n23061) );
  sky130_fd_sc_hd__a2bb2oi_1 U28283 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[51]), .B2(n26740), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[54]), .A2_N(n26736), .Y(n23060) );
  sky130_fd_sc_hd__nand2_1 U28284 ( .A(n23061), .B(n23060), .Y(n23064) );
  sky130_fd_sc_hd__a21oi_1 U28285 ( .A1(n25323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[55]), .B1(n23062), .Y(n23063) );
  sky130_fd_sc_hd__nand2_1 U28286 ( .A(n23064), .B(n23063), .Y(n23067) );
  sky130_fd_sc_hd__nand2_1 U28287 ( .A(n23067), .B(n23066), .Y(n23076) );
  sky130_fd_sc_hd__nand2_1 U28288 ( .A(n26742), .B(
        j202_soc_core_intc_core_00_rg_ipr[62]), .Y(n23069) );
  sky130_fd_sc_hd__o2bb2ai_1 U28289 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[60]), .B2(n26755), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[57]), .A2_N(n25488), .Y(n23068) );
  sky130_fd_sc_hd__o211ai_1 U28290 ( .A1(j202_soc_core_intc_core_00_rg_ipr[57]), .A2(n25488), .B1(n23069), .C1(n23068), .Y(n23071) );
  sky130_fd_sc_hd__a2bb2oi_1 U28291 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[59]), .B2(n26759), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[62]), .A2_N(n26742), .Y(n23070) );
  sky130_fd_sc_hd__nand2_1 U28292 ( .A(n23071), .B(n23070), .Y(n23075) );
  sky130_fd_sc_hd__a21oi_1 U28293 ( .A1(n26757), .A2(
        j202_soc_core_intc_core_00_rg_ipr[63]), .B1(n23072), .Y(n23074) );
  sky130_fd_sc_hd__inv_2 U28294 ( .A(n27325), .Y(n23080) );
  sky130_fd_sc_hd__mux2i_1 U28295 ( .A0(j202_soc_core_intc_core_00_rg_ipr[62]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[58]), .S(n23080), .Y(n23077) );
  sky130_fd_sc_hd__mux2_2 U28296 ( .A0(j202_soc_core_intc_core_00_rg_ipr[51]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[55]), .S(n27328), .X(n23142) );
  sky130_fd_sc_hd__mux2_2 U28297 ( .A0(j202_soc_core_intc_core_00_rg_ipr[57]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[61]), .S(n27325), .X(n23125) );
  sky130_fd_sc_hd__mux2i_1 U28298 ( .A0(j202_soc_core_intc_core_00_rg_ipr[53]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[49]), .S(n23076), .Y(n23124) );
  sky130_fd_sc_hd__mux2i_1 U28299 ( .A0(j202_soc_core_intc_core_00_rg_ipr[60]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[56]), .S(n23080), .Y(n23134) );
  sky130_fd_sc_hd__nand2_1 U28300 ( .A(n23085), .B(n23077), .Y(n23078) );
  sky130_fd_sc_hd__nand2_1 U28301 ( .A(n23079), .B(n23078), .Y(n23081) );
  sky130_fd_sc_hd__mux2i_1 U28302 ( .A0(j202_soc_core_intc_core_00_rg_ipr[63]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[59]), .S(n23080), .Y(n23143) );
  sky130_fd_sc_hd__o21ai_1 U28303 ( .A1(n23142), .A2(n23081), .B1(n23143), .Y(
        n23083) );
  sky130_fd_sc_hd__nand2_1 U28304 ( .A(n23081), .B(n23142), .Y(n23082) );
  sky130_fd_sc_hd__nand3_1 U28305 ( .A(n23083), .B(n23275), .C(n23082), .Y(
        n27327) );
  sky130_fd_sc_hd__nand2_1 U28306 ( .A(n27327), .B(n23141), .Y(n27326) );
  sky130_fd_sc_hd__mux2_2 U28307 ( .A0(n23085), .A1(n23084), .S(n27326), .X(
        n23150) );
  sky130_fd_sc_hd__nand2_1 U28308 ( .A(n26711), .B(
        j202_soc_core_intc_core_00_rg_ipr[38]), .Y(n23087) );
  sky130_fd_sc_hd__o2bb2ai_1 U28309 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[36]), .B2(n26727), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[33]), .A2_N(n26726), .Y(n23086) );
  sky130_fd_sc_hd__o211ai_1 U28310 ( .A1(j202_soc_core_intc_core_00_rg_ipr[33]), .A2(n26726), .B1(n23087), .C1(n23086), .Y(n23089) );
  sky130_fd_sc_hd__nand2_1 U28311 ( .A(n23089), .B(n23088), .Y(n23092) );
  sky130_fd_sc_hd__a21oi_1 U28312 ( .A1(n26729), .A2(
        j202_soc_core_intc_core_00_rg_ipr[39]), .B1(n23090), .Y(n23091) );
  sky130_fd_sc_hd__nand2_1 U28313 ( .A(n23092), .B(n23091), .Y(n23095) );
  sky130_fd_sc_hd__mux2i_1 U28314 ( .A0(j202_soc_core_intc_core_00_rg_ipr[38]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[34]), .S(n23104), .Y(n23120) );
  sky130_fd_sc_hd__nand2_1 U28315 ( .A(n25070), .B(
        j202_soc_core_intc_core_00_rg_ipr[46]), .Y(n23097) );
  sky130_fd_sc_hd__o2bb2ai_1 U28316 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[44]), .B2(n26734), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[41]), .A2_N(n25790), .Y(n23096) );
  sky130_fd_sc_hd__o211ai_1 U28317 ( .A1(j202_soc_core_intc_core_00_rg_ipr[41]), .A2(n25790), .B1(n23097), .C1(n23096), .Y(n23099) );
  sky130_fd_sc_hd__a2bb2oi_1 U28318 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[43]), .B2(n26122), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[46]), .A2_N(n25070), .Y(n23098) );
  sky130_fd_sc_hd__nand2_1 U28319 ( .A(n23099), .B(n23098), .Y(n23103) );
  sky130_fd_sc_hd__a21oi_1 U28320 ( .A1(n26735), .A2(
        j202_soc_core_intc_core_00_rg_ipr[47]), .B1(n23100), .Y(n23102) );
  sky130_fd_sc_hd__mux2_2 U28321 ( .A0(j202_soc_core_intc_core_00_rg_ipr[42]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[46]), .S(n27329), .X(n23113) );
  sky130_fd_sc_hd__mux2_2 U28322 ( .A0(j202_soc_core_intc_core_00_rg_ipr[35]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[39]), .S(n27332), .X(n23123) );
  sky130_fd_sc_hd__nand2_1 U28323 ( .A(n23113), .B(n23120), .Y(n23112) );
  sky130_fd_sc_hd__mux2_2 U28324 ( .A0(j202_soc_core_intc_core_00_rg_ipr[41]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[45]), .S(n27329), .X(n23107) );
  sky130_fd_sc_hd__nand2_1 U28325 ( .A(n23107), .B(n23127), .Y(n23106) );
  sky130_fd_sc_hd__inv_1 U28326 ( .A(n27329), .Y(n23114) );
  sky130_fd_sc_hd__mux2i_1 U28327 ( .A0(j202_soc_core_intc_core_00_rg_ipr[44]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[40]), .S(n23114), .Y(n23131) );
  sky130_fd_sc_hd__mux2i_1 U28328 ( .A0(n26728), .A1(n26727), .S(n23104), .Y(
        n23105) );
  sky130_fd_sc_hd__nand3_1 U28329 ( .A(n23106), .B(n23131), .C(n23105), .Y(
        n23110) );
  sky130_fd_sc_hd__inv_1 U28330 ( .A(n23127), .Y(n23108) );
  sky130_fd_sc_hd__nand2_1 U28331 ( .A(n23108), .B(n23128), .Y(n23109) );
  sky130_fd_sc_hd__nand2_1 U28332 ( .A(n23110), .B(n23109), .Y(n23111) );
  sky130_fd_sc_hd__o2bb2ai_1 U28333 ( .B1(n23113), .B2(n23120), .A1_N(n23112), 
        .A2_N(n23111), .Y(n23115) );
  sky130_fd_sc_hd__mux2i_1 U28334 ( .A0(j202_soc_core_intc_core_00_rg_ipr[47]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[43]), .S(n23114), .Y(n23121) );
  sky130_fd_sc_hd__o21ai_1 U28335 ( .A1(n23123), .A2(n23115), .B1(n23121), .Y(
        n23118) );
  sky130_fd_sc_hd__nand2_1 U28336 ( .A(n23115), .B(n23123), .Y(n23116) );
  sky130_fd_sc_hd__nand3_1 U28337 ( .A(n23118), .B(n23117), .C(n23116), .Y(
        n27331) );
  sky130_fd_sc_hd__mux2_2 U28338 ( .A0(n23123), .A1(n23122), .S(n27330), .X(
        n23268) );
  sky130_fd_sc_hd__mux2_2 U28339 ( .A0(n23126), .A1(n23125), .S(n27326), .X(
        n23259) );
  sky130_fd_sc_hd__nand2_1 U28340 ( .A(n27330), .B(n23128), .Y(n23129) );
  sky130_fd_sc_hd__nand2_1 U28341 ( .A(n23130), .B(n23129), .Y(n23136) );
  sky130_fd_sc_hd__mux2i_1 U28342 ( .A0(j202_soc_core_intc_core_00_rg_ipr[36]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[32]), .S(n23104), .Y(n23132) );
  sky130_fd_sc_hd__mux2i_1 U28343 ( .A0(n23132), .A1(n23131), .S(n27330), .Y(
        n23254) );
  sky130_fd_sc_hd__nand2_1 U28344 ( .A(n23149), .B(n23138), .Y(n23139) );
  sky130_fd_sc_hd__nand2_1 U28345 ( .A(n23140), .B(n23139), .Y(n23145) );
  sky130_fd_sc_hd__o2bb2ai_1 U28346 ( .B1(n23141), .B2(n23275), .A1_N(n23268), 
        .A2_N(n23145), .Y(n23148) );
  sky130_fd_sc_hd__mux2_2 U28347 ( .A0(n23144), .A1(n23143), .S(n27326), .X(
        n23267) );
  sky130_fd_sc_hd__o21a_1 U28348 ( .A1(n23268), .A2(n23145), .B1(n23267), .X(
        n23147) );
  sky130_fd_sc_hd__o21a_2 U28349 ( .A1(n23148), .A2(n23147), .B1(n23146), .X(
        n27333) );
  sky130_fd_sc_hd__mux2i_1 U28350 ( .A0(n23150), .A1(n23149), .S(n27333), .Y(
        n23281) );
  sky130_fd_sc_hd__nand2_1 U28351 ( .A(n25071), .B(
        j202_soc_core_intc_core_00_rg_ipr[14]), .Y(n23152) );
  sky130_fd_sc_hd__o211ai_1 U28352 ( .A1(j202_soc_core_intc_core_00_rg_ipr[9]), 
        .A2(n25162), .B1(n23152), .C1(n23151), .Y(n23154) );
  sky130_fd_sc_hd__nand2_1 U28353 ( .A(n25155), .B(
        j202_soc_core_intc_core_00_rg_ipr[10]), .Y(n23153) );
  sky130_fd_sc_hd__nand2_1 U28354 ( .A(n23154), .B(n23153), .Y(n23156) );
  sky130_fd_sc_hd__nand2_1 U28355 ( .A(n26672), .B(
        j202_soc_core_intc_core_00_rg_ipr[15]), .Y(n23155) );
  sky130_fd_sc_hd__a21oi_1 U28356 ( .A1(n26123), .A2(
        j202_soc_core_intc_core_00_rg_ipr[11]), .B1(n23157), .Y(n23159) );
  sky130_fd_sc_hd__mux2_2 U28357 ( .A0(n25155), .A1(n25071), .S(n27315), .X(
        n23176) );
  sky130_fd_sc_hd__nand2_1 U28358 ( .A(n25154), .B(
        j202_soc_core_intc_core_00_rg_ipr[2]), .Y(n23163) );
  sky130_fd_sc_hd__nand2_1 U28359 ( .A(n24809), .B(
        j202_soc_core_intc_core_00_rg_ipr[5]), .Y(n23161) );
  sky130_fd_sc_hd__nand3_1 U28360 ( .A(n23161), .B(
        j202_soc_core_intc_core_00_rg_ipr[0]), .C(n24827), .Y(n23162) );
  sky130_fd_sc_hd__o211ai_1 U28361 ( .A1(j202_soc_core_intc_core_00_rg_ipr[5]), 
        .A2(n24809), .B1(n23163), .C1(n23162), .Y(n23165) );
  sky130_fd_sc_hd__a2bb2oi_1 U28362 ( .B1(j202_soc_core_intc_core_00_rg_ipr[7]), .B2(n27574), .A1_N(j202_soc_core_intc_core_00_rg_ipr[2]), .A2_N(n25154), .Y(
        n23164) );
  sky130_fd_sc_hd__nand2_1 U28363 ( .A(n23165), .B(n23164), .Y(n23168) );
  sky130_fd_sc_hd__a21oi_1 U28364 ( .A1(n27150), .A2(
        j202_soc_core_intc_core_00_rg_ipr[3]), .B1(n23166), .Y(n23167) );
  sky130_fd_sc_hd__nand2_1 U28365 ( .A(n23168), .B(n23167), .Y(n23171) );
  sky130_fd_sc_hd__mux2_2 U28366 ( .A0(j202_soc_core_intc_core_00_rg_ipr[6]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[2]), .S(n23172), .X(n23183) );
  sky130_fd_sc_hd__mux2i_1 U28367 ( .A0(j202_soc_core_intc_core_00_rg_ipr[3]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[7]), .S(n27316), .Y(n23238) );
  sky130_fd_sc_hd__mux2_2 U28368 ( .A0(j202_soc_core_intc_core_00_rg_ipr[15]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[11]), .S(n27315), .X(n23240) );
  sky130_fd_sc_hd__o21ai_1 U28369 ( .A1(n23238), .A2(n23240), .B1(n23173), .Y(
        n23182) );
  sky130_fd_sc_hd__mux2i_1 U28370 ( .A0(j202_soc_core_intc_core_00_rg_ipr[0]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[4]), .S(n27316), .Y(n23227) );
  sky130_fd_sc_hd__mux2_2 U28371 ( .A0(j202_soc_core_intc_core_00_rg_ipr[12]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[8]), .S(n27315), .X(n23230) );
  sky130_fd_sc_hd__mux2_2 U28372 ( .A0(j202_soc_core_intc_core_00_rg_ipr[13]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[9]), .S(n27315), .X(n23221) );
  sky130_fd_sc_hd__mux2i_1 U28373 ( .A0(j202_soc_core_intc_core_00_rg_ipr[1]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[5]), .S(n27316), .Y(n23222) );
  sky130_fd_sc_hd__nand2_1 U28374 ( .A(n23221), .B(n23222), .Y(n23174) );
  sky130_fd_sc_hd__nand2_1 U28375 ( .A(n23175), .B(n23174), .Y(n23179) );
  sky130_fd_sc_hd__nand2_1 U28376 ( .A(n23176), .B(n23183), .Y(n23178) );
  sky130_fd_sc_hd__o2bb2ai_1 U28377 ( .B1(n23183), .B2(n23176), .A1_N(n23240), 
        .A2_N(n23238), .Y(n23177) );
  sky130_fd_sc_hd__a21oi_1 U28378 ( .A1(n23179), .A2(n23178), .B1(n23177), .Y(
        n23181) );
  sky130_fd_sc_hd__o21a_2 U28379 ( .A1(n23182), .A2(n23181), .B1(n23180), .X(
        n23228) );
  sky130_fd_sc_hd__mux2_2 U28380 ( .A0(n23184), .A1(n23183), .S(n23228), .X(
        n23220) );
  sky130_fd_sc_hd__nand2_1 U28381 ( .A(n30173), .B(
        j202_soc_core_intc_core_00_rg_ipr[22]), .Y(n23186) );
  sky130_fd_sc_hd__a2bb2oi_1 U28382 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[19]), .B2(n26688), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[22]), .A2_N(n30173), .Y(n23187) );
  sky130_fd_sc_hd__nand2_1 U28383 ( .A(n23188), .B(n23187), .Y(n23191) );
  sky130_fd_sc_hd__a21oi_1 U28384 ( .A1(n25324), .A2(
        j202_soc_core_intc_core_00_rg_ipr[23]), .B1(n23189), .Y(n23190) );
  sky130_fd_sc_hd__nand2_1 U28385 ( .A(n23191), .B(n23190), .Y(n23194) );
  sky130_fd_sc_hd__inv_2 U28387 ( .A(n23203), .Y(n27321) );
  sky130_fd_sc_hd__inv_1 U28389 ( .A(n23209), .Y(n23219) );
  sky130_fd_sc_hd__nand2_1 U28390 ( .A(n26690), .B(
        j202_soc_core_intc_core_00_rg_ipr[30]), .Y(n23196) );
  sky130_fd_sc_hd__o2bb2ai_1 U28391 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[28]), .B2(n26706), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[25]), .A2_N(n25490), .Y(n23195) );
  sky130_fd_sc_hd__o211ai_1 U28392 ( .A1(j202_soc_core_intc_core_00_rg_ipr[25]), .A2(n25490), .B1(n23196), .C1(n23195), .Y(n23198) );
  sky130_fd_sc_hd__a2bb2oi_1 U28393 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[27]), .B2(n26709), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[30]), .A2_N(n26690), .Y(n23197) );
  sky130_fd_sc_hd__nand2_1 U28394 ( .A(n23198), .B(n23197), .Y(n23202) );
  sky130_fd_sc_hd__a21oi_1 U28395 ( .A1(n26708), .A2(
        j202_soc_core_intc_core_00_rg_ipr[31]), .B1(n23199), .Y(n23201) );
  sky130_fd_sc_hd__mux2i_1 U28396 ( .A0(j202_soc_core_intc_core_00_rg_ipr[30]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[26]), .S(n23212), .Y(n23218) );
  sky130_fd_sc_hd__mux2_2 U28397 ( .A0(j202_soc_core_intc_core_00_rg_ipr[19]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[23]), .S(n27321), .X(n23242) );
  sky130_fd_sc_hd__mux2_2 U28398 ( .A0(j202_soc_core_intc_core_00_rg_ipr[25]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[29]), .S(n27318), .X(n23232) );
  sky130_fd_sc_hd__mux2i_1 U28399 ( .A0(j202_soc_core_intc_core_00_rg_ipr[21]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[17]), .S(n23203), .Y(n23231) );
  sky130_fd_sc_hd__nand2_1 U28400 ( .A(n23232), .B(n23231), .Y(n23204) );
  sky130_fd_sc_hd__mux2i_1 U28401 ( .A0(j202_soc_core_intc_core_00_rg_ipr[28]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[24]), .S(n23212), .Y(n23225) );
  sky130_fd_sc_hd__nand3_1 U28402 ( .A(n23204), .B(n23224), .C(n23225), .Y(
        n23205) );
  sky130_fd_sc_hd__o21ai_1 U28403 ( .A1(n23232), .A2(n23231), .B1(n23205), .Y(
        n23208) );
  sky130_fd_sc_hd__nand2_1 U28406 ( .A(n23208), .B(n30010), .Y(n23211) );
  sky130_fd_sc_hd__nand2_1 U28407 ( .A(n23209), .B(n23218), .Y(n23210) );
  sky130_fd_sc_hd__nand2_1 U28408 ( .A(n23211), .B(n23210), .Y(n23213) );
  sky130_fd_sc_hd__mux2i_1 U28409 ( .A0(j202_soc_core_intc_core_00_rg_ipr[31]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[27]), .S(n23212), .Y(n23243) );
  sky130_fd_sc_hd__o21ai_1 U28410 ( .A1(n23242), .A2(n23213), .B1(n23243), .Y(
        n23216) );
  sky130_fd_sc_hd__nand2_1 U28411 ( .A(n23213), .B(n23242), .Y(n23214) );
  sky130_fd_sc_hd__nand3_1 U28412 ( .A(n23216), .B(n23215), .C(n23214), .Y(
        n27320) );
  sky130_fd_sc_hd__nand2_1 U28413 ( .A(n27320), .B(n23217), .Y(n27319) );
  sky130_fd_sc_hd__mux2_2 U28414 ( .A0(n23219), .A1(n23218), .S(n30169), .X(
        n23251) );
  sky130_fd_sc_hd__nor2_1 U28415 ( .A(n23220), .B(n23251), .Y(n23236) );
  sky130_fd_sc_hd__mux2_2 U28416 ( .A0(n23223), .A1(n23222), .S(n23228), .X(
        n23262) );
  sky130_fd_sc_hd__mux2_2 U28417 ( .A0(n23226), .A1(n23225), .S(n27319), .X(
        n23357) );
  sky130_fd_sc_hd__mux2_2 U28418 ( .A0(n23230), .A1(n23229), .S(n23228), .X(
        n23352) );
  sky130_fd_sc_hd__nand2_1 U28419 ( .A(n23357), .B(n23352), .Y(n23234) );
  sky130_fd_sc_hd__maj3_2 U28420 ( .A(n23262), .B(n23234), .C(n23260), .X(
        n23235) );
  sky130_fd_sc_hd__mux2_2 U28421 ( .A0(n23240), .A1(n23239), .S(n23228), .X(
        n23264) );
  sky130_fd_sc_hd__a21oi_1 U28422 ( .A1(n23245), .A2(n23264), .B1(n23241), .Y(
        n23247) );
  sky130_fd_sc_hd__mux2_2 U28423 ( .A0(n23244), .A1(n23243), .S(n30169), .X(
        n23265) );
  sky130_fd_sc_hd__o21ai_1 U28424 ( .A1(n23264), .A2(n23245), .B1(n23265), .Y(
        n23246) );
  sky130_fd_sc_hd__nand2_1 U28425 ( .A(n23247), .B(n23246), .Y(n23250) );
  sky130_fd_sc_hd__nand2_4 U28426 ( .A(n23250), .B(n23249), .Y(n27322) );
  sky130_fd_sc_hd__mux2i_1 U28427 ( .A0(n23252), .A1(n23251), .S(n27322), .Y(
        n23270) );
  sky130_fd_sc_hd__mux2i_1 U28429 ( .A0(n23256), .A1(n23255), .S(n27333), .Y(
        n23353) );
  sky130_fd_sc_hd__nor2_1 U28430 ( .A(n23257), .B(n23353), .Y(n23263) );
  sky130_fd_sc_hd__mux2i_1 U28431 ( .A0(n23259), .A1(n23258), .S(n27333), .Y(
        n23349) );
  sky130_fd_sc_hd__inv_1 U28432 ( .A(n23260), .Y(n23261) );
  sky130_fd_sc_hd__mux2i_1 U28433 ( .A0(n23262), .A1(n23261), .S(n27322), .Y(
        n23350) );
  sky130_fd_sc_hd__mux2i_1 U28434 ( .A0(n23269), .A1(n23268), .S(n27333), .Y(
        n23273) );
  sky130_fd_sc_hd__o22a_1 U28435 ( .A1(n23281), .A2(n23270), .B1(n23368), .B2(
        n23273), .X(n23271) );
  sky130_fd_sc_hd__o22a_1 U28436 ( .A1(n23276), .A2(n23275), .B1(n23366), .B2(
        n23274), .X(n23277) );
  sky130_fd_sc_hd__nand2_1 U28437 ( .A(n23279), .B(n23278), .Y(n23354) );
  sky130_fd_sc_hd__inv_2 U28438 ( .A(n23354), .Y(n23365) );
  sky130_fd_sc_hd__mux2_2 U28439 ( .A0(n23281), .A1(n23280), .S(n23365), .X(
        n24383) );
  sky130_fd_sc_hd__o21ai_1 U28440 ( .A1(j202_soc_core_intc_core_00_rg_ipr[65]), 
        .A2(n27151), .B1(j202_soc_core_intc_core_00_rg_ipr[64]), .Y(n23282) );
  sky130_fd_sc_hd__o22ai_1 U28441 ( .A1(j202_soc_core_intc_core_00_rg_ipr[68]), 
        .A2(n23282), .B1(j202_soc_core_intc_core_00_rg_ipr[69]), .B2(n28552), 
        .Y(n23283) );
  sky130_fd_sc_hd__a222oi_1 U28442 ( .A1(j202_soc_core_intc_core_00_rg_ipr[66]), .A2(n26761), .B1(j202_soc_core_intc_core_00_rg_ipr[66]), .B2(n23283), .C1(
        n26761), .C2(n23283), .Y(n23284) );
  sky130_fd_sc_hd__maj3_1 U28443 ( .A(j202_soc_core_intc_core_00_rg_ipr[71]), 
        .B(n27684), .C(n23284), .X(n23288) );
  sky130_fd_sc_hd__nand2_1 U28444 ( .A(n27342), .B(
        j202_soc_core_intc_core_00_rg_ipr[66]), .Y(n23289) );
  sky130_fd_sc_hd__a21oi_1 U28446 ( .A1(j202_soc_core_intc_core_00_rg_ipr[77]), 
        .A2(n27936), .B1(j202_soc_core_intc_core_00_rg_ipr[76]), .Y(n23291) );
  sky130_fd_sc_hd__o22ai_1 U28447 ( .A1(j202_soc_core_intc_core_00_rg_ipr[77]), 
        .A2(n27936), .B1(j202_soc_core_intc_core_00_rg_ipr[78]), .B2(n25076), 
        .Y(n23290) );
  sky130_fd_sc_hd__a21oi_1 U28448 ( .A1(j202_soc_core_intc_core_00_rg_ipr[72]), 
        .A2(n23291), .B1(n23290), .Y(n23293) );
  sky130_fd_sc_hd__o22ai_1 U28449 ( .A1(j202_soc_core_intc_core_00_rg_ipr[75]), 
        .A2(n26124), .B1(j202_soc_core_intc_core_00_rg_ipr[74]), .B2(n26883), 
        .Y(n23292) );
  sky130_fd_sc_hd__o22ai_1 U28450 ( .A1(n23293), .A2(n23292), .B1(
        j202_soc_core_intc_core_00_rg_ipr[79]), .B2(n26767), .Y(n23297) );
  sky130_fd_sc_hd__nand2_1 U28451 ( .A(n27339), .B(n26883), .Y(n23298) );
  sky130_fd_sc_hd__o21ai_1 U28452 ( .A1(j202_soc_core_intc_core_00_rg_ipr[74]), 
        .A2(n27339), .B1(n23298), .Y(n23315) );
  sky130_fd_sc_hd__nand2_1 U28453 ( .A(n27342), .B(n28230), .Y(n23299) );
  sky130_fd_sc_hd__o21ai_1 U28454 ( .A1(j202_soc_core_intc_core_00_rg_ipr[68]), 
        .A2(n27342), .B1(n23299), .Y(n23324) );
  sky130_fd_sc_hd__nand2_1 U28455 ( .A(n27339), .B(n25791), .Y(n23300) );
  sky130_fd_sc_hd__nand2_1 U28457 ( .A(n27342), .B(
        j202_soc_core_intc_core_00_rg_ipr[65]), .Y(n23301) );
  sky130_fd_sc_hd__o21ai_1 U28458 ( .A1(n27151), .A2(n27342), .B1(n23301), .Y(
        n23328) );
  sky130_fd_sc_hd__nand2_1 U28459 ( .A(n27339), .B(n25192), .Y(n23302) );
  sky130_fd_sc_hd__o21ai_1 U28460 ( .A1(j202_soc_core_intc_core_00_rg_ipr[72]), 
        .A2(n27339), .B1(n23302), .Y(n23323) );
  sky130_fd_sc_hd__o2bb2ai_1 U28462 ( .B1(n23324), .B2(n23303), .A1_N(n23327), 
        .A2_N(n23328), .Y(n23304) );
  sky130_fd_sc_hd__nand2b_1 U28463 ( .A_N(n27339), .B(n26767), .Y(n23306) );
  sky130_fd_sc_hd__nand2_1 U28464 ( .A(n27339), .B(n26124), .Y(n23305) );
  sky130_fd_sc_hd__nand2_1 U28465 ( .A(n23306), .B(n23305), .Y(n23318) );
  sky130_fd_sc_hd__a21oi_1 U28466 ( .A1(n23310), .A2(n23318), .B1(n23308), .Y(
        n23312) );
  sky130_fd_sc_hd__nand2_1 U28467 ( .A(n27342), .B(
        j202_soc_core_intc_core_00_rg_ipr[67]), .Y(n23309) );
  sky130_fd_sc_hd__o21ai_1 U28468 ( .A1(n26766), .A2(n27342), .B1(n23309), .Y(
        n23319) );
  sky130_fd_sc_hd__o21ai_1 U28469 ( .A1(n23318), .A2(n23310), .B1(n23319), .Y(
        n23311) );
  sky130_fd_sc_hd__nand2_1 U28470 ( .A(n23312), .B(n23311), .Y(n23314) );
  sky130_fd_sc_hd__nand2_1 U28471 ( .A(n24392), .B(n23315), .Y(n23316) );
  sky130_fd_sc_hd__o21ai_1 U28472 ( .A1(n23317), .A2(n24392), .B1(n23316), .Y(
        n23334) );
  sky130_fd_sc_hd__nor2_1 U28473 ( .A(n23320), .B(n24392), .Y(n23321) );
  sky130_fd_sc_hd__a21oi_1 U28474 ( .A1(n23322), .A2(n24392), .B1(n23321), .Y(
        n23369) );
  sky130_fd_sc_hd__nor2_1 U28475 ( .A(n23324), .B(n24392), .Y(n23325) );
  sky130_fd_sc_hd__a21oi_1 U28476 ( .A1(n24392), .A2(n23326), .B1(n23325), .Y(
        n24372) );
  sky130_fd_sc_hd__nand2_1 U28477 ( .A(n24392), .B(n23327), .Y(n23331) );
  sky130_fd_sc_hd__nand2_1 U28478 ( .A(n27341), .B(n23329), .Y(n23330) );
  sky130_fd_sc_hd__nand2_1 U28479 ( .A(n23331), .B(n23330), .Y(n23348) );
  sky130_fd_sc_hd__o22ai_1 U28480 ( .A1(j202_soc_core_intc_core_00_rg_ipr[80]), 
        .A2(n24372), .B1(n23348), .B2(j202_soc_core_intc_core_00_rg_ipr[81]), 
        .Y(n23333) );
  sky130_fd_sc_hd__nand2_1 U28481 ( .A(n23348), .B(
        j202_soc_core_intc_core_00_rg_ipr[81]), .Y(n23332) );
  sky130_fd_sc_hd__nand2_1 U28482 ( .A(n23333), .B(n23332), .Y(n23335) );
  sky130_fd_sc_hd__o21ai_1 U28483 ( .A1(j202_soc_core_intc_core_00_rg_ipr[82]), 
        .A2(n23335), .B1(n23334), .Y(n23337) );
  sky130_fd_sc_hd__nand2_1 U28484 ( .A(n23335), .B(
        j202_soc_core_intc_core_00_rg_ipr[82]), .Y(n23336) );
  sky130_fd_sc_hd__nand2_1 U28485 ( .A(n23337), .B(n23336), .Y(n23338) );
  sky130_fd_sc_hd__nand2_1 U28487 ( .A(n23369), .B(
        j202_soc_core_intc_core_00_rg_ipr[83]), .Y(n23339) );
  sky130_fd_sc_hd__nand2_1 U28488 ( .A(n23340), .B(n23339), .Y(n23343) );
  sky130_fd_sc_hd__nand2_1 U28489 ( .A(n23343), .B(n23342), .Y(n23346) );
  sky130_fd_sc_hd__mux2_2 U28490 ( .A0(n23347), .A1(
        j202_soc_core_intc_core_00_rg_ipr[82]), .S(n24376), .X(n24382) );
  sky130_fd_sc_hd__nor2_1 U28491 ( .A(n24383), .B(n24382), .Y(n23364) );
  sky130_fd_sc_hd__mux2_2 U28492 ( .A0(n23348), .A1(n25747), .S(n24376), .X(
        n24381) );
  sky130_fd_sc_hd__mux2_2 U28493 ( .A0(n23351), .A1(n23350), .S(n23365), .X(
        n24379) );
  sky130_fd_sc_hd__nor2_1 U28494 ( .A(n23352), .B(n27322), .Y(n23356) );
  sky130_fd_sc_hd__buf_4 U28495 ( .A(n23354), .X(n27336) );
  sky130_fd_sc_hd__inv_1 U28497 ( .A(n27322), .Y(n24387) );
  sky130_fd_sc_hd__nand2_1 U28498 ( .A(n24391), .B(n23357), .Y(n23358) );
  sky130_fd_sc_hd__nand2_1 U28499 ( .A(n23359), .B(n23358), .Y(n24374) );
  sky130_fd_sc_hd__mux2i_1 U28500 ( .A0(n24372), .A1(n27098), .S(n24376), .Y(
        n23360) );
  sky130_fd_sc_hd__nor2_1 U28501 ( .A(n24374), .B(n23360), .Y(n23361) );
  sky130_fd_sc_hd__o21ai_1 U28502 ( .A1(n24381), .A2(n24379), .B1(n23361), .Y(
        n23363) );
  sky130_fd_sc_hd__nand2_1 U28503 ( .A(n24379), .B(n24381), .Y(n23362) );
  sky130_fd_sc_hd__buf_2 U28505 ( .A(n23365), .X(n27713) );
  sky130_fd_sc_hd__nor2_1 U28506 ( .A(n23273), .B(n27713), .Y(n23367) );
  sky130_fd_sc_hd__mux2_2 U28507 ( .A0(n23369), .A1(n25325), .S(n24376), .X(
        n24371) );
  sky130_fd_sc_hd__a2bb2oi_1 U28508 ( .B1(n24383), .B2(n24382), .A1_N(n12093), 
        .A2_N(n24371), .Y(n23370) );
  sky130_fd_sc_hd__nand2_1 U28509 ( .A(n23371), .B(n23370), .Y(n23375) );
  sky130_fd_sc_hd__a21oi_1 U28510 ( .A1(n24371), .A2(n12093), .B1(n23373), .Y(
        n23374) );
  sky130_fd_sc_hd__nand2_4 U28511 ( .A(n30088), .B(n12861), .Y(n23403) );
  sky130_fd_sc_hd__nand2_1 U28513 ( .A(n24546), .B(n24551), .Y(n23381) );
  sky130_fd_sc_hd__inv_2 U28514 ( .A(n29589), .Y(n23398) );
  sky130_fd_sc_hd__nand2b_4 U28515 ( .A_N(n12236), .B(n23394), .Y(n27730) );
  sky130_fd_sc_hd__buf_2 U28516 ( .A(n23396), .X(n24106) );
  sky130_fd_sc_hd__nand2_1 U28518 ( .A(n24593), .B(n23392), .Y(n23611) );
  sky130_fd_sc_hd__nand2_1 U28519 ( .A(n23604), .B(n10960), .Y(n23383) );
  sky130_fd_sc_hd__nand2_1 U28520 ( .A(n23392), .B(n11494), .Y(n23385) );
  sky130_fd_sc_hd__nor2_1 U28521 ( .A(n24616), .B(n24619), .Y(n24553) );
  sky130_fd_sc_hd__nor2_1 U28523 ( .A(n23389), .B(n12336), .Y(n24399) );
  sky130_fd_sc_hd__nor2_1 U28524 ( .A(n24628), .B(n28388), .Y(n23390) );
  sky130_fd_sc_hd__inv_1 U28525 ( .A(n10960), .Y(n24102) );
  sky130_fd_sc_hd__nand2_1 U28526 ( .A(n27901), .B(n24102), .Y(n23946) );
  sky130_fd_sc_hd__nor2_2 U28528 ( .A(n11395), .B(n27899), .Y(n23547) );
  sky130_fd_sc_hd__nor2_1 U28529 ( .A(n23608), .B(n23404), .Y(n23410) );
  sky130_fd_sc_hd__nand3_1 U28531 ( .A(n24406), .B(n24409), .C(n24111), .Y(
        n24654) );
  sky130_fd_sc_hd__nor2_1 U28532 ( .A(n12038), .B(n24654), .Y(n23409) );
  sky130_fd_sc_hd__nand2_1 U28533 ( .A(n28394), .B(n28379), .Y(n23411) );
  sky130_fd_sc_hd__nor2_1 U28534 ( .A(n28373), .B(n24394), .Y(n24416) );
  sky130_fd_sc_hd__nor2_1 U28535 ( .A(n23420), .B(n23412), .Y(n24585) );
  sky130_fd_sc_hd__and3_1 U28536 ( .A(n23414), .B(
        j202_soc_core_j22_cpu_opst[3]), .C(n23413), .X(n24417) );
  sky130_fd_sc_hd__nor2_1 U28537 ( .A(n24585), .B(n24417), .Y(n23415) );
  sky130_fd_sc_hd__nand3_1 U28538 ( .A(n23416), .B(n24540), .C(n23415), .Y(
        n24685) );
  sky130_fd_sc_hd__nand2_1 U28539 ( .A(n23417), .B(n28085), .Y(n24539) );
  sky130_fd_sc_hd__nand2_1 U28540 ( .A(n24539), .B(n28071), .Y(n24697) );
  sky130_fd_sc_hd__nand2b_1 U28541 ( .A_N(n24685), .B(n23418), .Y(n24603) );
  sky130_fd_sc_hd__nor2_1 U28542 ( .A(n23419), .B(n24603), .Y(n24109) );
  sky130_fd_sc_hd__nand2_1 U28544 ( .A(n28360), .B(n28403), .Y(n28127) );
  sky130_fd_sc_hd__nor2_1 U28545 ( .A(n23421), .B(n27743), .Y(n23424) );
  sky130_fd_sc_hd__nand2_1 U28546 ( .A(n22003), .B(n29490), .Y(n23422) );
  sky130_fd_sc_hd__o21ai_1 U28548 ( .A1(n23424), .A2(n12232), .B1(n30089), .Y(
        n23425) );
  sky130_fd_sc_hd__nand2_1 U28549 ( .A(n23425), .B(n12254), .Y(n23432) );
  sky130_fd_sc_hd__nand2_1 U28550 ( .A(n24560), .B(n23426), .Y(n23430) );
  sky130_fd_sc_hd__nand2_1 U28551 ( .A(n23427), .B(n29489), .Y(n23428) );
  sky130_fd_sc_hd__nand2_1 U28553 ( .A(n29587), .B(n23549), .Y(n23435) );
  sky130_fd_sc_hd__a21oi_1 U28554 ( .A1(n29490), .A2(n12317), .B1(n24591), .Y(
        n23440) );
  sky130_fd_sc_hd__nand3_1 U28555 ( .A(n11646), .B(n23444), .C(n12332), .Y(
        n24690) );
  sky130_fd_sc_hd__nand3_1 U28556 ( .A(n23445), .B(n30083), .C(n24690), .Y(
        n23450) );
  sky130_fd_sc_hd__nand2_1 U28558 ( .A(n12669), .B(n29587), .Y(n27726) );
  sky130_fd_sc_hd__nand2_1 U28559 ( .A(n28117), .B(n28127), .Y(n23453) );
  sky130_fd_sc_hd__nor2_1 U28560 ( .A(n23453), .B(n23452), .Y(n23454) );
  sky130_fd_sc_hd__nand2_1 U28561 ( .A(n24574), .B(n23550), .Y(n23457) );
  sky130_fd_sc_hd__nand3_1 U28562 ( .A(n23459), .B(n23458), .C(n12235), .Y(
        n23460) );
  sky130_fd_sc_hd__a21oi_1 U28563 ( .A1(n23460), .A2(n28417), .B1(n24696), .Y(
        n27894) );
  sky130_fd_sc_hd__nor2_1 U28564 ( .A(n23462), .B(n23461), .Y(n23467) );
  sky130_fd_sc_hd__nand2_1 U28565 ( .A(n23463), .B(n23471), .Y(n23465) );
  sky130_fd_sc_hd__nand4_1 U28566 ( .A(n23469), .B(n24855), .C(n23470), .D(
        n26032), .Y(n23464) );
  sky130_fd_sc_hd__nor2_1 U28567 ( .A(n23465), .B(n23464), .Y(n23466) );
  sky130_fd_sc_hd__nor2_1 U28568 ( .A(n26032), .B(n23469), .Y(n23474) );
  sky130_fd_sc_hd__nor2_1 U28569 ( .A(n24855), .B(n23470), .Y(n23473) );
  sky130_fd_sc_hd__nand4_1 U28570 ( .A(n23474), .B(n23473), .C(n25770), .D(
        n23472), .Y(n23475) );
  sky130_fd_sc_hd__inv_1 U28571 ( .A(n23475), .Y(n23491) );
  sky130_fd_sc_hd__nor2_1 U28572 ( .A(n23477), .B(n23476), .Y(n23481) );
  sky130_fd_sc_hd__nor2_1 U28573 ( .A(n23479), .B(n23478), .Y(n23480) );
  sky130_fd_sc_hd__nand2_1 U28574 ( .A(n23481), .B(n23480), .Y(n23482) );
  sky130_fd_sc_hd__nor2_1 U28576 ( .A(n23484), .B(n27362), .Y(n23488) );
  sky130_fd_sc_hd__nor2_1 U28577 ( .A(n25890), .B(n23485), .Y(n23486) );
  sky130_fd_sc_hd__nor2_1 U28578 ( .A(n23492), .B(n24854), .Y(n23563) );
  sky130_fd_sc_hd__buf_2 U28579 ( .A(n23494), .X(n25772) );
  sky130_fd_sc_hd__a21oi_1 U28580 ( .A1(n23495), .A2(n11146), .B1(n24853), .Y(
        n23496) );
  sky130_fd_sc_hd__nand2_4 U28581 ( .A(n25772), .B(n23496), .Y(n23588) );
  sky130_fd_sc_hd__nand2_1 U28582 ( .A(n27768), .B(n11392), .Y(n23497) );
  sky130_fd_sc_hd__o211ai_1 U28583 ( .A1(n25869), .A2(n27770), .B1(n23588), 
        .C1(n23497), .Y(j202_soc_core_j22_cpu_ml_maclj[18]) );
  sky130_fd_sc_hd__a211o_1 U28584 ( .A1(n23753), .A2(n23500), .B1(n23499), 
        .C1(n23498), .X(n23501) );
  sky130_fd_sc_hd__nand2b_1 U28585 ( .A_N(n23502), .B(
        j202_soc_core_j22_cpu_ma_M_MEM[0]), .Y(n23510) );
  sky130_fd_sc_hd__nand2b_1 U28587 ( .A_N(n26048), .B(n23517), .Y(n25638) );
  sky130_fd_sc_hd__nand2_1 U28588 ( .A(n27787), .B(n25397), .Y(n25636) );
  sky130_fd_sc_hd__o21ai_1 U28589 ( .A1(n25682), .A2(n26329), .B1(n25636), .Y(
        n23518) );
  sky130_fd_sc_hd__o211ai_1 U28590 ( .A1(n11123), .A2(n26329), .B1(n25638), 
        .C1(n23518), .Y(n23539) );
  sky130_fd_sc_hd__nand2_1 U28591 ( .A(n25385), .B(n27789), .Y(n23537) );
  sky130_fd_sc_hd__nor2_1 U28592 ( .A(n26268), .B(n26311), .Y(n23521) );
  sky130_fd_sc_hd__nand3_1 U28593 ( .A(n23520), .B(n26375), .C(n28489), .Y(
        n26049) );
  sky130_fd_sc_hd__nor2_1 U28594 ( .A(n27147), .B(n26049), .Y(n24883) );
  sky130_fd_sc_hd__a21o_1 U28595 ( .A1(n23522), .A2(n23521), .B1(n24883), .X(
        n25840) );
  sky130_fd_sc_hd__nand2_1 U28596 ( .A(n25840), .B(n26426), .Y(n27814) );
  sky130_fd_sc_hd__o22ai_1 U28597 ( .A1(n27383), .A2(n27795), .B1(n26324), 
        .B2(n27803), .Y(n23525) );
  sky130_fd_sc_hd__nand2b_1 U28598 ( .A_N(n23523), .B(n25999), .Y(n27797) );
  sky130_fd_sc_hd__o22ai_1 U28599 ( .A1(n26296), .A2(n26943), .B1(n11189), 
        .B2(n27797), .Y(n23524) );
  sky130_fd_sc_hd__nor2_1 U28600 ( .A(n23525), .B(n23524), .Y(n23529) );
  sky130_fd_sc_hd__xnor2_1 U28601 ( .A(n28499), .B(n26329), .Y(n26225) );
  sky130_fd_sc_hd__a2bb2oi_1 U28602 ( .B1(n25697), .B2(n27808), .A1_N(n25872), 
        .A2_N(n26225), .Y(n23528) );
  sky130_fd_sc_hd__nand2_1 U28603 ( .A(n25999), .B(n28509), .Y(n27799) );
  sky130_fd_sc_hd__o22ai_1 U28604 ( .A1(n28499), .A2(n27793), .B1(n26321), 
        .B2(n27799), .Y(n23526) );
  sky130_fd_sc_hd__a21oi_1 U28605 ( .A1(n27810), .A2(n25271), .B1(n23526), .Y(
        n23527) );
  sky130_fd_sc_hd__nand4_1 U28606 ( .A(n27814), .B(n23529), .C(n23528), .D(
        n23527), .Y(n23535) );
  sky130_fd_sc_hd__nand2_1 U28607 ( .A(n23531), .B(n24888), .Y(n25820) );
  sky130_fd_sc_hd__nand2_1 U28608 ( .A(n25820), .B(n26426), .Y(n27817) );
  sky130_fd_sc_hd__nand2b_1 U28609 ( .A_N(n23533), .B(n26424), .Y(n25821) );
  sky130_fd_sc_hd__nand2_1 U28610 ( .A(n25821), .B(n26426), .Y(n27815) );
  sky130_fd_sc_hd__o22ai_1 U28611 ( .A1(n26281), .A2(n27817), .B1(n26421), 
        .B2(n27815), .Y(n23534) );
  sky130_fd_sc_hd__nor2_1 U28612 ( .A(n23535), .B(n23534), .Y(n23536) );
  sky130_fd_sc_hd__nand2_1 U28613 ( .A(n23537), .B(n23536), .Y(n23538) );
  sky130_fd_sc_hd__nand2_1 U28614 ( .A(n28499), .B(n27791), .Y(n23540) );
  sky130_fd_sc_hd__nand2_1 U28615 ( .A(n23540), .B(n26919), .Y(n23541) );
  sky130_fd_sc_hd__nand2_1 U28616 ( .A(n23541), .B(n26329), .Y(n25558) );
  sky130_fd_sc_hd__and3_1 U28617 ( .A(n25377), .B(n27828), .C(n25376), .X(
        n23543) );
  sky130_fd_sc_hd__nand3_1 U28619 ( .A(n23469), .B(n25679), .C(n23545), .Y(
        n25560) );
  sky130_fd_sc_hd__o22ai_1 U28620 ( .A1(n25964), .A2(n25594), .B1(n27847), 
        .B2(n12267), .Y(j202_soc_core_j22_cpu_rf_N2702) );
  sky130_fd_sc_hd__nand2_1 U28621 ( .A(n24401), .B(n28387), .Y(n24627) );
  sky130_fd_sc_hd__nand2_1 U28622 ( .A(n28394), .B(n28367), .Y(n24960) );
  sky130_fd_sc_hd__nand2_1 U28623 ( .A(n12208), .B(n28417), .Y(n24959) );
  sky130_fd_sc_hd__nor2_1 U28624 ( .A(n24959), .B(n28121), .Y(n23558) );
  sky130_fd_sc_hd__nand2_1 U28625 ( .A(n23554), .B(n11007), .Y(n24126) );
  sky130_fd_sc_hd__nand2_1 U28626 ( .A(n24126), .B(n28417), .Y(n27990) );
  sky130_fd_sc_hd__nand3_1 U28627 ( .A(n25146), .B(n28417), .C(n29559), .Y(
        n23556) );
  sky130_fd_sc_hd__nor2_1 U28628 ( .A(n23558), .B(n13043), .Y(n23559) );
  sky130_fd_sc_hd__nand2_1 U28629 ( .A(n11689), .B(n23559), .Y(n10534) );
  sky130_fd_sc_hd__nand2_1 U28630 ( .A(n12234), .B(n23563), .Y(n25769) );
  sky130_fd_sc_hd__inv_2 U28631 ( .A(n25779), .Y(n26077) );
  sky130_fd_sc_hd__nand2_1 U28632 ( .A(n26077), .B(n23562), .Y(n23565) );
  sky130_fd_sc_hd__nand2_1 U28633 ( .A(n28056), .B(n27767), .Y(n23564) );
  sky130_fd_sc_hd__nand2_1 U28634 ( .A(n23565), .B(n13081), .Y(n29839) );
  sky130_fd_sc_hd__nand2_1 U28635 ( .A(n26077), .B(n23566), .Y(n23569) );
  sky130_fd_sc_hd__nand2_1 U28636 ( .A(n28056), .B(n23567), .Y(n23568) );
  sky130_fd_sc_hd__nand2_1 U28637 ( .A(n23569), .B(n13080), .Y(n29840) );
  sky130_fd_sc_hd__nand2_1 U28638 ( .A(n26077), .B(n23570), .Y(n23573) );
  sky130_fd_sc_hd__nand2_1 U28639 ( .A(n28056), .B(n23571), .Y(n23572) );
  sky130_fd_sc_hd__nand2_1 U28640 ( .A(n23573), .B(n13079), .Y(n29838) );
  sky130_fd_sc_hd__nand2_1 U28641 ( .A(n26077), .B(n23574), .Y(n23576) );
  sky130_fd_sc_hd__nand2_1 U28642 ( .A(n28056), .B(
        j202_soc_core_j22_cpu_ml_bufa[24]), .Y(n23575) );
  sky130_fd_sc_hd__nand2_1 U28643 ( .A(n23576), .B(n13095), .Y(n29841) );
  sky130_fd_sc_hd__o211ai_1 U28644 ( .A1(n24854), .A2(n23580), .B1(n23579), 
        .C1(n23578), .Y(n23581) );
  sky130_fd_sc_hd__nand2_1 U28645 ( .A(n26077), .B(n23581), .Y(n23584) );
  sky130_fd_sc_hd__nand2_1 U28646 ( .A(n28056), .B(n23582), .Y(n23583) );
  sky130_fd_sc_hd__nand2_1 U28647 ( .A(n23584), .B(n13078), .Y(n29837) );
  sky130_fd_sc_hd__nand2_1 U28648 ( .A(n26077), .B(n25665), .Y(n23586) );
  sky130_fd_sc_hd__nand2_1 U28649 ( .A(n28056), .B(n11474), .Y(n23585) );
  sky130_fd_sc_hd__nand2_1 U28650 ( .A(n23586), .B(n13077), .Y(n29843) );
  sky130_fd_sc_hd__nand2_1 U28651 ( .A(n12330), .B(
        j202_soc_core_j22_cpu_ml_macl[4]), .Y(n23592) );
  sky130_fd_sc_hd__a21oi_1 U28652 ( .A1(n27768), .A2(
        j202_soc_core_j22_cpu_ml_bufa[4]), .B1(n27766), .Y(n23591) );
  sky130_fd_sc_hd__inv_2 U28653 ( .A(n24312), .Y(n24325) );
  sky130_fd_sc_hd__nand2_1 U28654 ( .A(n24325), .B(n22317), .Y(n23590) );
  sky130_fd_sc_hd__nand3_1 U28655 ( .A(n23590), .B(n23592), .C(n23591), .Y(
        j202_soc_core_j22_cpu_ml_maclj[4]) );
  sky130_fd_sc_hd__nand2_1 U28656 ( .A(n12330), .B(
        j202_soc_core_j22_cpu_ml_macl[2]), .Y(n23596) );
  sky130_fd_sc_hd__a21oi_1 U28657 ( .A1(n27768), .A2(n12436), .B1(n27766), .Y(
        n23595) );
  sky130_fd_sc_hd__nand2_1 U28658 ( .A(n24325), .B(n22364), .Y(n23594) );
  sky130_fd_sc_hd__nand3_1 U28659 ( .A(n23594), .B(n23596), .C(n23595), .Y(
        j202_soc_core_j22_cpu_ml_maclj[2]) );
  sky130_fd_sc_hd__nand3_1 U28660 ( .A(n11098), .B(n24401), .C(n28344), .Y(
        n23620) );
  sky130_fd_sc_hd__nand3_1 U28662 ( .A(n24583), .B(n23599), .C(n24409), .Y(
        n23600) );
  sky130_fd_sc_hd__nand2b_1 U28663 ( .A_N(n12285), .B(n11728), .Y(n24124) );
  sky130_fd_sc_hd__nand3_1 U28664 ( .A(n27901), .B(n23603), .C(n12332), .Y(
        n23996) );
  sky130_fd_sc_hd__nand2b_1 U28665 ( .A_N(n30072), .B(n23604), .Y(n24572) );
  sky130_fd_sc_hd__nand4_1 U28666 ( .A(n23606), .B(n23996), .C(n23605), .D(
        n24572), .Y(n23607) );
  sky130_fd_sc_hd__nor2_1 U28667 ( .A(n23612), .B(n27981), .Y(n24579) );
  sky130_fd_sc_hd__nand3_1 U28668 ( .A(n12136), .B(n23614), .C(n29587), .Y(
        n24110) );
  sky130_fd_sc_hd__clkbuf_1 U28671 ( .A(la_data_out[16]), .X(io_out[36]) );
  sky130_fd_sc_hd__and3_1 U28672 ( .A(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[0]), .C(n23898), .X(io_oeb[12]) );
  sky130_fd_sc_hd__clkbuf_1 U28673 ( .A(la_data_out[15]), .X(io_out[35]) );
  sky130_fd_sc_hd__clkbuf_1 U28674 ( .A(io_oeb[12]), .X(io_oeb[10]) );
  sky130_fd_sc_hd__clkbuf_1 U28675 ( .A(la_data_out[14]), .X(io_out[34]) );
  sky130_fd_sc_hd__clkbuf_1 U28676 ( .A(la_data_out[13]), .X(io_out[33]) );
  sky130_fd_sc_hd__clkbuf_1 U28677 ( .A(la_data_out[12]), .X(io_out[32]) );
  sky130_fd_sc_hd__clkbuf_1 U28678 ( .A(la_data_out[0]), .X(io_out[0]) );
  sky130_fd_sc_hd__clkbuf_1 U28679 ( .A(la_data_out[10]), .X(io_out[30]) );
  sky130_fd_sc_hd__clkbuf_1 U28680 ( .A(la_data_out[1]), .X(io_out[1]) );
  sky130_fd_sc_hd__clkbuf_1 U28681 ( .A(la_data_out[9]), .X(io_out[29]) );
  sky130_fd_sc_hd__clkbuf_1 U28682 ( .A(la_data_out[8]), .X(io_out[28]) );
  sky130_fd_sc_hd__clkbuf_1 U28683 ( .A(la_data_out[7]), .X(io_out[27]) );
  sky130_fd_sc_hd__clkbuf_1 U28684 ( .A(la_data_out[6]), .X(io_out[26]) );
  sky130_fd_sc_hd__clkbuf_1 U28685 ( .A(la_data_out[3]), .X(io_out[3]) );
  sky130_fd_sc_hd__clkbuf_1 U28686 ( .A(la_data_out[5]), .X(io_out[7]) );
  sky130_fd_sc_hd__clkbuf_1 U28687 ( .A(la_data_out[4]), .X(io_out[4]) );
  sky130_fd_sc_hd__nor2_1 U28688 ( .A(n23626), .B(n23625), .Y(n28432) );
  sky130_fd_sc_hd__nand2_1 U28689 ( .A(n23627), .B(n28538), .Y(n28512) );
  sky130_fd_sc_hd__nand3_1 U28690 ( .A(n24428), .B(
        j202_soc_core_j22_cpu_macop_MAC_[3]), .C(n27763), .Y(n24430) );
  sky130_fd_sc_hd__nor2_1 U28691 ( .A(j202_soc_core_ahb2apb_02_state[2]), .B(
        j202_soc_core_ahb2apb_02_state[0]), .Y(n26899) );
  sky130_fd_sc_hd__nand4_1 U28692 ( .A(j202_soc_core_pstrb[1]), .B(
        j202_soc_core_pstrb[0]), .C(j202_soc_core_pstrb[3]), .D(
        j202_soc_core_pstrb[2]), .Y(n23628) );
  sky130_fd_sc_hd__nor2_1 U28693 ( .A(n23628), .B(n24296), .Y(n23629) );
  sky130_fd_sc_hd__nand3_1 U28694 ( .A(n26899), .B(n23629), .C(
        j202_soc_core_pwrite[2]), .Y(n26783) );
  sky130_fd_sc_hd__nor2_1 U28695 ( .A(j202_soc_core_gpio_core_00_reg_addr[4]), 
        .B(n26908), .Y(n26910) );
  sky130_fd_sc_hd__nor2_1 U28696 ( .A(j202_soc_core_gpio_core_00_reg_addr[7]), 
        .B(j202_soc_core_gpio_core_00_reg_addr[1]), .Y(n23631) );
  sky130_fd_sc_hd__nor2_1 U28697 ( .A(j202_soc_core_gpio_core_00_reg_addr[5]), 
        .B(j202_soc_core_gpio_core_00_reg_addr[6]), .Y(n23630) );
  sky130_fd_sc_hd__and3_1 U28698 ( .A(n23631), .B(n23630), .C(n26777), .X(
        n23882) );
  sky130_fd_sc_hd__nand2_1 U28699 ( .A(n23882), .B(n23856), .Y(n26903) );
  sky130_fd_sc_hd__nand3_1 U28700 ( .A(n26530), .B(n28739), .C(n27614), .Y(
        n27293) );
  sky130_fd_sc_hd__nand2_1 U28701 ( .A(j202_soc_core_qspi_wb_addr[24]), .B(
        j202_soc_core_ahb2wbqspi_00_stb_o), .Y(n23871) );
  sky130_fd_sc_hd__nand2_1 U28702 ( .A(n26543), .B(n27238), .Y(n27288) );
  sky130_fd_sc_hd__nor2_1 U28703 ( .A(j202_soc_core_wbqspiflash_00_state[4]), 
        .B(j202_soc_core_wbqspiflash_00_state[2]), .Y(n28840) );
  sky130_fd_sc_hd__nand2_1 U28704 ( .A(n28840), .B(n28647), .Y(n27210) );
  sky130_fd_sc_hd__nand2b_1 U28705 ( .A_N(n27210), .B(n28870), .Y(n28865) );
  sky130_fd_sc_hd__nor2_1 U28706 ( .A(n27288), .B(n28865), .Y(n28677) );
  sky130_fd_sc_hd__nor2_1 U28707 ( .A(j202_soc_core_wbqspiflash_00_state[1]), 
        .B(n27224), .Y(n27285) );
  sky130_fd_sc_hd__nor2_1 U28708 ( .A(j202_soc_core_wbqspiflash_00_state[4]), 
        .B(n26588), .Y(n27268) );
  sky130_fd_sc_hd__nand2_1 U28709 ( .A(n27268), .B(n28647), .Y(n27201) );
  sky130_fd_sc_hd__nand2_1 U28710 ( .A(n27285), .B(n28871), .Y(n26511) );
  sky130_fd_sc_hd__nor2_1 U28711 ( .A(j202_soc_core_wbqspiflash_00_spi_len[0]), 
        .B(j202_soc_core_wbqspiflash_00_spi_len[1]), .Y(n28708) );
  sky130_fd_sc_hd__nand2_1 U28712 ( .A(n27285), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n27280) );
  sky130_fd_sc_hd__nor2_1 U28713 ( .A(n23633), .B(n27280), .Y(n27431) );
  sky130_fd_sc_hd__a21oi_1 U28714 ( .A1(n23634), .A2(n28708), .B1(n27431), .Y(
        n23635) );
  sky130_fd_sc_hd__nand2_1 U28715 ( .A(n29133), .B(
        j202_soc_core_wbqspiflash_00_spi_valid), .Y(n26513) );
  sky130_fd_sc_hd__nand2_1 U28716 ( .A(n27285), .B(n28840), .Y(n28684) );
  sky130_fd_sc_hd__nor2_1 U28717 ( .A(n28647), .B(n28684), .Y(n26514) );
  sky130_fd_sc_hd__o22ai_1 U28718 ( .A1(n23635), .A2(n27307), .B1(n26513), 
        .B2(n26597), .Y(n26539) );
  sky130_fd_sc_hd__a21oi_1 U28719 ( .A1(n26544), .A2(n28677), .B1(n26539), .Y(
        n23637) );
  sky130_fd_sc_hd__nand2_1 U28720 ( .A(j202_soc_core_wbqspiflash_00_state[1]), 
        .B(j202_soc_core_wbqspiflash_00_state[3]), .Y(n25205) );
  sky130_fd_sc_hd__nor2_1 U28721 ( .A(n25205), .B(n27201), .Y(n27429) );
  sky130_fd_sc_hd__nand2_1 U28722 ( .A(n27429), .B(
        j202_soc_core_wbqspiflash_00_spi_valid), .Y(n25340) );
  sky130_fd_sc_hd__nand2_1 U28723 ( .A(n28870), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n27254) );
  sky130_fd_sc_hd__nor2_1 U28724 ( .A(n27284), .B(n27254), .Y(n23869) );
  sky130_fd_sc_hd__nand2_1 U28725 ( .A(n26530), .B(n28739), .Y(n23872) );
  sky130_fd_sc_hd__nor2_1 U28726 ( .A(n23872), .B(n27288), .Y(n23866) );
  sky130_fd_sc_hd__nand2_1 U28727 ( .A(n23869), .B(n23866), .Y(n26548) );
  sky130_fd_sc_hd__nor2_1 U28728 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[0]), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[1]), .Y(n29274) );
  sky130_fd_sc_hd__or3_1 U28729 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[2]), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[3]), .C(n26474), .X(n28645)
         );
  sky130_fd_sc_hd__nor2_1 U28730 ( .A(n28653), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[7]), .Y(n26469) );
  sky130_fd_sc_hd__nand2_1 U28731 ( .A(n26469), .B(n23638), .Y(n26471) );
  sky130_fd_sc_hd__nand2b_1 U28732 ( .A_N(n26471), .B(n26477), .Y(n26651) );
  sky130_fd_sc_hd__nand2_1 U28733 ( .A(n23639), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n26479) );
  sky130_fd_sc_hd__nand2_1 U28734 ( .A(n23640), .B(n27224), .Y(n26483) );
  sky130_fd_sc_hd__nor2_1 U28735 ( .A(n26483), .B(n27284), .Y(n26467) );
  sky130_fd_sc_hd__nand2_1 U28736 ( .A(n28367), .B(n29745), .Y(n24651) );
  sky130_fd_sc_hd__nand2_1 U28737 ( .A(n23641), .B(n24718), .Y(n23830) );
  sky130_fd_sc_hd__nor3_1 U28738 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__3_), 
        .B(n23830), .C(n28109), .Y(n23642) );
  sky130_fd_sc_hd__nand2_1 U28739 ( .A(n28870), .B(n26580), .Y(n27183) );
  sky130_fd_sc_hd__xor2_1 U28740 ( .A(j202_soc_core_qspi_wb_addr[8]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[8]), .X(n23659) );
  sky130_fd_sc_hd__nand2_1 U28741 ( .A(n23644), .B(
        j202_soc_core_ahb2wbqspi_00_stb_o), .Y(n27229) );
  sky130_fd_sc_hd__nor2_1 U28742 ( .A(n27238), .B(n27229), .Y(n27197) );
  sky130_fd_sc_hd__clkinv_1 U28743 ( .A(n27197), .Y(n23645) );
  sky130_fd_sc_hd__nor2_1 U28744 ( .A(n23659), .B(n23645), .Y(n23745) );
  sky130_fd_sc_hd__nor2_1 U28745 ( .A(j202_soc_core_qspi_wb_addr[23]), .B(
        n23646), .Y(n23744) );
  sky130_fd_sc_hd__xnor2_1 U28746 ( .A(n23648), .B(n13070), .Y(n23737) );
  sky130_fd_sc_hd__xor2_1 U28747 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]), .B(
        j202_soc_core_qspi_wb_addr[20]), .X(n23650) );
  sky130_fd_sc_hd__xnor2_1 U28748 ( .A(n23651), .B(n23650), .Y(n23730) );
  sky130_fd_sc_hd__xor2_1 U28749 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .B(
        j202_soc_core_qspi_wb_addr[18]), .X(n23653) );
  sky130_fd_sc_hd__xnor2_1 U28750 ( .A(n23654), .B(n23653), .Y(n23723) );
  sky130_fd_sc_hd__xnor2_1 U28751 ( .A(n23656), .B(n13068), .Y(n23716) );
  sky130_fd_sc_hd__xnor2_1 U28752 ( .A(n23658), .B(n13069), .Y(n23662) );
  sky130_fd_sc_hd__xnor2_1 U28753 ( .A(n23660), .B(n23659), .Y(n23661) );
  sky130_fd_sc_hd__nor2_1 U28754 ( .A(n23662), .B(n23661), .Y(n23672) );
  sky130_fd_sc_hd__xnor2_1 U28755 ( .A(j202_soc_core_qspi_wb_addr[7]), .B(
        n23663), .Y(n23664) );
  sky130_fd_sc_hd__xnor2_1 U28756 ( .A(n23665), .B(n23664), .Y(n23670) );
  sky130_fd_sc_hd__xnor2_1 U28757 ( .A(j202_soc_core_qspi_wb_addr[6]), .B(
        n23666), .Y(n23667) );
  sky130_fd_sc_hd__xnor2_1 U28758 ( .A(n23668), .B(n23667), .Y(n23669) );
  sky130_fd_sc_hd__nor2_1 U28759 ( .A(n23670), .B(n23669), .Y(n23671) );
  sky130_fd_sc_hd__nand2_1 U28760 ( .A(n23672), .B(n23671), .Y(n23687) );
  sky130_fd_sc_hd__xnor2_1 U28761 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .B(
        j202_soc_core_qspi_wb_addr[2]), .Y(n23675) );
  sky130_fd_sc_hd__xnor2_1 U28762 ( .A(j202_soc_core_qspi_wb_addr[3]), .B(
        n23860), .Y(n23673) );
  sky130_fd_sc_hd__xnor2_1 U28763 ( .A(n23862), .B(n23673), .Y(n23674) );
  sky130_fd_sc_hd__nor2_1 U28764 ( .A(n23675), .B(n23674), .Y(n23685) );
  sky130_fd_sc_hd__xnor2_1 U28765 ( .A(j202_soc_core_qspi_wb_addr[5]), .B(
        n23676), .Y(n23677) );
  sky130_fd_sc_hd__xnor2_1 U28766 ( .A(n23678), .B(n23677), .Y(n23683) );
  sky130_fd_sc_hd__xnor2_1 U28767 ( .A(j202_soc_core_qspi_wb_addr[4]), .B(
        n23679), .Y(n23681) );
  sky130_fd_sc_hd__xnor2_1 U28768 ( .A(n23681), .B(n23680), .Y(n23682) );
  sky130_fd_sc_hd__nor2_1 U28769 ( .A(n23683), .B(n23682), .Y(n23684) );
  sky130_fd_sc_hd__nand2_1 U28770 ( .A(n23685), .B(n23684), .Y(n23686) );
  sky130_fd_sc_hd__nor2_1 U28771 ( .A(n23687), .B(n23686), .Y(n23714) );
  sky130_fd_sc_hd__xor2_1 U28772 ( .A(j202_soc_core_qspi_wb_addr[14]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]), .X(n23689) );
  sky130_fd_sc_hd__xor2_1 U28773 ( .A(n23690), .B(n23689), .X(n23694) );
  sky130_fd_sc_hd__xor2_1 U28774 ( .A(n23692), .B(n13066), .X(n23693) );
  sky130_fd_sc_hd__nand2_1 U28775 ( .A(n23694), .B(n23693), .Y(n23712) );
  sky130_fd_sc_hd__xor2_1 U28776 ( .A(j202_soc_core_qspi_wb_addr[11]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[11]), .X(n23696) );
  sky130_fd_sc_hd__xnor2_1 U28777 ( .A(n23697), .B(n23696), .Y(n23701) );
  sky130_fd_sc_hd__xnor2_1 U28778 ( .A(n23699), .B(n13073), .Y(n23700) );
  sky130_fd_sc_hd__nor2_1 U28779 ( .A(n23701), .B(n23700), .Y(n23710) );
  sky130_fd_sc_hd__xor2_1 U28780 ( .A(j202_soc_core_qspi_wb_addr[13]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[13]), .X(n23703) );
  sky130_fd_sc_hd__xnor2_1 U28781 ( .A(n23704), .B(n23703), .Y(n23708) );
  sky130_fd_sc_hd__xnor2_1 U28782 ( .A(n23706), .B(n13052), .Y(n23707) );
  sky130_fd_sc_hd__nor2_1 U28783 ( .A(n23708), .B(n23707), .Y(n23709) );
  sky130_fd_sc_hd__nand2_1 U28784 ( .A(n23710), .B(n23709), .Y(n23711) );
  sky130_fd_sc_hd__nor2_1 U28785 ( .A(n23712), .B(n23711), .Y(n23713) );
  sky130_fd_sc_hd__nand2_1 U28786 ( .A(n23714), .B(n23713), .Y(n23715) );
  sky130_fd_sc_hd__nor2_1 U28787 ( .A(n23716), .B(n23715), .Y(n23721) );
  sky130_fd_sc_hd__xor2_1 U28788 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]), .B(
        j202_soc_core_qspi_wb_addr[17]), .X(n23718) );
  sky130_fd_sc_hd__xor2_1 U28789 ( .A(n23719), .B(n23718), .X(n23720) );
  sky130_fd_sc_hd__nand2_1 U28790 ( .A(n23721), .B(n23720), .Y(n23722) );
  sky130_fd_sc_hd__nor2_1 U28791 ( .A(n23723), .B(n23722), .Y(n23728) );
  sky130_fd_sc_hd__xor2_1 U28792 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .B(
        j202_soc_core_qspi_wb_addr[19]), .X(n23725) );
  sky130_fd_sc_hd__xor2_1 U28793 ( .A(n23726), .B(n23725), .X(n23727) );
  sky130_fd_sc_hd__nand2_1 U28794 ( .A(n23728), .B(n23727), .Y(n23729) );
  sky130_fd_sc_hd__nor2_1 U28795 ( .A(n23730), .B(n23729), .Y(n23735) );
  sky130_fd_sc_hd__xor2_1 U28796 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]), .B(
        j202_soc_core_qspi_wb_addr[21]), .X(n23732) );
  sky130_fd_sc_hd__xor2_1 U28797 ( .A(n23733), .B(n23732), .X(n23734) );
  sky130_fd_sc_hd__nand2_1 U28798 ( .A(n23735), .B(n23734), .Y(n23736) );
  sky130_fd_sc_hd__nor2_1 U28799 ( .A(n23737), .B(n23736), .Y(n23742) );
  sky130_fd_sc_hd__xor2_1 U28800 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]), .B(
        j202_soc_core_qspi_wb_addr[23]), .X(n23739) );
  sky130_fd_sc_hd__xor2_1 U28801 ( .A(n23740), .B(n23739), .X(n23741) );
  sky130_fd_sc_hd__nand2_1 U28802 ( .A(n23742), .B(n23741), .Y(n23743) );
  sky130_fd_sc_hd__nor2_1 U28803 ( .A(n23744), .B(n23743), .Y(n26629) );
  sky130_fd_sc_hd__and2_0 U28804 ( .A(n23745), .B(n26629), .X(n26554) );
  sky130_fd_sc_hd__nand2_1 U28805 ( .A(n26554), .B(n26558), .Y(n27225) );
  sky130_fd_sc_hd__nor3_1 U28806 ( .A(n27254), .B(n27226), .C(n27225), .Y(
        n26510) );
  sky130_fd_sc_hd__nor2_1 U28807 ( .A(j202_soc_core_wbqspiflash_00_state[2]), 
        .B(n26580), .Y(n27219) );
  sky130_fd_sc_hd__nor2_1 U28808 ( .A(n27219), .B(n27268), .Y(n26519) );
  sky130_fd_sc_hd__nand2_1 U28810 ( .A(n23892), .B(n23840), .Y(n24716) );
  sky130_fd_sc_hd__nand2_1 U28811 ( .A(n23746), .B(n24718), .Y(n23839) );
  sky130_fd_sc_hd__nor2_1 U28812 ( .A(n12347), .B(n24771), .Y(n23748) );
  sky130_fd_sc_hd__nor2_1 U28813 ( .A(j202_soc_core_j22_cpu_regop_We__3_), .B(
        j202_soc_core_j22_cpu_regop_We__2_), .Y(n23747) );
  sky130_fd_sc_hd__nand3_1 U28814 ( .A(n28109), .B(n23748), .C(n23747), .Y(
        n23749) );
  sky130_fd_sc_hd__nor2_1 U28815 ( .A(n23751), .B(n24673), .Y(n23786) );
  sky130_fd_sc_hd__nand3_1 U28816 ( .A(n23786), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__2_), .C(n23752), .Y(n23813) );
  sky130_fd_sc_hd__nand2_1 U28817 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__0_), 
        .B(j202_soc_core_j22_cpu_regop_M_Rn__1_), .Y(n23850) );
  sky130_fd_sc_hd__nand2b_1 U28818 ( .A_N(n23841), .B(n23754), .Y(n23759) );
  sky130_fd_sc_hd__nand2b_1 U28819 ( .A_N(n23826), .B(n23757), .Y(n23758) );
  sky130_fd_sc_hd__nand2_1 U28821 ( .A(n23786), .B(n23760), .Y(n23834) );
  sky130_fd_sc_hd__nand2b_1 U28822 ( .A_N(n23841), .B(n11200), .Y(n23764) );
  sky130_fd_sc_hd__nand2b_1 U28823 ( .A_N(n23826), .B(n23762), .Y(n23763) );
  sky130_fd_sc_hd__nand2_1 U28825 ( .A(n23765), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__1_), .Y(n23801) );
  sky130_fd_sc_hd__nand2b_1 U28826 ( .A_N(n23841), .B(n16507), .Y(n23769) );
  sky130_fd_sc_hd__nand2b_1 U28827 ( .A_N(n23826), .B(n23767), .Y(n23768) );
  sky130_fd_sc_hd__nand2_1 U28828 ( .A(n23770), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__0_), .Y(n23829) );
  sky130_fd_sc_hd__nand2b_1 U28829 ( .A_N(n23841), .B(n13566), .Y(n23774) );
  sky130_fd_sc_hd__nand2b_1 U28830 ( .A_N(n23826), .B(n23772), .Y(n23773) );
  sky130_fd_sc_hd__nand3_1 U28831 ( .A(n23786), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__3_), .C(n23775), .Y(n23818) );
  sky130_fd_sc_hd__nand2b_1 U28833 ( .A_N(n23826), .B(n23778), .Y(n23779) );
  sky130_fd_sc_hd__nand2b_1 U28835 ( .A_N(n23826), .B(n23783), .Y(n23784) );
  sky130_fd_sc_hd__nand2_1 U28836 ( .A(n23785), .B(n23784), .Y(n25982) );
  sky130_fd_sc_hd__inv_2 U28837 ( .A(n25982), .Y(n27837) );
  sky130_fd_sc_hd__nand3_1 U28838 ( .A(n23786), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__2_), .C(
        j202_soc_core_j22_cpu_regop_M_Rn__3_), .Y(n23849) );
  sky130_fd_sc_hd__nand2b_1 U28839 ( .A_N(n23841), .B(n23787), .Y(n23791) );
  sky130_fd_sc_hd__nand2b_1 U28840 ( .A_N(n23826), .B(n23789), .Y(n23790) );
  sky130_fd_sc_hd__nand2b_1 U28841 ( .A_N(n23841), .B(n23792), .Y(n23796) );
  sky130_fd_sc_hd__nand2b_1 U28842 ( .A_N(n23826), .B(n23794), .Y(n23795) );
  sky130_fd_sc_hd__nand2b_1 U28843 ( .A_N(n23841), .B(n15017), .Y(n23800) );
  sky130_fd_sc_hd__nand2b_1 U28844 ( .A_N(n23826), .B(n23798), .Y(n23799) );
  sky130_fd_sc_hd__nand2b_1 U28846 ( .A_N(n23841), .B(n23802), .Y(n23806) );
  sky130_fd_sc_hd__nand2b_1 U28847 ( .A_N(n23826), .B(n23804), .Y(n23805) );
  sky130_fd_sc_hd__nand2b_1 U28849 ( .A_N(n23841), .B(n23808), .Y(n23812) );
  sky130_fd_sc_hd__nand2b_1 U28850 ( .A_N(n23826), .B(n23810), .Y(n23811) );
  sky130_fd_sc_hd__nand2b_1 U28851 ( .A_N(n23841), .B(n14275), .Y(n23817) );
  sky130_fd_sc_hd__nand2b_1 U28852 ( .A_N(n23826), .B(n23815), .Y(n23816) );
  sky130_fd_sc_hd__nand2b_1 U28854 ( .A_N(n23841), .B(n15950), .Y(n23822) );
  sky130_fd_sc_hd__nand2b_1 U28855 ( .A_N(n23826), .B(n23820), .Y(n23821) );
  sky130_fd_sc_hd__nand2b_1 U28856 ( .A_N(n23841), .B(n23823), .Y(n23828) );
  sky130_fd_sc_hd__nand2b_1 U28857 ( .A_N(n23826), .B(n23825), .Y(n23827) );
  sky130_fd_sc_hd__nor3_1 U28858 ( .A(n23831), .B(n23830), .C(n24673), .Y(
        n24681) );
  sky130_fd_sc_hd__nand2_1 U28859 ( .A(n28109), .B(n12347), .Y(n23845) );
  sky130_fd_sc_hd__nand2_1 U28860 ( .A(n23892), .B(n23832), .Y(n23833) );
  sky130_fd_sc_hd__o211ai_2 U28861 ( .A1(n23835), .A2(n23834), .B1(n23833), 
        .C1(n27847), .Y(j202_soc_core_j22_cpu_rf_N2709) );
  sky130_fd_sc_hd__nand2_1 U28862 ( .A(n28109), .B(n23836), .Y(n23838) );
  sky130_fd_sc_hd__nor2_1 U28863 ( .A(j202_soc_core_j22_cpu_regop_We__0_), .B(
        n12347), .Y(n23837) );
  sky130_fd_sc_hd__nand4_1 U28864 ( .A(n23892), .B(
        j202_soc_core_j22_cpu_regop_M_Wm__2_), .C(n23840), .D(n24717), .Y(
        n23848) );
  sky130_fd_sc_hd__nand2b_1 U28865 ( .A_N(n23841), .B(n13820), .Y(n23847) );
  sky130_fd_sc_hd__a21oi_1 U28866 ( .A1(n23843), .A2(
        j202_soc_core_j22_cpu_regop_We__0_), .B1(n23842), .Y(n23844) );
  sky130_fd_sc_hd__nand2b_1 U28867 ( .A_N(n23845), .B(n23844), .Y(n23846) );
  sky130_fd_sc_hd__nor2_1 U28868 ( .A(n23852), .B(n23851), .Y(n26660) );
  sky130_fd_sc_hd__nand3_1 U28869 ( .A(n26568), .B(n23853), .C(
        j202_soc_core_wbqspiflash_00_lldriver_state[0]), .Y(n26661) );
  sky130_fd_sc_hd__nand3_1 U28870 ( .A(n26660), .B(n29183), .C(n26661), .Y(
        n26567) );
  sky130_fd_sc_hd__nand2_1 U28871 ( .A(n28895), .B(n26661), .Y(n23855) );
  sky130_fd_sc_hd__nand2_1 U28872 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B(n26569), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N423) );
  sky130_fd_sc_hd__nand3_1 U28874 ( .A(n23882), .B(
        j202_soc_core_gpio_core_00_reg_addr[2]), .C(n26910), .Y(n26905) );
  sky130_fd_sc_hd__o21ai_1 U28875 ( .A1(n26783), .A2(n26905), .B1(n29827), .Y(
        n10712) );
  sky130_fd_sc_hd__nor2_1 U28876 ( .A(j202_soc_core_gpio_core_00_reg_addr[4]), 
        .B(n23856), .Y(n23857) );
  sky130_fd_sc_hd__nand3_1 U28877 ( .A(n23882), .B(n23857), .C(n26908), .Y(
        n26907) );
  sky130_fd_sc_hd__o21ai_1 U28878 ( .A1(n26783), .A2(n26907), .B1(n29827), .Y(
        n10714) );
  sky130_fd_sc_hd__nand2_1 U28879 ( .A(n23898), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_cs_n), .Y(n23859) );
  sky130_fd_sc_hd__nand2_1 U28880 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .B(
        j202_soc_core_wbqspiflash_00_alt_cmd), .Y(n23858) );
  sky130_fd_sc_hd__nand2_1 U28881 ( .A(n23859), .B(n23858), .Y(io_out[8]) );
  sky130_fd_sc_hd__nand3_1 U28882 ( .A(n28669), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .C(
        j202_soc_core_wbqspiflash_00_state[2]), .Y(n26640) );
  sky130_fd_sc_hd__nand2_1 U28883 ( .A(j202_soc_core_wbqspiflash_00_state[2]), 
        .B(j202_soc_core_wbqspiflash_00_state[4]), .Y(n27264) );
  sky130_fd_sc_hd__nor2_1 U28884 ( .A(n27264), .B(n26483), .Y(n28861) );
  sky130_fd_sc_hd__nand2_1 U28885 ( .A(n26558), .B(n26623), .Y(n26612) );
  sky130_fd_sc_hd__nor3_1 U28886 ( .A(n26633), .B(n26588), .C(n26612), .Y(
        n23864) );
  sky130_fd_sc_hd__nand2_1 U28887 ( .A(n23860), .B(n23862), .Y(n27430) );
  sky130_fd_sc_hd__nand2_1 U28888 ( .A(j202_soc_core_wbqspiflash_00_spif_cmd), 
        .B(j202_soc_core_wbqspiflash_00_spif_ctrl), .Y(n26532) );
  sky130_fd_sc_hd__nand2_1 U28889 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .Y(n26485) );
  sky130_fd_sc_hd__nand3_1 U28890 ( .A(n27430), .B(n23861), .C(n26485), .Y(
        n27275) );
  sky130_fd_sc_hd__o211ai_1 U28891 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[31]), .B1(n23862), .C1(n23861), 
        .Y(n27233) );
  sky130_fd_sc_hd__nor2_1 U28892 ( .A(j202_soc_core_wbqspiflash_00_spif_cmd), 
        .B(n26481), .Y(n28837) );
  sky130_fd_sc_hd__nand2_1 U28893 ( .A(n28837), .B(n27430), .Y(n23863) );
  sky130_fd_sc_hd__and3_1 U28894 ( .A(n27275), .B(n27233), .C(n23863), .X(
        n26587) );
  sky130_fd_sc_hd__nand2_1 U28895 ( .A(n26481), .B(
        j202_soc_core_wbqspiflash_00_spif_cmd), .Y(n27251) );
  sky130_fd_sc_hd__nor2_1 U28896 ( .A(
        j202_soc_core_wbqspiflash_00_write_protect), .B(n27251), .Y(n27271) );
  sky130_fd_sc_hd__nand2_1 U28897 ( .A(n27271), .B(n27614), .Y(n27203) );
  sky130_fd_sc_hd__nand2_1 U28898 ( .A(n26587), .B(n27203), .Y(n26631) );
  sky130_fd_sc_hd__nand2_1 U28899 ( .A(n26623), .B(
        j202_soc_core_wbqspiflash_00_state[4]), .Y(n26634) );
  sky130_fd_sc_hd__a21oi_1 U28900 ( .A1(n23864), .A2(n26631), .B1(n23878), .Y(
        n23865) );
  sky130_fd_sc_hd__a21oi_1 U28901 ( .A1(n23865), .A2(n26479), .B1(n26483), .Y(
        n23868) );
  sky130_fd_sc_hd__nand2_1 U28902 ( .A(n28840), .B(
        j202_soc_core_ahb2wbqspi_00_stb_o), .Y(n23867) );
  sky130_fd_sc_hd__nor2_1 U28903 ( .A(j202_soc_core_qspi_wb_we), .B(n27229), 
        .Y(n28841) );
  sky130_fd_sc_hd__nor4_1 U28904 ( .A(n23867), .B(n27254), .C(n28841), .D(
        n23866), .Y(n26635) );
  sky130_fd_sc_hd__nor4_1 U28905 ( .A(n25344), .B(n28861), .C(n23868), .D(
        n26635), .Y(n23870) );
  sky130_fd_sc_hd__nand2_1 U28906 ( .A(n23869), .B(n28841), .Y(n28817) );
  sky130_fd_sc_hd__nor2_1 U28907 ( .A(n28647), .B(n26483), .Y(n28688) );
  sky130_fd_sc_hd__nand2_1 U28908 ( .A(n28688), .B(n27284), .Y(n27190) );
  sky130_fd_sc_hd__nand3_1 U28909 ( .A(n23870), .B(n28817), .C(n27190), .Y(
        n26502) );
  sky130_fd_sc_hd__nor2_1 U28910 ( .A(n27268), .B(n27280), .Y(n27208) );
  sky130_fd_sc_hd__nand2_1 U28911 ( .A(n26588), .B(n28647), .Y(n27181) );
  sky130_fd_sc_hd__nor2_1 U28912 ( .A(j202_soc_core_wbqspiflash_00_state[1]), 
        .B(n27181), .Y(n27211) );
  sky130_fd_sc_hd__nand2_1 U28913 ( .A(n27211), .B(
        j202_soc_core_wbqspiflash_00_state[3]), .Y(n25342) );
  sky130_fd_sc_hd__nand2_1 U28914 ( .A(n26588), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n27286) );
  sky130_fd_sc_hd__nand2_1 U28915 ( .A(n26486), .B(
        j202_soc_core_wbqspiflash_00_state[3]), .Y(n26506) );
  sky130_fd_sc_hd__nand2_1 U28916 ( .A(n25342), .B(n26506), .Y(n25206) );
  sky130_fd_sc_hd__nor2_1 U28917 ( .A(n27208), .B(n25206), .Y(n26583) );
  sky130_fd_sc_hd__nand3_1 U28918 ( .A(n27226), .B(n28866), .C(
        j202_soc_core_wbqspiflash_00_write_in_progress), .Y(n27289) );
  sky130_fd_sc_hd__nand2_1 U28919 ( .A(n27288), .B(n27289), .Y(n28842) );
  sky130_fd_sc_hd__nand2_1 U28920 ( .A(j202_soc_core_qspi_wb_addr[3]), .B(
        j202_soc_core_qspi_wb_addr[2]), .Y(n28867) );
  sky130_fd_sc_hd__nor2_1 U28921 ( .A(n27238), .B(n23871), .Y(n27193) );
  sky130_fd_sc_hd__nand2_1 U28922 ( .A(n27193), .B(n23872), .Y(n26546) );
  sky130_fd_sc_hd__nor2_1 U28923 ( .A(n26490), .B(n26546), .Y(n26585) );
  sky130_fd_sc_hd__a21oi_1 U28924 ( .A1(n28842), .A2(n27293), .B1(n26585), .Y(
        n23876) );
  sky130_fd_sc_hd__nand2_1 U28925 ( .A(n27193), .B(
        j202_soc_core_qspi_wb_wdat[31]), .Y(n27294) );
  sky130_fd_sc_hd__nand2_1 U28927 ( .A(n23873), .B(n27407), .Y(n23874) );
  sky130_fd_sc_hd__nand3_1 U28928 ( .A(n23874), .B(n23876), .C(n25345), .Y(
        n26616) );
  sky130_fd_sc_hd__a21oi_1 U28929 ( .A1(n23876), .A2(
        j202_soc_core_wbqspiflash_00_write_in_progress), .B1(n23875), .Y(
        n26497) );
  sky130_fd_sc_hd__nor2_1 U28930 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(n27183), .Y(n27298) );
  sky130_fd_sc_hd__a21oi_1 U28931 ( .A1(n26534), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .B1(n26481), .Y(n28859)
         );
  sky130_fd_sc_hd__nor2_1 U28932 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(j202_soc_core_wbqspiflash_00_state[3]), .Y(n23877) );
  sky130_fd_sc_hd__and3_1 U28933 ( .A(io_out[8]), .B(n23878), .C(n23877), .X(
        n26482) );
  sky130_fd_sc_hd__nand2_1 U28934 ( .A(n26482), .B(
        j202_soc_core_wbqspiflash_00_state[1]), .Y(n26504) );
  sky130_fd_sc_hd__nand2_1 U28935 ( .A(n28647), .B(
        j202_soc_core_wbqspiflash_00_state[2]), .Y(n27279) );
  sky130_fd_sc_hd__nand2_1 U28936 ( .A(n26484), .B(n28870), .Y(n27257) );
  sky130_fd_sc_hd__o21ai_1 U28937 ( .A1(n28859), .A2(n26504), .B1(n27257), .Y(
        n23879) );
  sky130_fd_sc_hd__a21oi_1 U28938 ( .A1(n26497), .A2(n27298), .B1(n23879), .Y(
        n26649) );
  sky130_fd_sc_hd__nand2_1 U28939 ( .A(n26908), .B(
        j202_soc_core_gpio_core_00_reg_addr[4]), .Y(n26904) );
  sky130_fd_sc_hd__nand3_1 U28940 ( .A(n23882), .B(n23881), .C(
        j202_soc_core_gpio_core_00_reg_addr[2]), .Y(n26901) );
  sky130_fd_sc_hd__o21ai_1 U28941 ( .A1(n26783), .A2(n26901), .B1(n29830), .Y(
        n10711) );
  sky130_fd_sc_hd__nor2_1 U28942 ( .A(j202_soc_core_j22_cpu_rte4), .B(n23887), 
        .Y(n23884) );
  sky130_fd_sc_hd__and3_1 U28943 ( .A(n23885), .B(n23884), .C(n23883), .X(
        n23886) );
  sky130_fd_sc_hd__nand3_1 U28944 ( .A(n24710), .B(n23886), .C(n24704), .Y(
        n24039) );
  sky130_fd_sc_hd__nor2_1 U28945 ( .A(n29088), .B(n23887), .Y(n24032) );
  sky130_fd_sc_hd__nand2_1 U28946 ( .A(n24176), .B(n23888), .Y(n23890) );
  sky130_fd_sc_hd__nand3_1 U28947 ( .A(n28109), .B(
        j202_soc_core_j22_cpu_regop_We__2_), .C(n23889), .Y(n27364) );
  sky130_fd_sc_hd__nand2_1 U28948 ( .A(n23890), .B(n27364), .Y(n24040) );
  sky130_fd_sc_hd__o22ai_1 U28949 ( .A1(n23892), .A2(n27855), .B1(n23891), 
        .B2(n24040), .Y(n23893) );
  sky130_fd_sc_hd__nand2_1 U28950 ( .A(j202_soc_core_uart_TOP_rx_go), .B(
        j202_soc_core_uart_TOP_rx_sio_ce), .Y(n28593) );
  sky130_fd_sc_hd__nor2_1 U28952 ( .A(j202_soc_core_uart_TOP_rx_valid_r), .B(
        n23897), .Y(n27958) );
  sky130_fd_sc_hd__and3_1 U28953 ( .A(n27958), .B(
        j202_soc_core_uart_TOP_rx_fifo_wp[0]), .C(
        j202_soc_core_uart_TOP_rx_fifo_wp[1]), .X(n29723) );
  sky130_fd_sc_hd__nand2_1 U28954 ( .A(n27958), .B(
        j202_soc_core_uart_TOP_rx_fifo_wp[0]), .Y(n27954) );
  sky130_fd_sc_hd__nor2_1 U28955 ( .A(j202_soc_core_uart_TOP_rx_fifo_wp[1]), 
        .B(n27954), .Y(n29870) );
  sky130_fd_sc_hd__nor2b_1 U28956 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[25]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N28) );
  sky130_fd_sc_hd__nor2b_1 U28957 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[31]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N34) );
  sky130_fd_sc_hd__nor2b_1 U28958 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[23]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N26) );
  sky130_fd_sc_hd__nor2b_1 U28959 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[26]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N29) );
  sky130_fd_sc_hd__nor2b_1 U28960 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[21]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N24) );
  sky130_fd_sc_hd__nor2b_1 U28961 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[10]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N13) );
  sky130_fd_sc_hd__nor2b_1 U28962 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[14]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N17) );
  sky130_fd_sc_hd__nor2b_1 U28963 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[29]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N32) );
  sky130_fd_sc_hd__nor2b_1 U28964 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[6]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N9) );
  sky130_fd_sc_hd__nand3_1 U28965 ( .A(n28910), .B(
        j202_soc_core_uart_TOP_tx_fifo_wp[0]), .C(j202_soc_core_uart_WRTXD1), 
        .Y(n27922) );
  sky130_fd_sc_hd__nor2_1 U28966 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[1]), 
        .B(n27922), .Y(n29880) );
  sky130_fd_sc_hd__nor2b_1 U28967 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[11]), .A(n29088), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N14) );
  sky130_fd_sc_hd__nor2b_1 U28968 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[1]), .A(n29088), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N4) );
  sky130_fd_sc_hd__nor2b_1 U28969 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[7]), .A(n29088), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N10) );
  sky130_fd_sc_hd__nor2b_1 U28970 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[20]), .A(n29088), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N23) );
  sky130_fd_sc_hd__nor2b_1 U28971 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[8]), .A(n29088), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N11) );
  sky130_fd_sc_hd__nor2b_1 U28972 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[15]), .A(n29088), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N18) );
  sky130_fd_sc_hd__nor2b_1 U28973 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[13]), .A(n29088), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N16) );
  sky130_fd_sc_hd__nor2b_1 U28974 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[3]), .A(n29088), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N6) );
  sky130_fd_sc_hd__nor2b_1 U28975 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[19]), .A(n29088), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N22) );
  sky130_fd_sc_hd__nor2b_1 U28976 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[2]), .A(n29088), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N5) );
  sky130_fd_sc_hd__nor2b_1 U28977 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[5]), .A(n29088), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N8) );
  sky130_fd_sc_hd__nor2b_1 U28978 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[12]), .A(n29088), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N15) );
  sky130_fd_sc_hd__nor2b_1 U28979 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[16]), .A(n29088), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N19) );
  sky130_fd_sc_hd__nor2b_1 U28980 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[0]), .A(n29088), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N3) );
  sky130_fd_sc_hd__nor2b_1 U28981 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[4]), .A(n29088), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N7) );
  sky130_fd_sc_hd__nor2b_1 U28982 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[17]), .A(n29088), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N20) );
  sky130_fd_sc_hd__nor2b_1 U28983 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[22]), .A(n29088), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N25) );
  sky130_fd_sc_hd__nor2b_1 U28984 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[18]), .A(n29088), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N21) );
  sky130_fd_sc_hd__nor2b_1 U28985 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[9]), .A(n29088), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N12) );
  sky130_fd_sc_hd__nor2b_1 U28986 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[30]), .A(n29088), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N33) );
  sky130_fd_sc_hd__nor2b_1 U28987 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[27]), .A(n29088), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N30) );
  sky130_fd_sc_hd__nor2b_1 U28988 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[24]), .A(n29088), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N27) );
  sky130_fd_sc_hd__nor2b_1 U28989 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[28]), .A(n29088), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N31) );
  sky130_fd_sc_hd__nand3_1 U28990 ( .A(n23899), .B(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[1]), .C(
        j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_2), .Y(n24022) );
  sky130_fd_sc_hd__nor2_1 U28991 ( .A(j202_soc_core_cmt_core_00_reg_addr[1]), 
        .B(j202_soc_core_cmt_core_00_reg_addr[7]), .Y(n23902) );
  sky130_fd_sc_hd__nand3_1 U28992 ( .A(n23902), .B(n23901), .C(n23900), .Y(
        n24020) );
  sky130_fd_sc_hd__nand3_1 U28993 ( .A(n23903), .B(
        j202_soc_core_cmt_core_00_reg_addr[4]), .C(n24019), .Y(n24750) );
  sky130_fd_sc_hd__nor2_1 U28994 ( .A(n24022), .B(n24750), .Y(n24736) );
  sky130_fd_sc_hd__nand3_1 U28995 ( .A(n28222), .B(n28221), .C(n24736), .Y(
        n27530) );
  sky130_fd_sc_hd__nor2_1 U28996 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[2]), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[8]), .Y(n23905) );
  sky130_fd_sc_hd__and3_1 U28997 ( .A(n23905), .B(n23904), .C(n28566), .X(
        n23916) );
  sky130_fd_sc_hd__nor2_1 U28998 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[4]), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[6]), .Y(n23915) );
  sky130_fd_sc_hd__a22oi_1 U28999 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[9]), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[5]), .B1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[7]), .B2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[3]), .Y(n23912) );
  sky130_fd_sc_hd__nand3_1 U29000 ( .A(n23906), .B(n28575), .C(n28571), .Y(
        n23911) );
  sky130_fd_sc_hd__nand3_1 U29001 ( .A(n23907), .B(n28580), .C(
        j202_soc_core_cmt_core_00_cks1[1]), .Y(n23910) );
  sky130_fd_sc_hd__and4_1 U29003 ( .A(n23912), .B(n23911), .C(n23910), .D(
        n23909), .X(n23914) );
  sky130_fd_sc_hd__nand4_1 U29005 ( .A(n23916), .B(n23915), .C(n23914), .D(
        n23913), .Y(n23943) );
  sky130_fd_sc_hd__nor2_1 U29006 ( .A(n27544), .B(n23943), .Y(n27514) );
  sky130_fd_sc_hd__xor2_1 U29007 ( .A(j202_soc_core_cmt_core_00_const1[7]), 
        .B(j202_soc_core_cmt_core_00_cnt1[7]), .X(n23934) );
  sky130_fd_sc_hd__xnor2_1 U29008 ( .A(j202_soc_core_cmt_core_00_const1[15]), 
        .B(j202_soc_core_cmt_core_00_cnt1[15]), .Y(n23919) );
  sky130_fd_sc_hd__xnor2_1 U29009 ( .A(j202_soc_core_cmt_core_00_const1[11]), 
        .B(j202_soc_core_cmt_core_00_cnt1[11]), .Y(n23918) );
  sky130_fd_sc_hd__xnor2_1 U29010 ( .A(j202_soc_core_cmt_core_00_const1[2]), 
        .B(j202_soc_core_cmt_core_00_cnt1[2]), .Y(n23917) );
  sky130_fd_sc_hd__nand3_1 U29011 ( .A(n23919), .B(n23918), .C(n23917), .Y(
        n23933) );
  sky130_fd_sc_hd__xor2_1 U29012 ( .A(j202_soc_core_cmt_core_00_const1[14]), 
        .B(j202_soc_core_cmt_core_00_cnt1[14]), .X(n23921) );
  sky130_fd_sc_hd__xor2_1 U29013 ( .A(j202_soc_core_cmt_core_00_const1[0]), 
        .B(j202_soc_core_cmt_core_00_cnt1[0]), .X(n23920) );
  sky130_fd_sc_hd__nor2_1 U29014 ( .A(n23921), .B(n23920), .Y(n23931) );
  sky130_fd_sc_hd__xnor2_1 U29015 ( .A(j202_soc_core_cmt_core_00_const1[10]), 
        .B(j202_soc_core_cmt_core_00_cnt1[10]), .Y(n23923) );
  sky130_fd_sc_hd__xnor2_1 U29016 ( .A(j202_soc_core_cmt_core_00_const1[5]), 
        .B(j202_soc_core_cmt_core_00_cnt1[5]), .Y(n23922) );
  sky130_fd_sc_hd__xnor2_1 U29017 ( .A(j202_soc_core_cmt_core_00_const1[3]), 
        .B(j202_soc_core_cmt_core_00_cnt1[3]), .Y(n23925) );
  sky130_fd_sc_hd__xnor2_1 U29018 ( .A(j202_soc_core_cmt_core_00_const1[4]), 
        .B(j202_soc_core_cmt_core_00_cnt1[4]), .Y(n23924) );
  sky130_fd_sc_hd__xnor2_1 U29019 ( .A(j202_soc_core_cmt_core_00_const1[12]), 
        .B(j202_soc_core_cmt_core_00_cnt1[12]), .Y(n23927) );
  sky130_fd_sc_hd__xnor2_1 U29020 ( .A(j202_soc_core_cmt_core_00_const1[1]), 
        .B(j202_soc_core_cmt_core_00_cnt1[1]), .Y(n23926) );
  sky130_fd_sc_hd__nand4_1 U29021 ( .A(n23931), .B(n23930), .C(n23929), .D(
        n23928), .Y(n23932) );
  sky130_fd_sc_hd__nor3_1 U29022 ( .A(n23934), .B(n23933), .C(n23932), .Y(
        n23940) );
  sky130_fd_sc_hd__xor2_1 U29023 ( .A(j202_soc_core_cmt_core_00_const1[13]), 
        .B(j202_soc_core_cmt_core_00_cnt1[13]), .X(n23936) );
  sky130_fd_sc_hd__xor2_1 U29024 ( .A(j202_soc_core_cmt_core_00_const1[6]), 
        .B(j202_soc_core_cmt_core_00_cnt1[6]), .X(n23935) );
  sky130_fd_sc_hd__nor2_1 U29025 ( .A(n23936), .B(n23935), .Y(n23939) );
  sky130_fd_sc_hd__xnor2_1 U29026 ( .A(j202_soc_core_cmt_core_00_const1[9]), 
        .B(j202_soc_core_cmt_core_00_cnt1[9]), .Y(n23938) );
  sky130_fd_sc_hd__xnor2_1 U29027 ( .A(j202_soc_core_cmt_core_00_const1[8]), 
        .B(j202_soc_core_cmt_core_00_cnt1[8]), .Y(n23937) );
  sky130_fd_sc_hd__nand4_1 U29028 ( .A(n23940), .B(n23939), .C(n23938), .D(
        n23937), .Y(n29170) );
  sky130_fd_sc_hd__nand2_1 U29029 ( .A(j202_soc_core_cmt_core_00_cnt1[3]), .B(
        j202_soc_core_cmt_core_00_cnt1[2]), .Y(n23941) );
  sky130_fd_sc_hd__nand2_1 U29030 ( .A(j202_soc_core_cmt_core_00_cnt1[0]), .B(
        j202_soc_core_cmt_core_00_cnt1[1]), .Y(n27523) );
  sky130_fd_sc_hd__nor2_1 U29031 ( .A(n23941), .B(n27523), .Y(n27537) );
  sky130_fd_sc_hd__nand3_1 U29032 ( .A(n27537), .B(
        j202_soc_core_cmt_core_00_cnt1[4]), .C(
        j202_soc_core_cmt_core_00_cnt1[5]), .Y(n27536) );
  sky130_fd_sc_hd__o21ai_1 U29033 ( .A1(n27540), .A2(n27536), .B1(n23942), .Y(
        n23944) );
  sky130_fd_sc_hd__nor2_1 U29034 ( .A(n23942), .B(n27536), .Y(n24971) );
  sky130_fd_sc_hd__nand2_1 U29035 ( .A(n27530), .B(n23943), .Y(n28583) );
  sky130_fd_sc_hd__o2bb2ai_1 U29037 ( .B1(n27530), .B2(n27465), .A1_N(n23944), 
        .A2_N(n27545), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[6])
         );
  sky130_fd_sc_hd__nand2_1 U29038 ( .A(n29745), .B(
        j202_soc_core_wbqspiflash_00_spi_valid), .Y(n27306) );
  sky130_fd_sc_hd__nand2_1 U29039 ( .A(n26559), .B(
        j202_soc_core_wbqspiflash_00_spi_wr), .Y(n27246) );
  sky130_fd_sc_hd__o31ai_2 U29040 ( .A1(n27306), .A2(n26597), .A3(n27246), 
        .B1(n23945), .Y(n29630) );
  sky130_fd_sc_hd__nand2b_1 U29041 ( .A_N(n28155), .B(
        j202_soc_core_j22_cpu_opst[2]), .Y(n24686) );
  sky130_fd_sc_hd__nor2_1 U29042 ( .A(n23947), .B(n23946), .Y(n23953) );
  sky130_fd_sc_hd__nor2_1 U29043 ( .A(n23949), .B(n23948), .Y(n23952) );
  sky130_fd_sc_hd__nand3_1 U29044 ( .A(n23952), .B(n11172), .C(n23951), .Y(
        n24576) );
  sky130_fd_sc_hd__nor2_1 U29045 ( .A(n23953), .B(n24576), .Y(n28142) );
  sky130_fd_sc_hd__nand2_1 U29046 ( .A(n12669), .B(n24574), .Y(n23954) );
  sky130_fd_sc_hd__nor2_1 U29047 ( .A(n23954), .B(n24573), .Y(n23958) );
  sky130_fd_sc_hd__a21oi_1 U29048 ( .A1(n11729), .A2(n28133), .B1(n28091), .Y(
        n23956) );
  sky130_fd_sc_hd__nand4_1 U29049 ( .A(n23956), .B(n27729), .C(n28259), .D(
        n27736), .Y(n23957) );
  sky130_fd_sc_hd__nor2_1 U29050 ( .A(n23958), .B(n23957), .Y(n23959) );
  sky130_fd_sc_hd__o2bb2ai_1 U29051 ( .B1(n28355), .B2(n24686), .A1_N(n28417), 
        .A2_N(n23960), .Y(n10636) );
  sky130_fd_sc_hd__nor2_1 U29052 ( .A(n12040), .B(n24587), .Y(n23970) );
  sky130_fd_sc_hd__nand3_1 U29053 ( .A(n23961), .B(n12040), .C(n24587), .Y(
        n23972) );
  sky130_fd_sc_hd__o22ai_1 U29054 ( .A1(n23970), .A2(n23962), .B1(
        j202_soc_core_j22_cpu_memop_MEM__1_), .B2(n29581), .Y(n23964) );
  sky130_fd_sc_hd__nand2_1 U29055 ( .A(n23964), .B(n23963), .Y(n25480) );
  sky130_fd_sc_hd__o21a_1 U29056 ( .A1(n29565), .A2(n29581), .B1(n25480), .X(
        n23965) );
  sky130_fd_sc_hd__o21a_1 U29057 ( .A1(n27090), .A2(n29581), .B1(n25480), .X(
        n23967) );
  sky130_fd_sc_hd__nor2_1 U29059 ( .A(n23970), .B(n23969), .Y(n23971) );
  sky130_fd_sc_hd__a21oi_1 U29061 ( .A1(n29581), .A2(n23973), .B1(n24302), .Y(
        n23974) );
  sky130_fd_sc_hd__nand2_1 U29062 ( .A(n23975), .B(n23974), .Y(n27914) );
  sky130_fd_sc_hd__a21oi_1 U29063 ( .A1(n27090), .A2(n29581), .B1(n27914), .Y(
        n23976) );
  sky130_fd_sc_hd__a21oi_1 U29064 ( .A1(n29581), .A2(n29565), .B1(n27914), .Y(
        n23978) );
  sky130_fd_sc_hd__nand2_1 U29066 ( .A(n29879), .B(n28109), .Y(n23990) );
  sky130_fd_sc_hd__nor2b_1 U29067 ( .B_N(j202_soc_core_j22_cpu_regop_Wm__1_), 
        .A(n23990), .Y(j202_soc_core_j22_cpu_id_idec_N957) );
  sky130_fd_sc_hd__nor2b_1 U29068 ( .B_N(j202_soc_core_j22_cpu_regop_Wm__3_), 
        .A(n23990), .Y(j202_soc_core_j22_cpu_id_idec_N959) );
  sky130_fd_sc_hd__nor2b_1 U29069 ( .B_N(j202_soc_core_j22_cpu_regop_Wm__0_), 
        .A(n23990), .Y(j202_soc_core_j22_cpu_id_idec_N956) );
  sky130_fd_sc_hd__nor2b_1 U29070 ( .B_N(j202_soc_core_j22_cpu_regop_Wm__2_), 
        .A(n23990), .Y(j202_soc_core_j22_cpu_id_idec_N958) );
  sky130_fd_sc_hd__nand2_1 U29071 ( .A(n27219), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n27231) );
  sky130_fd_sc_hd__nor2_1 U29072 ( .A(n25205), .B(n27231), .Y(n28814) );
  sky130_fd_sc_hd__nand2_1 U29073 ( .A(n23991), .B(n29827), .Y(
        j202_soc_core_wbqspiflash_00_N710) );
  sky130_fd_sc_hd__nand2_1 U29074 ( .A(n29485), .B(n29828), .Y(n23992) );
  sky130_fd_sc_hd__nor2b_1 U29075 ( .B_N(j202_soc_core_prdata[8]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N136) );
  sky130_fd_sc_hd__nor2b_1 U29076 ( .B_N(j202_soc_core_prdata[0]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N128) );
  sky130_fd_sc_hd__nor2b_1 U29077 ( .B_N(j202_soc_core_prdata[3]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N131) );
  sky130_fd_sc_hd__nor2b_1 U29078 ( .B_N(j202_soc_core_prdata[7]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N135) );
  sky130_fd_sc_hd__nor2b_1 U29079 ( .B_N(j202_soc_core_prdata[11]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N139) );
  sky130_fd_sc_hd__nor2b_1 U29080 ( .B_N(j202_soc_core_prdata[14]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N142) );
  sky130_fd_sc_hd__nor2b_1 U29081 ( .B_N(j202_soc_core_prdata[10]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N138) );
  sky130_fd_sc_hd__nor2b_1 U29082 ( .B_N(j202_soc_core_prdata[1]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N129) );
  sky130_fd_sc_hd__nor2b_1 U29083 ( .B_N(j202_soc_core_prdata[4]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N132) );
  sky130_fd_sc_hd__nor2b_1 U29084 ( .B_N(j202_soc_core_prdata[12]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N140) );
  sky130_fd_sc_hd__nor2b_1 U29085 ( .B_N(j202_soc_core_prdata[2]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N130) );
  sky130_fd_sc_hd__nor2b_1 U29086 ( .B_N(j202_soc_core_prdata[15]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N143) );
  sky130_fd_sc_hd__nor2b_1 U29087 ( .B_N(j202_soc_core_prdata[13]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N141) );
  sky130_fd_sc_hd__nor2b_1 U29088 ( .B_N(j202_soc_core_prdata[5]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N133) );
  sky130_fd_sc_hd__nor2b_1 U29089 ( .B_N(j202_soc_core_prdata[6]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N134) );
  sky130_fd_sc_hd__nor2b_1 U29090 ( .B_N(j202_soc_core_prdata[9]), .A(n23992), 
        .Y(j202_soc_core_ahb2apb_00_N137) );
  sky130_fd_sc_hd__inv_1 U29091 ( .A(n24400), .Y(n23993) );
  sky130_fd_sc_hd__nand3_1 U29092 ( .A(n12232), .B(n12254), .C(n11423), .Y(
        n23995) );
  sky130_fd_sc_hd__nand4_1 U29093 ( .A(n28029), .B(n12399), .C(n23996), .D(
        n23995), .Y(n23997) );
  sky130_fd_sc_hd__o2bb2ai_1 U29094 ( .B1(n23998), .B2(n28405), .A1_N(n28417), 
        .A2_N(n23997), .Y(n10542) );
  sky130_fd_sc_hd__nor2_1 U29096 ( .A(n29088), .B(
        j202_soc_core_ahb2aqu_00_aqu_st_0_), .Y(n25030) );
  sky130_fd_sc_hd__nand2b_1 U29097 ( .A_N(n25478), .B(n25030), .Y(
        j202_soc_core_ahb2aqu_00_N95) );
  sky130_fd_sc_hd__nor2_1 U29098 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[1]), 
        .B(n29172), .Y(n28589) );
  sky130_fd_sc_hd__nor2b_1 U29099 ( .B_N(j202_soc_core_uart_TOP_rx_bit_cnt[3]), 
        .A(j202_soc_core_uart_TOP_rx_bit_cnt[2]), .Y(n29173) );
  sky130_fd_sc_hd__nor2_1 U29100 ( .A(n29172), .B(n24000), .Y(n24001) );
  sky130_fd_sc_hd__nor2_1 U29101 ( .A(j202_soc_core_rst), .B(n28593), .Y(
        n24273) );
  sky130_fd_sc_hd__nand2_1 U29102 ( .A(n24001), .B(
        j202_soc_core_uart_TOP_rx_bit_cnt[2]), .Y(n28591) );
  sky130_fd_sc_hd__o211a_2 U29103 ( .A1(j202_soc_core_uart_TOP_rx_bit_cnt[2]), 
        .A2(n24001), .B1(n24273), .C1(n28591), .X(j202_soc_core_uart_TOP_N88)
         );
  sky130_fd_sc_hd__nand2_1 U29104 ( .A(j202_soc_core_uart_sio_ce), .B(
        j202_soc_core_uart_TOP_load), .Y(n29301) );
  sky130_fd_sc_hd__nand3_1 U29105 ( .A(j202_soc_core_uart_sio_ce), .B(
        j202_soc_core_uart_TOP_shift_en), .C(n29301), .Y(n28595) );
  sky130_fd_sc_hd__nand3_1 U29106 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[2]), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .C(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .Y(n24520) );
  sky130_fd_sc_hd__nor2_1 U29107 ( .A(n24521), .B(n24520), .Y(n24522) );
  sky130_fd_sc_hd__nand2_1 U29108 ( .A(n24522), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[4]), .Y(n24524) );
  sky130_fd_sc_hd__nor2_1 U29109 ( .A(n24525), .B(n24524), .Y(n24527) );
  sky130_fd_sc_hd__nand2_1 U29110 ( .A(n24527), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .Y(n24530) );
  sky130_fd_sc_hd__o211a_2 U29111 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .A2(n24527), .B1(
        n28547), .C1(n24530), .X(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[6]) );
  sky130_fd_sc_hd__nand2_1 U29112 ( .A(n27958), .B(n27955), .Y(n27953) );
  sky130_fd_sc_hd__nor2_1 U29113 ( .A(j202_soc_core_uart_TOP_rx_fifo_wp[1]), 
        .B(n27953), .Y(n29868) );
  sky130_fd_sc_hd__nor2_1 U29114 ( .A(n24002), .B(n27953), .Y(n29869) );
  sky130_fd_sc_hd__nand3_1 U29115 ( .A(n28910), .B(j202_soc_core_uart_WRTXD1), 
        .C(n27921), .Y(n24003) );
  sky130_fd_sc_hd__nor2_1 U29116 ( .A(n24004), .B(n24003), .Y(n29863) );
  sky130_fd_sc_hd__nor2_1 U29117 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[1]), 
        .B(n24003), .Y(n29865) );
  sky130_fd_sc_hd__nand2_1 U29118 ( .A(j202_soc_core_cmt_core_00_str1), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[0]), .Y(n28567) );
  sky130_fd_sc_hd__nor2_1 U29119 ( .A(n28566), .B(n28567), .Y(n28568) );
  sky130_fd_sc_hd__nand2_1 U29120 ( .A(n28568), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[2]), .Y(n28570) );
  sky130_fd_sc_hd__nor2_1 U29121 ( .A(n28571), .B(n28570), .Y(n28572) );
  sky130_fd_sc_hd__nand2_1 U29122 ( .A(n28572), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[4]), .Y(n28574) );
  sky130_fd_sc_hd__nor2_1 U29123 ( .A(n28575), .B(n28574), .Y(n28576) );
  sky130_fd_sc_hd__nand2_1 U29124 ( .A(n28576), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[6]), .Y(n28579) );
  sky130_fd_sc_hd__nor2_1 U29125 ( .A(n28580), .B(n28579), .Y(n28578) );
  sky130_fd_sc_hd__nand2_1 U29126 ( .A(n28578), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[8]), .Y(n28581) );
  sky130_fd_sc_hd__o211a_2 U29127 ( .A1(n28578), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[8]), .B1(n29171), .C1(
        n28581), .X(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[8]) );
  sky130_fd_sc_hd__nor2_1 U29128 ( .A(n24004), .B(n27922), .Y(n29864) );
  sky130_fd_sc_hd__nand2_1 U29129 ( .A(j202_soc_core_cmt_core_00_str0), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[0]), .Y(n28554) );
  sky130_fd_sc_hd__nor2_1 U29130 ( .A(n24269), .B(n28554), .Y(n24268) );
  sky130_fd_sc_hd__nand2_1 U29131 ( .A(n24268), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[2]), .Y(n24265) );
  sky130_fd_sc_hd__nor2_1 U29132 ( .A(n24266), .B(n24265), .Y(n24264) );
  sky130_fd_sc_hd__nand2_1 U29133 ( .A(n24264), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[4]), .Y(n28557) );
  sky130_fd_sc_hd__nor2_1 U29134 ( .A(n28558), .B(n28557), .Y(n28556) );
  sky130_fd_sc_hd__nand2_1 U29135 ( .A(n28556), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[6]), .Y(n28560) );
  sky130_fd_sc_hd__nor2_1 U29136 ( .A(n28561), .B(n28560), .Y(n28559) );
  sky130_fd_sc_hd__nor2_1 U29137 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[2]), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[8]), .Y(n24006) );
  sky130_fd_sc_hd__and3_1 U29138 ( .A(n24006), .B(n24005), .C(n24269), .X(
        n24017) );
  sky130_fd_sc_hd__nor2_1 U29139 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[4]), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[6]), .Y(n24016) );
  sky130_fd_sc_hd__a22oi_1 U29140 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[9]), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[5]), .B1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[7]), .B2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[3]), .Y(n24013) );
  sky130_fd_sc_hd__nand3_1 U29141 ( .A(n24007), .B(n28558), .C(n24266), .Y(
        n24012) );
  sky130_fd_sc_hd__nand3_1 U29142 ( .A(n24008), .B(n28561), .C(
        j202_soc_core_cmt_core_00_cks0[1]), .Y(n24011) );
  sky130_fd_sc_hd__and4_1 U29144 ( .A(n24013), .B(n24012), .C(n24011), .D(
        n24010), .X(n24015) );
  sky130_fd_sc_hd__nand4_1 U29146 ( .A(n24017), .B(n24016), .C(n24015), .D(
        n24014), .Y(n24979) );
  sky130_fd_sc_hd__nand2_1 U29147 ( .A(j202_soc_core_cmt_core_00_reg_addr[2]), 
        .B(j202_soc_core_cmt_core_00_reg_addr[3]), .Y(n24755) );
  sky130_fd_sc_hd__nand2_1 U29148 ( .A(n24019), .B(n24018), .Y(n24021) );
  sky130_fd_sc_hd__nor2_1 U29149 ( .A(n24021), .B(n24020), .Y(n24754) );
  sky130_fd_sc_hd__nand2_1 U29150 ( .A(n24754), .B(n24023), .Y(n28210) );
  sky130_fd_sc_hd__nor2_1 U29151 ( .A(n24024), .B(n27486), .Y(n29169) );
  sky130_fd_sc_hd__nand2_1 U29152 ( .A(n28559), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[8]), .Y(n28562) );
  sky130_fd_sc_hd__o211a_2 U29153 ( .A1(n28559), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[8]), .B1(n29169), .C1(
        n28562), .X(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[8]) );
  sky130_fd_sc_hd__nand2_1 U29154 ( .A(n24026), .B(n12069), .Y(
        j202_soc_core_ahb2apb_00_N127) );
  sky130_fd_sc_hd__nand2_1 U29155 ( .A(n24912), .B(n12069), .Y(n10603) );
  sky130_fd_sc_hd__nand2_1 U29156 ( .A(n24028), .B(n28367), .Y(n10601) );
  sky130_fd_sc_hd__nand2_1 U29157 ( .A(n24029), .B(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .Y(n26666) );
  sky130_fd_sc_hd__nand2_1 U29158 ( .A(n26666), .B(n29745), .Y(n29266) );
  sky130_fd_sc_hd__nand2_1 U29159 ( .A(n29267), .B(n26570), .Y(n29166) );
  sky130_fd_sc_hd__nand2_1 U29160 ( .A(n24031), .B(n24030), .Y(n26667) );
  sky130_fd_sc_hd__nand2_1 U29161 ( .A(n26667), .B(n26661), .Y(n29270) );
  sky130_fd_sc_hd__nand2_1 U29162 ( .A(n29166), .B(n28702), .Y(n26662) );
  sky130_fd_sc_hd__nand3_1 U29163 ( .A(n27219), .B(
        j202_soc_core_wbqspiflash_00_spi_valid), .C(n28780), .Y(n26557) );
  sky130_fd_sc_hd__nor2_1 U29164 ( .A(n26557), .B(n27267), .Y(n26576) );
  sky130_fd_sc_hd__nand2_1 U29165 ( .A(n28849), .B(
        j202_soc_core_wbqspiflash_00_state[4]), .Y(n27240) );
  sky130_fd_sc_hd__nor2_1 U29166 ( .A(n26612), .B(n27240), .Y(n26641) );
  sky130_fd_sc_hd__a211oi_1 U29167 ( .A1(n26467), .A2(n28647), .B1(n26576), 
        .C1(n26641), .Y(n27223) );
  sky130_fd_sc_hd__o22ai_1 U29168 ( .A1(n26516), .A2(n27306), .B1(n29088), 
        .B2(n27223), .Y(j202_soc_core_wbqspiflash_00_N749) );
  sky130_fd_sc_hd__nor2_1 U29169 ( .A(n28726), .B(n26661), .Y(n29184) );
  sky130_fd_sc_hd__nand2_1 U29170 ( .A(n29267), .B(
        j202_soc_core_wbqspiflash_00_spi_spd), .Y(n29196) );
  sky130_fd_sc_hd__nand2_1 U29171 ( .A(n28508), .B(n25724), .Y(n24043) );
  sky130_fd_sc_hd__nand2_1 U29172 ( .A(n24040), .B(n24032), .Y(n24037) );
  sky130_fd_sc_hd__a22oi_1 U29173 ( .A1(n26070), .A2(n28509), .B1(n24035), 
        .B2(n26068), .Y(n24042) );
  sky130_fd_sc_hd__nand2b_1 U29174 ( .A_N(n24037), .B(n24036), .Y(n24038) );
  sky130_fd_sc_hd__nand2_1 U29175 ( .A(n26071), .B(n27507), .Y(n24041) );
  sky130_fd_sc_hd__nand3_1 U29176 ( .A(n24043), .B(n24042), .C(n24041), .Y(
        j202_soc_core_j22_cpu_rf_N302) );
  sky130_fd_sc_hd__nand2_1 U29177 ( .A(n28501), .B(n25724), .Y(n24047) );
  sky130_fd_sc_hd__a22oi_1 U29178 ( .A1(n26070), .A2(n28502), .B1(n24044), 
        .B2(n26068), .Y(n24046) );
  sky130_fd_sc_hd__nand2_1 U29179 ( .A(n26071), .B(n24803), .Y(n24045) );
  sky130_fd_sc_hd__nand3_1 U29180 ( .A(n24047), .B(n24046), .C(n24045), .Y(
        j202_soc_core_j22_cpu_rf_N303) );
  sky130_fd_sc_hd__a22oi_1 U29181 ( .A1(n26070), .A2(n28521), .B1(n24048), 
        .B2(n26068), .Y(n24050) );
  sky130_fd_sc_hd__nand2_1 U29182 ( .A(n26071), .B(n27125), .Y(n24049) );
  sky130_fd_sc_hd__nand3_1 U29183 ( .A(n24051), .B(n24050), .C(n24049), .Y(
        j202_soc_core_j22_cpu_rf_N300) );
  sky130_fd_sc_hd__nand2_1 U29184 ( .A(n12431), .B(n25724), .Y(n24055) );
  sky130_fd_sc_hd__a22oi_1 U29185 ( .A1(n26070), .A2(n12354), .B1(n24052), 
        .B2(n26068), .Y(n24054) );
  sky130_fd_sc_hd__nand2_1 U29186 ( .A(n26071), .B(n24792), .Y(n24053) );
  sky130_fd_sc_hd__nand3_1 U29187 ( .A(n24055), .B(n24054), .C(n24053), .Y(
        j202_soc_core_j22_cpu_rf_N299) );
  sky130_fd_sc_hd__nand2_1 U29188 ( .A(n12402), .B(n25724), .Y(n24059) );
  sky130_fd_sc_hd__a22oi_1 U29189 ( .A1(n26070), .A2(n28495), .B1(n24056), 
        .B2(n26068), .Y(n24058) );
  sky130_fd_sc_hd__nand2_1 U29190 ( .A(n26071), .B(n25152), .Y(n24057) );
  sky130_fd_sc_hd__nand3_1 U29191 ( .A(n24059), .B(n24058), .C(n24057), .Y(
        j202_soc_core_j22_cpu_rf_N304) );
  sky130_fd_sc_hd__nand2_1 U29192 ( .A(n29486), .B(n25392), .Y(n24061) );
  sky130_fd_sc_hd__nand2_1 U29193 ( .A(n26191), .B(n25938), .Y(n24060) );
  sky130_fd_sc_hd__nand2_1 U29194 ( .A(n24061), .B(n24060), .Y(n24953) );
  sky130_fd_sc_hd__nand2_1 U29196 ( .A(n28483), .B(n25724), .Y(n24064) );
  sky130_fd_sc_hd__a22oi_1 U29197 ( .A1(n26070), .A2(n28484), .B1(n24947), 
        .B2(n26068), .Y(n24063) );
  sky130_fd_sc_hd__nand2_1 U29198 ( .A(n26071), .B(n26974), .Y(n24062) );
  sky130_fd_sc_hd__nand3_1 U29199 ( .A(n24064), .B(n24063), .C(n24062), .Y(
        j202_soc_core_j22_cpu_rf_N306) );
  sky130_fd_sc_hd__nand2_1 U29200 ( .A(n28459), .B(n25724), .Y(n24067) );
  sky130_fd_sc_hd__a22oi_1 U29201 ( .A1(n26070), .A2(n28460), .B1(n26016), 
        .B2(n26068), .Y(n24066) );
  sky130_fd_sc_hd__nand2_1 U29202 ( .A(n26071), .B(n26026), .Y(n24065) );
  sky130_fd_sc_hd__nand3_1 U29203 ( .A(n24067), .B(n24066), .C(n24065), .Y(
        j202_soc_core_j22_cpu_rf_N310) );
  sky130_fd_sc_hd__o22a_1 U29204 ( .A1(n24069), .A2(n12423), .B1(n25940), .B2(
        n12409), .X(n26187) );
  sky130_fd_sc_hd__nand2_1 U29205 ( .A(n28466), .B(n25724), .Y(n24073) );
  sky130_fd_sc_hd__a22oi_1 U29206 ( .A1(n26070), .A2(n28467), .B1(n25926), 
        .B2(n26068), .Y(n24072) );
  sky130_fd_sc_hd__nand2_1 U29207 ( .A(n26071), .B(n24070), .Y(n24071) );
  sky130_fd_sc_hd__nand3_1 U29208 ( .A(n24073), .B(n24072), .C(n24071), .Y(
        j202_soc_core_j22_cpu_rf_N309) );
  sky130_fd_sc_hd__nor2_1 U29209 ( .A(n26192), .B(n12361), .Y(n24869) );
  sky130_fd_sc_hd__inv_2 U29210 ( .A(n24869), .Y(n24901) );
  sky130_fd_sc_hd__a22oi_1 U29211 ( .A1(n26070), .A2(n28478), .B1(n24873), 
        .B2(n26068), .Y(n24077) );
  sky130_fd_sc_hd__nand2_1 U29212 ( .A(n26071), .B(n24075), .Y(n24076) );
  sky130_fd_sc_hd__o211ai_1 U29213 ( .A1(n27855), .A2(n28480), .B1(n24077), 
        .C1(n24076), .Y(j202_soc_core_j22_cpu_rf_N307) );
  sky130_fd_sc_hd__buf_2 U29214 ( .A(n12212), .X(n24629) );
  sky130_fd_sc_hd__nand2_1 U29215 ( .A(n24629), .B(n28417), .Y(n24648) );
  sky130_fd_sc_hd__nor2_1 U29216 ( .A(n11178), .B(n24648), .Y(
        j202_soc_core_j22_cpu_id_idec_N900) );
  sky130_fd_sc_hd__nand2_1 U29217 ( .A(n11442), .B(n25724), .Y(n24081) );
  sky130_fd_sc_hd__a22oi_1 U29218 ( .A1(n26070), .A2(n28541), .B1(n24078), 
        .B2(n26068), .Y(n24080) );
  sky130_fd_sc_hd__nand2_1 U29219 ( .A(n26071), .B(j202_soc_core_j22_cpu_pc[0]), .Y(n24079) );
  sky130_fd_sc_hd__nand3_1 U29220 ( .A(n24081), .B(n24080), .C(n24079), .Y(
        j202_soc_core_j22_cpu_rf_N298) );
  sky130_fd_sc_hd__a22oi_1 U29221 ( .A1(n26070), .A2(n28515), .B1(n24082), 
        .B2(n26068), .Y(n24084) );
  sky130_fd_sc_hd__nand2_1 U29222 ( .A(n26071), .B(n24773), .Y(n24083) );
  sky130_fd_sc_hd__nand3_1 U29223 ( .A(n24085), .B(n24084), .C(n24083), .Y(
        j202_soc_core_j22_cpu_rf_N301) );
  sky130_fd_sc_hd__nor2_1 U29224 ( .A(n26195), .B(n12360), .Y(n24680) );
  sky130_fd_sc_hd__a22oi_1 U29225 ( .A1(n26070), .A2(n28489), .B1(n24086), 
        .B2(n26068), .Y(n24088) );
  sky130_fd_sc_hd__nand2_1 U29226 ( .A(n26071), .B(n24713), .Y(n24087) );
  sky130_fd_sc_hd__o211ai_1 U29227 ( .A1(n27855), .A2(n11180), .B1(n24088), 
        .C1(n24087), .Y(j202_soc_core_j22_cpu_rf_N305) );
  sky130_fd_sc_hd__nand2_1 U29228 ( .A(n26158), .B(n25938), .Y(n24089) );
  sky130_fd_sc_hd__o21a_1 U29229 ( .A1(n25940), .A2(n24090), .B1(n24089), .X(
        n26174) );
  sky130_fd_sc_hd__nor2_1 U29230 ( .A(n24091), .B(n12360), .Y(n26917) );
  sky130_fd_sc_hd__a22oi_1 U29231 ( .A1(n26070), .A2(n28473), .B1(n26956), 
        .B2(n26068), .Y(n24094) );
  sky130_fd_sc_hd__nand2_1 U29232 ( .A(n26071), .B(n24092), .Y(n24093) );
  sky130_fd_sc_hd__o211ai_1 U29233 ( .A1(n27855), .A2(n26965), .B1(n24094), 
        .C1(n24093), .Y(j202_soc_core_j22_cpu_rf_N308) );
  sky130_fd_sc_hd__inv_1 U29234 ( .A(n28091), .Y(n24096) );
  sky130_fd_sc_hd__nand2_1 U29235 ( .A(n24629), .B(n11423), .Y(n24095) );
  sky130_fd_sc_hd__nand4_1 U29236 ( .A(n11449), .B(n24096), .C(n25904), .D(
        n24095), .Y(n24100) );
  sky130_fd_sc_hd__inv_1 U29237 ( .A(n24097), .Y(n24098) );
  sky130_fd_sc_hd__nor2_1 U29238 ( .A(n24099), .B(n28090), .Y(n24692) );
  sky130_fd_sc_hd__inv_1 U29239 ( .A(n28387), .Y(n24101) );
  sky130_fd_sc_hd__nor2_1 U29240 ( .A(n24423), .B(n24101), .Y(n24103) );
  sky130_fd_sc_hd__a22oi_1 U29241 ( .A1(n27885), .A2(n29587), .B1(n24112), 
        .B2(n24102), .Y(n27909) );
  sky130_fd_sc_hd__nand2_1 U29242 ( .A(n12064), .B(n28130), .Y(n24104) );
  sky130_fd_sc_hd__nand2_1 U29243 ( .A(n11646), .B(n24634), .Y(n24105) );
  sky130_fd_sc_hd__o211a_1 U29244 ( .A1(n27899), .A2(n27739), .B1(n24406), 
        .C1(n24105), .X(n28147) );
  sky130_fd_sc_hd__nand3_1 U29245 ( .A(n24547), .B(n11110), .C(n28147), .Y(
        n24107) );
  sky130_fd_sc_hd__nor2_1 U29246 ( .A(n24107), .B(n28151), .Y(n24108) );
  sky130_fd_sc_hd__nand2_1 U29247 ( .A(n24109), .B(n28072), .Y(n24396) );
  sky130_fd_sc_hd__nand2_1 U29248 ( .A(n28360), .B(n24396), .Y(n24119) );
  sky130_fd_sc_hd__nand4_1 U29249 ( .A(n12287), .B(n12399), .C(n24111), .D(
        n24110), .Y(n24114) );
  sky130_fd_sc_hd__nor2_1 U29250 ( .A(n24114), .B(n24113), .Y(n28150) );
  sky130_fd_sc_hd__nand2_1 U29251 ( .A(n24117), .B(n28417), .Y(n24118) );
  sky130_fd_sc_hd__nor2_1 U29252 ( .A(n11669), .B(n27885), .Y(n24120) );
  sky130_fd_sc_hd__nand2_1 U29253 ( .A(n24958), .B(n24120), .Y(n24122) );
  sky130_fd_sc_hd__nand2b_1 U29254 ( .A_N(n24124), .B(n11545), .Y(n24125) );
  sky130_fd_sc_hd__nand2_1 U29255 ( .A(n28033), .B(n11395), .Y(n24130) );
  sky130_fd_sc_hd__a21o_1 U29256 ( .A1(n11141), .A2(n24127), .B1(n24126), .X(
        n28030) );
  sky130_fd_sc_hd__nand2_1 U29257 ( .A(n28030), .B(n12417), .Y(n24129) );
  sky130_fd_sc_hd__nand3_1 U29258 ( .A(n24131), .B(n24130), .C(n24129), .Y(
        n24132) );
  sky130_fd_sc_hd__nand2_1 U29259 ( .A(n28030), .B(n29491), .Y(n24136) );
  sky130_fd_sc_hd__nand2_1 U29260 ( .A(n24133), .B(n29560), .Y(n24135) );
  sky130_fd_sc_hd__nand2_1 U29261 ( .A(n25146), .B(n11520), .Y(n24134) );
  sky130_fd_sc_hd__nand3_1 U29262 ( .A(n24136), .B(n24135), .C(n24134), .Y(
        n24137) );
  sky130_fd_sc_hd__nand2_1 U29263 ( .A(n28030), .B(n11395), .Y(n24140) );
  sky130_fd_sc_hd__nand2_1 U29264 ( .A(n24133), .B(n11520), .Y(n24139) );
  sky130_fd_sc_hd__nand2_1 U29265 ( .A(n28033), .B(n29491), .Y(n24138) );
  sky130_fd_sc_hd__nand3_1 U29266 ( .A(n24140), .B(n24139), .C(n24138), .Y(
        n24142) );
  sky130_fd_sc_hd__and4_1 U29267 ( .A(n24146), .B(n12421), .C(n29745), .D(
        n24143), .X(n29633) );
  sky130_fd_sc_hd__and3_1 U29268 ( .A(n24146), .B(n24145), .C(n29827), .X(
        n29634) );
  sky130_fd_sc_hd__and4_1 U29269 ( .A(n24149), .B(n27052), .C(n24148), .D(
        n24154), .X(n24150) );
  sky130_fd_sc_hd__a21oi_1 U29270 ( .A1(n24151), .A2(n24150), .B1(n26926), .Y(
        n24173) );
  sky130_fd_sc_hd__nand2_1 U29271 ( .A(n24152), .B(n24173), .Y(n24175) );
  sky130_fd_sc_hd__nand3_1 U29272 ( .A(n24155), .B(n27828), .C(n24154), .Y(
        n24172) );
  sky130_fd_sc_hd__nor2_1 U29274 ( .A(n24156), .B(n12351), .Y(n24165) );
  sky130_fd_sc_hd__nand2_1 U29275 ( .A(n24165), .B(n26916), .Y(n24157) );
  sky130_fd_sc_hd__o22ai_1 U29276 ( .A1(n24929), .A2(n27793), .B1(n26317), 
        .B2(n27797), .Y(n24159) );
  sky130_fd_sc_hd__o22ai_1 U29277 ( .A1(n26322), .A2(n27799), .B1(n27796), 
        .B2(n27803), .Y(n24158) );
  sky130_fd_sc_hd__nor2_1 U29278 ( .A(n24159), .B(n24158), .Y(n24162) );
  sky130_fd_sc_hd__xnor2_1 U29279 ( .A(n24929), .B(n27807), .Y(n26233) );
  sky130_fd_sc_hd__o22a_1 U29280 ( .A1(n26431), .A2(n27795), .B1(n25872), .B2(
        n26233), .X(n24161) );
  sky130_fd_sc_hd__a22oi_1 U29281 ( .A1(n27810), .A2(n27788), .B1(n27808), 
        .B2(n25642), .Y(n24160) );
  sky130_fd_sc_hd__nand4_1 U29282 ( .A(n27814), .B(n24162), .C(n24161), .D(
        n24160), .Y(n24164) );
  sky130_fd_sc_hd__o22ai_1 U29283 ( .A1(n28481), .A2(n27817), .B1(n24931), 
        .B2(n27815), .Y(n24163) );
  sky130_fd_sc_hd__nor2_1 U29284 ( .A(n24164), .B(n24163), .Y(n24170) );
  sky130_fd_sc_hd__o211ai_1 U29286 ( .A1(n11123), .A2(n27807), .B1(n25638), 
        .C1(n24166), .Y(n24167) );
  sky130_fd_sc_hd__nand2_1 U29287 ( .A(n25209), .B(n24167), .Y(n24169) );
  sky130_fd_sc_hd__nand2_1 U29288 ( .A(n26461), .B(n27789), .Y(n24168) );
  sky130_fd_sc_hd__nand3_1 U29289 ( .A(n24176), .B(
        j202_soc_core_j22_cpu_regop_We__0_), .C(
        j202_soc_core_j22_cpu_regop_We__3_), .Y(n27644) );
  sky130_fd_sc_hd__nor2_1 U29290 ( .A(j202_soc_core_ahb2apb_00_state[2]), .B(
        n24177), .Y(n24178) );
  sky130_fd_sc_hd__a22oi_1 U29291 ( .A1(n26070), .A2(n28431), .B1(n26417), 
        .B2(n26068), .Y(n24180) );
  sky130_fd_sc_hd__and3_1 U29293 ( .A(n28109), .B(n29882), .C(n24183), .X(
        n29649) );
  sky130_fd_sc_hd__nand2_1 U29294 ( .A(n26467), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n29276) );
  sky130_fd_sc_hd__and3_1 U29295 ( .A(n24184), .B(la_data_in[31]), .C(n29830), 
        .X(n29652) );
  sky130_fd_sc_hd__and3_1 U29296 ( .A(n24185), .B(la_data_in[30]), .C(n29830), 
        .X(n29653) );
  sky130_fd_sc_hd__and3_1 U29297 ( .A(n24186), .B(la_data_in[29]), .C(n29828), 
        .X(n29654) );
  sky130_fd_sc_hd__and3_1 U29298 ( .A(n24187), .B(la_data_in[28]), .C(n12069), 
        .X(n29655) );
  sky130_fd_sc_hd__and3_1 U29299 ( .A(n24188), .B(la_data_in[27]), .C(n29830), 
        .X(n29656) );
  sky130_fd_sc_hd__and3_1 U29300 ( .A(n24189), .B(la_data_in[26]), .C(n12069), 
        .X(n29657) );
  sky130_fd_sc_hd__and3_1 U29301 ( .A(n24190), .B(la_data_in[25]), .C(n12069), 
        .X(n29658) );
  sky130_fd_sc_hd__and3_1 U29302 ( .A(n24191), .B(la_data_in[24]), .C(n29827), 
        .X(n29659) );
  sky130_fd_sc_hd__and3_1 U29303 ( .A(n24192), .B(la_data_in[23]), .C(n12069), 
        .X(n29660) );
  sky130_fd_sc_hd__and3_1 U29304 ( .A(n24193), .B(la_data_in[22]), .C(n29745), 
        .X(n29661) );
  sky130_fd_sc_hd__and3_1 U29305 ( .A(n24194), .B(la_data_in[21]), .C(n12069), 
        .X(n29662) );
  sky130_fd_sc_hd__and3_1 U29306 ( .A(n24195), .B(la_data_in[20]), .C(n29827), 
        .X(n29663) );
  sky130_fd_sc_hd__and3_1 U29307 ( .A(n24196), .B(la_data_in[19]), .C(n29827), 
        .X(n29664) );
  sky130_fd_sc_hd__and3_1 U29308 ( .A(n24197), .B(la_data_in[18]), .C(n12069), 
        .X(n29665) );
  sky130_fd_sc_hd__and3_1 U29309 ( .A(n24198), .B(la_data_in[17]), .C(n29828), 
        .X(n29666) );
  sky130_fd_sc_hd__nand2b_1 U29310 ( .A_N(n26514), .B(n26511), .Y(n28026) );
  sky130_fd_sc_hd__o22ai_1 U29311 ( .A1(n29115), .A2(n24200), .B1(n24199), 
        .B2(n29493), .Y(n24201) );
  sky130_fd_sc_hd__nand2_1 U29312 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[27]), .Y(n24203) );
  sky130_fd_sc_hd__nand2_1 U29313 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[24]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24202) );
  sky130_fd_sc_hd__nand2_1 U29314 ( .A(n24203), .B(n24202), .Y(n25552) );
  sky130_fd_sc_hd__nand2_1 U29315 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[23]), .Y(n24205) );
  sky130_fd_sc_hd__nand2_1 U29316 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[20]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24204) );
  sky130_fd_sc_hd__nand2_1 U29317 ( .A(n24205), .B(n24204), .Y(n25544) );
  sky130_fd_sc_hd__nand2_1 U29318 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[22]), .Y(n24207) );
  sky130_fd_sc_hd__nand2_1 U29319 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[19]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24206) );
  sky130_fd_sc_hd__nand2_1 U29320 ( .A(n24207), .B(n24206), .Y(n25542) );
  sky130_fd_sc_hd__nand2_1 U29321 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[21]), .Y(n24209) );
  sky130_fd_sc_hd__nand2_1 U29322 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[18]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24208) );
  sky130_fd_sc_hd__nand2_1 U29323 ( .A(n24209), .B(n24208), .Y(n25540) );
  sky130_fd_sc_hd__nand2_1 U29324 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[20]), .Y(n24211) );
  sky130_fd_sc_hd__nand2_1 U29325 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[17]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24210) );
  sky130_fd_sc_hd__nand2_1 U29326 ( .A(n24211), .B(n24210), .Y(n25538) );
  sky130_fd_sc_hd__nand2_1 U29327 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[19]), .Y(n24213) );
  sky130_fd_sc_hd__nand2_1 U29328 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[16]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24212) );
  sky130_fd_sc_hd__nand2_1 U29329 ( .A(n24213), .B(n24212), .Y(n25536) );
  sky130_fd_sc_hd__nand2_1 U29330 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[9]), .Y(n24215) );
  sky130_fd_sc_hd__nand2_1 U29331 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[6]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24214) );
  sky130_fd_sc_hd__nand2_1 U29332 ( .A(n24215), .B(n24214), .Y(n25516) );
  sky130_fd_sc_hd__nand2_1 U29333 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[3]), .Y(n24217) );
  sky130_fd_sc_hd__nand2_1 U29334 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[0]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24216) );
  sky130_fd_sc_hd__nand2_1 U29335 ( .A(n24217), .B(n24216), .Y(n25504) );
  sky130_fd_sc_hd__nand2_1 U29336 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[25]), .Y(n24219) );
  sky130_fd_sc_hd__nand2_1 U29337 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[22]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24218) );
  sky130_fd_sc_hd__nand2_1 U29338 ( .A(n24219), .B(n24218), .Y(n25548) );
  sky130_fd_sc_hd__nand2_1 U29339 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[18]), .Y(n24221) );
  sky130_fd_sc_hd__nand2_1 U29340 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[15]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24220) );
  sky130_fd_sc_hd__nand2_1 U29341 ( .A(n24221), .B(n24220), .Y(n25534) );
  sky130_fd_sc_hd__nand2_1 U29342 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[7]), .Y(n24223) );
  sky130_fd_sc_hd__nand2_1 U29343 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[4]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24222) );
  sky130_fd_sc_hd__nand2_1 U29344 ( .A(n24223), .B(n24222), .Y(n25512) );
  sky130_fd_sc_hd__nand2_1 U29345 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[29]), .Y(n24225) );
  sky130_fd_sc_hd__nand2_1 U29346 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[26]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24224) );
  sky130_fd_sc_hd__nand2_1 U29347 ( .A(n24225), .B(n24224), .Y(n28893) );
  sky130_fd_sc_hd__nand2_1 U29348 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[28]), .Y(n24227) );
  sky130_fd_sc_hd__nand2_1 U29349 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[25]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24226) );
  sky130_fd_sc_hd__nand2_1 U29350 ( .A(n24227), .B(n24226), .Y(n28023) );
  sky130_fd_sc_hd__nand2_1 U29351 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[26]), .Y(n24229) );
  sky130_fd_sc_hd__nand2_1 U29352 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[23]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24228) );
  sky130_fd_sc_hd__nand2_1 U29353 ( .A(n24229), .B(n24228), .Y(n25550) );
  sky130_fd_sc_hd__nand2_1 U29354 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[16]), .Y(n24231) );
  sky130_fd_sc_hd__nand2_1 U29355 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[13]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24230) );
  sky130_fd_sc_hd__nand2_1 U29356 ( .A(n24231), .B(n24230), .Y(n25530) );
  sky130_fd_sc_hd__nand2_1 U29357 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[14]), .Y(n24233) );
  sky130_fd_sc_hd__nand2_1 U29358 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[11]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24232) );
  sky130_fd_sc_hd__nand2_1 U29359 ( .A(n24233), .B(n24232), .Y(n25526) );
  sky130_fd_sc_hd__nand2_1 U29360 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[12]), .Y(n24235) );
  sky130_fd_sc_hd__nand2_1 U29361 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[9]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24234) );
  sky130_fd_sc_hd__nand2_1 U29362 ( .A(n24235), .B(n24234), .Y(n25522) );
  sky130_fd_sc_hd__nand2_1 U29363 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[10]), .Y(n24237) );
  sky130_fd_sc_hd__nand2_1 U29364 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[7]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24236) );
  sky130_fd_sc_hd__nand2_1 U29365 ( .A(n24237), .B(n24236), .Y(n25518) );
  sky130_fd_sc_hd__nand2_1 U29366 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[8]), .Y(n24239) );
  sky130_fd_sc_hd__nand2_1 U29367 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[5]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24238) );
  sky130_fd_sc_hd__nand2_1 U29368 ( .A(n24239), .B(n24238), .Y(n25514) );
  sky130_fd_sc_hd__nand2_1 U29369 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[6]), .Y(n24241) );
  sky130_fd_sc_hd__nand2_1 U29370 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[3]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24240) );
  sky130_fd_sc_hd__nand2_1 U29371 ( .A(n24241), .B(n24240), .Y(n25510) );
  sky130_fd_sc_hd__nand2_1 U29372 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[4]), .Y(n24243) );
  sky130_fd_sc_hd__nand2_1 U29373 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[1]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24242) );
  sky130_fd_sc_hd__nand2_1 U29374 ( .A(n24243), .B(n24242), .Y(n25506) );
  sky130_fd_sc_hd__nand2_1 U29375 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[24]), .Y(n24245) );
  sky130_fd_sc_hd__nand2_1 U29376 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[21]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24244) );
  sky130_fd_sc_hd__nand2_1 U29377 ( .A(n24245), .B(n24244), .Y(n25546) );
  sky130_fd_sc_hd__nand2_1 U29378 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[17]), .Y(n24247) );
  sky130_fd_sc_hd__nand2_1 U29379 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[14]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24246) );
  sky130_fd_sc_hd__nand2_1 U29380 ( .A(n24247), .B(n24246), .Y(n25532) );
  sky130_fd_sc_hd__nand2_1 U29381 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[13]), .Y(n24249) );
  sky130_fd_sc_hd__nand2_1 U29382 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[10]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24248) );
  sky130_fd_sc_hd__nand2_1 U29383 ( .A(n24249), .B(n24248), .Y(n25524) );
  sky130_fd_sc_hd__nand2_1 U29384 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[5]), .Y(n24251) );
  sky130_fd_sc_hd__nand2_1 U29385 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[2]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24250) );
  sky130_fd_sc_hd__nand2_1 U29386 ( .A(n24251), .B(n24250), .Y(n25508) );
  sky130_fd_sc_hd__nand2_1 U29387 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[15]), .Y(n24253) );
  sky130_fd_sc_hd__nand2_1 U29388 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[12]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24252) );
  sky130_fd_sc_hd__nand2_1 U29389 ( .A(n24253), .B(n24252), .Y(n25528) );
  sky130_fd_sc_hd__nand2_1 U29390 ( .A(n28896), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[11]), .Y(n24255) );
  sky130_fd_sc_hd__nand2_1 U29391 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[8]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24254) );
  sky130_fd_sc_hd__nand2_1 U29392 ( .A(n24255), .B(n24254), .Y(n25520) );
  sky130_fd_sc_hd__nand3_1 U29393 ( .A(j202_soc_core_cmt_core_00_cmf0), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[6]), .C(n29830), .Y(
        n26764) );
  sky130_fd_sc_hd__nand3_1 U29394 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[4]), .B(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[6]), .C(j202_soc_core_intc_core_00_cp_intack_all_0_), .Y(n25735) );
  sky130_fd_sc_hd__nor2_1 U29395 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .B(n25735), .Y(n26853) );
  sky130_fd_sc_hd__and3_1 U29396 ( .A(n26853), .B(n25736), .C(n29072), .X(
        n27310) );
  sky130_fd_sc_hd__nor2_1 U29397 ( .A(j202_soc_core_intc_core_00_rg_irqc[16]), 
        .B(n29088), .Y(n24256) );
  sky130_fd_sc_hd__o211ai_1 U29398 ( .A1(n24257), .A2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]), .B1(j202_soc_core_intc_core_00_in_intreq[16]), .C1(n24256), .Y(n24258) );
  sky130_fd_sc_hd__o21ai_1 U29399 ( .A1(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[16]), 
        .A2(n26764), .B1(n24258), .Y(n24259) );
  sky130_fd_sc_hd__o211a_2 U29400 ( .A1(n24264), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[4]), .B1(n28557), .C1(
        n29169), .X(n29724) );
  sky130_fd_sc_hd__o211a_2 U29401 ( .A1(n24268), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[2]), .B1(n24265), .C1(
        n29169), .X(n29725) );
  sky130_fd_sc_hd__o211a_2 U29402 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[6]), .A2(n28556), .B1(
        n29169), .C1(n28560), .X(n29726) );
  sky130_fd_sc_hd__nor2_1 U29403 ( .A(j202_soc_core_ahb2apb_02_state[2]), .B(
        n24260), .Y(n24274) );
  sky130_fd_sc_hd__and3_1 U29404 ( .A(n24274), .B(n24296), .C(n12069), .X(
        n29730) );
  sky130_fd_sc_hd__nand3_1 U29405 ( .A(j202_soc_core_uart_TOP_tx_bit_cnt[0]), 
        .B(j202_soc_core_uart_TOP_tx_bit_cnt[1]), .C(
        j202_soc_core_uart_TOP_tx_bit_cnt[2]), .Y(n28594) );
  sky130_fd_sc_hd__nor2_1 U29406 ( .A(n24261), .B(j202_soc_core_uart_TOP_load), 
        .Y(n24262) );
  sky130_fd_sc_hd__o211a_2 U29407 ( .A1(n24263), .A2(
        j202_soc_core_uart_TOP_tx_bit_cnt[2]), .B1(n24262), .C1(n29494), .X(
        n29731) );
  sky130_fd_sc_hd__a21oi_1 U29408 ( .A1(n24266), .A2(n24265), .B1(n24264), .Y(
        n24267) );
  sky130_fd_sc_hd__a21oi_1 U29409 ( .A1(n28554), .A2(n24269), .B1(n24268), .Y(
        n24270) );
  sky130_fd_sc_hd__xor2_1 U29410 ( .A(j202_soc_core_uart_TOP_tx_bit_cnt[0]), 
        .B(j202_soc_core_uart_TOP_tx_bit_cnt[1]), .X(n24272) );
  sky130_fd_sc_hd__and3_1 U29411 ( .A(n24272), .B(n29494), .C(n24271), .X(
        n29740) );
  sky130_fd_sc_hd__nor2_1 U29412 ( .A(j202_soc_core_rst), .B(
        j202_soc_core_ahb2apb_00_state[2]), .Y(n24276) );
  sky130_fd_sc_hd__and3_1 U29413 ( .A(n24276), .B(
        j202_soc_core_ahb2apb_00_state[0]), .C(
        j202_soc_core_ahb2apb_00_state[1]), .X(n29741) );
  sky130_fd_sc_hd__nor2_1 U29414 ( .A(n29088), .B(n24296), .Y(n26900) );
  sky130_fd_sc_hd__nand2_1 U29415 ( .A(n24728), .B(
        j202_soc_core_ahb2apb_00_state[1]), .Y(n24275) );
  sky130_fd_sc_hd__mux2i_1 U29416 ( .A0(n24275), .A1(
        j202_soc_core_ahb2apb_00_state[1]), .S(
        j202_soc_core_ahb2apb_00_state[0]), .Y(n24277) );
  sky130_fd_sc_hd__nand2_1 U29417 ( .A(n29270), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[1]), .Y(n28696) );
  sky130_fd_sc_hd__nand2_1 U29418 ( .A(n29270), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[0]), .Y(n28700) );
  sky130_fd_sc_hd__nand2_1 U29419 ( .A(n29603), .B(n28727), .Y(n24279) );
  sky130_fd_sc_hd__nor2_1 U29420 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd), .B(n26667), .Y(n26653)
         );
  sky130_fd_sc_hd__o211ai_1 U29421 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd), .A2(n26661), .B1(n24279), 
        .C1(n24278), .Y(n28701) );
  sky130_fd_sc_hd__nand2_1 U29422 ( .A(n28700), .B(n28701), .Y(n28698) );
  sky130_fd_sc_hd__nand2_1 U29423 ( .A(n28696), .B(n24280), .Y(
        DP_OP_1508J1_126_2326_n4) );
  sky130_fd_sc_hd__buf_2 U29424 ( .A(n25696), .X(n25720) );
  sky130_fd_sc_hd__nor2_1 U29425 ( .A(n24285), .B(n24284), .Y(n24291) );
  sky130_fd_sc_hd__or4_1 U29426 ( .A(j202_soc_core_j22_cpu_macop_MAC_[2]), .B(
        n28053), .C(n24286), .D(n24287), .X(n28428) );
  sky130_fd_sc_hd__nand2_1 U29427 ( .A(n27764), .B(n25697), .Y(n24293) );
  sky130_fd_sc_hd__nand2_1 U29428 ( .A(j202_soc_core_j22_cpu_macop_MAC_[3]), 
        .B(j202_soc_core_j22_cpu_macop_MAC_[1]), .Y(n24667) );
  sky130_fd_sc_hd__nor3_1 U29429 ( .A(j202_soc_core_j22_cpu_macop_MAC_[2]), 
        .B(n27052), .C(n24667), .Y(n28438) );
  sky130_fd_sc_hd__and3_1 U29430 ( .A(n26064), .B(n28438), .C(n27615), .X(
        n24290) );
  sky130_fd_sc_hd__o211ai_1 U29431 ( .A1(n25720), .A2(n27388), .B1(n24293), 
        .C1(n24292), .Y(j202_soc_core_j22_cpu_ml_N322) );
  sky130_fd_sc_hd__nand2_1 U29432 ( .A(n27764), .B(n27033), .Y(n24295) );
  sky130_fd_sc_hd__o211ai_1 U29433 ( .A1(n27642), .A2(n27388), .B1(n24295), 
        .C1(n24292), .Y(j202_soc_core_j22_cpu_ml_N333) );
  sky130_fd_sc_hd__nand2_1 U29434 ( .A(n26899), .B(n24296), .Y(n24298) );
  sky130_fd_sc_hd__nor2_1 U29435 ( .A(n24298), .B(n24307), .Y(
        j202_soc_core_ahb2apb_02_N89) );
  sky130_fd_sc_hd__nor2_1 U29436 ( .A(n24818), .B(n24307), .Y(
        j202_soc_core_ahb2apb_02_N26) );
  sky130_fd_sc_hd__nor2_1 U29437 ( .A(n25053), .B(n24307), .Y(
        j202_soc_core_ahb2apb_02_N27) );
  sky130_fd_sc_hd__nor2_1 U29438 ( .A(n24817), .B(n24307), .Y(
        j202_soc_core_ahb2apb_02_N25) );
  sky130_fd_sc_hd__nor2_1 U29439 ( .A(n25054), .B(n24307), .Y(
        j202_soc_core_ahb2apb_02_N28) );
  sky130_fd_sc_hd__nor2_1 U29440 ( .A(n25036), .B(n24307), .Y(
        j202_soc_core_ahb2apb_02_N29) );
  sky130_fd_sc_hd__nor2_1 U29441 ( .A(n25035), .B(n24307), .Y(
        j202_soc_core_ahb2apb_02_N30) );
  sky130_fd_sc_hd__nor2_1 U29442 ( .A(n27919), .B(n24307), .Y(
        j202_soc_core_ahb2apb_02_N24) );
  sky130_fd_sc_hd__nor2_1 U29443 ( .A(n27090), .B(n24307), .Y(
        j202_soc_core_ahb2apb_02_N23) );
  sky130_fd_sc_hd__nor2_1 U29445 ( .A(n27091), .B(n24307), .Y(
        j202_soc_core_ahb2apb_02_N56) );
  sky130_fd_sc_hd__nand3_1 U29446 ( .A(n24305), .B(n24304), .C(n24303), .Y(
        n24306) );
  sky130_fd_sc_hd__o21ba_2 U29447 ( .A1(n28103), .A2(n29581), .B1_N(n24306), 
        .X(n25476) );
  sky130_fd_sc_hd__nor2_1 U29448 ( .A(n25476), .B(n24307), .Y(
        j202_soc_core_ahb2apb_02_N57) );
  sky130_fd_sc_hd__nor2_1 U29449 ( .A(n12842), .B(n24307), .Y(
        j202_soc_core_ahb2apb_02_N55) );
  sky130_fd_sc_hd__nand2_1 U29450 ( .A(n12330), .B(
        j202_soc_core_j22_cpu_ml_macl[6]), .Y(n24311) );
  sky130_fd_sc_hd__inv_2 U29451 ( .A(n24312), .Y(n24365) );
  sky130_fd_sc_hd__nand2_1 U29452 ( .A(n24365), .B(n24308), .Y(n24310) );
  sky130_fd_sc_hd__a21oi_1 U29453 ( .A1(n27768), .A2(
        j202_soc_core_j22_cpu_ml_bufa[6]), .B1(n27766), .Y(n24309) );
  sky130_fd_sc_hd__nand3_1 U29454 ( .A(n24310), .B(n24311), .C(n24309), .Y(
        j202_soc_core_j22_cpu_ml_maclj[6]) );
  sky130_fd_sc_hd__inv_2 U29455 ( .A(n24312), .Y(n26967) );
  sky130_fd_sc_hd__nand2_1 U29456 ( .A(n26967), .B(n24313), .Y(n24316) );
  sky130_fd_sc_hd__nand2_1 U29457 ( .A(n24363), .B(
        j202_soc_core_j22_cpu_ml_macl[10]), .Y(n24315) );
  sky130_fd_sc_hd__a21oi_1 U29458 ( .A1(n27768), .A2(n30145), .B1(n27766), .Y(
        n24314) );
  sky130_fd_sc_hd__nand3_1 U29459 ( .A(n24316), .B(n24315), .C(n24314), .Y(
        j202_soc_core_j22_cpu_ml_maclj[10]) );
  sky130_fd_sc_hd__nand2_1 U29460 ( .A(n26967), .B(n24462), .Y(n24319) );
  sky130_fd_sc_hd__nand2_1 U29461 ( .A(n24363), .B(
        j202_soc_core_j22_cpu_ml_macl[14]), .Y(n24318) );
  sky130_fd_sc_hd__a21oi_1 U29462 ( .A1(n27768), .A2(n24454), .B1(n27766), .Y(
        n24317) );
  sky130_fd_sc_hd__nand3_1 U29463 ( .A(n24319), .B(n24318), .C(n24317), .Y(
        j202_soc_core_j22_cpu_ml_maclj[14]) );
  sky130_fd_sc_hd__nand2_1 U29464 ( .A(n24325), .B(n24320), .Y(n24323) );
  sky130_fd_sc_hd__nand2_1 U29465 ( .A(n12330), .B(
        j202_soc_core_j22_cpu_ml_macl[1]), .Y(n24322) );
  sky130_fd_sc_hd__a21oi_1 U29466 ( .A1(n27768), .A2(n21943), .B1(n27766), .Y(
        n24321) );
  sky130_fd_sc_hd__nand3_1 U29467 ( .A(n24323), .B(n24322), .C(n24321), .Y(
        j202_soc_core_j22_cpu_ml_maclj[1]) );
  sky130_fd_sc_hd__nand2_1 U29468 ( .A(n12330), .B(
        j202_soc_core_j22_cpu_ml_macl[7]), .Y(n24328) );
  sky130_fd_sc_hd__nand2_1 U29469 ( .A(n24325), .B(n24324), .Y(n24327) );
  sky130_fd_sc_hd__a21oi_1 U29470 ( .A1(n27768), .A2(n27618), .B1(n27766), .Y(
        n24326) );
  sky130_fd_sc_hd__nand3_1 U29471 ( .A(n24328), .B(n24326), .C(n24327), .Y(
        j202_soc_core_j22_cpu_ml_maclj[7]) );
  sky130_fd_sc_hd__nand2_1 U29472 ( .A(n24325), .B(n24329), .Y(n24332) );
  sky130_fd_sc_hd__nand2_1 U29473 ( .A(n24363), .B(
        j202_soc_core_j22_cpu_ml_macl[3]), .Y(n24331) );
  sky130_fd_sc_hd__a21oi_1 U29474 ( .A1(n27768), .A2(n21219), .B1(n27766), .Y(
        n24330) );
  sky130_fd_sc_hd__nand3_1 U29475 ( .A(n24332), .B(n24331), .C(n24330), .Y(
        j202_soc_core_j22_cpu_ml_maclj[3]) );
  sky130_fd_sc_hd__nand2_1 U29476 ( .A(n26967), .B(n24333), .Y(n24336) );
  sky130_fd_sc_hd__nand2_1 U29477 ( .A(n24363), .B(
        j202_soc_core_j22_cpu_ml_macl[9]), .Y(n24335) );
  sky130_fd_sc_hd__a21oi_1 U29478 ( .A1(n27768), .A2(n24799), .B1(n27766), .Y(
        n24334) );
  sky130_fd_sc_hd__nand3_1 U29479 ( .A(n24336), .B(n24335), .C(n24334), .Y(
        j202_soc_core_j22_cpu_ml_maclj[9]) );
  sky130_fd_sc_hd__nand2_1 U29480 ( .A(n24365), .B(n24337), .Y(n24340) );
  sky130_fd_sc_hd__nand2_1 U29481 ( .A(n24363), .B(
        j202_soc_core_j22_cpu_ml_macl[15]), .Y(n24339) );
  sky130_fd_sc_hd__a21oi_1 U29482 ( .A1(n27768), .A2(n18887), .B1(n27766), .Y(
        n24338) );
  sky130_fd_sc_hd__nand3_1 U29483 ( .A(n24340), .B(n24339), .C(n24338), .Y(
        j202_soc_core_j22_cpu_ml_maclj[15]) );
  sky130_fd_sc_hd__nand2_1 U29484 ( .A(n12330), .B(
        j202_soc_core_j22_cpu_ml_macl[11]), .Y(n24344) );
  sky130_fd_sc_hd__nand2_1 U29485 ( .A(n24365), .B(n24341), .Y(n24343) );
  sky130_fd_sc_hd__a21oi_1 U29486 ( .A1(n27768), .A2(n21280), .B1(n27766), .Y(
        n24342) );
  sky130_fd_sc_hd__nand3_1 U29487 ( .A(n24344), .B(n24342), .C(n24343), .Y(
        j202_soc_core_j22_cpu_ml_maclj[11]) );
  sky130_fd_sc_hd__nand2_1 U29488 ( .A(n12330), .B(
        j202_soc_core_j22_cpu_ml_macl[13]), .Y(n24348) );
  sky130_fd_sc_hd__nand2_1 U29489 ( .A(n24365), .B(n24444), .Y(n24347) );
  sky130_fd_sc_hd__a21oi_1 U29490 ( .A1(n27768), .A2(n24345), .B1(n27766), .Y(
        n24346) );
  sky130_fd_sc_hd__nand3_1 U29491 ( .A(n24347), .B(n24348), .C(n24346), .Y(
        j202_soc_core_j22_cpu_ml_maclj[13]) );
  sky130_fd_sc_hd__nand2_1 U29492 ( .A(n26967), .B(n24349), .Y(n24352) );
  sky130_fd_sc_hd__nand2_1 U29493 ( .A(n24363), .B(
        j202_soc_core_j22_cpu_ml_macl[12]), .Y(n24351) );
  sky130_fd_sc_hd__a21oi_1 U29494 ( .A1(n27768), .A2(
        j202_soc_core_j22_cpu_ml_bufa[12]), .B1(n27766), .Y(n24350) );
  sky130_fd_sc_hd__nand3_1 U29495 ( .A(n24352), .B(n24351), .C(n24350), .Y(
        j202_soc_core_j22_cpu_ml_maclj[12]) );
  sky130_fd_sc_hd__nand2_1 U29496 ( .A(n26967), .B(n24353), .Y(n24356) );
  sky130_fd_sc_hd__nand2_1 U29497 ( .A(n24363), .B(
        j202_soc_core_j22_cpu_ml_macl[0]), .Y(n24355) );
  sky130_fd_sc_hd__a21oi_1 U29498 ( .A1(n27768), .A2(
        j202_soc_core_j22_cpu_ml_bufa[0]), .B1(n27766), .Y(n24354) );
  sky130_fd_sc_hd__nand3_1 U29499 ( .A(n24356), .B(n24355), .C(n24354), .Y(
        j202_soc_core_j22_cpu_ml_maclj[0]) );
  sky130_fd_sc_hd__nand2_1 U29500 ( .A(n27764), .B(n27032), .Y(n24359) );
  sky130_fd_sc_hd__o211ai_1 U29501 ( .A1(n27388), .A2(n28477), .B1(n24359), 
        .C1(n24292), .Y(j202_soc_core_j22_cpu_ml_N329) );
  sky130_fd_sc_hd__nand2_1 U29502 ( .A(n28055), .B(n27153), .Y(n24362) );
  sky130_fd_sc_hd__nand2_1 U29503 ( .A(n28056), .B(n24366), .Y(n24361) );
  sky130_fd_sc_hd__nand3_1 U29504 ( .A(n24362), .B(n12203), .C(n24361), .Y(
        j202_soc_core_j22_cpu_ml_machj[5]) );
  sky130_fd_sc_hd__nand2_1 U29505 ( .A(n12330), .B(
        j202_soc_core_j22_cpu_ml_macl[5]), .Y(n24369) );
  sky130_fd_sc_hd__nand2_1 U29506 ( .A(n24365), .B(n24364), .Y(n24368) );
  sky130_fd_sc_hd__a21oi_1 U29507 ( .A1(n27768), .A2(n24366), .B1(n27766), .Y(
        n24367) );
  sky130_fd_sc_hd__nand3_1 U29508 ( .A(n24369), .B(n24367), .C(n24368), .Y(
        j202_soc_core_j22_cpu_ml_maclj[5]) );
  sky130_fd_sc_hd__o22ai_1 U29509 ( .A1(n24371), .A2(n24384), .B1(n24370), 
        .B2(n27712), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N6) );
  sky130_fd_sc_hd__mux2i_1 U29510 ( .A0(n24373), .A1(
        j202_soc_core_intc_core_00_rg_ipr[80]), .S(n24376), .Y(n24375) );
  sky130_fd_sc_hd__o22ai_1 U29511 ( .A1(n24375), .A2(n24384), .B1(n24374), 
        .B2(n27712), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N3) );
  sky130_fd_sc_hd__a21oi_1 U29512 ( .A1(n24377), .A2(n27336), .B1(n24391), .Y(
        n24378) );
  sky130_fd_sc_hd__o22ai_1 U29513 ( .A1(n27344), .A2(n24384), .B1(n24378), 
        .B2(n27712), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N5) );
  sky130_fd_sc_hd__inv_1 U29514 ( .A(n24379), .Y(n24380) );
  sky130_fd_sc_hd__o22ai_1 U29515 ( .A1(n24381), .A2(n24384), .B1(n24380), 
        .B2(n27712), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N4) );
  sky130_fd_sc_hd__o22ai_1 U29516 ( .A1(n24385), .A2(n24384), .B1(n24383), 
        .B2(n27712), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N5) );
  sky130_fd_sc_hd__nand2_1 U29517 ( .A(n24387), .B(n24386), .Y(n24389) );
  sky130_fd_sc_hd__mux2i_1 U29518 ( .A0(n27326), .A1(n27330), .S(n27333), .Y(
        n24388) );
  sky130_fd_sc_hd__mux2i_1 U29519 ( .A0(n24389), .A1(n24388), .S(n27336), .Y(
        n24390) );
  sky130_fd_sc_hd__a21oi_1 U29520 ( .A1(n24391), .A2(n30169), .B1(n24390), .Y(
        n24393) );
  sky130_fd_sc_hd__nor3_1 U29521 ( .A(j202_soc_core_j22_cpu_opst[3]), .B(
        n28373), .C(n24395), .Y(n24397) );
  sky130_fd_sc_hd__nor3_1 U29522 ( .A(n28359), .B(n24397), .C(n24396), .Y(
        n24398) );
  sky130_fd_sc_hd__nand2_1 U29523 ( .A(n28379), .B(n28367), .Y(n28125) );
  sky130_fd_sc_hd__o21ai_1 U29524 ( .A1(n24398), .A2(n24613), .B1(n24412), .Y(
        n10609) );
  sky130_fd_sc_hd__nor2_1 U29525 ( .A(j202_soc_core_j22_cpu_opst[2]), .B(
        n28155), .Y(n24411) );
  sky130_fd_sc_hd__nand2_1 U29526 ( .A(n24413), .B(n24412), .Y(n24414) );
  sky130_fd_sc_hd__nand2_1 U29527 ( .A(n28360), .B(n24416), .Y(n28352) );
  sky130_fd_sc_hd__nand2_1 U29528 ( .A(n28394), .B(n28352), .Y(n24419) );
  sky130_fd_sc_hd__nand2_1 U29529 ( .A(n28360), .B(n24417), .Y(n27892) );
  sky130_fd_sc_hd__nand2b_1 U29530 ( .A_N(n27892), .B(
        j202_soc_core_j22_cpu_opst[0]), .Y(n24649) );
  sky130_fd_sc_hd__nand2_1 U29531 ( .A(n28360), .B(n24418), .Y(n28082) );
  sky130_fd_sc_hd__nand2b_1 U29532 ( .A_N(n28082), .B(
        j202_soc_core_j22_cpu_opst[1]), .Y(n28361) );
  sky130_fd_sc_hd__nand2_1 U29533 ( .A(n24649), .B(n28361), .Y(n24653) );
  sky130_fd_sc_hd__nor2_1 U29534 ( .A(n24419), .B(n24653), .Y(n24420) );
  sky130_fd_sc_hd__nand3_1 U29535 ( .A(n27644), .B(n29828), .C(n27364), .Y(
        j202_soc_core_j22_cpu_rf_N2668) );
  sky130_fd_sc_hd__nand3_1 U29536 ( .A(n24428), .B(
        j202_soc_core_j22_cpu_macop_MAC_[2]), .C(n27763), .Y(n24429) );
  sky130_fd_sc_hd__nand3_1 U29537 ( .A(n27615), .B(n24430), .C(n24429), .Y(
        n29750) );
  sky130_fd_sc_hd__nand3_1 U29538 ( .A(n25038), .B(n24431), .C(
        j202_soc_core_ahb2apb_01_state[1]), .Y(n24785) );
  sky130_fd_sc_hd__nand2_1 U29539 ( .A(n24785), .B(n12069), .Y(n29751) );
  sky130_fd_sc_hd__inv_2 U29540 ( .A(n24432), .Y(n24433) );
  sky130_fd_sc_hd__buf_6 U29541 ( .A(n24433), .X(n29762) );
  sky130_fd_sc_hd__buf_6 U29542 ( .A(n24433), .X(n29763) );
  sky130_fd_sc_hd__buf_6 U29544 ( .A(n24435), .X(n29764) );
  sky130_fd_sc_hd__buf_6 U29545 ( .A(n24435), .X(n29765) );
  sky130_fd_sc_hd__inv_2 U29546 ( .A(n24436), .Y(n24437) );
  sky130_fd_sc_hd__buf_6 U29547 ( .A(n24437), .X(n29766) );
  sky130_fd_sc_hd__buf_6 U29548 ( .A(n24437), .X(n29767) );
  sky130_fd_sc_hd__nand2_1 U29549 ( .A(n24438), .B(n24450), .Y(n27720) );
  sky130_fd_sc_hd__nand2_1 U29550 ( .A(n24439), .B(n24452), .Y(n24443) );
  sky130_fd_sc_hd__o22ai_1 U29551 ( .A1(n24456), .A2(n17994), .B1(n24440), 
        .B2(n28045), .Y(n24441) );
  sky130_fd_sc_hd__a21oi_1 U29552 ( .A1(n25442), .A2(n25679), .B1(n24441), .Y(
        n24442) );
  sky130_fd_sc_hd__nand2_1 U29553 ( .A(n24443), .B(n24442), .Y(n25421) );
  sky130_fd_sc_hd__nand2_1 U29554 ( .A(n25421), .B(n27828), .Y(n27716) );
  sky130_fd_sc_hd__nand2_1 U29555 ( .A(n24444), .B(n24461), .Y(n27714) );
  sky130_fd_sc_hd__o22ai_1 U29556 ( .A1(n17994), .A2(n26001), .B1(n24445), 
        .B2(n24463), .Y(n25406) );
  sky130_fd_sc_hd__and3_1 U29557 ( .A(n27714), .B(n27715), .C(n27720), .X(
        n24446) );
  sky130_fd_sc_hd__buf_6 U29558 ( .A(n30014), .X(n29768) );
  sky130_fd_sc_hd__buf_6 U29559 ( .A(n30014), .X(n29769) );
  sky130_fd_sc_hd__nand2_1 U29560 ( .A(n24451), .B(n24450), .Y(n26871) );
  sky130_fd_sc_hd__o22ai_1 U29561 ( .A1(n24456), .A2(n24465), .B1(n24455), 
        .B2(n28045), .Y(n24457) );
  sky130_fd_sc_hd__a21oi_1 U29562 ( .A1(n24458), .A2(n22940), .B1(n24457), .Y(
        n24459) );
  sky130_fd_sc_hd__nand2_1 U29563 ( .A(n24460), .B(n24459), .Y(n25965) );
  sky130_fd_sc_hd__nand2_1 U29564 ( .A(n25965), .B(n27828), .Y(n26868) );
  sky130_fd_sc_hd__nand2_1 U29565 ( .A(n24462), .B(n24461), .Y(n26866) );
  sky130_fd_sc_hd__o22ai_1 U29566 ( .A1(n24465), .A2(n26001), .B1(n24464), 
        .B2(n24463), .Y(n25945) );
  sky130_fd_sc_hd__and3_1 U29567 ( .A(n26866), .B(n26867), .C(n26871), .X(
        n24466) );
  sky130_fd_sc_hd__a22oi_1 U29568 ( .A1(n24467), .A2(n26871), .B1(n26868), 
        .B2(n24466), .Y(n24468) );
  sky130_fd_sc_hd__buf_4 U29569 ( .A(n24472), .X(n29772) );
  sky130_fd_sc_hd__nand2_1 U29570 ( .A(n29503), .B(n12214), .Y(n24473) );
  sky130_fd_sc_hd__inv_2 U29571 ( .A(n24473), .Y(n24474) );
  sky130_fd_sc_hd__buf_6 U29572 ( .A(n24474), .X(n29774) );
  sky130_fd_sc_hd__buf_6 U29573 ( .A(n24474), .X(n29775) );
  sky130_fd_sc_hd__buf_6 U29574 ( .A(n30193), .X(n29776) );
  sky130_fd_sc_hd__buf_6 U29575 ( .A(n30193), .X(n29777) );
  sky130_fd_sc_hd__nand2_1 U29576 ( .A(n29505), .B(n11853), .Y(n24477) );
  sky130_fd_sc_hd__buf_6 U29577 ( .A(n24478), .X(n29778) );
  sky130_fd_sc_hd__buf_6 U29578 ( .A(n24478), .X(n29779) );
  sky130_fd_sc_hd__buf_6 U29579 ( .A(n24480), .X(n29780) );
  sky130_fd_sc_hd__nand2_1 U29580 ( .A(n29507), .B(n11853), .Y(n24481) );
  sky130_fd_sc_hd__buf_6 U29581 ( .A(n24482), .X(n29781) );
  sky130_fd_sc_hd__buf_6 U29582 ( .A(n24482), .X(n29782) );
  sky130_fd_sc_hd__nand2_1 U29583 ( .A(n29508), .B(n11853), .Y(n24483) );
  sky130_fd_sc_hd__buf_6 U29584 ( .A(n24484), .X(n29783) );
  sky130_fd_sc_hd__buf_6 U29585 ( .A(n24484), .X(n29784) );
  sky130_fd_sc_hd__buf_6 U29587 ( .A(n30195), .X(n29785) );
  sky130_fd_sc_hd__buf_6 U29588 ( .A(n30195), .X(n29786) );
  sky130_fd_sc_hd__buf_4 U29590 ( .A(n30192), .X(n29787) );
  sky130_fd_sc_hd__buf_4 U29591 ( .A(n30192), .X(n29788) );
  sky130_fd_sc_hd__nand2_1 U29592 ( .A(n29511), .B(n11853), .Y(n24489) );
  sky130_fd_sc_hd__buf_6 U29593 ( .A(n24490), .X(n29789) );
  sky130_fd_sc_hd__buf_6 U29594 ( .A(n24490), .X(n29790) );
  sky130_fd_sc_hd__inv_2 U29595 ( .A(n24491), .Y(n24492) );
  sky130_fd_sc_hd__buf_6 U29596 ( .A(n24492), .X(n29791) );
  sky130_fd_sc_hd__buf_6 U29597 ( .A(n24492), .X(n29792) );
  sky130_fd_sc_hd__inv_2 U29598 ( .A(n24493), .Y(n24494) );
  sky130_fd_sc_hd__buf_6 U29599 ( .A(n24494), .X(n29793) );
  sky130_fd_sc_hd__buf_6 U29600 ( .A(n24494), .X(n29794) );
  sky130_fd_sc_hd__buf_6 U29601 ( .A(n24496), .X(n29795) );
  sky130_fd_sc_hd__buf_6 U29602 ( .A(n24496), .X(n29796) );
  sky130_fd_sc_hd__nand2_1 U29603 ( .A(n29515), .B(n12214), .Y(n24497) );
  sky130_fd_sc_hd__buf_6 U29604 ( .A(n24498), .X(n29797) );
  sky130_fd_sc_hd__buf_6 U29605 ( .A(n24498), .X(n29798) );
  sky130_fd_sc_hd__buf_6 U29606 ( .A(n24499), .X(n29799) );
  sky130_fd_sc_hd__buf_6 U29607 ( .A(n24499), .X(n29800) );
  sky130_fd_sc_hd__nand2_1 U29608 ( .A(n29518), .B(n11853), .Y(n24500) );
  sky130_fd_sc_hd__buf_6 U29609 ( .A(n24501), .X(n29801) );
  sky130_fd_sc_hd__buf_6 U29610 ( .A(n24501), .X(n29802) );
  sky130_fd_sc_hd__buf_6 U29611 ( .A(n30197), .X(n29803) );
  sky130_fd_sc_hd__buf_6 U29612 ( .A(n30197), .X(n29804) );
  sky130_fd_sc_hd__buf_6 U29613 ( .A(n24504), .X(n29805) );
  sky130_fd_sc_hd__buf_6 U29614 ( .A(n24504), .X(n29806) );
  sky130_fd_sc_hd__nand2_1 U29615 ( .A(n29521), .B(n12214), .Y(n24505) );
  sky130_fd_sc_hd__buf_6 U29616 ( .A(n24506), .X(n29807) );
  sky130_fd_sc_hd__buf_6 U29617 ( .A(n24506), .X(n29808) );
  sky130_fd_sc_hd__nand2_1 U29618 ( .A(n29522), .B(n11853), .Y(n24507) );
  sky130_fd_sc_hd__buf_6 U29619 ( .A(n24508), .X(n29809) );
  sky130_fd_sc_hd__buf_6 U29620 ( .A(n24508), .X(n29810) );
  sky130_fd_sc_hd__buf_6 U29622 ( .A(n30196), .X(n29811) );
  sky130_fd_sc_hd__buf_6 U29623 ( .A(n30196), .X(n29812) );
  sky130_fd_sc_hd__buf_4 U29625 ( .A(n30191), .X(n29813) );
  sky130_fd_sc_hd__buf_4 U29626 ( .A(n30191), .X(n29814) );
  sky130_fd_sc_hd__nand2_1 U29627 ( .A(n29525), .B(n12214), .Y(n24513) );
  sky130_fd_sc_hd__buf_6 U29628 ( .A(n24514), .X(n29815) );
  sky130_fd_sc_hd__buf_6 U29629 ( .A(n24514), .X(n29816) );
  sky130_fd_sc_hd__buf_6 U29630 ( .A(n11151), .X(n29817) );
  sky130_fd_sc_hd__buf_6 U29631 ( .A(n11151), .X(n29818) );
  sky130_fd_sc_hd__nand2_1 U29632 ( .A(n29301), .B(n24518), .Y(
        j202_soc_core_uart_TOP_N24) );
  sky130_fd_sc_hd__xnor2_1 U29633 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .Y(n24519) );
  sky130_fd_sc_hd__nor2_1 U29634 ( .A(n24519), .B(n29115), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[1]) );
  sky130_fd_sc_hd__a211oi_1 U29635 ( .A1(n24521), .A2(n24520), .B1(n24522), 
        .C1(n29115), .Y(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[3])
         );
  sky130_fd_sc_hd__nor2_1 U29637 ( .A(n24523), .B(n29115), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[4]) );
  sky130_fd_sc_hd__a21o_1 U29638 ( .A1(n24525), .A2(n24524), .B1(n29115), .X(
        n24526) );
  sky130_fd_sc_hd__nor2_1 U29639 ( .A(n24527), .B(n24526), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[5]) );
  sky130_fd_sc_hd__nand2b_1 U29640 ( .A_N(n29115), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]), .Y(n24528) );
  sky130_fd_sc_hd__nor2_1 U29641 ( .A(n24528), .B(n24530), .Y(n24535) );
  sky130_fd_sc_hd__nor2_1 U29642 ( .A(n29115), .B(n24535), .Y(n24532) );
  sky130_fd_sc_hd__a21oi_1 U29643 ( .A1(n24531), .A2(n24530), .B1(n24529), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[7]) );
  sky130_fd_sc_hd__nand2_1 U29644 ( .A(n24532), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .Y(n24533) );
  sky130_fd_sc_hd__o21ai_1 U29645 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .A2(n24534), .B1(
        n24533), .Y(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[8]) );
  sky130_fd_sc_hd__a22oi_1 U29646 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]), .A2(n28547), .B1(
        n24535), .B2(j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .Y(
        n24536) );
  sky130_fd_sc_hd__and3_1 U29647 ( .A(n24535), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .C(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]), .X(n28548) );
  sky130_fd_sc_hd__nor2_1 U29648 ( .A(n24536), .B(n28548), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[9]) );
  sky130_fd_sc_hd__nand3_1 U29649 ( .A(n24538), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .C(n28547), .Y(
        n24537) );
  sky130_fd_sc_hd__o21ai_1 U29650 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .A2(n24538), .B1(
        n24537), .Y(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[10]) );
  sky130_fd_sc_hd__inv_1 U29651 ( .A(n29528), .Y(n10585) );
  sky130_fd_sc_hd__inv_1 U29652 ( .A(n29529), .Y(n10587) );
  sky130_fd_sc_hd__inv_1 U29653 ( .A(n29530), .Y(n10588) );
  sky130_fd_sc_hd__inv_1 U29654 ( .A(n29531), .Y(n10584) );
  sky130_fd_sc_hd__inv_1 U29655 ( .A(n29532), .Y(n10581) );
  sky130_fd_sc_hd__inv_1 U29656 ( .A(n29533), .Y(n10582) );
  sky130_fd_sc_hd__inv_1 U29657 ( .A(n29534), .Y(n10596) );
  sky130_fd_sc_hd__inv_1 U29658 ( .A(n29535), .Y(n10593) );
  sky130_fd_sc_hd__inv_1 U29659 ( .A(n29536), .Y(n10594) );
  sky130_fd_sc_hd__inv_1 U29660 ( .A(n29537), .Y(n10595) );
  sky130_fd_sc_hd__inv_1 U29661 ( .A(n29538), .Y(n10592) );
  sky130_fd_sc_hd__inv_1 U29662 ( .A(n29539), .Y(n10589) );
  sky130_fd_sc_hd__nand4_1 U29663 ( .A(n24542), .B(n24541), .C(n24540), .D(
        n24539), .Y(n10574) );
  sky130_fd_sc_hd__nand2_1 U29664 ( .A(n24583), .B(n24547), .Y(n24548) );
  sky130_fd_sc_hd__nor2_1 U29665 ( .A(n24549), .B(n24548), .Y(n24555) );
  sky130_fd_sc_hd__nand4_1 U29666 ( .A(n24553), .B(n24555), .C(n24554), .D(
        n12350), .Y(n24556) );
  sky130_fd_sc_hd__o21ai_1 U29667 ( .A1(n24557), .A2(n24556), .B1(n28417), .Y(
        n24558) );
  sky130_fd_sc_hd__nand2_1 U29668 ( .A(n24558), .B(n28394), .Y(n10644) );
  sky130_fd_sc_hd__nand3_1 U29669 ( .A(n28133), .B(n12228), .C(n28267), .Y(
        n24561) );
  sky130_fd_sc_hd__nor2_1 U29670 ( .A(n24564), .B(n10960), .Y(n27740) );
  sky130_fd_sc_hd__nand2_1 U29671 ( .A(n27740), .B(n11646), .Y(n24565) );
  sky130_fd_sc_hd__nor2_1 U29672 ( .A(n11929), .B(n24565), .Y(n27980) );
  sky130_fd_sc_hd__nand3_1 U29673 ( .A(n24568), .B(n24567), .C(n24566), .Y(
        n24569) );
  sky130_fd_sc_hd__nand2_1 U29674 ( .A(n24569), .B(n28417), .Y(n24571) );
  sky130_fd_sc_hd__nand2_1 U29675 ( .A(n24571), .B(n24570), .Y(n10624) );
  sky130_fd_sc_hd__o22a_1 U29676 ( .A1(n24574), .A2(n24573), .B1(n11494), .B2(
        n24572), .X(n24575) );
  sky130_fd_sc_hd__nor2_1 U29677 ( .A(n24577), .B(n24576), .Y(n28270) );
  sky130_fd_sc_hd__nand4_1 U29678 ( .A(n24578), .B(n24579), .C(n11449), .D(
        n12219), .Y(n24580) );
  sky130_fd_sc_hd__nor2_1 U29679 ( .A(n24581), .B(n24580), .Y(n24582) );
  sky130_fd_sc_hd__nand3_1 U29680 ( .A(n28270), .B(n24583), .C(n24582), .Y(
        n24584) );
  sky130_fd_sc_hd__nand2_1 U29681 ( .A(n24584), .B(n28417), .Y(n24586) );
  sky130_fd_sc_hd__nand2_1 U29682 ( .A(n28360), .B(n24585), .Y(n27986) );
  sky130_fd_sc_hd__nand2b_1 U29683 ( .A_N(n27892), .B(n28355), .Y(n28145) );
  sky130_fd_sc_hd__nand2_1 U29684 ( .A(n24686), .B(n28145), .Y(n27751) );
  sky130_fd_sc_hd__nand2_1 U29685 ( .A(n27751), .B(n28355), .Y(n28272) );
  sky130_fd_sc_hd__nand3_1 U29686 ( .A(n24586), .B(n27986), .C(n28272), .Y(
        n10634) );
  sky130_fd_sc_hd__o21ai_1 U29687 ( .A1(n24588), .A2(n24587), .B1(n24589), .Y(
        j202_soc_core_j22_cpu_ma_N53) );
  sky130_fd_sc_hd__nand2_1 U29688 ( .A(n24589), .B(n29882), .Y(n24646) );
  sky130_fd_sc_hd__nor2_1 U29689 ( .A(n24590), .B(n24646), .Y(
        j202_soc_core_j22_cpu_ma_N54) );
  sky130_fd_sc_hd__nand2_1 U29690 ( .A(n28033), .B(n11659), .Y(n24595) );
  sky130_fd_sc_hd__nor2_1 U29691 ( .A(n27737), .B(n23950), .Y(n24600) );
  sky130_fd_sc_hd__nand2_1 U29692 ( .A(n30083), .B(n11449), .Y(n24598) );
  sky130_fd_sc_hd__nor2_1 U29693 ( .A(n24598), .B(n25146), .Y(n24599) );
  sky130_fd_sc_hd__o21ai_1 U29694 ( .A1(n24601), .A2(n12237), .B1(n28417), .Y(
        n24605) );
  sky130_fd_sc_hd__a21oi_1 U29695 ( .A1(n28360), .A2(n24603), .B1(n24602), .Y(
        n24604) );
  sky130_fd_sc_hd__nand2_1 U29696 ( .A(n24607), .B(n24606), .Y(n24608) );
  sky130_fd_sc_hd__a31oi_1 U29697 ( .A1(n24609), .A2(n27730), .A3(n24608), 
        .B1(n28379), .Y(j202_soc_core_j22_cpu_id_idec_N917) );
  sky130_fd_sc_hd__a21oi_1 U29698 ( .A1(n24610), .A2(n28417), .B1(n13072), .Y(
        n24611) );
  sky130_fd_sc_hd__nand2_1 U29700 ( .A(n24613), .B(n28367), .Y(n10645) );
  sky130_fd_sc_hd__nand2_1 U29701 ( .A(n24615), .B(n24614), .Y(n24637) );
  sky130_fd_sc_hd__o21ai_1 U29702 ( .A1(n24626), .A2(n24623), .B1(n28417), .Y(
        n24625) );
  sky130_fd_sc_hd__nand2_1 U29703 ( .A(n28083), .B(n24649), .Y(n24624) );
  sky130_fd_sc_hd__nand4_1 U29704 ( .A(n24625), .B(n25147), .C(n28078), .D(
        n12061), .Y(n10617) );
  sky130_fd_sc_hd__nand2_1 U29705 ( .A(n24629), .B(n24634), .Y(n24630) );
  sky130_fd_sc_hd__nand2_1 U29706 ( .A(n12064), .B(n24634), .Y(n24635) );
  sky130_fd_sc_hd__o211ai_1 U29707 ( .A1(n11142), .A2(n25904), .B1(n24636), 
        .C1(n24635), .Y(n24638) );
  sky130_fd_sc_hd__nor2_1 U29708 ( .A(n24637), .B(n24638), .Y(n24639) );
  sky130_fd_sc_hd__nand2_1 U29709 ( .A(n24641), .B(n28367), .Y(n10616) );
  sky130_fd_sc_hd__nand2_1 U29710 ( .A(n29587), .B(n28417), .Y(n24642) );
  sky130_fd_sc_hd__nand2_1 U29711 ( .A(n24642), .B(n28405), .Y(n10614) );
  sky130_fd_sc_hd__nand2_1 U29712 ( .A(n23549), .B(n28417), .Y(n24643) );
  sky130_fd_sc_hd__nand2_1 U29713 ( .A(n24643), .B(n28405), .Y(n10615) );
  sky130_fd_sc_hd__nand2_1 U29714 ( .A(n12669), .B(n28417), .Y(n24644) );
  sky130_fd_sc_hd__nand2_1 U29715 ( .A(n24644), .B(n28405), .Y(n10613) );
  sky130_fd_sc_hd__nand2_1 U29716 ( .A(n29593), .B(n28417), .Y(n24645) );
  sky130_fd_sc_hd__nand2_1 U29717 ( .A(n24645), .B(n28405), .Y(n10612) );
  sky130_fd_sc_hd__nor2_1 U29718 ( .A(n12041), .B(n24646), .Y(
        j202_soc_core_j22_cpu_ma_N55) );
  sky130_fd_sc_hd__nor2_1 U29719 ( .A(n24647), .B(n24646), .Y(
        j202_soc_core_j22_cpu_ma_N56) );
  sky130_fd_sc_hd__nor2_1 U29720 ( .A(n28036), .B(n24648), .Y(n24657) );
  sky130_fd_sc_hd__nand2_1 U29721 ( .A(n24649), .B(n28352), .Y(n28031) );
  sky130_fd_sc_hd__a31oi_1 U29722 ( .A1(n11389), .A2(n28417), .A3(n12326), 
        .B1(n28031), .Y(n24650) );
  sky130_fd_sc_hd__nand2b_1 U29723 ( .A_N(n24657), .B(n24650), .Y(n10638) );
  sky130_fd_sc_hd__nand2_1 U29724 ( .A(n24652), .B(n28346), .Y(n10599) );
  sky130_fd_sc_hd__nand2_1 U29725 ( .A(n28083), .B(n28357), .Y(n28342) );
  sky130_fd_sc_hd__inv_1 U29726 ( .A(n24654), .Y(n24656) );
  sky130_fd_sc_hd__nand3_1 U29727 ( .A(n11389), .B(n10957), .C(n12326), .Y(
        n24655) );
  sky130_fd_sc_hd__nand3_1 U29728 ( .A(n24656), .B(n27886), .C(n24655), .Y(
        n24661) );
  sky130_fd_sc_hd__a21oi_1 U29729 ( .A1(n24661), .A2(n28417), .B1(n24657), .Y(
        n24658) );
  sky130_fd_sc_hd__nand2_1 U29730 ( .A(n24659), .B(n24658), .Y(n10639) );
  sky130_fd_sc_hd__nand3_1 U29731 ( .A(n28148), .B(n24660), .C(n12287), .Y(
        n24662) );
  sky130_fd_sc_hd__o21ai_1 U29732 ( .A1(n24662), .A2(n24661), .B1(n28417), .Y(
        n24664) );
  sky130_fd_sc_hd__nand2_1 U29733 ( .A(n24664), .B(n24663), .Y(n10640) );
  sky130_fd_sc_hd__nand3_1 U29734 ( .A(n24666), .B(n27052), .C(
        j202_soc_core_j22_cpu_rfuo_sr__s_), .Y(n27754) );
  sky130_fd_sc_hd__nand4_1 U29735 ( .A(n27757), .B(n29746), .C(n27756), .D(
        n27754), .Y(n28423) );
  sky130_fd_sc_hd__nor3_1 U29736 ( .A(n27052), .B(n24668), .C(n24667), .Y(
        n24669) );
  sky130_fd_sc_hd__nand3_1 U29737 ( .A(n29746), .B(n24670), .C(n24669), .Y(
        n28422) );
  sky130_fd_sc_hd__o21ai_1 U29738 ( .A1(n27828), .A2(n28423), .B1(n28422), .Y(
        j202_soc_core_j22_cpu_ml_N191) );
  sky130_fd_sc_hd__nand2_1 U29739 ( .A(n28109), .B(n24671), .Y(n28052) );
  sky130_fd_sc_hd__nor2_1 U29740 ( .A(n13325), .B(n27760), .Y(n28050) );
  sky130_fd_sc_hd__nand2_1 U29741 ( .A(n24676), .B(n24675), .Y(n28048) );
  sky130_fd_sc_hd__o21ai_1 U29742 ( .A1(n28047), .A2(n24677), .B1(n28048), .Y(
        n24678) );
  sky130_fd_sc_hd__a21oi_1 U29743 ( .A1(n28050), .A2(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]), .B1(n24678), .Y(n24679) );
  sky130_fd_sc_hd__o22ai_1 U29745 ( .A1(n11180), .A2(n27859), .B1(n27858), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N3317) );
  sky130_fd_sc_hd__nand2_1 U29746 ( .A(n28360), .B(n24685), .Y(n28154) );
  sky130_fd_sc_hd__o211ai_1 U29747 ( .A1(j202_soc_core_j22_cpu_opst[0]), .A2(
        n28394), .B1(n28154), .C1(n24686), .Y(n24687) );
  sky130_fd_sc_hd__a21oi_1 U29748 ( .A1(n24688), .A2(n28417), .B1(n24687), .Y(
        n24689) );
  sky130_fd_sc_hd__nand2_1 U29749 ( .A(n28083), .B(n24689), .Y(n10526) );
  sky130_fd_sc_hd__nor2_1 U29751 ( .A(n28198), .B(n27751), .Y(n28074) );
  sky130_fd_sc_hd__nand4_1 U29752 ( .A(n24694), .B(n28074), .C(n28352), .D(
        n28361), .Y(n10527) );
  sky130_fd_sc_hd__a21oi_1 U29753 ( .A1(n28360), .A2(n24697), .B1(n24696), .Y(
        n24698) );
  sky130_fd_sc_hd__o21ai_1 U29754 ( .A1(n24699), .A2(n24700), .B1(n28417), .Y(
        n24701) );
  sky130_fd_sc_hd__nand2_1 U29755 ( .A(n24701), .B(n28394), .Y(n10643) );
  sky130_fd_sc_hd__mux2i_1 U29756 ( .A0(n27988), .A1(n11180), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3278) );
  sky130_fd_sc_hd__a21oi_1 U29757 ( .A1(n24703), .A2(n24702), .B1(n28084), .Y(
        n24706) );
  sky130_fd_sc_hd__or4_1 U29758 ( .A(n24708), .B(n24707), .C(n24706), .D(
        n24705), .X(n24709) );
  sky130_fd_sc_hd__o21ai_1 U29759 ( .A1(n24710), .A2(n24709), .B1(n29827), .Y(
        n10597) );
  sky130_fd_sc_hd__nand2_1 U29760 ( .A(n28383), .B(n24711), .Y(n10646) );
  sky130_fd_sc_hd__nor2_1 U29761 ( .A(n27644), .B(n27988), .Y(
        j202_soc_core_j22_cpu_rf_N2649) );
  sky130_fd_sc_hd__o22ai_1 U29762 ( .A1(n11180), .A2(n27841), .B1(n24712), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N3241) );
  sky130_fd_sc_hd__o22ai_1 U29763 ( .A1(n11180), .A2(n25964), .B1(n27847), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N2686) );
  sky130_fd_sc_hd__a2bb2oi_1 U29764 ( .B1(n24713), .B2(n27862), .A1_N(n27774), 
        .A2_N(n11180), .Y(n24714) );
  sky130_fd_sc_hd__o21ai_0 U29765 ( .A1(n27648), .A2(n27988), .B1(n24714), .Y(
        j202_soc_core_j22_cpu_rf_N3352) );
  sky130_fd_sc_hd__nor2_1 U29766 ( .A(n24771), .B(n24715), .Y(n26157) );
  sky130_fd_sc_hd__nand2_1 U29767 ( .A(n28109), .B(n26157), .Y(n27753) );
  sky130_fd_sc_hd__o31ai_1 U29768 ( .A1(n24718), .A2(n24717), .A3(n24716), 
        .B1(n27753), .Y(j202_soc_core_j22_cpu_rf_N2627) );
  sky130_fd_sc_hd__nand2_1 U29769 ( .A(n24721), .B(j202_soc_core_uart_RDRXD1), 
        .Y(n27961) );
  sky130_fd_sc_hd__nor2_1 U29770 ( .A(n27957), .B(n27961), .Y(n27952) );
  sky130_fd_sc_hd__o22ai_1 U29771 ( .A1(n24723), .A2(n27961), .B1(n24722), 
        .B2(n27952), .Y(n104) );
  sky130_fd_sc_hd__nand3_1 U29772 ( .A(n24725), .B(n24724), .C(
        j202_soc_core_ahb2apb_00_state[0]), .Y(n24751) );
  sky130_fd_sc_hd__o22ai_1 U29773 ( .A1(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[0]), .A2(n24751), .B1(
        n24728), .B2(n24727), .Y(
        j202_soc_core_cmt_core_00_cmt_apb_00_nxt_state_0_) );
  sky130_fd_sc_hd__nor2_1 U29774 ( .A(n24729), .B(n24751), .Y(
        j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen) );
  sky130_fd_sc_hd__nand2_1 U29775 ( .A(n28222), .B(
        j202_soc_core_cmt_core_00_reg_addr[3]), .Y(n24758) );
  sky130_fd_sc_hd__nand2_1 U29776 ( .A(n24739), .B(n24732), .Y(n28287) );
  sky130_fd_sc_hd__nand2_1 U29778 ( .A(n24731), .B(n24730), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_nxt_latch_status_0_) );
  sky130_fd_sc_hd__nand2_1 U29779 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[7]), .Y(n24733) );
  sky130_fd_sc_hd__o21ai_1 U29780 ( .A1(n27550), .A2(n28289), .B1(n24733), .Y(
        n114) );
  sky130_fd_sc_hd__nand2_1 U29781 ( .A(n28287), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[4]), .Y(n24734) );
  sky130_fd_sc_hd__o21ai_1 U29782 ( .A1(n24741), .A2(n28287), .B1(n24734), .Y(
        n73) );
  sky130_fd_sc_hd__nand2_1 U29783 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[4]), .Y(n24735) );
  sky130_fd_sc_hd__o21ai_1 U29784 ( .A1(n24741), .A2(n28289), .B1(n24735), .Y(
        n75) );
  sky130_fd_sc_hd__nand2_1 U29785 ( .A(n28221), .B(
        j202_soc_core_cmt_core_00_reg_addr[2]), .Y(n24757) );
  sky130_fd_sc_hd__nand2_1 U29786 ( .A(n24738), .B(n24736), .Y(n28291) );
  sky130_fd_sc_hd__nand2_1 U29787 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[4]), .Y(n24737) );
  sky130_fd_sc_hd__o21ai_1 U29788 ( .A1(n24741), .A2(n28291), .B1(n24737), .Y(
        n74) );
  sky130_fd_sc_hd__nand2_1 U29789 ( .A(n24739), .B(n24738), .Y(n28293) );
  sky130_fd_sc_hd__nand2_1 U29790 ( .A(n28293), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[4]), .Y(n24740) );
  sky130_fd_sc_hd__nand2_1 U29792 ( .A(n28287), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[6]), .Y(n24742) );
  sky130_fd_sc_hd__o21ai_1 U29793 ( .A1(n27465), .A2(n28287), .B1(n24742), .Y(
        n110) );
  sky130_fd_sc_hd__nand2_1 U29794 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[6]), .Y(n24743) );
  sky130_fd_sc_hd__o21ai_1 U29795 ( .A1(n27465), .A2(n28289), .B1(n24743), .Y(
        n112) );
  sky130_fd_sc_hd__nand2_1 U29796 ( .A(n28293), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[6]), .Y(n24744) );
  sky130_fd_sc_hd__o21ai_1 U29797 ( .A1(n27465), .A2(n28293), .B1(n24744), .Y(
        n134) );
  sky130_fd_sc_hd__nand2_1 U29798 ( .A(n28287), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[5]), .Y(n24745) );
  sky130_fd_sc_hd__o21ai_1 U29799 ( .A1(n24749), .A2(n28287), .B1(n24745), .Y(
        n107) );
  sky130_fd_sc_hd__nand2_1 U29800 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[5]), .Y(n24746) );
  sky130_fd_sc_hd__o21ai_1 U29801 ( .A1(n24749), .A2(n28289), .B1(n24746), .Y(
        n109) );
  sky130_fd_sc_hd__nand2_1 U29802 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[5]), .Y(n24747) );
  sky130_fd_sc_hd__o21ai_1 U29803 ( .A1(n24749), .A2(n28291), .B1(n24747), .Y(
        n108) );
  sky130_fd_sc_hd__nand2_1 U29804 ( .A(n28293), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[5]), .Y(n24748) );
  sky130_fd_sc_hd__o21ai_1 U29805 ( .A1(n24749), .A2(n28293), .B1(n24748), .Y(
        n106) );
  sky130_fd_sc_hd__nor2_1 U29806 ( .A(j202_soc_core_pwrite[0]), .B(n24751), 
        .Y(n24753) );
  sky130_fd_sc_hd__nand2_1 U29807 ( .A(n24752), .B(n24753), .Y(n24756) );
  sky130_fd_sc_hd__nor2_1 U29808 ( .A(n24758), .B(n24756), .Y(n28296) );
  sky130_fd_sc_hd__nand2_1 U29809 ( .A(n28222), .B(n28221), .Y(n28211) );
  sky130_fd_sc_hd__a22oi_1 U29810 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[5]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[5]), .Y(
        n24762) );
  sky130_fd_sc_hd__nand2_1 U29811 ( .A(n24754), .B(n24753), .Y(n28219) );
  sky130_fd_sc_hd__nor2_1 U29812 ( .A(n28219), .B(n24755), .Y(n28297) );
  sky130_fd_sc_hd__nor2_1 U29813 ( .A(n28219), .B(n24757), .Y(n28299) );
  sky130_fd_sc_hd__a22oi_1 U29814 ( .A1(n28297), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[5]), 
        .B1(n28299), .B2(j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[5]), .Y(
        n24761) );
  sky130_fd_sc_hd__nor2_1 U29815 ( .A(n24757), .B(n24756), .Y(n28301) );
  sky130_fd_sc_hd__nand2_1 U29816 ( .A(n28301), .B(
        j202_soc_core_cmt_core_00_const0[5]), .Y(n24760) );
  sky130_fd_sc_hd__nor2_1 U29817 ( .A(n28219), .B(n24758), .Y(n28300) );
  sky130_fd_sc_hd__nand2_1 U29818 ( .A(n28300), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[5]), .Y(n24759) );
  sky130_fd_sc_hd__nand4_1 U29819 ( .A(n24762), .B(n24761), .C(n24760), .D(
        n24759), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[5]) );
  sky130_fd_sc_hd__a21oi_1 U29820 ( .A1(n24765), .A2(n24764), .B1(n24763), .Y(
        n24766) );
  sky130_fd_sc_hd__inv_2 U29821 ( .A(n27766), .Y(n25374) );
  sky130_fd_sc_hd__o21ai_1 U29822 ( .A1(n24766), .A2(n27770), .B1(n25374), .Y(
        j202_soc_core_j22_cpu_ml_maclj[28]) );
  sky130_fd_sc_hd__mux2i_1 U29823 ( .A0(n24779), .A1(n11190), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N306) );
  sky130_fd_sc_hd__nand2_1 U29824 ( .A(n28055), .B(n24772), .Y(n24768) );
  sky130_fd_sc_hd__nand2_1 U29825 ( .A(n28056), .B(n21219), .Y(n24767) );
  sky130_fd_sc_hd__nand3_1 U29826 ( .A(n24768), .B(n12203), .C(n24767), .Y(
        j202_soc_core_j22_cpu_ml_machj[3]) );
  sky130_fd_sc_hd__inv_1 U29827 ( .A(n24769), .Y(n24774) );
  sky130_fd_sc_hd__o22ai_1 U29828 ( .A1(n24779), .A2(n27859), .B1(n27858), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N3313) );
  sky130_fd_sc_hd__mux2i_1 U29829 ( .A0(n24778), .A1(n24779), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3273) );
  sky130_fd_sc_hd__o22ai_1 U29830 ( .A1(n24771), .A2(n27364), .B1(n27644), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N2645) );
  sky130_fd_sc_hd__o22ai_1 U29831 ( .A1(n24779), .A2(n27841), .B1(n24712), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N3236) );
  sky130_fd_sc_hd__o22ai_1 U29832 ( .A1(n24779), .A2(n25964), .B1(n27847), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N2681) );
  sky130_fd_sc_hd__nor2_1 U29833 ( .A(n27355), .B(n27648), .Y(n27772) );
  sky130_fd_sc_hd__nand2_1 U29834 ( .A(n24772), .B(n27772), .Y(n24777) );
  sky130_fd_sc_hd__nand2_1 U29835 ( .A(n24774), .B(n27860), .Y(n24775) );
  sky130_fd_sc_hd__nand3_1 U29836 ( .A(n24777), .B(n24776), .C(n24775), .Y(
        j202_soc_core_j22_cpu_rf_N3348) );
  sky130_fd_sc_hd__o22ai_1 U29837 ( .A1(n24779), .A2(n25977), .B1(n28061), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N2866) );
  sky130_fd_sc_hd__o22ai_1 U29838 ( .A1(n24779), .A2(n25978), .B1(n27834), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N2940) );
  sky130_fd_sc_hd__o22ai_1 U29839 ( .A1(n24779), .A2(n25979), .B1(n28112), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N3199) );
  sky130_fd_sc_hd__o22ai_1 U29840 ( .A1(n24779), .A2(n25980), .B1(n27835), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N2792) );
  sky130_fd_sc_hd__o22ai_1 U29841 ( .A1(n24779), .A2(n25981), .B1(n27836), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N3162) );
  sky130_fd_sc_hd__o22ai_1 U29842 ( .A1(n24779), .A2(n25982), .B1(n27837), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N3014) );
  sky130_fd_sc_hd__o22ai_1 U29843 ( .A1(n24779), .A2(n25983), .B1(n27838), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N3051) );
  sky130_fd_sc_hd__o22ai_1 U29844 ( .A1(n24779), .A2(n26894), .B1(n27839), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N2903) );
  sky130_fd_sc_hd__o22ai_1 U29845 ( .A1(n24779), .A2(n25984), .B1(n27840), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N2718) );
  sky130_fd_sc_hd__o22ai_1 U29846 ( .A1(n24779), .A2(n25985), .B1(n27842), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N3088) );
  sky130_fd_sc_hd__o22ai_1 U29847 ( .A1(n24779), .A2(n25986), .B1(n27843), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N2977) );
  sky130_fd_sc_hd__o22ai_1 U29848 ( .A1(n24779), .A2(n25987), .B1(n27844), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N3125) );
  sky130_fd_sc_hd__o22ai_1 U29849 ( .A1(n24779), .A2(n25988), .B1(n27845), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N2829) );
  sky130_fd_sc_hd__o22ai_1 U29850 ( .A1(n24779), .A2(n25989), .B1(n27846), 
        .B2(n24778), .Y(j202_soc_core_j22_cpu_rf_N2755) );
  sky130_fd_sc_hd__nor4_1 U29851 ( .A(j202_soc_core_intc_core_00_bs_addr[5]), 
        .B(j202_soc_core_intc_core_00_bs_addr[4]), .C(
        j202_soc_core_intc_core_00_bs_addr[9]), .D(n24780), .Y(n24786) );
  sky130_fd_sc_hd__nor2_1 U29852 ( .A(j202_soc_core_intc_core_00_bs_addr[11]), 
        .B(j202_soc_core_intc_core_00_bs_addr[10]), .Y(n24783) );
  sky130_fd_sc_hd__nand4_1 U29853 ( .A(j202_soc_core_pstrb[5]), .B(
        j202_soc_core_pstrb[4]), .C(j202_soc_core_pstrb[6]), .D(
        j202_soc_core_pstrb[7]), .Y(n24781) );
  sky130_fd_sc_hd__nand2_1 U29854 ( .A(j202_soc_core_pwrite[1]), .B(n24781), 
        .Y(n24782) );
  sky130_fd_sc_hd__nand2_1 U29855 ( .A(n24783), .B(n24782), .Y(n24784) );
  sky130_fd_sc_hd__nor2_1 U29856 ( .A(n24785), .B(n24784), .Y(n27416) );
  sky130_fd_sc_hd__nor2_1 U29857 ( .A(j202_soc_core_intc_core_00_bs_addr[1]), 
        .B(j202_soc_core_intc_core_00_bs_addr[0]), .Y(n25073) );
  sky130_fd_sc_hd__nand3_1 U29858 ( .A(n25073), .B(n25072), .C(n29403), .Y(
        n25090) );
  sky130_fd_sc_hd__nand3_1 U29859 ( .A(n24786), .B(n27416), .C(n29406), .Y(
        n25081) );
  sky130_fd_sc_hd__nor3_1 U29860 ( .A(j202_soc_core_intc_core_00_bs_addr[6]), 
        .B(n25061), .C(n25081), .Y(n29143) );
  sky130_fd_sc_hd__nand2_1 U29861 ( .A(n28064), .B(n29827), .Y(n28063) );
  sky130_fd_sc_hd__o22ai_1 U29862 ( .A1(n29161), .A2(n28064), .B1(n27352), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U29863 ( .A1(n29152), .A2(n28064), .B1(n27312), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__nand2_1 U29864 ( .A(n28109), .B(
        j202_soc_core_j22_cpu_intack), .Y(n26860) );
  sky130_fd_sc_hd__nand2_1 U29865 ( .A(n26860), .B(n29827), .Y(n29073) );
  sky130_fd_sc_hd__o22ai_1 U29866 ( .A1(n29073), .A2(n26674), .B1(n24787), 
        .B2(n29070), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N5) );
  sky130_fd_sc_hd__o22ai_1 U29867 ( .A1(n24788), .A2(n27859), .B1(n27858), 
        .B2(n24791), .Y(j202_soc_core_j22_cpu_rf_N3309) );
  sky130_fd_sc_hd__nor2_1 U29868 ( .A(n27644), .B(n24791), .Y(
        j202_soc_core_j22_cpu_rf_N2643) );
  sky130_fd_sc_hd__o22ai_1 U29869 ( .A1(n24788), .A2(n27841), .B1(n24712), 
        .B2(n11164), .Y(j202_soc_core_j22_cpu_rf_N3234) );
  sky130_fd_sc_hd__o22ai_1 U29870 ( .A1(n24788), .A2(n25977), .B1(n28061), 
        .B2(n24791), .Y(j202_soc_core_j22_cpu_rf_N2864) );
  sky130_fd_sc_hd__o22ai_1 U29871 ( .A1(n24788), .A2(n25978), .B1(n27834), 
        .B2(n11164), .Y(j202_soc_core_j22_cpu_rf_N2938) );
  sky130_fd_sc_hd__o22ai_1 U29872 ( .A1(n24788), .A2(n25979), .B1(n28112), 
        .B2(n11164), .Y(j202_soc_core_j22_cpu_rf_N3197) );
  sky130_fd_sc_hd__o22ai_1 U29873 ( .A1(n24788), .A2(n25980), .B1(n27835), 
        .B2(n11164), .Y(j202_soc_core_j22_cpu_rf_N2790) );
  sky130_fd_sc_hd__o22ai_1 U29874 ( .A1(n24788), .A2(n25981), .B1(n27836), 
        .B2(n11164), .Y(j202_soc_core_j22_cpu_rf_N3160) );
  sky130_fd_sc_hd__o22ai_1 U29875 ( .A1(n24788), .A2(n25982), .B1(n27837), 
        .B2(n11164), .Y(j202_soc_core_j22_cpu_rf_N3012) );
  sky130_fd_sc_hd__o22ai_1 U29876 ( .A1(n24788), .A2(n25983), .B1(n27838), 
        .B2(n11164), .Y(j202_soc_core_j22_cpu_rf_N3049) );
  sky130_fd_sc_hd__o22ai_1 U29877 ( .A1(n24788), .A2(n26894), .B1(n27839), 
        .B2(n24791), .Y(j202_soc_core_j22_cpu_rf_N2901) );
  sky130_fd_sc_hd__o22ai_1 U29878 ( .A1(n24788), .A2(n25984), .B1(n27840), 
        .B2(n24791), .Y(j202_soc_core_j22_cpu_rf_N2716) );
  sky130_fd_sc_hd__o22ai_1 U29879 ( .A1(n24788), .A2(n25985), .B1(n27842), 
        .B2(n24791), .Y(j202_soc_core_j22_cpu_rf_N3086) );
  sky130_fd_sc_hd__o22ai_1 U29880 ( .A1(n24788), .A2(n25986), .B1(n27843), 
        .B2(n11164), .Y(j202_soc_core_j22_cpu_rf_N2975) );
  sky130_fd_sc_hd__o22ai_1 U29881 ( .A1(n24788), .A2(n25987), .B1(n27844), 
        .B2(n11164), .Y(j202_soc_core_j22_cpu_rf_N3123) );
  sky130_fd_sc_hd__o22ai_1 U29882 ( .A1(n24788), .A2(n25988), .B1(n27845), 
        .B2(n11164), .Y(j202_soc_core_j22_cpu_rf_N2827) );
  sky130_fd_sc_hd__o22ai_1 U29883 ( .A1(n24788), .A2(n25989), .B1(n27846), 
        .B2(n24791), .Y(j202_soc_core_j22_cpu_rf_N2753) );
  sky130_fd_sc_hd__o22ai_1 U29884 ( .A1(n24788), .A2(n25964), .B1(n27847), 
        .B2(n11164), .Y(j202_soc_core_j22_cpu_rf_N2679) );
  sky130_fd_sc_hd__a22oi_1 U29885 ( .A1(n27862), .A2(n24792), .B1(n12431), 
        .B2(n27861), .Y(n24793) );
  sky130_fd_sc_hd__o21ai_0 U29886 ( .A1(n27648), .A2(n11164), .B1(n24793), .Y(
        j202_soc_core_j22_cpu_rf_N3346) );
  sky130_fd_sc_hd__mux2i_1 U29887 ( .A0(n24788), .A1(n26284), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N304) );
  sky130_fd_sc_hd__nand2_1 U29888 ( .A(n28055), .B(n24794), .Y(n24795) );
  sky130_fd_sc_hd__nand2_1 U29889 ( .A(n24795), .B(n12203), .Y(
        j202_soc_core_j22_cpu_ml_machj[1]) );
  sky130_fd_sc_hd__mux2i_1 U29890 ( .A0(n28480), .A1(n26944), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N312) );
  sky130_fd_sc_hd__nand2_1 U29891 ( .A(n28055), .B(n24904), .Y(n24801) );
  sky130_fd_sc_hd__nand2_1 U29892 ( .A(n28056), .B(n24799), .Y(n24800) );
  sky130_fd_sc_hd__nand3_1 U29893 ( .A(n24801), .B(n12203), .C(n24800), .Y(
        j202_soc_core_j22_cpu_ml_machj[9]) );
  sky130_fd_sc_hd__buf_2 U29894 ( .A(n24802), .X(n27159) );
  sky130_fd_sc_hd__o22ai_1 U29895 ( .A1(n27433), .A2(n25977), .B1(n28061), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N2868) );
  sky130_fd_sc_hd__o22ai_1 U29896 ( .A1(n27433), .A2(n25978), .B1(n27834), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N2942) );
  sky130_fd_sc_hd__o22ai_1 U29897 ( .A1(n27433), .A2(n25979), .B1(n28112), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N3201) );
  sky130_fd_sc_hd__o22ai_1 U29898 ( .A1(n27433), .A2(n25980), .B1(n27835), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N2794) );
  sky130_fd_sc_hd__o22ai_1 U29899 ( .A1(n27433), .A2(n25981), .B1(n27836), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N3164) );
  sky130_fd_sc_hd__o22ai_1 U29900 ( .A1(n27433), .A2(n25982), .B1(n27837), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N3016) );
  sky130_fd_sc_hd__o22ai_1 U29901 ( .A1(n27433), .A2(n25983), .B1(n27838), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N3053) );
  sky130_fd_sc_hd__o22ai_1 U29902 ( .A1(n27433), .A2(n26894), .B1(n27839), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N2905) );
  sky130_fd_sc_hd__o22ai_1 U29903 ( .A1(n27433), .A2(n25984), .B1(n27840), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N2720) );
  sky130_fd_sc_hd__o22ai_1 U29904 ( .A1(n27433), .A2(n27841), .B1(n24712), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N3238) );
  sky130_fd_sc_hd__o22ai_1 U29905 ( .A1(n27433), .A2(n25985), .B1(n27842), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N3090) );
  sky130_fd_sc_hd__o22ai_1 U29906 ( .A1(n27433), .A2(n25986), .B1(n27843), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N2979) );
  sky130_fd_sc_hd__o22ai_1 U29907 ( .A1(n27433), .A2(n25987), .B1(n27844), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N3127) );
  sky130_fd_sc_hd__o22ai_1 U29908 ( .A1(n27433), .A2(n25988), .B1(n27845), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N2831) );
  sky130_fd_sc_hd__o22ai_1 U29909 ( .A1(n27433), .A2(n25989), .B1(n27846), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N2757) );
  sky130_fd_sc_hd__o22ai_1 U29910 ( .A1(n27433), .A2(n25964), .B1(n27847), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N2683) );
  sky130_fd_sc_hd__mux2i_1 U29911 ( .A0(n24805), .A1(n27433), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3275) );
  sky130_fd_sc_hd__o22ai_1 U29912 ( .A1(n27433), .A2(n27859), .B1(n27858), 
        .B2(n24805), .Y(j202_soc_core_j22_cpu_rf_N3315) );
  sky130_fd_sc_hd__nor2_1 U29913 ( .A(n27644), .B(n24805), .Y(
        j202_soc_core_j22_cpu_rf_N2647) );
  sky130_fd_sc_hd__a22oi_1 U29914 ( .A1(n24803), .A2(n27862), .B1(n28501), 
        .B2(n27861), .Y(n24804) );
  sky130_fd_sc_hd__o21ai_0 U29915 ( .A1(n27648), .A2(n24805), .B1(n24804), .Y(
        j202_soc_core_j22_cpu_rf_N3350) );
  sky130_fd_sc_hd__nor2_1 U29916 ( .A(j202_soc_core_intc_core_00_bs_addr[5]), 
        .B(j202_soc_core_intc_core_00_bs_addr[4]), .Y(n24807) );
  sky130_fd_sc_hd__nor3_1 U29917 ( .A(j202_soc_core_intc_core_00_bs_addr[7]), 
        .B(j202_soc_core_intc_core_00_bs_addr[6]), .C(n27414), .Y(n24806) );
  sky130_fd_sc_hd__nand3_1 U29918 ( .A(n27416), .B(n24807), .C(n24806), .Y(
        n25088) );
  sky130_fd_sc_hd__nor2_1 U29919 ( .A(j202_soc_core_intc_core_00_bs_addr[8]), 
        .B(n25088), .Y(n25074) );
  sky130_fd_sc_hd__nand2_1 U29920 ( .A(n25074), .B(n29406), .Y(n25096) );
  sky130_fd_sc_hd__nand2_1 U29921 ( .A(n24808), .B(j202_soc_core_pwrite[1]), 
        .Y(n27575) );
  sky130_fd_sc_hd__nand2_1 U29922 ( .A(n27575), .B(n12069), .Y(n27573) );
  sky130_fd_sc_hd__o22ai_1 U29923 ( .A1(n29163), .A2(n27575), .B1(n24809), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U29924 ( .A1(n29159), .A2(n27575), .B1(n24810), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__mux2i_1 U29925 ( .A0(n27668), .A1(n11188), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N303) );
  sky130_fd_sc_hd__nand2_1 U29926 ( .A(n28055), .B(n27645), .Y(n24811) );
  sky130_fd_sc_hd__o22ai_1 U29927 ( .A1(n29165), .A2(n28064), .B1(n24816), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__nand4_1 U29928 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[6]), .B(j202_soc_core_intc_core_00_cp_intack_all_0_), .C(n25736), .D(n29069), .Y(
        n24820) );
  sky130_fd_sc_hd__nor2_1 U29929 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .B(n24820), .Y(n26719) );
  sky130_fd_sc_hd__nor2_1 U29930 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]), .B(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[3]), .Y(n27350) );
  sky130_fd_sc_hd__a21oi_1 U29931 ( .A1(n26719), .A2(n27350), .B1(
        j202_soc_core_intc_core_00_rg_irqc[0]), .Y(n24814) );
  sky130_fd_sc_hd__nor2_1 U29932 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[0]), 
        .B(n24812), .Y(n24813) );
  sky130_fd_sc_hd__a31oi_1 U29933 ( .A1(n24814), .A2(
        j202_soc_core_intc_core_00_in_intreq[0]), .A3(n29827), .B1(n24813), 
        .Y(n24815) );
  sky130_fd_sc_hd__nor2_1 U29934 ( .A(n24816), .B(n24815), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N3) );
  sky130_fd_sc_hd__nand3_1 U29935 ( .A(n25063), .B(j202_soc_core_pwrite[1]), 
        .C(j202_soc_core_intc_core_00_bs_addr[8]), .Y(n25077) );
  sky130_fd_sc_hd__nor2_1 U29936 ( .A(n25090), .B(n25077), .Y(n26704) );
  sky130_fd_sc_hd__nor2_1 U29937 ( .A(n29088), .B(
        j202_soc_core_qspi_wb_wdat[0]), .Y(n28246) );
  sky130_fd_sc_hd__o22ai_1 U29938 ( .A1(n26704), .A2(n24819), .B1(n28246), 
        .B2(n26702), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U29939 ( .A1(n29163), .A2(n28064), .B1(n24822), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__nor2_1 U29940 ( .A(n24820), .B(n27349), .Y(n26713) );
  sky130_fd_sc_hd__nand2_1 U29941 ( .A(n26713), .B(n27350), .Y(n24821) );
  sky130_fd_sc_hd__nand4b_1 U29942 ( .A_N(
        j202_soc_core_intc_core_00_rg_irqc[1]), .B(n24821), .C(
        j202_soc_core_intc_core_00_in_intreq[1]), .D(n12069), .Y(n24824) );
  sky130_fd_sc_hd__nand2b_1 U29943 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[1]), 
        .B(n29544), .Y(n24823) );
  sky130_fd_sc_hd__a21oi_1 U29944 ( .A1(n24824), .A2(n24823), .B1(n24822), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N4) );
  sky130_fd_sc_hd__nor2_1 U29945 ( .A(n29088), .B(
        j202_soc_core_qspi_wb_wdat[4]), .Y(n28931) );
  sky130_fd_sc_hd__o22ai_1 U29946 ( .A1(n26704), .A2(n24825), .B1(n28931), 
        .B2(n26702), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__nor2_1 U29947 ( .A(n25061), .B(n29165), .Y(n29405) );
  sky130_fd_sc_hd__o22ai_1 U29948 ( .A1(n25096), .A2(n29399), .B1(n24826), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U29949 ( .A1(n29160), .A2(n27575), .B1(n24827), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__a21oi_1 U29951 ( .A1(n24829), .A2(n28056), .B1(n25776), .Y(
        n24830) );
  sky130_fd_sc_hd__o21ai_1 U29952 ( .A1(n24831), .A2(n25779), .B1(n24830), .Y(
        n29833) );
  sky130_fd_sc_hd__nand2_4 U29953 ( .A(n24833), .B(n30076), .Y(n28537) );
  sky130_fd_sc_hd__nand2_1 U29954 ( .A(n26414), .B(n27052), .Y(n25658) );
  sky130_fd_sc_hd__o22ai_1 U29955 ( .A1(n26317), .A2(n27799), .B1(n11188), 
        .B2(n27797), .Y(n24843) );
  sky130_fd_sc_hd__o22ai_1 U29956 ( .A1(n26430), .A2(n27795), .B1(n26323), 
        .B2(n26943), .Y(n24842) );
  sky130_fd_sc_hd__xor2_1 U29957 ( .A(n27111), .B(n28532), .X(n26226) );
  sky130_fd_sc_hd__nand2_1 U29958 ( .A(n27810), .B(n27115), .Y(n24834) );
  sky130_fd_sc_hd__o22a_1 U29960 ( .A1(n26926), .A2(n24837), .B1(n27355), .B2(
        n24836), .X(n24838) );
  sky130_fd_sc_hd__o21ai_0 U29961 ( .A1(n26320), .A2(n27803), .B1(n24838), .Y(
        n24839) );
  sky130_fd_sc_hd__a211o_1 U29962 ( .A1(n27808), .A2(n26009), .B1(n24840), 
        .C1(n24839), .X(n24841) );
  sky130_fd_sc_hd__nor3_1 U29963 ( .A(n24843), .B(n24842), .C(n24841), .Y(
        n24846) );
  sky130_fd_sc_hd__mux2_2 U29964 ( .A0(n27817), .A1(n27793), .S(n28532), .X(
        n24845) );
  sky130_fd_sc_hd__nand2_1 U29965 ( .A(n25648), .B(n28541), .Y(n24844) );
  sky130_fd_sc_hd__nand4_1 U29966 ( .A(n27814), .B(n24846), .C(n24845), .D(
        n24844), .Y(n24847) );
  sky130_fd_sc_hd__a21oi_1 U29967 ( .A1(n24865), .A2(n27789), .B1(n24847), .Y(
        n24850) );
  sky130_fd_sc_hd__nand2_1 U29968 ( .A(n27111), .B(n27785), .Y(n24848) );
  sky130_fd_sc_hd__o211ai_1 U29969 ( .A1(n11123), .A2(n27111), .B1(n26922), 
        .C1(n24848), .Y(n24849) );
  sky130_fd_sc_hd__nor2_1 U29970 ( .A(n27355), .B(n24852), .Y(n27361) );
  sky130_fd_sc_hd__nand2_1 U29971 ( .A(n24853), .B(n27361), .Y(n24857) );
  sky130_fd_sc_hd__nor2_1 U29972 ( .A(n24854), .B(n27355), .Y(n25889) );
  sky130_fd_sc_hd__nand2_1 U29973 ( .A(n24855), .B(n25889), .Y(n24856) );
  sky130_fd_sc_hd__nand2_1 U29974 ( .A(n24861), .B(n24832), .Y(n24858) );
  sky130_fd_sc_hd__o21ai_0 U29975 ( .A1(n24832), .A2(n28537), .B1(n24858), .Y(
        j202_soc_core_j22_cpu_rf_N3288) );
  sky130_fd_sc_hd__a22oi_1 U29976 ( .A1(n27862), .A2(n24862), .B1(n24859), 
        .B2(n27861), .Y(n24860) );
  sky130_fd_sc_hd__o22ai_1 U29978 ( .A1(n27841), .A2(n28537), .B1(n24712), 
        .B2(n12256), .Y(j202_soc_core_j22_cpu_rf_N3251) );
  sky130_fd_sc_hd__o22ai_1 U29979 ( .A1(n28532), .A2(n27850), .B1(n24863), 
        .B2(n27848), .Y(n24864) );
  sky130_fd_sc_hd__a21oi_1 U29980 ( .A1(n24865), .A2(n26068), .B1(n24864), .Y(
        n24866) );
  sky130_fd_sc_hd__o21ai_0 U29981 ( .A1(n27855), .A2(n28537), .B1(n24866), .Y(
        j202_soc_core_j22_cpu_rf_N314) );
  sky130_fd_sc_hd__o22ai_1 U29982 ( .A1(n27859), .A2(n28537), .B1(n27858), 
        .B2(n28060), .Y(j202_soc_core_j22_cpu_rf_N3327) );
  sky130_fd_sc_hd__o22ai_1 U29983 ( .A1(n25964), .A2(n28537), .B1(n27847), 
        .B2(n12256), .Y(j202_soc_core_j22_cpu_rf_N2696) );
  sky130_fd_sc_hd__nand2_1 U29985 ( .A(n27764), .B(n27042), .Y(n24867) );
  sky130_fd_sc_hd__o211ai_1 U29986 ( .A1(n27388), .A2(n27019), .B1(n24867), 
        .C1(n24292), .Y(j202_soc_core_j22_cpu_ml_N331) );
  sky130_fd_sc_hd__o21ai_1 U29987 ( .A1(n27021), .A2(n27770), .B1(n25374), .Y(
        j202_soc_core_j22_cpu_ml_maclj[27]) );
  sky130_fd_sc_hd__nand2_1 U29988 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[11]), .Y(n24868) );
  sky130_fd_sc_hd__o21ai_1 U29989 ( .A1(n26996), .A2(n28289), .B1(n24868), .Y(
        n125) );
  sky130_fd_sc_hd__nand2_1 U29990 ( .A(n24869), .B(n26916), .Y(n24870) );
  sky130_fd_sc_hd__nand2_1 U29991 ( .A(n25916), .B(n28478), .Y(n26292) );
  sky130_fd_sc_hd__nand2_1 U29992 ( .A(n26292), .B(n27806), .Y(n24891) );
  sky130_fd_sc_hd__nand3_1 U29993 ( .A(n24870), .B(n26919), .C(n24891), .Y(
        n24871) );
  sky130_fd_sc_hd__nand2_1 U29994 ( .A(n24871), .B(n25916), .Y(n24903) );
  sky130_fd_sc_hd__nand2_1 U29995 ( .A(n25916), .B(n27785), .Y(n24872) );
  sky130_fd_sc_hd__o211ai_1 U29996 ( .A1(n11123), .A2(n25916), .B1(n26922), 
        .C1(n24872), .Y(n24900) );
  sky130_fd_sc_hd__nand2_1 U29997 ( .A(n24873), .B(n27789), .Y(n24896) );
  sky130_fd_sc_hd__o22ai_1 U29998 ( .A1(n26926), .A2(n24874), .B1(n27793), 
        .B2(n28478), .Y(n24875) );
  sky130_fd_sc_hd__a21oi_1 U29999 ( .A1(n26003), .A2(n27032), .B1(n24875), .Y(
        n24878) );
  sky130_fd_sc_hd__o22a_1 U30000 ( .A1(n26926), .A2(n24876), .B1(n26939), .B2(
        n26292), .X(n24877) );
  sky130_fd_sc_hd__o211ai_1 U30001 ( .A1(n27798), .A2(n27803), .B1(n24878), 
        .C1(n24877), .Y(n24882) );
  sky130_fd_sc_hd__o22ai_1 U30003 ( .A1(n11144), .A2(n26936), .B1(n26276), 
        .B2(n26932), .Y(n24880) );
  sky130_fd_sc_hd__nor3_1 U30004 ( .A(n24882), .B(n24881), .C(n24880), .Y(
        n24895) );
  sky130_fd_sc_hd__o22ai_1 U30005 ( .A1(n26284), .A2(n27799), .B1(n26320), 
        .B2(n26943), .Y(n24886) );
  sky130_fd_sc_hd__o22ai_1 U30006 ( .A1(n26317), .A2(n27795), .B1(n27796), 
        .B2(n25996), .Y(n24885) );
  sky130_fd_sc_hd__nand2_1 U30007 ( .A(n24883), .B(n26426), .Y(n26933) );
  sky130_fd_sc_hd__nor3_1 U30008 ( .A(n24886), .B(n24885), .C(n24884), .Y(
        n24894) );
  sky130_fd_sc_hd__nand2_1 U30009 ( .A(n26332), .B(n24887), .Y(n24889) );
  sky130_fd_sc_hd__nand2_1 U30010 ( .A(n24889), .B(n24888), .Y(n24890) );
  sky130_fd_sc_hd__nand2_1 U30011 ( .A(n24890), .B(n26426), .Y(n26934) );
  sky130_fd_sc_hd__nand2_1 U30012 ( .A(n26934), .B(n24891), .Y(n24892) );
  sky130_fd_sc_hd__nand2_1 U30013 ( .A(n24892), .B(n28478), .Y(n24893) );
  sky130_fd_sc_hd__nand4_1 U30014 ( .A(n24896), .B(n24895), .C(n24894), .D(
        n24893), .Y(n24897) );
  sky130_fd_sc_hd__o21bai_1 U30015 ( .A1(n26926), .A2(n24898), .B1_N(n24897), 
        .Y(n24899) );
  sky130_fd_sc_hd__a21oi_1 U30016 ( .A1(n24901), .A2(n24900), .B1(n24899), .Y(
        n24902) );
  sky130_fd_sc_hd__nand2_1 U30017 ( .A(n24903), .B(n24902), .Y(n24907) );
  sky130_fd_sc_hd__o22ai_1 U30018 ( .A1(n28480), .A2(n25977), .B1(n28061), 
        .B2(n27162), .Y(j202_soc_core_j22_cpu_rf_N2873) );
  sky130_fd_sc_hd__o22ai_1 U30019 ( .A1(n28480), .A2(n25978), .B1(n27834), 
        .B2(n27162), .Y(j202_soc_core_j22_cpu_rf_N2947) );
  sky130_fd_sc_hd__o22ai_1 U30020 ( .A1(n28480), .A2(n25979), .B1(n28112), 
        .B2(n27162), .Y(j202_soc_core_j22_cpu_rf_N3206) );
  sky130_fd_sc_hd__o22ai_1 U30021 ( .A1(n28480), .A2(n25980), .B1(n27835), 
        .B2(n27162), .Y(j202_soc_core_j22_cpu_rf_N2799) );
  sky130_fd_sc_hd__o22ai_1 U30022 ( .A1(n28480), .A2(n25981), .B1(n27836), 
        .B2(n12225), .Y(j202_soc_core_j22_cpu_rf_N3169) );
  sky130_fd_sc_hd__o22ai_1 U30023 ( .A1(n28480), .A2(n25982), .B1(n27837), 
        .B2(n27162), .Y(j202_soc_core_j22_cpu_rf_N3021) );
  sky130_fd_sc_hd__o22ai_1 U30024 ( .A1(n28480), .A2(n26894), .B1(n27839), 
        .B2(n12225), .Y(j202_soc_core_j22_cpu_rf_N2910) );
  sky130_fd_sc_hd__o22ai_1 U30025 ( .A1(n28480), .A2(n25984), .B1(n27840), 
        .B2(n27162), .Y(j202_soc_core_j22_cpu_rf_N2725) );
  sky130_fd_sc_hd__o22ai_1 U30026 ( .A1(n28480), .A2(n27841), .B1(n24712), 
        .B2(n12225), .Y(j202_soc_core_j22_cpu_rf_N3243) );
  sky130_fd_sc_hd__o22ai_1 U30027 ( .A1(n28480), .A2(n25985), .B1(n27842), 
        .B2(n27162), .Y(j202_soc_core_j22_cpu_rf_N3095) );
  sky130_fd_sc_hd__o22ai_1 U30028 ( .A1(n28480), .A2(n25986), .B1(n27843), 
        .B2(n12225), .Y(j202_soc_core_j22_cpu_rf_N2984) );
  sky130_fd_sc_hd__o22ai_1 U30029 ( .A1(n28480), .A2(n25987), .B1(n27844), 
        .B2(n27162), .Y(j202_soc_core_j22_cpu_rf_N3132) );
  sky130_fd_sc_hd__o22ai_1 U30030 ( .A1(n28480), .A2(n25988), .B1(n27845), 
        .B2(n27162), .Y(j202_soc_core_j22_cpu_rf_N2836) );
  sky130_fd_sc_hd__o22ai_1 U30031 ( .A1(n28480), .A2(n25989), .B1(n27846), 
        .B2(n27162), .Y(j202_soc_core_j22_cpu_rf_N2762) );
  sky130_fd_sc_hd__o22ai_1 U30032 ( .A1(n28480), .A2(n25964), .B1(n27847), 
        .B2(n12225), .Y(j202_soc_core_j22_cpu_rf_N2688) );
  sky130_fd_sc_hd__o22ai_1 U30033 ( .A1(n28480), .A2(n27859), .B1(n27858), 
        .B2(n27162), .Y(j202_soc_core_j22_cpu_rf_N3319) );
  sky130_fd_sc_hd__mux2i_1 U30034 ( .A0(n27162), .A1(n28480), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3280) );
  sky130_fd_sc_hd__nor2_1 U30035 ( .A(n27644), .B(n12225), .Y(
        j202_soc_core_j22_cpu_rf_N2652) );
  sky130_fd_sc_hd__o22ai_1 U30036 ( .A1(n24905), .A2(n27775), .B1(n27774), 
        .B2(n28480), .Y(n24906) );
  sky130_fd_sc_hd__a21oi_1 U30037 ( .A1(n24907), .A2(n27860), .B1(n24906), .Y(
        n24908) );
  sky130_fd_sc_hd__nand2_1 U30039 ( .A(n26149), .B(n24910), .Y(n24914) );
  sky130_fd_sc_hd__a21oi_1 U30040 ( .A1(n24911), .A2(n24914), .B1(n24912), .Y(
        n24918) );
  sky130_fd_sc_hd__nor2_1 U30041 ( .A(n24914), .B(n24912), .Y(n24919) );
  sky130_fd_sc_hd__nand3_1 U30042 ( .A(n24919), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[0]), .C(n28431), .Y(n24917) );
  sky130_fd_sc_hd__inv_1 U30043 ( .A(n24913), .Y(n24915) );
  sky130_fd_sc_hd__nand4_1 U30044 ( .A(n24915), .B(n28109), .C(n26157), .D(
        n24914), .Y(n24916) );
  sky130_fd_sc_hd__o211ai_1 U30045 ( .A1(n28480), .A2(n24918), .B1(n24917), 
        .C1(n24916), .Y(j202_soc_core_j22_cpu_rf_N2640) );
  sky130_fd_sc_hd__nand2_1 U30046 ( .A(n26865), .B(n24920), .Y(
        j202_soc_core_j22_cpu_rf_N2639) );
  sky130_fd_sc_hd__a21oi_1 U30047 ( .A1(j202_soc_core_j22_cpu_ml_bufa[8]), 
        .A2(n28056), .B1(n24921), .Y(n24923) );
  sky130_fd_sc_hd__nand3_2 U30048 ( .A(n24924), .B(n24923), .C(n24922), .Y(
        n26973) );
  sky130_fd_sc_hd__o21ai_0 U30049 ( .A1(n11123), .A2(n26945), .B1(n26922), .Y(
        n24925) );
  sky130_fd_sc_hd__nand2_1 U30050 ( .A(n28483), .B(n24925), .Y(n24956) );
  sky130_fd_sc_hd__mux2i_1 U30051 ( .A0(n26934), .A1(n27793), .S(n24931), .Y(
        n24945) );
  sky130_fd_sc_hd__nand2_1 U30052 ( .A(n26935), .B(n27807), .Y(n24926) );
  sky130_fd_sc_hd__o211ai_1 U30053 ( .A1(n26265), .A2(n26936), .B1(n24926), 
        .C1(n26933), .Y(n24944) );
  sky130_fd_sc_hd__o22ai_1 U30054 ( .A1(n11188), .A2(n27799), .B1(n27616), 
        .B2(n27795), .Y(n24928) );
  sky130_fd_sc_hd__o22ai_1 U30055 ( .A1(n26322), .A2(n26943), .B1(n26944), 
        .B2(n27803), .Y(n24927) );
  sky130_fd_sc_hd__nor2_1 U30056 ( .A(n24928), .B(n24927), .Y(n24942) );
  sky130_fd_sc_hd__nand2_1 U30057 ( .A(n24930), .B(n24929), .Y(n24941) );
  sky130_fd_sc_hd__nand2b_1 U30058 ( .A_N(n24931), .B(n26945), .Y(n26308) );
  sky130_fd_sc_hd__o21a_1 U30059 ( .A1(n28484), .A2(n26945), .B1(n26308), .X(
        n26211) );
  sky130_fd_sc_hd__nor2_1 U30060 ( .A(n11116), .B(n26001), .Y(n24934) );
  sky130_fd_sc_hd__nand2_1 U30062 ( .A(n24935), .B(n27791), .Y(n24936) );
  sky130_fd_sc_hd__o211ai_1 U30063 ( .A1(n26317), .A2(n26919), .B1(n24937), 
        .C1(n24936), .Y(n24938) );
  sky130_fd_sc_hd__a21oi_1 U30064 ( .A1(n26211), .A2(n27806), .B1(n24938), .Y(
        n24940) );
  sky130_fd_sc_hd__a22oi_1 U30065 ( .A1(n27810), .A2(n26923), .B1(n27808), 
        .B2(n26378), .Y(n24939) );
  sky130_fd_sc_hd__nand4_1 U30066 ( .A(n24942), .B(n24941), .C(n24940), .D(
        n24939), .Y(n24943) );
  sky130_fd_sc_hd__nor3_1 U30067 ( .A(n24945), .B(n24944), .C(n24943), .Y(
        n24946) );
  sky130_fd_sc_hd__nand2_1 U30068 ( .A(n24953), .B(n24952), .Y(n24948) );
  sky130_fd_sc_hd__a21oi_2 U30072 ( .A1(n26973), .A2(n27152), .B1(n26978), .Y(
        n24957) );
  sky130_fd_sc_hd__o22ai_1 U30074 ( .A1(n26975), .A2(n26894), .B1(n27839), 
        .B2(n26972), .Y(j202_soc_core_j22_cpu_rf_N2909) );
  sky130_fd_sc_hd__o22ai_1 U30075 ( .A1(n26975), .A2(n25986), .B1(n27843), 
        .B2(n30071), .Y(j202_soc_core_j22_cpu_rf_N2983) );
  sky130_fd_sc_hd__o22ai_1 U30076 ( .A1(n26975), .A2(n25982), .B1(n27837), 
        .B2(n26972), .Y(j202_soc_core_j22_cpu_rf_N3020) );
  sky130_fd_sc_hd__o22ai_1 U30077 ( .A1(n26975), .A2(n25964), .B1(n27847), 
        .B2(n26972), .Y(j202_soc_core_j22_cpu_rf_N2687) );
  sky130_fd_sc_hd__o22ai_1 U30078 ( .A1(n26975), .A2(n25985), .B1(n27842), 
        .B2(n26972), .Y(j202_soc_core_j22_cpu_rf_N3094) );
  sky130_fd_sc_hd__nor2_1 U30079 ( .A(n27644), .B(n30071), .Y(
        j202_soc_core_j22_cpu_rf_N2651) );
  sky130_fd_sc_hd__o22ai_1 U30080 ( .A1(n26975), .A2(n25984), .B1(n27840), 
        .B2(n30071), .Y(j202_soc_core_j22_cpu_rf_N2724) );
  sky130_fd_sc_hd__o22ai_1 U30081 ( .A1(n26975), .A2(n27841), .B1(n24712), 
        .B2(n30071), .Y(j202_soc_core_j22_cpu_rf_N3242) );
  sky130_fd_sc_hd__nand2_1 U30082 ( .A(n25146), .B(n25901), .Y(n24967) );
  sky130_fd_sc_hd__nor2_1 U30083 ( .A(n24959), .B(n24958), .Y(n24963) );
  sky130_fd_sc_hd__o21ai_0 U30084 ( .A1(n28379), .A2(n28387), .B1(n24961), .Y(
        n24962) );
  sky130_fd_sc_hd__nor2_1 U30085 ( .A(n24963), .B(n24962), .Y(n24965) );
  sky130_fd_sc_hd__inv_1 U30086 ( .A(n25902), .Y(n24966) );
  sky130_fd_sc_hd__o211ai_1 U30087 ( .A1(n24968), .A2(n27990), .B1(n24967), 
        .C1(n24966), .Y(n10533) );
  sky130_fd_sc_hd__o22ai_1 U30088 ( .A1(n26975), .A2(n25980), .B1(n27835), 
        .B2(n30071), .Y(j202_soc_core_j22_cpu_rf_N2798) );
  sky130_fd_sc_hd__o22ai_1 U30089 ( .A1(n26975), .A2(n25983), .B1(n27838), 
        .B2(n30071), .Y(j202_soc_core_j22_cpu_rf_N3057) );
  sky130_fd_sc_hd__o22ai_1 U30090 ( .A1(n26975), .A2(n25979), .B1(n28112), 
        .B2(n30071), .Y(j202_soc_core_j22_cpu_rf_N3205) );
  sky130_fd_sc_hd__o22ai_1 U30091 ( .A1(n26975), .A2(n25981), .B1(n27836), 
        .B2(n30071), .Y(j202_soc_core_j22_cpu_rf_N3168) );
  sky130_fd_sc_hd__o22ai_1 U30092 ( .A1(n26975), .A2(n25987), .B1(n27844), 
        .B2(n30071), .Y(j202_soc_core_j22_cpu_rf_N3131) );
  sky130_fd_sc_hd__o22ai_1 U30093 ( .A1(n26975), .A2(n25989), .B1(n27846), 
        .B2(n30071), .Y(j202_soc_core_j22_cpu_rf_N2761) );
  sky130_fd_sc_hd__o22ai_1 U30094 ( .A1(n26975), .A2(n25988), .B1(n27845), 
        .B2(n30071), .Y(j202_soc_core_j22_cpu_rf_N2835) );
  sky130_fd_sc_hd__o22ai_1 U30095 ( .A1(n26975), .A2(n25978), .B1(n27834), 
        .B2(n30071), .Y(j202_soc_core_j22_cpu_rf_N2946) );
  sky130_fd_sc_hd__nand2_1 U30096 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[10]), .Y(n24969) );
  sky130_fd_sc_hd__o21ai_1 U30097 ( .A1(n24976), .A2(n28289), .B1(n24969), .Y(
        n124) );
  sky130_fd_sc_hd__nand2_1 U30098 ( .A(j202_soc_core_cmt_core_00_cnt1[7]), .B(
        j202_soc_core_cmt_core_00_cnt1[8]), .Y(n26984) );
  sky130_fd_sc_hd__nand4_1 U30099 ( .A(n24971), .B(n24972), .C(
        j202_soc_core_cmt_core_00_cnt1[9]), .D(
        j202_soc_core_cmt_core_00_cnt1[10]), .Y(n25166) );
  sky130_fd_sc_hd__nand2_1 U30100 ( .A(n25166), .B(n26990), .Y(n24970) );
  sky130_fd_sc_hd__nand2_1 U30101 ( .A(n24970), .B(n28583), .Y(n26992) );
  sky130_fd_sc_hd__nand2_1 U30102 ( .A(n24971), .B(n26990), .Y(n27548) );
  sky130_fd_sc_hd__a31oi_1 U30103 ( .A1(n26982), .A2(
        j202_soc_core_cmt_core_00_cnt1[9]), .A3(n24972), .B1(
        j202_soc_core_cmt_core_00_cnt1[10]), .Y(n24973) );
  sky130_fd_sc_hd__o22ai_1 U30104 ( .A1(n24976), .A2(n27530), .B1(n24974), 
        .B2(n24973), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[10])
         );
  sky130_fd_sc_hd__nand2_1 U30105 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[10]), .Y(n24975) );
  sky130_fd_sc_hd__o21ai_1 U30106 ( .A1(n24976), .A2(n28291), .B1(n24975), .Y(
        n130) );
  sky130_fd_sc_hd__nand2_1 U30107 ( .A(n27472), .B(
        j202_soc_core_cmt_core_00_cnt0[2]), .Y(n27476) );
  sky130_fd_sc_hd__nor2_1 U30108 ( .A(n24977), .B(n27476), .Y(n27479) );
  sky130_fd_sc_hd__nand3_1 U30109 ( .A(n27479), .B(
        j202_soc_core_cmt_core_00_cnt0[4]), .C(
        j202_soc_core_cmt_core_00_cnt0[5]), .Y(n27434) );
  sky130_fd_sc_hd__nor2_1 U30110 ( .A(n24978), .B(n27434), .Y(n25009) );
  sky130_fd_sc_hd__nor2_1 U30111 ( .A(n24979), .B(n27486), .Y(n27467) );
  sky130_fd_sc_hd__xnor2_1 U30112 ( .A(j202_soc_core_cmt_core_00_cnt0[15]), 
        .B(j202_soc_core_cmt_core_00_const0[15]), .Y(n24981) );
  sky130_fd_sc_hd__xnor2_1 U30113 ( .A(j202_soc_core_cmt_core_00_cnt0[5]), .B(
        j202_soc_core_cmt_core_00_const0[5]), .Y(n24980) );
  sky130_fd_sc_hd__nand2_1 U30114 ( .A(n24981), .B(n24980), .Y(n24998) );
  sky130_fd_sc_hd__xnor2_1 U30115 ( .A(j202_soc_core_cmt_core_00_const0[0]), 
        .B(j202_soc_core_cmt_core_00_cnt0[0]), .Y(n24983) );
  sky130_fd_sc_hd__xnor2_1 U30116 ( .A(j202_soc_core_cmt_core_00_cnt0[2]), .B(
        j202_soc_core_cmt_core_00_const0[2]), .Y(n24982) );
  sky130_fd_sc_hd__nand2_1 U30117 ( .A(n24983), .B(n24982), .Y(n24997) );
  sky130_fd_sc_hd__xnor2_1 U30118 ( .A(j202_soc_core_cmt_core_00_const0[10]), 
        .B(j202_soc_core_cmt_core_00_cnt0[10]), .Y(n24985) );
  sky130_fd_sc_hd__xnor2_1 U30119 ( .A(j202_soc_core_cmt_core_00_const0[1]), 
        .B(j202_soc_core_cmt_core_00_cnt0[1]), .Y(n24984) );
  sky130_fd_sc_hd__xnor2_1 U30120 ( .A(j202_soc_core_cmt_core_00_const0[9]), 
        .B(j202_soc_core_cmt_core_00_cnt0[9]), .Y(n24987) );
  sky130_fd_sc_hd__xnor2_1 U30121 ( .A(j202_soc_core_cmt_core_00_const0[11]), 
        .B(j202_soc_core_cmt_core_00_cnt0[11]), .Y(n24986) );
  sky130_fd_sc_hd__xnor2_1 U30122 ( .A(j202_soc_core_cmt_core_00_const0[3]), 
        .B(j202_soc_core_cmt_core_00_cnt0[3]), .Y(n24989) );
  sky130_fd_sc_hd__xnor2_1 U30123 ( .A(j202_soc_core_cmt_core_00_const0[8]), 
        .B(j202_soc_core_cmt_core_00_cnt0[8]), .Y(n24988) );
  sky130_fd_sc_hd__xnor2_1 U30124 ( .A(j202_soc_core_cmt_core_00_const0[7]), 
        .B(j202_soc_core_cmt_core_00_cnt0[7]), .Y(n24991) );
  sky130_fd_sc_hd__xnor2_1 U30125 ( .A(j202_soc_core_cmt_core_00_const0[12]), 
        .B(j202_soc_core_cmt_core_00_cnt0[12]), .Y(n24990) );
  sky130_fd_sc_hd__nand4_1 U30126 ( .A(n24995), .B(n24994), .C(n24993), .D(
        n24992), .Y(n24996) );
  sky130_fd_sc_hd__nor3_1 U30127 ( .A(n24998), .B(n24997), .C(n24996), .Y(
        n25004) );
  sky130_fd_sc_hd__xor2_1 U30128 ( .A(j202_soc_core_cmt_core_00_const0[13]), 
        .B(j202_soc_core_cmt_core_00_cnt0[13]), .X(n25000) );
  sky130_fd_sc_hd__xor2_1 U30129 ( .A(j202_soc_core_cmt_core_00_const0[6]), 
        .B(j202_soc_core_cmt_core_00_cnt0[6]), .X(n24999) );
  sky130_fd_sc_hd__nor2_1 U30130 ( .A(n25000), .B(n24999), .Y(n25003) );
  sky130_fd_sc_hd__xnor2_1 U30131 ( .A(j202_soc_core_cmt_core_00_const0[4]), 
        .B(j202_soc_core_cmt_core_00_cnt0[4]), .Y(n25002) );
  sky130_fd_sc_hd__xnor2_1 U30132 ( .A(j202_soc_core_cmt_core_00_const0[14]), 
        .B(j202_soc_core_cmt_core_00_cnt0[14]), .Y(n25001) );
  sky130_fd_sc_hd__nand4_1 U30133 ( .A(n25004), .B(n25003), .C(n25002), .D(
        n25001), .Y(n29168) );
  sky130_fd_sc_hd__nand2_1 U30134 ( .A(n27467), .B(n29168), .Y(n27484) );
  sky130_fd_sc_hd__nor2_1 U30135 ( .A(n27477), .B(n29169), .Y(n25013) );
  sky130_fd_sc_hd__nor3_1 U30137 ( .A(n27484), .B(
        j202_soc_core_cmt_core_00_cnt0[7]), .C(n25005), .Y(n25006) );
  sky130_fd_sc_hd__a21oi_1 U30138 ( .A1(n27486), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[7]), .B1(n25006), .Y(n25007) );
  sky130_fd_sc_hd__o21ai_1 U30139 ( .A1(n25008), .A2(n27438), .B1(n25007), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[7]) );
  sky130_fd_sc_hd__nand3_1 U30140 ( .A(n25009), .B(
        j202_soc_core_cmt_core_00_cnt0[7]), .C(
        j202_soc_core_cmt_core_00_cnt0[8]), .Y(n25015) );
  sky130_fd_sc_hd__a21oi_1 U30141 ( .A1(n25009), .A2(
        j202_soc_core_cmt_core_00_cnt0[7]), .B1(
        j202_soc_core_cmt_core_00_cnt0[8]), .Y(n25011) );
  sky130_fd_sc_hd__a22oi_1 U30142 ( .A1(n27486), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[8]), .B1(n29169), .B2(
        j202_soc_core_cmt_core_00_cnt0[8]), .Y(n25010) );
  sky130_fd_sc_hd__o31ai_1 U30143 ( .A1(n27484), .A2(n25012), .A3(n25011), 
        .B1(n25010), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[8])
         );
  sky130_fd_sc_hd__nor2_1 U30144 ( .A(n25014), .B(n25015), .Y(n25017) );
  sky130_fd_sc_hd__a21oi_1 U30145 ( .A1(n25017), .A2(n28564), .B1(n25013), .Y(
        n25171) );
  sky130_fd_sc_hd__a22o_1 U30147 ( .A1(n27486), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[9]), .B1(n25171), .B2(n25016), 
        .X(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[9]) );
  sky130_fd_sc_hd__nand2_1 U30148 ( .A(n25017), .B(n27477), .Y(n26104) );
  sky130_fd_sc_hd__a22oi_1 U30149 ( .A1(n27486), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[10]), .B1(n26095), .B2(n25019), 
        .Y(n25018) );
  sky130_fd_sc_hd__o21ai_1 U30150 ( .A1(n25019), .A2(n26097), .B1(n25018), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[10]) );
  sky130_fd_sc_hd__a22oi_1 U30151 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[10]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[10]), 
        .Y(n25021) );
  sky130_fd_sc_hd__a22oi_1 U30152 ( .A1(n28297), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[10]), 
        .B1(n28301), .B2(j202_soc_core_cmt_core_00_const0[10]), .Y(n25020) );
  sky130_fd_sc_hd__nand2_1 U30153 ( .A(n25021), .B(n25020), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[10]) );
  sky130_fd_sc_hd__nand2_1 U30154 ( .A(n25022), .B(n28385), .Y(n27915) );
  sky130_fd_sc_hd__nand2b_4 U30156 ( .A_N(n27915), .B(n25023), .Y(n27093) );
  sky130_fd_sc_hd__nand2_1 U30157 ( .A(n12466), .B(n28385), .Y(n28274) );
  sky130_fd_sc_hd__nand2_1 U30158 ( .A(n28274), .B(n25025), .Y(n25026) );
  sky130_fd_sc_hd__nand2_1 U30159 ( .A(n25026), .B(n12359), .Y(
        j202_soc_core_ahb2aqu_00_N128) );
  sky130_fd_sc_hd__nor2_1 U30160 ( .A(n29547), .B(n29546), .Y(n25028) );
  sky130_fd_sc_hd__nor3_1 U30161 ( .A(n29550), .B(n29549), .C(n29548), .Y(
        n25027) );
  sky130_fd_sc_hd__nor2_1 U30163 ( .A(n29552), .B(n27950), .Y(
        j202_soc_core_ahb2aqu_00_N97) );
  sky130_fd_sc_hd__nand2_1 U30164 ( .A(n12359), .B(n25031), .Y(
        j202_soc_core_ahb2aqu_00_N93) );
  sky130_fd_sc_hd__nor2_1 U30165 ( .A(n25034), .B(n25033), .Y(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_nxt_state_1_) );
  sky130_fd_sc_hd__nand2_1 U30166 ( .A(n25038), .B(
        j202_soc_core_ahb2apb_01_state[0]), .Y(n25041) );
  sky130_fd_sc_hd__nor3_1 U30167 ( .A(j202_soc_core_rst), .B(n25037), .C(
        n25041), .Y(j202_soc_core_ahb2apb_01_N91) );
  sky130_fd_sc_hd__nand2_1 U30168 ( .A(n25039), .B(n25038), .Y(n25040) );
  sky130_fd_sc_hd__nor3_1 U30169 ( .A(j202_soc_core_ahb2apb_01_state[1]), .B(
        n29088), .C(n25041), .Y(j202_soc_core_ahb2apb_01_N90) );
  sky130_fd_sc_hd__nand2_1 U30170 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[0]), 
        .B(j202_soc_core_ahb2apb_01_hsize_buf[1]), .Y(
        j202_soc_core_ahb2apb_01_N123) );
  sky130_fd_sc_hd__clkinv_1 U30171 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[0]), 
        .Y(n25044) );
  sky130_fd_sc_hd__nor2_1 U30172 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[1]), 
        .B(n25044), .Y(n25047) );
  sky130_fd_sc_hd__clkinv_1 U30173 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[1]), 
        .Y(n25042) );
  sky130_fd_sc_hd__nor2_1 U30174 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[0]), 
        .B(n25042), .Y(n25045) );
  sky130_fd_sc_hd__a21oi_1 U30175 ( .A1(j202_soc_core_intc_core_00_bs_addr[1]), 
        .A2(n25047), .B1(n25045), .Y(n25043) );
  sky130_fd_sc_hd__o31ai_1 U30176 ( .A1(j202_soc_core_intc_core_00_bs_addr[1]), 
        .A2(j202_soc_core_ahb2apb_01_hsize_buf[0]), .A3(n25050), .B1(n25043), 
        .Y(n10785) );
  sky130_fd_sc_hd__o21ai_0 U30177 ( .A1(j202_soc_core_ahb2apb_01_hsize_buf[0]), 
        .A2(n25066), .B1(n25043), .Y(n10786) );
  sky130_fd_sc_hd__nand2_1 U30178 ( .A(j202_soc_core_intc_core_00_bs_addr[1]), 
        .B(n25044), .Y(n25049) );
  sky130_fd_sc_hd__a21oi_1 U30179 ( .A1(n25047), .A2(n25046), .B1(n25045), .Y(
        n25048) );
  sky130_fd_sc_hd__o21ai_0 U30180 ( .A1(j202_soc_core_intc_core_00_bs_addr[0]), 
        .A2(n25049), .B1(n25048), .Y(n10784) );
  sky130_fd_sc_hd__o21ai_0 U30181 ( .A1(n25050), .A2(n25049), .B1(n25048), .Y(
        n10783) );
  sky130_fd_sc_hd__o22ai_1 U30182 ( .A1(n29156), .A2(n28064), .B1(n25059), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__nor2_1 U30183 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]), .B(n29072), .Y(n28065) );
  sky130_fd_sc_hd__nand4_1 U30184 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[1]), .B(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[6]), .C(j202_soc_core_intc_core_00_cp_intack_all_0_), .D(n29069), .Y(n26114) );
  sky130_fd_sc_hd__nor2_1 U30185 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .B(n26114), .Y(n26747) );
  sky130_fd_sc_hd__a21oi_1 U30186 ( .A1(n28065), .A2(n26747), .B1(
        j202_soc_core_intc_core_00_rg_irqc[10]), .Y(n25057) );
  sky130_fd_sc_hd__nor2_1 U30187 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[10]), 
        .B(n25055), .Y(n25056) );
  sky130_fd_sc_hd__a31oi_1 U30188 ( .A1(n25057), .A2(
        j202_soc_core_intc_core_00_in_intreq[10]), .A3(n29827), .B1(n25056), 
        .Y(n25058) );
  sky130_fd_sc_hd__nor2_1 U30189 ( .A(n25059), .B(n25058), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N13) );
  sky130_fd_sc_hd__o22ai_1 U30190 ( .A1(n29156), .A2(n28310), .B1(n25060), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__nor2_1 U30191 ( .A(j202_soc_core_intc_core_00_bs_addr[3]), 
        .B(n25061), .Y(n25068) );
  sky130_fd_sc_hd__nand3_1 U30192 ( .A(n25063), .B(n25073), .C(n25062), .Y(
        n25095) );
  sky130_fd_sc_hd__nor2_1 U30193 ( .A(n25064), .B(n25095), .Y(n26746) );
  sky130_fd_sc_hd__o22ai_1 U30194 ( .A1(n29156), .A2(n28313), .B1(n25065), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__nand2_1 U30195 ( .A(j202_soc_core_pwrite[1]), .B(
        j202_soc_core_intc_core_00_bs_addr[3]), .Y(n25079) );
  sky130_fd_sc_hd__nor2_1 U30196 ( .A(n25072), .B(n25066), .Y(n29398) );
  sky130_fd_sc_hd__nand2_1 U30197 ( .A(n25074), .B(n29398), .Y(n25097) );
  sky130_fd_sc_hd__o22ai_1 U30198 ( .A1(n29156), .A2(n28316), .B1(n25067), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__nand2_1 U30199 ( .A(n26760), .B(n29827), .Y(n26758) );
  sky130_fd_sc_hd__o22ai_1 U30200 ( .A1(n29156), .A2(n26760), .B1(n25070), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o22ai_1 U30201 ( .A1(n29156), .A2(n27575), .B1(n25071), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__nand3_1 U30202 ( .A(n25073), .B(
        j202_soc_core_intc_core_00_bs_addr[3]), .C(n25072), .Y(n25086) );
  sky130_fd_sc_hd__nand2_1 U30203 ( .A(n25074), .B(n29402), .Y(n28231) );
  sky130_fd_sc_hd__nand2_1 U30204 ( .A(n25075), .B(j202_soc_core_pwrite[1]), 
        .Y(n28553) );
  sky130_fd_sc_hd__nand2_1 U30205 ( .A(n28553), .B(n29745), .Y(n28551) );
  sky130_fd_sc_hd__o22ai_1 U30206 ( .A1(n29156), .A2(n28553), .B1(n25076), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__nor2_1 U30207 ( .A(n25086), .B(n25077), .Y(n27658) );
  sky130_fd_sc_hd__o22ai_1 U30208 ( .A1(n29156), .A2(n29082), .B1(n25078), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__nor2_1 U30209 ( .A(n25079), .B(n25095), .Y(n28235) );
  sky130_fd_sc_hd__o22ai_1 U30210 ( .A1(n29156), .A2(n29076), .B1(n25080), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__nand2_1 U30211 ( .A(n29828), .B(
        j202_soc_core_intc_core_00_bs_addr[3]), .Y(n25094) );
  sky130_fd_sc_hd__nor4_1 U30212 ( .A(n29088), .B(
        j202_soc_core_intc_core_00_bs_addr[7]), .C(
        j202_soc_core_intc_core_00_bs_addr[6]), .D(n25081), .Y(n28318) );
  sky130_fd_sc_hd__nand3_1 U30213 ( .A(n25082), .B(
        j202_soc_core_intc_core_00_bs_addr[6]), .C(n29745), .Y(n25083) );
  sky130_fd_sc_hd__a22oi_1 U30214 ( .A1(n28318), .A2(
        j202_soc_core_intc_core_00_rg_ie[10]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[10]), .Y(n25092) );
  sky130_fd_sc_hd__nand2_1 U30215 ( .A(n29828), .B(
        j202_soc_core_intc_core_00_bs_addr[8]), .Y(n25089) );
  sky130_fd_sc_hd__nand2b_1 U30216 ( .A_N(n25086), .B(n25085), .Y(n25087) );
  sky130_fd_sc_hd__nor2_1 U30217 ( .A(n25087), .B(n25088), .Y(n28322) );
  sky130_fd_sc_hd__nor3_1 U30218 ( .A(n25090), .B(n25089), .C(n25088), .Y(
        n27398) );
  sky130_fd_sc_hd__a22oi_1 U30219 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[82]), .B1(n27398), .B2(
        j202_soc_core_intc_core_00_rg_itgt[66]), .Y(n25091) );
  sky130_fd_sc_hd__nand3_1 U30220 ( .A(n25092), .B(n28238), .C(n25091), .Y(
        n25093) );
  sky130_fd_sc_hd__a21oi_1 U30221 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[106]), .B1(n25093), .Y(n25102) );
  sky130_fd_sc_hd__nand2_1 U30222 ( .A(n29403), .B(n29828), .Y(n25098) );
  sky130_fd_sc_hd__a22oi_1 U30223 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[90]), .B1(n28331), .B2(
        j202_soc_core_intc_core_00_rg_itgt[74]), .Y(n25101) );
  sky130_fd_sc_hd__a22oi_1 U30224 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[10]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[42]), .B2(n28330), .Y(n25100) );
  sky130_fd_sc_hd__nand2_1 U30225 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[74]), .Y(n25099) );
  sky130_fd_sc_hd__nand4_1 U30226 ( .A(n25102), .B(n25101), .C(n25100), .D(
        n25099), .Y(j202_soc_core_ahb2apb_01_N138) );
  sky130_fd_sc_hd__nand2b_1 U30227 ( .A_N(n12279), .B(n12366), .Y(n25103) );
  sky130_fd_sc_hd__nand2_1 U30228 ( .A(n27764), .B(n26330), .Y(n25104) );
  sky130_fd_sc_hd__o211ai_1 U30229 ( .A1(n27388), .A2(n28448), .B1(n25104), 
        .C1(n24292), .Y(j202_soc_core_j22_cpu_ml_N334) );
  sky130_fd_sc_hd__a21oi_1 U30230 ( .A1(n12425), .A2(n28056), .B1(n25776), .Y(
        n25105) );
  sky130_fd_sc_hd__o21ai_1 U30231 ( .A1(n25106), .A2(n25779), .B1(n25105), .Y(
        n29835) );
  sky130_fd_sc_hd__nand2_1 U30232 ( .A(n11114), .B(n25682), .Y(n25126) );
  sky130_fd_sc_hd__nand2_1 U30233 ( .A(n26330), .B(n25263), .Y(n25107) );
  sky130_fd_sc_hd__a22o_1 U30234 ( .A1(n27785), .A2(n26330), .B1(n25107), .B2(
        n27786), .X(n25108) );
  sky130_fd_sc_hd__nand2_1 U30235 ( .A(n11114), .B(n25108), .Y(n25125) );
  sky130_fd_sc_hd__o22a_1 U30236 ( .A1(n26275), .A2(n27817), .B1(n25973), .B2(
        n27815), .X(n25122) );
  sky130_fd_sc_hd__nand2_1 U30237 ( .A(n28446), .B(n27791), .Y(n25110) );
  sky130_fd_sc_hd__nand2_1 U30238 ( .A(n25110), .B(n25266), .Y(n25115) );
  sky130_fd_sc_hd__a2bb2oi_1 U30239 ( .B1(n25868), .B2(n25112), .A1_N(n26926), 
        .A2_N(n25111), .Y(n25113) );
  sky130_fd_sc_hd__o21ai_1 U30240 ( .A1(n27793), .A2(n28446), .B1(n25113), .Y(
        n25114) );
  sky130_fd_sc_hd__a21oi_1 U30241 ( .A1(n26330), .A2(n25115), .B1(n25114), .Y(
        n25116) );
  sky130_fd_sc_hd__o21ai_1 U30242 ( .A1(n26324), .A2(n27799), .B1(n25116), .Y(
        n25117) );
  sky130_fd_sc_hd__a21oi_1 U30243 ( .A1(n27808), .A2(n27809), .B1(n25117), .Y(
        n25121) );
  sky130_fd_sc_hd__o22ai_1 U30244 ( .A1(n26296), .A2(n27795), .B1(n28429), 
        .B2(n27803), .Y(n25119) );
  sky130_fd_sc_hd__xnor2_1 U30245 ( .A(n28446), .B(n26330), .Y(n26235) );
  sky130_fd_sc_hd__o22ai_1 U30246 ( .A1(n26319), .A2(n27797), .B1(n25872), 
        .B2(n26235), .Y(n25118) );
  sky130_fd_sc_hd__nor2_1 U30247 ( .A(n25119), .B(n25118), .Y(n25120) );
  sky130_fd_sc_hd__nand4_1 U30248 ( .A(n25122), .B(n25121), .C(n25120), .D(
        n27814), .Y(n25123) );
  sky130_fd_sc_hd__a21oi_1 U30249 ( .A1(n25141), .A2(n27789), .B1(n25123), .Y(
        n25124) );
  sky130_fd_sc_hd__nand2_1 U30250 ( .A(n25129), .B(n25868), .Y(n25130) );
  sky130_fd_sc_hd__nand2_1 U30251 ( .A(n25135), .B(n24832), .Y(n25134) );
  sky130_fd_sc_hd__o21ai_0 U30252 ( .A1(n24832), .A2(n28448), .B1(n25134), .Y(
        j202_soc_core_j22_cpu_rf_N3304) );
  sky130_fd_sc_hd__o22ai_1 U30253 ( .A1(n27859), .A2(n28448), .B1(n27858), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N3342) );
  sky130_fd_sc_hd__o22ai_1 U30254 ( .A1(n27841), .A2(n28448), .B1(n24712), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N3267) );
  sky130_fd_sc_hd__o22ai_1 U30255 ( .A1(n25964), .A2(n28448), .B1(n27847), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N2712) );
  sky130_fd_sc_hd__nand2_1 U30256 ( .A(n25135), .B(n27860), .Y(n25137) );
  sky130_fd_sc_hd__nand2_1 U30257 ( .A(n25137), .B(n25136), .Y(
        j202_soc_core_j22_cpu_rf_N3378) );
  sky130_fd_sc_hd__o22ai_1 U30258 ( .A1(n26275), .A2(n27850), .B1(n25139), 
        .B2(n27848), .Y(n25140) );
  sky130_fd_sc_hd__a21oi_1 U30259 ( .A1(n25141), .A2(n26068), .B1(n25140), .Y(
        n25142) );
  sky130_fd_sc_hd__o21ai_0 U30260 ( .A1(n27855), .A2(n28448), .B1(n25142), .Y(
        j202_soc_core_j22_cpu_rf_N328) );
  sky130_fd_sc_hd__o22ai_1 U30261 ( .A1(n25978), .A2(n28448), .B1(n27834), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N2971) );
  sky130_fd_sc_hd__o22ai_1 U30262 ( .A1(n25979), .A2(n28448), .B1(n28112), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N3230) );
  sky130_fd_sc_hd__o22ai_1 U30263 ( .A1(n25980), .A2(n28448), .B1(n27835), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N2823) );
  sky130_fd_sc_hd__o22ai_1 U30264 ( .A1(n25981), .A2(n28448), .B1(n27836), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N3193) );
  sky130_fd_sc_hd__o22ai_1 U30265 ( .A1(n25982), .A2(n28448), .B1(n27837), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N3045) );
  sky130_fd_sc_hd__o22ai_1 U30266 ( .A1(n25983), .A2(n28448), .B1(n27838), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N3082) );
  sky130_fd_sc_hd__o22ai_1 U30267 ( .A1(n26894), .A2(n28448), .B1(n27839), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N2934) );
  sky130_fd_sc_hd__o22ai_1 U30268 ( .A1(n25984), .A2(n28448), .B1(n27840), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N2749) );
  sky130_fd_sc_hd__o22ai_1 U30269 ( .A1(n25985), .A2(n28448), .B1(n27842), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N3119) );
  sky130_fd_sc_hd__o22ai_1 U30270 ( .A1(n25986), .A2(n28448), .B1(n27843), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N3008) );
  sky130_fd_sc_hd__o22ai_1 U30271 ( .A1(n25987), .A2(n28448), .B1(n27844), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N3156) );
  sky130_fd_sc_hd__o22ai_1 U30272 ( .A1(n25988), .A2(n28448), .B1(n27845), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N2860) );
  sky130_fd_sc_hd__o22ai_1 U30273 ( .A1(n25989), .A2(n28448), .B1(n27846), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N2786) );
  sky130_fd_sc_hd__a21oi_1 U30274 ( .A1(n27768), .A2(n12425), .B1(n27766), .Y(
        n25143) );
  sky130_fd_sc_hd__o22ai_1 U30276 ( .A1(n27461), .A2(n27859), .B1(n27858), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N3316) );
  sky130_fd_sc_hd__mux2i_1 U30277 ( .A0(n12471), .A1(n27461), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3276) );
  sky130_fd_sc_hd__a22oi_1 U30278 ( .A1(n25146), .A2(n29560), .B1(n29559), 
        .B2(n24133), .Y(n25151) );
  sky130_fd_sc_hd__o211ai_1 U30279 ( .A1(n25151), .A2(n28379), .B1(n25150), 
        .C1(n12061), .Y(n10535) );
  sky130_fd_sc_hd__nor2_1 U30280 ( .A(n27644), .B(n12471), .Y(
        j202_soc_core_j22_cpu_rf_N2648) );
  sky130_fd_sc_hd__o22ai_1 U30281 ( .A1(n27461), .A2(n27841), .B1(n24712), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N3239) );
  sky130_fd_sc_hd__o22ai_1 U30282 ( .A1(n27461), .A2(n25964), .B1(n27847), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N2684) );
  sky130_fd_sc_hd__a22oi_1 U30283 ( .A1(n25152), .A2(n27862), .B1(n12402), 
        .B2(n27861), .Y(n25153) );
  sky130_fd_sc_hd__o21ai_0 U30284 ( .A1(n27648), .A2(n12471), .B1(n25153), .Y(
        j202_soc_core_j22_cpu_rf_N3351) );
  sky130_fd_sc_hd__o22ai_1 U30285 ( .A1(n29158), .A2(n27575), .B1(n25154), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U30286 ( .A1(n29144), .A2(n27575), .B1(n25155), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U30287 ( .A1(n29162), .A2(n28064), .B1(n25160), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__a21oi_1 U30288 ( .A1(n26747), .A2(n27350), .B1(
        j202_soc_core_intc_core_00_rg_irqc[2]), .Y(n25158) );
  sky130_fd_sc_hd__nor2_1 U30289 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[2]), 
        .B(n25156), .Y(n25157) );
  sky130_fd_sc_hd__a31oi_1 U30290 ( .A1(n25158), .A2(
        j202_soc_core_intc_core_00_in_intreq[2]), .A3(n29830), .B1(n25157), 
        .Y(n25159) );
  sky130_fd_sc_hd__nor2_1 U30291 ( .A(n25160), .B(n25159), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N5) );
  sky130_fd_sc_hd__nor2_1 U30292 ( .A(j202_soc_core_rst), .B(
        j202_soc_core_qspi_wb_wdat[8]), .Y(n28959) );
  sky130_fd_sc_hd__o22ai_1 U30293 ( .A1(n26704), .A2(n25161), .B1(n28959), 
        .B2(n26702), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U30294 ( .A1(n29145), .A2(n27575), .B1(n25162), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U30295 ( .A1(n29148), .A2(n27575), .B1(n25163), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U30296 ( .A1(n29146), .A2(n27575), .B1(n25164), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__nand2_1 U30297 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[12]), .Y(n25165) );
  sky130_fd_sc_hd__o21ai_1 U30298 ( .A1(n25170), .A2(n28289), .B1(n25165), .Y(
        n121) );
  sky130_fd_sc_hd__a31oi_1 U30299 ( .A1(n26991), .A2(
        j202_soc_core_cmt_core_00_cnt1[11]), .A3(n26990), .B1(
        j202_soc_core_cmt_core_00_cnt1[12]), .Y(n25168) );
  sky130_fd_sc_hd__a21oi_1 U30300 ( .A1(j202_soc_core_cmt_core_00_cnt1[12]), 
        .A2(j202_soc_core_cmt_core_00_cnt1[11]), .B1(n27540), .Y(n25167) );
  sky130_fd_sc_hd__nor2_1 U30301 ( .A(n25167), .B(n26992), .Y(n26082) );
  sky130_fd_sc_hd__o22ai_1 U30302 ( .A1(n25170), .A2(n27530), .B1(n25168), 
        .B2(n26082), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[12])
         );
  sky130_fd_sc_hd__nand2_1 U30303 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[12]), .Y(n25169) );
  sky130_fd_sc_hd__o21ai_1 U30304 ( .A1(n25170), .A2(n28291), .B1(n25169), .Y(
        n120) );
  sky130_fd_sc_hd__a21oi_1 U30305 ( .A1(n26095), .A2(
        j202_soc_core_cmt_core_00_cnt0[10]), .B1(
        j202_soc_core_cmt_core_00_cnt0[11]), .Y(n25172) );
  sky130_fd_sc_hd__nand2_1 U30306 ( .A(j202_soc_core_cmt_core_00_cnt0[10]), 
        .B(j202_soc_core_cmt_core_00_cnt0[11]), .Y(n26094) );
  sky130_fd_sc_hd__a21oi_1 U30307 ( .A1(n27477), .A2(n26094), .B1(n25171), .Y(
        n25175) );
  sky130_fd_sc_hd__o22ai_1 U30308 ( .A1(n27482), .A2(n26996), .B1(n25172), 
        .B2(n25175), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[11])
         );
  sky130_fd_sc_hd__nor3_1 U30309 ( .A(j202_soc_core_cmt_core_00_cnt0[12]), .B(
        n26094), .C(n26104), .Y(n25173) );
  sky130_fd_sc_hd__a21oi_1 U30310 ( .A1(n27486), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[12]), .B1(n25173), .Y(n25174) );
  sky130_fd_sc_hd__o21ai_1 U30311 ( .A1(n25176), .A2(n25175), .B1(n25174), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[12]) );
  sky130_fd_sc_hd__a22oi_1 U30312 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[12]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[12]), 
        .Y(n25178) );
  sky130_fd_sc_hd__a22oi_1 U30313 ( .A1(n28297), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[12]), 
        .B1(n28301), .B2(j202_soc_core_cmt_core_00_const0[12]), .Y(n25177) );
  sky130_fd_sc_hd__nand2_1 U30314 ( .A(n25178), .B(n25177), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[12]) );
  sky130_fd_sc_hd__nand2_1 U30315 ( .A(n28201), .B(n25179), .Y(n25180) );
  sky130_fd_sc_hd__nand2_1 U30316 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[12]), .Y(n25181) );
  sky130_fd_sc_hd__o21ai_1 U30317 ( .A1(n25182), .A2(n28545), .B1(n25181), .Y(
        n58) );
  sky130_fd_sc_hd__o22ai_1 U30318 ( .A1(n29147), .A2(n28064), .B1(n25187), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__nor2_1 U30319 ( .A(n26674), .B(n29072), .Y(n26748) );
  sky130_fd_sc_hd__a21oi_1 U30320 ( .A1(n26748), .A2(n26719), .B1(
        j202_soc_core_intc_core_00_rg_irqc[12]), .Y(n25185) );
  sky130_fd_sc_hd__nor2_1 U30321 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[12]), 
        .B(n25183), .Y(n25184) );
  sky130_fd_sc_hd__a31oi_1 U30322 ( .A1(n25185), .A2(
        j202_soc_core_intc_core_00_in_intreq[12]), .A3(n29745), .B1(n25184), 
        .Y(n25186) );
  sky130_fd_sc_hd__nor2_1 U30323 ( .A(n25187), .B(n25186), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N15) );
  sky130_fd_sc_hd__nor2_1 U30324 ( .A(n29088), .B(
        j202_soc_core_qspi_wb_wdat[12]), .Y(n28984) );
  sky130_fd_sc_hd__o22ai_1 U30325 ( .A1(n26704), .A2(n25188), .B1(n28984), 
        .B2(n26702), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U30326 ( .A1(n26746), .A2(n25189), .B1(n28984), 
        .B2(n26744), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U30327 ( .A1(n29147), .A2(n28316), .B1(n25190), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U30328 ( .A1(n29147), .A2(n26760), .B1(n25191), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U30329 ( .A1(n29147), .A2(n28553), .B1(n25192), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U30330 ( .A1(n27658), .A2(n25193), .B1(n28984), 
        .B2(n27656), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U30331 ( .A1(n28235), .A2(n25194), .B1(n28984), 
        .B2(n28233), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__clkbuf_1 U30332 ( .A(n28318), .X(n28236) );
  sky130_fd_sc_hd__a22oi_1 U30333 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[12]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[12]), .Y(n25196) );
  sky130_fd_sc_hd__a22oi_1 U30334 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[19]), .B1(n27398), .B2(
        j202_soc_core_intc_core_00_rg_itgt[3]), .Y(n25195) );
  sky130_fd_sc_hd__nand3_1 U30335 ( .A(n25196), .B(n28238), .C(n25195), .Y(
        n25197) );
  sky130_fd_sc_hd__a21oi_1 U30336 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[108]), .B1(n25197), .Y(n25201) );
  sky130_fd_sc_hd__a22oi_1 U30337 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[27]), .B1(
        j202_soc_core_intc_core_00_rg_itgt[11]), .B2(n28331), .Y(n25200) );
  sky130_fd_sc_hd__a22oi_1 U30338 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[12]), .B1(n28330), .B2(
        j202_soc_core_intc_core_00_rg_ipr[44]), .Y(n25199) );
  sky130_fd_sc_hd__nand2_1 U30339 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[76]), .Y(n25198) );
  sky130_fd_sc_hd__nand4_1 U30340 ( .A(n25201), .B(n25200), .C(n25199), .D(
        n25198), .Y(j202_soc_core_ahb2apb_01_N140) );
  sky130_fd_sc_hd__nand2_1 U30341 ( .A(n25203), .B(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .Y(n26571) );
  sky130_fd_sc_hd__nand2_1 U30342 ( .A(n26571), .B(n29828), .Y(n26464) );
  sky130_fd_sc_hd__nand3_1 U30343 ( .A(n25204), .B(n26463), .C(n26567), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N312) );
  sky130_fd_sc_hd__o22ai_1 U30344 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(io_in[11]), .B1(
        n28896), .B2(io_in[10]), .Y(n25338) );
  sky130_fd_sc_hd__nor2_1 U30345 ( .A(n28898), .B(n25338), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N358) );
  sky130_fd_sc_hd__nor2_1 U30346 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(n27264), .Y(n26564) );
  sky130_fd_sc_hd__nand2_1 U30347 ( .A(n26564), .B(n27287), .Y(n28685) );
  sky130_fd_sc_hd__nand2_1 U30348 ( .A(n26516), .B(n28685), .Y(n26574) );
  sky130_fd_sc_hd__nand2_1 U30349 ( .A(n26574), .B(
        j202_soc_core_wbqspiflash_00_spi_out[0]), .Y(n25208) );
  sky130_fd_sc_hd__nor2_1 U30350 ( .A(n27264), .B(n27254), .Y(n26594) );
  sky130_fd_sc_hd__a21oi_1 U30351 ( .A1(n25206), .A2(
        j202_soc_core_wbqspiflash_00_state[4]), .B1(n26594), .Y(n25207) );
  sky130_fd_sc_hd__a21oi_1 U30352 ( .A1(n25208), .A2(n25207), .B1(n29088), .Y(
        j202_soc_core_wbqspiflash_00_N709) );
  sky130_fd_sc_hd__o22ai_1 U30353 ( .A1(n26894), .A2(n26456), .B1(n27839), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N2927) );
  sky130_fd_sc_hd__o22ai_1 U30354 ( .A1(n25980), .A2(n26456), .B1(n27835), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N2816) );
  sky130_fd_sc_hd__o22ai_1 U30355 ( .A1(n25986), .A2(n26456), .B1(n27843), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N3001) );
  sky130_fd_sc_hd__o22ai_1 U30356 ( .A1(n25982), .A2(n26456), .B1(n27837), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N3038) );
  sky130_fd_sc_hd__o22ai_1 U30357 ( .A1(n25985), .A2(n26456), .B1(n27842), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N3112) );
  sky130_fd_sc_hd__o22ai_1 U30358 ( .A1(n25987), .A2(n26456), .B1(n27844), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N3149) );
  sky130_fd_sc_hd__o22ai_1 U30359 ( .A1(n25984), .A2(n26456), .B1(n27840), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N2742) );
  sky130_fd_sc_hd__o22ai_1 U30360 ( .A1(n25978), .A2(n26456), .B1(n27834), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N2964) );
  sky130_fd_sc_hd__o22ai_1 U30361 ( .A1(n25983), .A2(n26456), .B1(n27838), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N3075) );
  sky130_fd_sc_hd__o22ai_1 U30362 ( .A1(n25977), .A2(n26456), .B1(n28061), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N2890) );
  sky130_fd_sc_hd__o22ai_1 U30363 ( .A1(n25979), .A2(n26456), .B1(n28112), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N3223) );
  sky130_fd_sc_hd__o22ai_1 U30364 ( .A1(n25981), .A2(n26456), .B1(n27836), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N3186) );
  sky130_fd_sc_hd__o22ai_1 U30365 ( .A1(n25964), .A2(n26456), .B1(n27847), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N2705) );
  sky130_fd_sc_hd__o22ai_1 U30366 ( .A1(n25989), .A2(n26456), .B1(n27846), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N2779) );
  sky130_fd_sc_hd__o22ai_1 U30367 ( .A1(n25988), .A2(n26456), .B1(n27845), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N2853) );
  sky130_fd_sc_hd__o22ai_1 U30368 ( .A1(n27841), .A2(n26456), .B1(n24712), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N3260) );
  sky130_fd_sc_hd__nand2_1 U30369 ( .A(n27764), .B(n27807), .Y(n25210) );
  sky130_fd_sc_hd__o211ai_1 U30370 ( .A1(n26456), .A2(n27388), .B1(n25210), 
        .C1(n24292), .Y(j202_soc_core_j22_cpu_ml_N328) );
  sky130_fd_sc_hd__a21oi_1 U30371 ( .A1(n27768), .A2(
        j202_soc_core_j22_cpu_ml_bufa[24]), .B1(n27766), .Y(n25212) );
  sky130_fd_sc_hd__o21ai_1 U30372 ( .A1(n25213), .A2(n27770), .B1(n25212), .Y(
        j202_soc_core_j22_cpu_ml_maclj[24]) );
  sky130_fd_sc_hd__nor2_1 U30373 ( .A(n25214), .B(n12279), .Y(n25240) );
  sky130_fd_sc_hd__nand2_1 U30374 ( .A(n27764), .B(n25271), .Y(n25215) );
  sky130_fd_sc_hd__o211ai_1 U30375 ( .A1(n25245), .A2(n27388), .B1(n25215), 
        .C1(n24292), .Y(j202_soc_core_j22_cpu_ml_N327) );
  sky130_fd_sc_hd__nand4_1 U30376 ( .A(n25222), .B(n25220), .C(n25219), .D(
        n25218), .Y(n25216) );
  sky130_fd_sc_hd__nand2_1 U30377 ( .A(n26077), .B(n25216), .Y(n25217) );
  sky130_fd_sc_hd__nand2_1 U30378 ( .A(n25217), .B(n27119), .Y(
        j202_soc_core_j22_cpu_ml_machj[23]) );
  sky130_fd_sc_hd__o21ai_1 U30379 ( .A1(n25224), .A2(n27770), .B1(n25374), .Y(
        j202_soc_core_j22_cpu_ml_maclj[23]) );
  sky130_fd_sc_hd__nand4_1 U30380 ( .A(n25220), .B(n27828), .C(n25219), .D(
        n25218), .Y(n25221) );
  sky130_fd_sc_hd__a21oi_1 U30381 ( .A1(n25224), .A2(n27052), .B1(n26926), .Y(
        n25225) );
  sky130_fd_sc_hd__nand3_1 U30382 ( .A(n25240), .B(n27786), .C(n25271), .Y(
        n25226) );
  sky130_fd_sc_hd__o21a_1 U30383 ( .A1(n25240), .A2(n27787), .B1(n25226), .X(
        n25243) );
  sky130_fd_sc_hd__nand2_1 U30384 ( .A(n25271), .B(n27785), .Y(n25227) );
  sky130_fd_sc_hd__o21a_1 U30385 ( .A1(n26411), .A2(n25271), .B1(n25227), .X(
        n25241) );
  sky130_fd_sc_hd__o22ai_1 U30386 ( .A1(n26430), .A2(n27799), .B1(n28429), 
        .B2(n26943), .Y(n25235) );
  sky130_fd_sc_hd__o22ai_1 U30387 ( .A1(n26324), .A2(n27795), .B1(n27616), 
        .B2(n27797), .Y(n25234) );
  sky130_fd_sc_hd__a21oi_1 U30388 ( .A1(n25230), .A2(n27791), .B1(n27790), .Y(
        n25228) );
  sky130_fd_sc_hd__o22ai_1 U30389 ( .A1(n27793), .A2(n25230), .B1(n26431), 
        .B2(n25228), .Y(n25229) );
  sky130_fd_sc_hd__a21oi_1 U30390 ( .A1(n26942), .A2(n27807), .B1(n25229), .Y(
        n25232) );
  sky130_fd_sc_hd__xor2_1 U30391 ( .A(n25230), .B(n25271), .X(n26228) );
  sky130_fd_sc_hd__a22oi_1 U30392 ( .A1(n26228), .A2(n27806), .B1(n27808), 
        .B2(n26329), .Y(n25231) );
  sky130_fd_sc_hd__o211ai_1 U30393 ( .A1(n27796), .A2(n25688), .B1(n25232), 
        .C1(n25231), .Y(n25233) );
  sky130_fd_sc_hd__nor3_1 U30394 ( .A(n25235), .B(n25234), .C(n25233), .Y(
        n25237) );
  sky130_fd_sc_hd__o22a_1 U30395 ( .A1(n28487), .A2(n27817), .B1(n26309), .B2(
        n27815), .X(n25236) );
  sky130_fd_sc_hd__nand3_1 U30396 ( .A(n25237), .B(n25236), .C(n27814), .Y(
        n25238) );
  sky130_fd_sc_hd__a21oi_1 U30397 ( .A1(n25252), .A2(n27789), .B1(n25238), .Y(
        n25239) );
  sky130_fd_sc_hd__o21a_1 U30398 ( .A1(n25241), .A2(n25240), .B1(n25239), .X(
        n25242) );
  sky130_fd_sc_hd__nand2_1 U30399 ( .A(n25246), .B(n24832), .Y(n25244) );
  sky130_fd_sc_hd__o21ai_0 U30400 ( .A1(n24832), .A2(n25245), .B1(n25244), .Y(
        j202_soc_core_j22_cpu_rf_N3296) );
  sky130_fd_sc_hd__o22ai_1 U30401 ( .A1(n25245), .A2(n27859), .B1(n27858), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N3335) );
  sky130_fd_sc_hd__o22ai_1 U30402 ( .A1(n27841), .A2(n25245), .B1(n24712), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N3259) );
  sky130_fd_sc_hd__o22ai_1 U30403 ( .A1(n25964), .A2(n25245), .B1(n27847), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N2704) );
  sky130_fd_sc_hd__nand2_1 U30404 ( .A(n25246), .B(n27860), .Y(n25249) );
  sky130_fd_sc_hd__o22a_1 U30405 ( .A1(n25250), .A2(n27775), .B1(n27774), .B2(
        n25245), .X(n25248) );
  sky130_fd_sc_hd__nand2_1 U30406 ( .A(n25249), .B(n25248), .Y(
        j202_soc_core_j22_cpu_rf_N3370) );
  sky130_fd_sc_hd__o22ai_1 U30407 ( .A1(n28487), .A2(n27850), .B1(n25250), 
        .B2(n27848), .Y(n25251) );
  sky130_fd_sc_hd__a21oi_1 U30408 ( .A1(n25252), .A2(n26068), .B1(n25251), .Y(
        n25253) );
  sky130_fd_sc_hd__o21ai_0 U30409 ( .A1(n27855), .A2(n25245), .B1(n25253), .Y(
        j202_soc_core_j22_cpu_rf_N321) );
  sky130_fd_sc_hd__o22ai_1 U30410 ( .A1(n25977), .A2(n25245), .B1(n28061), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N2889) );
  sky130_fd_sc_hd__o22ai_1 U30411 ( .A1(n25978), .A2(n25245), .B1(n27834), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N2963) );
  sky130_fd_sc_hd__o22ai_1 U30412 ( .A1(n25979), .A2(n25245), .B1(n28112), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N3222) );
  sky130_fd_sc_hd__o22ai_1 U30413 ( .A1(n25980), .A2(n25245), .B1(n27835), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N2815) );
  sky130_fd_sc_hd__o22ai_1 U30414 ( .A1(n25981), .A2(n25245), .B1(n27836), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N3185) );
  sky130_fd_sc_hd__o22ai_1 U30415 ( .A1(n25982), .A2(n25245), .B1(n27837), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N3037) );
  sky130_fd_sc_hd__o22ai_1 U30416 ( .A1(n26894), .A2(n25245), .B1(n27839), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N2926) );
  sky130_fd_sc_hd__o22ai_1 U30417 ( .A1(n25984), .A2(n25245), .B1(n27840), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N2741) );
  sky130_fd_sc_hd__o22ai_1 U30418 ( .A1(n25985), .A2(n25245), .B1(n27842), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N3111) );
  sky130_fd_sc_hd__o22ai_1 U30419 ( .A1(n25986), .A2(n25245), .B1(n27843), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N3000) );
  sky130_fd_sc_hd__o22ai_1 U30420 ( .A1(n25987), .A2(n25245), .B1(n27844), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N3148) );
  sky130_fd_sc_hd__o22ai_1 U30421 ( .A1(n25988), .A2(n25245), .B1(n27845), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N2852) );
  sky130_fd_sc_hd__o22ai_1 U30422 ( .A1(n25989), .A2(n25245), .B1(n27846), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N2778) );
  sky130_fd_sc_hd__a21oi_1 U30423 ( .A1(n27768), .A2(
        j202_soc_core_j22_cpu_ml_bufa[25]), .B1(n27766), .Y(n25254) );
  sky130_fd_sc_hd__nand2_1 U30425 ( .A(n25255), .B(n27828), .Y(n25257) );
  sky130_fd_sc_hd__nor2_1 U30426 ( .A(n25257), .B(n25256), .Y(n25258) );
  sky130_fd_sc_hd__a31oi_1 U30427 ( .A1(n25262), .A2(n27052), .A3(n25261), 
        .B1(n26926), .Y(n25280) );
  sky130_fd_sc_hd__nand3_1 U30428 ( .A(n28477), .B(n27786), .C(n27032), .Y(
        n25279) );
  sky130_fd_sc_hd__nand2_1 U30429 ( .A(n27032), .B(n25263), .Y(n25264) );
  sky130_fd_sc_hd__a22o_1 U30430 ( .A1(n27785), .A2(n27032), .B1(n25264), .B2(
        n27786), .X(n25265) );
  sky130_fd_sc_hd__inv_2 U30431 ( .A(n28477), .Y(n25282) );
  sky130_fd_sc_hd__o21a_1 U30432 ( .A1(n26939), .A2(n26276), .B1(n25266), .X(
        n25267) );
  sky130_fd_sc_hd__o22a_1 U30433 ( .A1(n28475), .A2(n27793), .B1(n27796), .B2(
        n25267), .X(n25268) );
  sky130_fd_sc_hd__o21ai_1 U30434 ( .A1(n26323), .A2(n27795), .B1(n25268), .Y(
        n25270) );
  sky130_fd_sc_hd__o22ai_1 U30435 ( .A1(n26320), .A2(n27799), .B1(n26944), 
        .B2(n27797), .Y(n25269) );
  sky130_fd_sc_hd__nor2_1 U30436 ( .A(n25270), .B(n25269), .Y(n25274) );
  sky130_fd_sc_hd__xor2_1 U30437 ( .A(n27032), .B(n26276), .X(n26236) );
  sky130_fd_sc_hd__o22a_1 U30438 ( .A1(n27825), .A2(n27803), .B1(n25872), .B2(
        n26236), .X(n25273) );
  sky130_fd_sc_hd__a22oi_1 U30439 ( .A1(n27810), .A2(n27042), .B1(n27808), 
        .B2(n25271), .Y(n25272) );
  sky130_fd_sc_hd__nand4_1 U30440 ( .A(n27814), .B(n25274), .C(n25273), .D(
        n25272), .Y(n25276) );
  sky130_fd_sc_hd__o22ai_1 U30441 ( .A1(n26276), .A2(n27817), .B1(n26215), 
        .B2(n27815), .Y(n25275) );
  sky130_fd_sc_hd__nor2_1 U30442 ( .A(n25276), .B(n25275), .Y(n25278) );
  sky130_fd_sc_hd__nand2_1 U30443 ( .A(n25288), .B(n27789), .Y(n25277) );
  sky130_fd_sc_hd__buf_6 U30444 ( .A(n25284), .X(n25290) );
  sky130_fd_sc_hd__nand2_1 U30445 ( .A(n25282), .B(n23749), .Y(n25283) );
  sky130_fd_sc_hd__buf_4 U30446 ( .A(n25284), .X(n25766) );
  sky130_fd_sc_hd__o22ai_1 U30447 ( .A1(n27859), .A2(n28477), .B1(n27858), 
        .B2(n25766), .Y(j202_soc_core_j22_cpu_rf_N3337) );
  sky130_fd_sc_hd__nor2_1 U30448 ( .A(n27644), .B(n25290), .Y(
        j202_soc_core_j22_cpu_rf_N2670) );
  sky130_fd_sc_hd__o22ai_1 U30449 ( .A1(n27841), .A2(n28477), .B1(n24712), 
        .B2(n25290), .Y(j202_soc_core_j22_cpu_rf_N3261) );
  sky130_fd_sc_hd__o22ai_1 U30450 ( .A1(n25964), .A2(n28477), .B1(n27847), 
        .B2(n25290), .Y(j202_soc_core_j22_cpu_rf_N2706) );
  sky130_fd_sc_hd__o22ai_1 U30451 ( .A1(n25286), .A2(n27775), .B1(n27774), 
        .B2(n28477), .Y(n25285) );
  sky130_fd_sc_hd__o22ai_1 U30452 ( .A1(n26276), .A2(n27850), .B1(n25286), 
        .B2(n27848), .Y(n25287) );
  sky130_fd_sc_hd__a21oi_1 U30453 ( .A1(n25288), .A2(n26068), .B1(n25287), .Y(
        n25289) );
  sky130_fd_sc_hd__o22ai_1 U30455 ( .A1(n25977), .A2(n28477), .B1(n28061), 
        .B2(n25290), .Y(j202_soc_core_j22_cpu_rf_N2891) );
  sky130_fd_sc_hd__o22ai_1 U30456 ( .A1(n25978), .A2(n28477), .B1(n27834), 
        .B2(n25290), .Y(j202_soc_core_j22_cpu_rf_N2965) );
  sky130_fd_sc_hd__o22ai_1 U30457 ( .A1(n25979), .A2(n28477), .B1(n28112), 
        .B2(n25766), .Y(j202_soc_core_j22_cpu_rf_N3224) );
  sky130_fd_sc_hd__o22ai_1 U30458 ( .A1(n25980), .A2(n28477), .B1(n27835), 
        .B2(n25290), .Y(j202_soc_core_j22_cpu_rf_N2817) );
  sky130_fd_sc_hd__o22ai_1 U30459 ( .A1(n25981), .A2(n28477), .B1(n27836), 
        .B2(n25766), .Y(j202_soc_core_j22_cpu_rf_N3187) );
  sky130_fd_sc_hd__o22ai_1 U30460 ( .A1(n25982), .A2(n28477), .B1(n27837), 
        .B2(n25290), .Y(j202_soc_core_j22_cpu_rf_N3039) );
  sky130_fd_sc_hd__o22ai_1 U30461 ( .A1(n25983), .A2(n28477), .B1(n27838), 
        .B2(n25766), .Y(j202_soc_core_j22_cpu_rf_N3076) );
  sky130_fd_sc_hd__o22ai_1 U30462 ( .A1(n25984), .A2(n28477), .B1(n27840), 
        .B2(n25290), .Y(j202_soc_core_j22_cpu_rf_N2743) );
  sky130_fd_sc_hd__o22ai_1 U30463 ( .A1(n25985), .A2(n28477), .B1(n27842), 
        .B2(n25290), .Y(j202_soc_core_j22_cpu_rf_N3113) );
  sky130_fd_sc_hd__o22ai_1 U30464 ( .A1(n25986), .A2(n28477), .B1(n27843), 
        .B2(n25290), .Y(j202_soc_core_j22_cpu_rf_N3002) );
  sky130_fd_sc_hd__o22ai_1 U30465 ( .A1(n25987), .A2(n28477), .B1(n27844), 
        .B2(n25290), .Y(j202_soc_core_j22_cpu_rf_N3150) );
  sky130_fd_sc_hd__o22ai_1 U30466 ( .A1(n25988), .A2(n28477), .B1(n27845), 
        .B2(n25766), .Y(j202_soc_core_j22_cpu_rf_N2854) );
  sky130_fd_sc_hd__o22ai_1 U30467 ( .A1(n25989), .A2(n28477), .B1(n27846), 
        .B2(n25290), .Y(j202_soc_core_j22_cpu_rf_N2780) );
  sky130_fd_sc_hd__nand2_1 U30469 ( .A(n26177), .B(n26189), .Y(n25291) );
  sky130_fd_sc_hd__o22ai_1 U30470 ( .A1(n26944), .A2(n27799), .B1(n27796), 
        .B2(n26943), .Y(n25293) );
  sky130_fd_sc_hd__o22ai_1 U30471 ( .A1(n26322), .A2(n27795), .B1(n26284), 
        .B2(n27797), .Y(n25292) );
  sky130_fd_sc_hd__nor2_1 U30472 ( .A(n25293), .B(n25292), .Y(n25299) );
  sky130_fd_sc_hd__xor2_1 U30473 ( .A(n26051), .B(n26285), .X(n26230) );
  sky130_fd_sc_hd__a22oi_1 U30474 ( .A1(n26414), .A2(n25294), .B1(n26285), 
        .B2(n26034), .Y(n25295) );
  sky130_fd_sc_hd__o21ai_0 U30475 ( .A1(n27800), .A2(n27803), .B1(n25295), .Y(
        n25296) );
  sky130_fd_sc_hd__a21oi_1 U30476 ( .A1(n27808), .A2(n26064), .B1(n25296), .Y(
        n25297) );
  sky130_fd_sc_hd__nand4_1 U30477 ( .A(n27814), .B(n25299), .C(n25298), .D(
        n25297), .Y(n25301) );
  sky130_fd_sc_hd__o22ai_1 U30478 ( .A1(n26285), .A2(n27817), .B1(n11144), 
        .B2(n27815), .Y(n25300) );
  sky130_fd_sc_hd__nor2_1 U30479 ( .A(n25301), .B(n25300), .Y(n25302) );
  sky130_fd_sc_hd__nand2_1 U30480 ( .A(n26051), .B(n27785), .Y(n25303) );
  sky130_fd_sc_hd__o211ai_1 U30481 ( .A1(n11123), .A2(n26051), .B1(n26922), 
        .C1(n25303), .Y(n25304) );
  sky130_fd_sc_hd__nand2_1 U30482 ( .A(n28525), .B(n25304), .Y(n25305) );
  sky130_fd_sc_hd__o211ai_1 U30483 ( .A1(n25658), .A2(n25307), .B1(n25306), 
        .C1(n25305), .Y(n25308) );
  sky130_fd_sc_hd__a21oi_2 U30484 ( .A1(n25309), .A2(n26051), .B1(n25308), .Y(
        n25722) );
  sky130_fd_sc_hd__o22ai_1 U30485 ( .A1(n25977), .A2(n25765), .B1(n28061), 
        .B2(n12056), .Y(j202_soc_core_j22_cpu_rf_N2882) );
  sky130_fd_sc_hd__o22ai_1 U30486 ( .A1(n25978), .A2(n25765), .B1(n27834), 
        .B2(n12056), .Y(j202_soc_core_j22_cpu_rf_N2956) );
  sky130_fd_sc_hd__o22ai_1 U30487 ( .A1(n25979), .A2(n25765), .B1(n28112), 
        .B2(n12056), .Y(j202_soc_core_j22_cpu_rf_N3215) );
  sky130_fd_sc_hd__o22ai_1 U30488 ( .A1(n25980), .A2(n25765), .B1(n27835), 
        .B2(n12056), .Y(j202_soc_core_j22_cpu_rf_N2808) );
  sky130_fd_sc_hd__o22ai_1 U30489 ( .A1(n25981), .A2(n25765), .B1(n27836), 
        .B2(n12057), .Y(j202_soc_core_j22_cpu_rf_N3178) );
  sky130_fd_sc_hd__o22ai_1 U30490 ( .A1(n25982), .A2(n25765), .B1(n27837), 
        .B2(n12057), .Y(j202_soc_core_j22_cpu_rf_N3030) );
  sky130_fd_sc_hd__o22ai_1 U30491 ( .A1(n25983), .A2(n25765), .B1(n27838), 
        .B2(n12056), .Y(j202_soc_core_j22_cpu_rf_N3067) );
  sky130_fd_sc_hd__o22ai_1 U30492 ( .A1(n25984), .A2(n25765), .B1(n27840), 
        .B2(n12057), .Y(j202_soc_core_j22_cpu_rf_N2734) );
  sky130_fd_sc_hd__o22ai_1 U30493 ( .A1(n27841), .A2(n25765), .B1(n24712), 
        .B2(n12057), .Y(j202_soc_core_j22_cpu_rf_N3252) );
  sky130_fd_sc_hd__o22ai_1 U30494 ( .A1(n25985), .A2(n25765), .B1(n27842), 
        .B2(n12056), .Y(j202_soc_core_j22_cpu_rf_N3104) );
  sky130_fd_sc_hd__o22ai_1 U30495 ( .A1(n25986), .A2(n25765), .B1(n27843), 
        .B2(n12056), .Y(j202_soc_core_j22_cpu_rf_N2993) );
  sky130_fd_sc_hd__o22ai_1 U30496 ( .A1(n25987), .A2(n25765), .B1(n27844), 
        .B2(n12056), .Y(j202_soc_core_j22_cpu_rf_N3141) );
  sky130_fd_sc_hd__o22ai_1 U30497 ( .A1(n25988), .A2(n25765), .B1(n27845), 
        .B2(n12057), .Y(j202_soc_core_j22_cpu_rf_N2845) );
  sky130_fd_sc_hd__o22ai_1 U30498 ( .A1(n25989), .A2(n25765), .B1(n27846), 
        .B2(n12056), .Y(j202_soc_core_j22_cpu_rf_N2771) );
  sky130_fd_sc_hd__o22ai_1 U30499 ( .A1(n25964), .A2(n25765), .B1(n27847), 
        .B2(n12057), .Y(j202_soc_core_j22_cpu_rf_N2697) );
  sky130_fd_sc_hd__nand2_1 U30500 ( .A(n25313), .B(n24832), .Y(n25312) );
  sky130_fd_sc_hd__nand2_1 U30501 ( .A(n28525), .B(n23749), .Y(n25311) );
  sky130_fd_sc_hd__nand2_1 U30502 ( .A(n25312), .B(n25311), .Y(
        j202_soc_core_j22_cpu_rf_N3289) );
  sky130_fd_sc_hd__o22ai_1 U30503 ( .A1(n25765), .A2(n27859), .B1(n27858), 
        .B2(n12057), .Y(j202_soc_core_j22_cpu_rf_N3328) );
  sky130_fd_sc_hd__o21ai_1 U30504 ( .A1(n25677), .A2(n27770), .B1(n25374), .Y(
        j202_soc_core_j22_cpu_ml_maclj[19]) );
  sky130_fd_sc_hd__nand2_1 U30505 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[19]), .Y(n25314) );
  sky130_fd_sc_hd__o21ai_1 U30506 ( .A1(n25315), .A2(n28545), .B1(n25314), .Y(
        n36) );
  sky130_fd_sc_hd__nand2_1 U30507 ( .A(n25317), .B(j202_soc_core_aquc_SEL__2_), 
        .Y(n27624) );
  sky130_fd_sc_hd__nand2_1 U30508 ( .A(n27624), .B(j202_soc_core_uart_div1[3]), 
        .Y(n25318) );
  sky130_fd_sc_hd__o22ai_1 U30510 ( .A1(n29150), .A2(n28310), .B1(n25320), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U30511 ( .A1(n29150), .A2(n28313), .B1(n25321), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U30512 ( .A1(n29150), .A2(n28316), .B1(n25322), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U30513 ( .A1(n29150), .A2(n26760), .B1(n25323), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U30514 ( .A1(n29150), .A2(n27575), .B1(n25324), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U30515 ( .A1(n29150), .A2(n28553), .B1(n25325), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U30516 ( .A1(n29150), .A2(n29082), .B1(n25326), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U30517 ( .A1(n29150), .A2(n29076), .B1(n25327), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__a22oi_1 U30518 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[19]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[19]), .Y(n25329) );
  sky130_fd_sc_hd__a22oi_1 U30519 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[116]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[100]), .Y(n25328) );
  sky130_fd_sc_hd__nand3_1 U30520 ( .A(n25329), .B(n28238), .C(n25328), .Y(
        n25330) );
  sky130_fd_sc_hd__a21oi_1 U30521 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[115]), .B1(n25330), .Y(n25334) );
  sky130_fd_sc_hd__a22oi_1 U30522 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[124]), .B1(n28331), .B2(
        j202_soc_core_intc_core_00_rg_itgt[108]), .Y(n25333) );
  sky130_fd_sc_hd__a22oi_1 U30523 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[19]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[51]), .B2(n28330), .Y(n25332) );
  sky130_fd_sc_hd__nand2_1 U30524 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[83]), .Y(n25331) );
  sky130_fd_sc_hd__nand4_1 U30525 ( .A(n25334), .B(n25333), .C(n25332), .D(
        n25331), .Y(j202_soc_core_ahb2apb_01_N147) );
  sky130_fd_sc_hd__nand2_1 U30526 ( .A(n26543), .B(n28914), .Y(n25335) );
  sky130_fd_sc_hd__nand2b_1 U30527 ( .A_N(n27183), .B(n26588), .Y(n27613) );
  sky130_fd_sc_hd__nor2_1 U30528 ( .A(n25335), .B(n27613), .Y(
        j202_soc_core_wbqspiflash_00_N744) );
  sky130_fd_sc_hd__nand2_1 U30529 ( .A(n25336), .B(n29827), .Y(
        j202_soc_core_wbqspiflash_00_N743) );
  sky130_fd_sc_hd__o31ai_1 U30530 ( .A1(n27238), .A2(n27232), .A3(n27284), 
        .B1(n25337), .Y(j202_soc_core_wbqspiflash_00_N663) );
  sky130_fd_sc_hd__nor2_1 U30531 ( .A(n28895), .B(n25338), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N323) );
  sky130_fd_sc_hd__mux2i_1 U30532 ( .A0(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[0]), .A1(io_in[11]), .S(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n25503) );
  sky130_fd_sc_hd__nor2_1 U30533 ( .A(n28898), .B(n25503), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N359) );
  sky130_fd_sc_hd__nor2_1 U30534 ( .A(n26575), .B(n27280), .Y(n28848) );
  sky130_fd_sc_hd__nand2_1 U30535 ( .A(n28848), .B(
        j202_soc_core_wbqspiflash_00_spif_data[1]), .Y(n28753) );
  sky130_fd_sc_hd__nand2_1 U30536 ( .A(n27429), .B(
        j202_soc_core_wbqspiflash_00_spi_out[1]), .Y(n25339) );
  sky130_fd_sc_hd__a21oi_1 U30537 ( .A1(n28753), .A2(n25339), .B1(
        j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N739) );
  sky130_fd_sc_hd__o211ai_1 U30538 ( .A1(n26612), .A2(n26512), .B1(n29830), 
        .C1(n25340), .Y(j202_soc_core_wbqspiflash_00_N738) );
  sky130_fd_sc_hd__nand2_1 U30539 ( .A(n28655), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .Y(n27261) );
  sky130_fd_sc_hd__nor2_1 U30540 ( .A(n26483), .B(n27201), .Y(n28836) );
  sky130_fd_sc_hd__o22ai_1 U30541 ( .A1(n27261), .A2(n26529), .B1(n28867), 
        .B2(n25341), .Y(n25343) );
  sky130_fd_sc_hd__nand2_1 U30542 ( .A(n28870), .B(n28647), .Y(n26498) );
  sky130_fd_sc_hd__nor2_1 U30543 ( .A(n26575), .B(n26498), .Y(n28730) );
  sky130_fd_sc_hd__nor2_1 U30544 ( .A(j202_soc_core_wbqspiflash_00_state[4]), 
        .B(n25342), .Y(n28878) );
  sky130_fd_sc_hd__nor2_1 U30545 ( .A(n28814), .B(n28878), .Y(n28666) );
  sky130_fd_sc_hd__o21ai_1 U30546 ( .A1(n28857), .A2(n27261), .B1(n28666), .Y(
        n28654) );
  sky130_fd_sc_hd__nor2_1 U30547 ( .A(n25343), .B(n28654), .Y(n28892) );
  sky130_fd_sc_hd__nand2b_1 U30548 ( .A_N(n26498), .B(n26521), .Y(n28724) );
  sky130_fd_sc_hd__nand2b_1 U30549 ( .A_N(n27183), .B(n26484), .Y(n28734) );
  sky130_fd_sc_hd__a22oi_1 U30550 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[31]), .B1(n28887), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]), .Y(n25347) );
  sky130_fd_sc_hd__nor2_1 U30551 ( .A(j202_soc_core_wbqspiflash_00_spif_ctrl), 
        .B(j202_soc_core_wbqspiflash_00_spif_cmd), .Y(n28729) );
  sky130_fd_sc_hd__nand2_1 U30552 ( .A(n27614), .B(n28841), .Y(n27297) );
  sky130_fd_sc_hd__nand2_1 U30553 ( .A(n27298), .B(n26489), .Y(n28747) );
  sky130_fd_sc_hd__nor2_1 U30554 ( .A(j202_soc_core_wbqspiflash_00_state[2]), 
        .B(n28747), .Y(n28847) );
  sky130_fd_sc_hd__a21oi_1 U30555 ( .A1(n28730), .A2(n28729), .B1(n28847), .Y(
        n28884) );
  sky130_fd_sc_hd__nor2_1 U30556 ( .A(n28884), .B(n27296), .Y(n28662) );
  sky130_fd_sc_hd__nor2_1 U30557 ( .A(n28662), .B(n25344), .Y(n28667) );
  sky130_fd_sc_hd__nand2b_1 U30558 ( .A_N(n27183), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n26507) );
  sky130_fd_sc_hd__nor2_1 U30559 ( .A(n25345), .B(n26507), .Y(n28675) );
  sky130_fd_sc_hd__nand2_1 U30560 ( .A(n28675), .B(
        j202_soc_core_qspi_wb_addr[23]), .Y(n25346) );
  sky130_fd_sc_hd__nand4_1 U30561 ( .A(n28892), .B(n25347), .C(n28667), .D(
        n25346), .Y(n10544) );
  sky130_fd_sc_hd__a21oi_1 U30562 ( .A1(n27768), .A2(n25627), .B1(n27766), .Y(
        n25348) );
  sky130_fd_sc_hd__o21ai_1 U30563 ( .A1(n25371), .A2(n27770), .B1(n25348), .Y(
        j202_soc_core_j22_cpu_ml_maclj[22]) );
  sky130_fd_sc_hd__nand2_1 U30564 ( .A(n26190), .B(n26189), .Y(n25350) );
  sky130_fd_sc_hd__nand2_1 U30565 ( .A(n25626), .B(n27152), .Y(n25373) );
  sky130_fd_sc_hd__o21a_1 U30566 ( .A1(n26277), .A2(n26939), .B1(n26919), .X(
        n25351) );
  sky130_fd_sc_hd__nand2_1 U30567 ( .A(n25352), .B(n25351), .Y(n25370) );
  sky130_fd_sc_hd__nand2_1 U30568 ( .A(n26324), .B(n26916), .Y(n25354) );
  sky130_fd_sc_hd__nand2_1 U30569 ( .A(n25642), .B(n27785), .Y(n25353) );
  sky130_fd_sc_hd__nand4_1 U30570 ( .A(n25354), .B(n27787), .C(n25353), .D(
        n25638), .Y(n25355) );
  sky130_fd_sc_hd__nand2_1 U30571 ( .A(n28492), .B(n25355), .Y(n25368) );
  sky130_fd_sc_hd__o22ai_1 U30572 ( .A1(n26280), .A2(n27795), .B1(n26435), 
        .B2(n26943), .Y(n25357) );
  sky130_fd_sc_hd__o22ai_1 U30573 ( .A1(n26431), .A2(n27803), .B1(n11191), 
        .B2(n27797), .Y(n25356) );
  sky130_fd_sc_hd__nor2_1 U30574 ( .A(n25357), .B(n25356), .Y(n25363) );
  sky130_fd_sc_hd__xor2_1 U30575 ( .A(n28493), .B(n25642), .X(n26227) );
  sky130_fd_sc_hd__a22oi_1 U30576 ( .A1(n26227), .A2(n27806), .B1(n27808), 
        .B2(n26331), .Y(n25362) );
  sky130_fd_sc_hd__o22ai_1 U30577 ( .A1(n26926), .A2(n25358), .B1(n27793), 
        .B2(n28493), .Y(n25360) );
  sky130_fd_sc_hd__nor2_1 U30578 ( .A(n26319), .B(n27799), .Y(n25359) );
  sky130_fd_sc_hd__a211oi_1 U30579 ( .A1(n27810), .A2(n27807), .B1(n25360), 
        .C1(n25359), .Y(n25361) );
  sky130_fd_sc_hd__nand4_1 U30580 ( .A(n27814), .B(n25363), .C(n25362), .D(
        n25361), .Y(n25365) );
  sky130_fd_sc_hd__o22ai_1 U30581 ( .A1(n26277), .A2(n27817), .B1(n25944), 
        .B2(n27815), .Y(n25364) );
  sky130_fd_sc_hd__nor2_1 U30582 ( .A(n25365), .B(n25364), .Y(n25367) );
  sky130_fd_sc_hd__nand2_1 U30583 ( .A(n25601), .B(n27789), .Y(n25366) );
  sky130_fd_sc_hd__o22ai_1 U30584 ( .A1(n26894), .A2(n25632), .B1(n27839), 
        .B2(n12059), .Y(j202_soc_core_j22_cpu_rf_N2925) );
  sky130_fd_sc_hd__o22ai_1 U30585 ( .A1(n25980), .A2(n25632), .B1(n27835), 
        .B2(n12058), .Y(j202_soc_core_j22_cpu_rf_N2814) );
  sky130_fd_sc_hd__o22ai_1 U30586 ( .A1(n25983), .A2(n25632), .B1(n27838), 
        .B2(n12059), .Y(j202_soc_core_j22_cpu_rf_N3073) );
  sky130_fd_sc_hd__o22ai_1 U30587 ( .A1(n25977), .A2(n25632), .B1(n28061), 
        .B2(n12058), .Y(j202_soc_core_j22_cpu_rf_N2888) );
  sky130_fd_sc_hd__o22ai_1 U30588 ( .A1(n25979), .A2(n25632), .B1(n28112), 
        .B2(n12059), .Y(j202_soc_core_j22_cpu_rf_N3221) );
  sky130_fd_sc_hd__o22ai_1 U30589 ( .A1(n25981), .A2(n25632), .B1(n27836), 
        .B2(n25604), .Y(j202_soc_core_j22_cpu_rf_N3184) );
  sky130_fd_sc_hd__o22ai_1 U30590 ( .A1(n25986), .A2(n25632), .B1(n27843), 
        .B2(n12058), .Y(j202_soc_core_j22_cpu_rf_N2999) );
  sky130_fd_sc_hd__o22ai_1 U30591 ( .A1(n25982), .A2(n25632), .B1(n27837), 
        .B2(n25604), .Y(j202_soc_core_j22_cpu_rf_N3036) );
  sky130_fd_sc_hd__o22ai_1 U30592 ( .A1(n25964), .A2(n25632), .B1(n27847), 
        .B2(n25604), .Y(j202_soc_core_j22_cpu_rf_N2703) );
  sky130_fd_sc_hd__o22ai_1 U30593 ( .A1(n25985), .A2(n25632), .B1(n27842), 
        .B2(n12059), .Y(j202_soc_core_j22_cpu_rf_N3110) );
  sky130_fd_sc_hd__o22ai_1 U30594 ( .A1(n25987), .A2(n25632), .B1(n27844), 
        .B2(n12058), .Y(j202_soc_core_j22_cpu_rf_N3147) );
  sky130_fd_sc_hd__o22ai_1 U30595 ( .A1(n25989), .A2(n25632), .B1(n27846), 
        .B2(n12059), .Y(j202_soc_core_j22_cpu_rf_N2777) );
  sky130_fd_sc_hd__o22ai_1 U30596 ( .A1(n25984), .A2(n25632), .B1(n27840), 
        .B2(n12058), .Y(j202_soc_core_j22_cpu_rf_N2740) );
  sky130_fd_sc_hd__o22ai_1 U30597 ( .A1(n25988), .A2(n25632), .B1(n27845), 
        .B2(n12059), .Y(j202_soc_core_j22_cpu_rf_N2851) );
  sky130_fd_sc_hd__o22ai_1 U30598 ( .A1(n25978), .A2(n25632), .B1(n27834), 
        .B2(n12058), .Y(j202_soc_core_j22_cpu_rf_N2962) );
  sky130_fd_sc_hd__o22ai_1 U30599 ( .A1(n27841), .A2(n25632), .B1(n24712), 
        .B2(n25604), .Y(j202_soc_core_j22_cpu_rf_N3258) );
  sky130_fd_sc_hd__nand4_1 U30601 ( .A(n25378), .B(n25379), .C(n25377), .D(
        n25376), .Y(n25380) );
  sky130_fd_sc_hd__nand2_1 U30602 ( .A(n25383), .B(n24832), .Y(n25382) );
  sky130_fd_sc_hd__o21ai_0 U30603 ( .A1(n24832), .A2(n25594), .B1(n25382), .Y(
        j202_soc_core_j22_cpu_rf_N3294) );
  sky130_fd_sc_hd__o22ai_1 U30604 ( .A1(n27841), .A2(n25594), .B1(n24712), 
        .B2(n12266), .Y(j202_soc_core_j22_cpu_rf_N3257) );
  sky130_fd_sc_hd__o22ai_1 U30605 ( .A1(n26281), .A2(n27850), .B1(n13047), 
        .B2(n27848), .Y(n25384) );
  sky130_fd_sc_hd__a21oi_1 U30606 ( .A1(n25385), .A2(n26068), .B1(n25384), .Y(
        n25386) );
  sky130_fd_sc_hd__o21ai_0 U30607 ( .A1(n27855), .A2(n25594), .B1(n25386), .Y(
        j202_soc_core_j22_cpu_rf_N319) );
  sky130_fd_sc_hd__o22ai_1 U30608 ( .A1(n25977), .A2(n25594), .B1(n28061), 
        .B2(n12266), .Y(j202_soc_core_j22_cpu_rf_N2887) );
  sky130_fd_sc_hd__o22ai_1 U30609 ( .A1(n25978), .A2(n25594), .B1(n27834), 
        .B2(n12267), .Y(j202_soc_core_j22_cpu_rf_N2961) );
  sky130_fd_sc_hd__o22ai_1 U30610 ( .A1(n25979), .A2(n25594), .B1(n28112), 
        .B2(n12267), .Y(j202_soc_core_j22_cpu_rf_N3220) );
  sky130_fd_sc_hd__o22ai_1 U30611 ( .A1(n25981), .A2(n25594), .B1(n27836), 
        .B2(n12266), .Y(j202_soc_core_j22_cpu_rf_N3183) );
  sky130_fd_sc_hd__o22ai_1 U30612 ( .A1(n25982), .A2(n25594), .B1(n27837), 
        .B2(n12266), .Y(j202_soc_core_j22_cpu_rf_N3035) );
  sky130_fd_sc_hd__o22ai_1 U30613 ( .A1(n25983), .A2(n25594), .B1(n27838), 
        .B2(n12266), .Y(j202_soc_core_j22_cpu_rf_N3072) );
  sky130_fd_sc_hd__o22ai_1 U30614 ( .A1(n26894), .A2(n25594), .B1(n27839), 
        .B2(n12267), .Y(j202_soc_core_j22_cpu_rf_N2924) );
  sky130_fd_sc_hd__o22ai_1 U30615 ( .A1(n25984), .A2(n25594), .B1(n27840), 
        .B2(n12267), .Y(j202_soc_core_j22_cpu_rf_N2739) );
  sky130_fd_sc_hd__o22ai_1 U30616 ( .A1(n25985), .A2(n25594), .B1(n27842), 
        .B2(n12266), .Y(j202_soc_core_j22_cpu_rf_N3109) );
  sky130_fd_sc_hd__o22ai_1 U30617 ( .A1(n25986), .A2(n25594), .B1(n27843), 
        .B2(n12266), .Y(j202_soc_core_j22_cpu_rf_N2998) );
  sky130_fd_sc_hd__o22ai_1 U30618 ( .A1(n25987), .A2(n25594), .B1(n27844), 
        .B2(n12267), .Y(j202_soc_core_j22_cpu_rf_N3146) );
  sky130_fd_sc_hd__o22ai_1 U30619 ( .A1(n25988), .A2(n25594), .B1(n27845), 
        .B2(n12266), .Y(j202_soc_core_j22_cpu_rf_N2850) );
  sky130_fd_sc_hd__o22ai_1 U30620 ( .A1(n25989), .A2(n25594), .B1(n27846), 
        .B2(n12267), .Y(j202_soc_core_j22_cpu_rf_N2776) );
  sky130_fd_sc_hd__nand2_1 U30621 ( .A(n12203), .B(n25464), .Y(n25388) );
  sky130_fd_sc_hd__nand2_1 U30622 ( .A(n28056), .B(n25389), .Y(n25387) );
  sky130_fd_sc_hd__nand3_1 U30623 ( .A(n25388), .B(n27119), .C(n25387), .Y(
        n29836) );
  sky130_fd_sc_hd__a21oi_1 U30624 ( .A1(n27768), .A2(n25389), .B1(n27766), .Y(
        n25390) );
  sky130_fd_sc_hd__o21ai_1 U30625 ( .A1(n25391), .A2(n27770), .B1(n25390), .Y(
        j202_soc_core_j22_cpu_ml_maclj[29]) );
  sky130_fd_sc_hd__nand2_1 U30626 ( .A(n29564), .B(n25392), .Y(n25396) );
  sky130_fd_sc_hd__nand3_2 U30627 ( .A(n11139), .B(n25396), .C(n25393), .Y(
        n28453) );
  sky130_fd_sc_hd__nand4_1 U30628 ( .A(n11139), .B(n26916), .C(n25396), .D(
        n25393), .Y(n25400) );
  sky130_fd_sc_hd__o21a_1 U30630 ( .A1(n25397), .A2(n25396), .B1(n25395), .X(
        n25399) );
  sky130_fd_sc_hd__nand2_1 U30631 ( .A(n12360), .B(n27785), .Y(n25398) );
  sky130_fd_sc_hd__nand3_1 U30632 ( .A(n25400), .B(n25399), .C(n25398), .Y(
        n25419) );
  sky130_fd_sc_hd__nand2_1 U30634 ( .A(n28453), .B(n25401), .Y(n25417) );
  sky130_fd_sc_hd__o21ai_1 U30635 ( .A1(n25451), .A2(n26934), .B1(n26933), .Y(
        n25413) );
  sky130_fd_sc_hd__nor2_1 U30636 ( .A(n26319), .B(n27803), .Y(n25405) );
  sky130_fd_sc_hd__nand2b_1 U30637 ( .A_N(n25451), .B(n26050), .Y(n26300) );
  sky130_fd_sc_hd__o22ai_1 U30638 ( .A1(n27793), .A2(n28454), .B1(n26939), 
        .B2(n26300), .Y(n25404) );
  sky130_fd_sc_hd__o22ai_1 U30639 ( .A1(n11189), .A2(n27799), .B1(n26280), 
        .B2(n26943), .Y(n25403) );
  sky130_fd_sc_hd__or4_1 U30641 ( .A(n25405), .B(n25404), .C(n25403), .D(
        n25402), .X(n25412) );
  sky130_fd_sc_hd__nand2_1 U30642 ( .A(n25406), .B(n26414), .Y(n25408) );
  sky130_fd_sc_hd__nand2_1 U30643 ( .A(n26321), .B(n25451), .Y(n26212) );
  sky130_fd_sc_hd__nand3_1 U30644 ( .A(n26300), .B(n26212), .C(n27806), .Y(
        n25407) );
  sky130_fd_sc_hd__o211a_2 U30645 ( .A1(n26318), .A2(n27795), .B1(n25408), 
        .C1(n25407), .X(n25410) );
  sky130_fd_sc_hd__a2bb2oi_1 U30646 ( .B1(n27033), .B2(n26935), .A1_N(n26421), 
        .A2_N(n26936), .Y(n25409) );
  sky130_fd_sc_hd__o211ai_1 U30647 ( .A1(n28451), .A2(n26932), .B1(n25410), 
        .C1(n25409), .Y(n25411) );
  sky130_fd_sc_hd__or3_1 U30648 ( .A(n25413), .B(n25412), .C(n25411), .X(
        n25414) );
  sky130_fd_sc_hd__a21oi_1 U30649 ( .A1(n25430), .A2(n27789), .B1(n25414), .Y(
        n25415) );
  sky130_fd_sc_hd__o21a_1 U30650 ( .A1(n26926), .A2(n27714), .B1(n25415), .X(
        n25416) );
  sky130_fd_sc_hd__a21oi_2 U30651 ( .A1(n26050), .A2(n25419), .B1(n25418), .Y(
        n25425) );
  sky130_fd_sc_hd__mux2i_1 U30653 ( .A0(n25420), .A1(n25556), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3284) );
  sky130_fd_sc_hd__nor2_1 U30654 ( .A(n27644), .B(n25420), .Y(
        j202_soc_core_j22_cpu_rf_N2656) );
  sky130_fd_sc_hd__mux2i_1 U30655 ( .A0(n25556), .A1(n26321), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N316) );
  sky130_fd_sc_hd__nand2_1 U30656 ( .A(n28055), .B(n25421), .Y(n25422) );
  sky130_fd_sc_hd__nand2_1 U30657 ( .A(n25422), .B(n12203), .Y(
        j202_soc_core_j22_cpu_ml_machj[13]) );
  sky130_fd_sc_hd__a22oi_1 U30658 ( .A1(n25423), .A2(n27862), .B1(n28453), 
        .B2(n27861), .Y(n25424) );
  sky130_fd_sc_hd__o21ai_0 U30659 ( .A1(n27648), .A2(n25427), .B1(n25426), .Y(
        j202_soc_core_j22_cpu_rf_N3359) );
  sky130_fd_sc_hd__nand2_1 U30660 ( .A(n28453), .B(n25724), .Y(n25432) );
  sky130_fd_sc_hd__o22ai_1 U30661 ( .A1(n25451), .A2(n27850), .B1(n25428), 
        .B2(n27848), .Y(n25429) );
  sky130_fd_sc_hd__a21oi_1 U30662 ( .A1(n25430), .A2(n26068), .B1(n25429), .Y(
        n25431) );
  sky130_fd_sc_hd__nand2_1 U30663 ( .A(n25432), .B(n25431), .Y(
        j202_soc_core_j22_cpu_rf_N311) );
  sky130_fd_sc_hd__nand2_1 U30664 ( .A(n25464), .B(n27152), .Y(n25462) );
  sky130_fd_sc_hd__nand2_1 U30665 ( .A(n25466), .B(n27785), .Y(n25436) );
  sky130_fd_sc_hd__o21a_1 U30666 ( .A1(n28451), .A2(n26939), .B1(n26919), .X(
        n25435) );
  sky130_fd_sc_hd__nand2_1 U30667 ( .A(n25433), .B(n26916), .Y(n25434) );
  sky130_fd_sc_hd__nand2_1 U30668 ( .A(n25437), .B(n27033), .Y(n25460) );
  sky130_fd_sc_hd__a31oi_1 U30669 ( .A1(n25440), .A2(n25439), .A3(n25438), 
        .B1(n25658), .Y(n25441) );
  sky130_fd_sc_hd__o21ai_1 U30671 ( .A1(n11123), .A2(n27033), .B1(n26922), .Y(
        n25457) );
  sky130_fd_sc_hd__nand2_1 U30672 ( .A(n25473), .B(n27789), .Y(n25455) );
  sky130_fd_sc_hd__o22ai_1 U30674 ( .A1(n26280), .A2(n27799), .B1(n26321), 
        .B2(n27797), .Y(n25446) );
  sky130_fd_sc_hd__nor2_1 U30675 ( .A(n25447), .B(n25446), .Y(n25450) );
  sky130_fd_sc_hd__xor2_1 U30676 ( .A(n27033), .B(n28451), .X(n26237) );
  sky130_fd_sc_hd__o22a_1 U30677 ( .A1(n27026), .A2(n27795), .B1(n25872), .B2(
        n26237), .X(n25449) );
  sky130_fd_sc_hd__a22oi_1 U30678 ( .A1(n27810), .A2(n26416), .B1(n27808), 
        .B2(n27042), .Y(n25448) );
  sky130_fd_sc_hd__nand4_1 U30679 ( .A(n27814), .B(n25450), .C(n25449), .D(
        n25448), .Y(n25453) );
  sky130_fd_sc_hd__o22ai_1 U30680 ( .A1(n28451), .A2(n27817), .B1(n25451), 
        .B2(n27815), .Y(n25452) );
  sky130_fd_sc_hd__nor2_1 U30681 ( .A(n25453), .B(n25452), .Y(n25454) );
  sky130_fd_sc_hd__nand2_1 U30682 ( .A(n25455), .B(n25454), .Y(n25456) );
  sky130_fd_sc_hd__a21oi_1 U30683 ( .A1(n25466), .A2(n25457), .B1(n25456), .Y(
        n25458) );
  sky130_fd_sc_hd__nand2_2 U30684 ( .A(n25462), .B(n25461), .Y(n25475) );
  sky130_fd_sc_hd__nand2_1 U30685 ( .A(n25475), .B(n24832), .Y(n25463) );
  sky130_fd_sc_hd__o21ai_0 U30686 ( .A1(n24832), .A2(n27642), .B1(n25463), .Y(
        j202_soc_core_j22_cpu_rf_N3303) );
  sky130_fd_sc_hd__nand2_1 U30687 ( .A(n25464), .B(n27772), .Y(n25470) );
  sky130_fd_sc_hd__o22ai_1 U30688 ( .A1(n25471), .A2(n27775), .B1(n27774), 
        .B2(n27642), .Y(n25467) );
  sky130_fd_sc_hd__a21oi_1 U30689 ( .A1(n25468), .A2(n27860), .B1(n25467), .Y(
        n25469) );
  sky130_fd_sc_hd__nand2_1 U30690 ( .A(n25470), .B(n25469), .Y(
        j202_soc_core_j22_cpu_rf_N3377) );
  sky130_fd_sc_hd__o22ai_1 U30691 ( .A1(n28451), .A2(n27850), .B1(n25471), 
        .B2(n27848), .Y(n25472) );
  sky130_fd_sc_hd__a21oi_1 U30692 ( .A1(n25473), .A2(n26068), .B1(n25472), .Y(
        n25474) );
  sky130_fd_sc_hd__o21ai_0 U30693 ( .A1(n27855), .A2(n27642), .B1(n25474), .Y(
        j202_soc_core_j22_cpu_rf_N327) );
  sky130_fd_sc_hd__o22ai_1 U30694 ( .A1(n27642), .A2(n27859), .B1(n27858), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N3341) );
  sky130_fd_sc_hd__o22ai_1 U30695 ( .A1(n25964), .A2(n27642), .B1(n27847), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N2711) );
  sky130_fd_sc_hd__o22ai_1 U30696 ( .A1(n27841), .A2(n27642), .B1(n24712), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N3266) );
  sky130_fd_sc_hd__nand2_1 U30698 ( .A(n25478), .B(n25477), .Y(n27916) );
  sky130_fd_sc_hd__o21a_1 U30699 ( .A1(n25480), .A2(n25479), .B1(n27916), .X(
        n27094) );
  sky130_fd_sc_hd__a21oi_1 U30700 ( .A1(n27091), .A2(n29565), .B1(n29581), .Y(
        n25481) );
  sky130_fd_sc_hd__nand2_1 U30701 ( .A(n27093), .B(n25481), .Y(n25482) );
  sky130_fd_sc_hd__nand2_1 U30702 ( .A(n27094), .B(n25482), .Y(
        j202_soc_core_ahb2aqu_00_N164) );
  sky130_fd_sc_hd__nand3_1 U30703 ( .A(j202_soc_core_aquc_WE_), .B(
        j202_soc_core_aquc_SEL__3_), .C(j202_soc_core_aquc_CE__1_), .Y(n27994)
         );
  sky130_fd_sc_hd__nand2_1 U30704 ( .A(n27994), .B(j202_soc_core_uart_div0[5]), 
        .Y(n25483) );
  sky130_fd_sc_hd__o22ai_1 U30706 ( .A1(n25494), .A2(n28310), .B1(n25485), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U30707 ( .A1(n25494), .A2(n28313), .B1(n25486), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U30708 ( .A1(n25494), .A2(n28316), .B1(n25487), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U30709 ( .A1(n25494), .A2(n26760), .B1(n25488), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U30710 ( .A1(n25494), .A2(n28064), .B1(n25489), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U30711 ( .A1(n25494), .A2(n27575), .B1(n25490), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U30712 ( .A1(n25494), .A2(n28553), .B1(n25491), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U30713 ( .A1(n25494), .A2(n29082), .B1(n25492), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U30714 ( .A1(n25494), .A2(n29076), .B1(n25493), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__a21oi_1 U30715 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[63]), .B1(n28326), .Y(n25502) );
  sky130_fd_sc_hd__nand2_1 U30716 ( .A(n28318), .B(
        j202_soc_core_intc_core_00_rg_ie[29]), .Y(n25497) );
  sky130_fd_sc_hd__a22oi_1 U30717 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[55]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[39]), .Y(n25496) );
  sky130_fd_sc_hd__nand2_1 U30718 ( .A(n28331), .B(
        j202_soc_core_intc_core_00_rg_itgt[47]), .Y(n25495) );
  sky130_fd_sc_hd__nand3_1 U30719 ( .A(n25497), .B(n25496), .C(n25495), .Y(
        n25498) );
  sky130_fd_sc_hd__a21oi_1 U30720 ( .A1(j202_soc_core_intc_core_00_rg_ipr[61]), 
        .A2(n28330), .B1(n25498), .Y(n25501) );
  sky130_fd_sc_hd__a22oi_1 U30721 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[29]), .B1(n28329), .B2(
        j202_soc_core_intc_core_00_rg_ipr[125]), .Y(n25500) );
  sky130_fd_sc_hd__nand2_1 U30722 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[93]), .Y(n25499) );
  sky130_fd_sc_hd__nand4_1 U30723 ( .A(n25502), .B(n25501), .C(n25500), .D(
        n25499), .Y(j202_soc_core_ahb2apb_01_N157) );
  sky130_fd_sc_hd__nor2_1 U30724 ( .A(n28895), .B(n25503), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N324) );
  sky130_fd_sc_hd__mux2i_1 U30725 ( .A0(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[1]), .A1(io_in[12]), .S(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n28193) );
  sky130_fd_sc_hd__nor2_1 U30726 ( .A(n28895), .B(n28193), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N325) );
  sky130_fd_sc_hd__mux2i_1 U30727 ( .A0(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[2]), .A1(io_in[13]), .S(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n27695) );
  sky130_fd_sc_hd__nor2_1 U30728 ( .A(n28895), .B(n27695), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N326) );
  sky130_fd_sc_hd__nor2_1 U30729 ( .A(n28895), .B(n25505), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N327) );
  sky130_fd_sc_hd__nor2_1 U30730 ( .A(n28895), .B(n25507), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N328) );
  sky130_fd_sc_hd__nor2_1 U30731 ( .A(n28895), .B(n25509), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N329) );
  sky130_fd_sc_hd__nor2_1 U30732 ( .A(n28895), .B(n25511), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N330) );
  sky130_fd_sc_hd__nor2_1 U30733 ( .A(n28895), .B(n25513), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N331) );
  sky130_fd_sc_hd__nor2_1 U30734 ( .A(n28895), .B(n25515), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N332) );
  sky130_fd_sc_hd__nor2_1 U30735 ( .A(n28895), .B(n25517), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N333) );
  sky130_fd_sc_hd__nor2_1 U30736 ( .A(n28895), .B(n25519), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N334) );
  sky130_fd_sc_hd__nor2_1 U30737 ( .A(n28895), .B(n25521), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N335) );
  sky130_fd_sc_hd__nor2_1 U30738 ( .A(n28895), .B(n25523), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N336) );
  sky130_fd_sc_hd__nor2_1 U30739 ( .A(n28895), .B(n25525), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N337) );
  sky130_fd_sc_hd__nor2_1 U30740 ( .A(n28895), .B(n25527), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N338) );
  sky130_fd_sc_hd__nor2_1 U30741 ( .A(n28895), .B(n25529), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N339) );
  sky130_fd_sc_hd__nor2_1 U30742 ( .A(n28895), .B(n25531), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N340) );
  sky130_fd_sc_hd__nor2_1 U30743 ( .A(n28895), .B(n25533), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N341) );
  sky130_fd_sc_hd__nor2_1 U30744 ( .A(n28895), .B(n25535), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N342) );
  sky130_fd_sc_hd__nor2_1 U30745 ( .A(n28895), .B(n25537), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N343) );
  sky130_fd_sc_hd__nor2_1 U30746 ( .A(n28895), .B(n25539), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N344) );
  sky130_fd_sc_hd__nor2_1 U30747 ( .A(n28895), .B(n25541), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N345) );
  sky130_fd_sc_hd__nor2_1 U30748 ( .A(n28895), .B(n25543), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N346) );
  sky130_fd_sc_hd__nor2_1 U30749 ( .A(n28895), .B(n25545), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N347) );
  sky130_fd_sc_hd__nor2_1 U30750 ( .A(n28895), .B(n25547), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N348) );
  sky130_fd_sc_hd__nor2_1 U30751 ( .A(n28895), .B(n25549), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N349) );
  sky130_fd_sc_hd__nor2_1 U30752 ( .A(n28895), .B(n25551), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N350) );
  sky130_fd_sc_hd__nor2_1 U30753 ( .A(n28895), .B(n25553), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N351) );
  sky130_fd_sc_hd__nand2_1 U30754 ( .A(n27431), .B(n25554), .Y(n27610) );
  sky130_fd_sc_hd__nand2_1 U30755 ( .A(n27610), .B(n27613), .Y(n28025) );
  sky130_fd_sc_hd__a22o_1 U30756 ( .A1(n28026), .A2(
        j202_soc_core_wbqspiflash_00_spi_out[29]), .B1(n28025), .B2(
        j202_soc_core_wbqspiflash_00_spi_busy), .X(
        j202_soc_core_wbqspiflash_00_N696) );
  sky130_fd_sc_hd__nand4_1 U30757 ( .A(n25561), .B(n25560), .C(n25559), .D(
        n25558), .Y(n25562) );
  sky130_fd_sc_hd__nand2_1 U30758 ( .A(n25562), .B(n27860), .Y(n25568) );
  sky130_fd_sc_hd__nand2_1 U30759 ( .A(n25564), .B(n25563), .Y(n25566) );
  sky130_fd_sc_hd__o22ai_1 U30760 ( .A1(n13047), .A2(n27775), .B1(n27774), 
        .B2(n25594), .Y(n25565) );
  sky130_fd_sc_hd__a21oi_1 U30761 ( .A1(n25566), .A2(n27860), .B1(n25565), .Y(
        n25567) );
  sky130_fd_sc_hd__nand2_1 U30762 ( .A(n25568), .B(n25567), .Y(
        j202_soc_core_j22_cpu_rf_N3368) );
  sky130_fd_sc_hd__nand2_1 U30763 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[21]), .Y(n25569) );
  sky130_fd_sc_hd__o21ai_1 U30764 ( .A1(n25570), .A2(n28545), .B1(n25569), .Y(
        n64) );
  sky130_fd_sc_hd__nand2_1 U30765 ( .A(n27624), .B(j202_soc_core_uart_div1[5]), 
        .Y(n25571) );
  sky130_fd_sc_hd__o21ai_1 U30766 ( .A1(n25572), .A2(n27624), .B1(n25571), .Y(
        n95) );
  sky130_fd_sc_hd__o22ai_1 U30767 ( .A1(n25582), .A2(n28310), .B1(n25573), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30768 ( .A1(n25582), .A2(n28313), .B1(n25574), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30769 ( .A1(n25582), .A2(n28316), .B1(n25575), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30770 ( .A1(n25582), .A2(n26760), .B1(n25576), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30771 ( .A1(n25582), .A2(n28064), .B1(n25577), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30772 ( .A1(n25582), .A2(n27575), .B1(n25578), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30773 ( .A1(n25582), .A2(n28553), .B1(n25579), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30774 ( .A1(n25582), .A2(n29082), .B1(n25580), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30775 ( .A1(n25582), .A2(n29076), .B1(n25581), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__a21oi_1 U30776 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[61]), .B1(n28326), .Y(n25590) );
  sky130_fd_sc_hd__nand2_1 U30777 ( .A(n28236), .B(
        j202_soc_core_intc_core_00_rg_ie[21]), .Y(n25585) );
  sky130_fd_sc_hd__a22oi_1 U30778 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[53]), .B1(n27398), .B2(
        j202_soc_core_intc_core_00_rg_itgt[37]), .Y(n25584) );
  sky130_fd_sc_hd__nand2_1 U30779 ( .A(n28331), .B(
        j202_soc_core_intc_core_00_rg_itgt[45]), .Y(n25583) );
  sky130_fd_sc_hd__nand3_1 U30780 ( .A(n25585), .B(n25584), .C(n25583), .Y(
        n25586) );
  sky130_fd_sc_hd__a21oi_1 U30781 ( .A1(j202_soc_core_intc_core_00_rg_ipr[53]), 
        .A2(n28330), .B1(n25586), .Y(n25589) );
  sky130_fd_sc_hd__a22oi_1 U30782 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[21]), .B1(n28329), .B2(
        j202_soc_core_intc_core_00_rg_ipr[117]), .Y(n25588) );
  sky130_fd_sc_hd__nand2_1 U30783 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[85]), .Y(n25587) );
  sky130_fd_sc_hd__nand4_1 U30784 ( .A(n25590), .B(n25589), .C(n25588), .D(
        n25587), .Y(j202_soc_core_ahb2apb_01_N149) );
  sky130_fd_sc_hd__nor2_1 U30785 ( .A(j202_soc_core_rst), .B(n25591), .Y(
        j202_soc_core_wbqspiflash_00_N718) );
  sky130_fd_sc_hd__a22o_1 U30786 ( .A1(n28026), .A2(
        j202_soc_core_wbqspiflash_00_spi_out[21]), .B1(n28025), .B2(
        j202_soc_core_wbqspiflash_00_erased_sector[7]), .X(
        j202_soc_core_wbqspiflash_00_N688) );
  sky130_fd_sc_hd__a22oi_1 U30787 ( .A1(n26329), .A2(n27764), .B1(n12222), 
        .B2(n28425), .Y(n25592) );
  sky130_fd_sc_hd__nand2_1 U30788 ( .A(n24292), .B(n25592), .Y(
        j202_soc_core_j22_cpu_ml_N325) );
  sky130_fd_sc_hd__o22ai_1 U30789 ( .A1(n25980), .A2(n25594), .B1(n27835), 
        .B2(n12266), .Y(j202_soc_core_j22_cpu_rf_N2813) );
  sky130_fd_sc_hd__nand2_1 U30790 ( .A(n25626), .B(n27772), .Y(n25598) );
  sky130_fd_sc_hd__o22ai_1 U30791 ( .A1(n25599), .A2(n27775), .B1(n27774), 
        .B2(n25632), .Y(n25596) );
  sky130_fd_sc_hd__a21oi_1 U30792 ( .A1(n30084), .A2(n27860), .B1(n25596), .Y(
        n25597) );
  sky130_fd_sc_hd__nand2_1 U30793 ( .A(n25598), .B(n25597), .Y(
        j202_soc_core_j22_cpu_rf_N3369) );
  sky130_fd_sc_hd__nand2_1 U30794 ( .A(n12396), .B(n25724), .Y(n25603) );
  sky130_fd_sc_hd__o22ai_1 U30795 ( .A1(n26277), .A2(n27850), .B1(n25599), 
        .B2(n27848), .Y(n25600) );
  sky130_fd_sc_hd__a21oi_1 U30796 ( .A1(n25601), .A2(n26068), .B1(n25600), .Y(
        n25602) );
  sky130_fd_sc_hd__nand2_1 U30797 ( .A(n25603), .B(n25602), .Y(
        j202_soc_core_j22_cpu_rf_N320) );
  sky130_fd_sc_hd__o22ai_1 U30798 ( .A1(n25632), .A2(n27859), .B1(n27858), 
        .B2(n25604), .Y(j202_soc_core_j22_cpu_rf_N3334) );
  sky130_fd_sc_hd__nand2_1 U30799 ( .A(n27624), .B(j202_soc_core_uart_div1[6]), 
        .Y(n25605) );
  sky130_fd_sc_hd__o21ai_1 U30800 ( .A1(n26834), .A2(n27624), .B1(n25605), .Y(
        n96) );
  sky130_fd_sc_hd__o22ai_1 U30801 ( .A1(n25614), .A2(n28310), .B1(n25606), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U30802 ( .A1(n25614), .A2(n28313), .B1(n25607), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U30803 ( .A1(n25614), .A2(n28316), .B1(n25608), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U30804 ( .A1(n25614), .A2(n26760), .B1(n12697), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U30805 ( .A1(n25614), .A2(n28064), .B1(n25609), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U30806 ( .A1(n25614), .A2(n27575), .B1(n25610), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U30807 ( .A1(n25614), .A2(n28553), .B1(n25611), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U30808 ( .A1(n25614), .A2(n29082), .B1(n25612), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U30809 ( .A1(n25614), .A2(n29076), .B1(n25613), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__a21oi_1 U30810 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[93]), .B1(n28326), .Y(n25622) );
  sky130_fd_sc_hd__nand2_1 U30811 ( .A(n28236), .B(
        j202_soc_core_intc_core_00_rg_ie[22]), .Y(n25617) );
  sky130_fd_sc_hd__a22oi_1 U30812 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[85]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[69]), .Y(n25616) );
  sky130_fd_sc_hd__nand2_1 U30813 ( .A(n28331), .B(
        j202_soc_core_intc_core_00_rg_itgt[77]), .Y(n25615) );
  sky130_fd_sc_hd__nand3_1 U30814 ( .A(n25617), .B(n25616), .C(n25615), .Y(
        n25618) );
  sky130_fd_sc_hd__a21oi_1 U30815 ( .A1(j202_soc_core_intc_core_00_rg_ipr[54]), 
        .A2(n28330), .B1(n25618), .Y(n25621) );
  sky130_fd_sc_hd__a22oi_1 U30816 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[22]), .B1(n28329), .B2(
        j202_soc_core_intc_core_00_rg_ipr[118]), .Y(n25620) );
  sky130_fd_sc_hd__nand2_1 U30817 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[86]), .Y(n25619) );
  sky130_fd_sc_hd__nand4_1 U30818 ( .A(n25622), .B(n25621), .C(n25620), .D(
        n25619), .Y(j202_soc_core_ahb2apb_01_N150) );
  sky130_fd_sc_hd__nand2_1 U30819 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[22]), .Y(n25623) );
  sky130_fd_sc_hd__o21ai_1 U30820 ( .A1(n25624), .A2(n28545), .B1(n25623), .Y(
        n65) );
  sky130_fd_sc_hd__a22oi_1 U30821 ( .A1(n25642), .A2(n27764), .B1(n12396), 
        .B2(n28425), .Y(n25625) );
  sky130_fd_sc_hd__nand2_1 U30822 ( .A(n24292), .B(n25625), .Y(
        j202_soc_core_j22_cpu_ml_N326) );
  sky130_fd_sc_hd__nand2_1 U30823 ( .A(n12203), .B(n25626), .Y(n25629) );
  sky130_fd_sc_hd__nand2_1 U30824 ( .A(n28056), .B(n25627), .Y(n25628) );
  sky130_fd_sc_hd__nand3_1 U30825 ( .A(n25629), .B(n27119), .C(n25628), .Y(
        n29842) );
  sky130_fd_sc_hd__nand2_1 U30826 ( .A(n25630), .B(n24832), .Y(n25631) );
  sky130_fd_sc_hd__nor2_1 U30828 ( .A(n26196), .B(n12351), .Y(n25634) );
  sky130_fd_sc_hd__nand2_1 U30830 ( .A(n25665), .B(n27152), .Y(n25659) );
  sky130_fd_sc_hd__nand2_1 U30831 ( .A(n25634), .B(n26916), .Y(n25635) );
  sky130_fd_sc_hd__o211ai_1 U30832 ( .A1(n28506), .A2(n26939), .B1(n26919), 
        .C1(n25635), .Y(n25656) );
  sky130_fd_sc_hd__o211ai_1 U30834 ( .A1(n11123), .A2(n26331), .B1(n25638), 
        .C1(n25637), .Y(n25639) );
  sky130_fd_sc_hd__nand2_1 U30835 ( .A(n25660), .B(n25639), .Y(n25654) );
  sky130_fd_sc_hd__o22ai_1 U30836 ( .A1(n26318), .A2(n27799), .B1(n27026), 
        .B2(n26943), .Y(n25647) );
  sky130_fd_sc_hd__o22ai_1 U30837 ( .A1(n27027), .A2(n27795), .B1(n27365), 
        .B2(n27797), .Y(n25646) );
  sky130_fd_sc_hd__xor2_1 U30838 ( .A(n26331), .B(n28506), .X(n26229) );
  sky130_fd_sc_hd__nand2_1 U30839 ( .A(n27808), .B(n27115), .Y(n25644) );
  sky130_fd_sc_hd__o22ai_1 U30840 ( .A1(n25640), .A2(n26926), .B1(n26280), 
        .B2(n27803), .Y(n25641) );
  sky130_fd_sc_hd__a21oi_1 U30841 ( .A1(n27810), .A2(n25642), .B1(n25641), .Y(
        n25643) );
  sky130_fd_sc_hd__o211ai_1 U30842 ( .A1(n26229), .A2(n25872), .B1(n25644), 
        .C1(n25643), .Y(n25645) );
  sky130_fd_sc_hd__nor3_1 U30843 ( .A(n25647), .B(n25646), .C(n25645), .Y(
        n25651) );
  sky130_fd_sc_hd__nand2_1 U30844 ( .A(n25648), .B(n28509), .Y(n25650) );
  sky130_fd_sc_hd__mux2_2 U30845 ( .A0(n27817), .A1(n27793), .S(n28506), .X(
        n25649) );
  sky130_fd_sc_hd__nand4_1 U30846 ( .A(n25651), .B(n25650), .C(n27814), .D(
        n25649), .Y(n25652) );
  sky130_fd_sc_hd__a21oi_1 U30847 ( .A1(n25674), .A2(n27789), .B1(n25652), .Y(
        n25653) );
  sky130_fd_sc_hd__nand2_1 U30848 ( .A(n25654), .B(n25653), .Y(n25655) );
  sky130_fd_sc_hd__a21oi_1 U30849 ( .A1(n25656), .A2(n26331), .B1(n25655), .Y(
        n25657) );
  sky130_fd_sc_hd__o22ai_1 U30850 ( .A1(n25977), .A2(n28505), .B1(n28061), 
        .B2(n27385), .Y(j202_soc_core_j22_cpu_rf_N2885) );
  sky130_fd_sc_hd__o22ai_1 U30851 ( .A1(n25978), .A2(n28505), .B1(n27834), 
        .B2(n27385), .Y(j202_soc_core_j22_cpu_rf_N2959) );
  sky130_fd_sc_hd__o22ai_1 U30852 ( .A1(n25979), .A2(n28505), .B1(n28112), 
        .B2(n27385), .Y(j202_soc_core_j22_cpu_rf_N3218) );
  sky130_fd_sc_hd__o22ai_1 U30853 ( .A1(n25980), .A2(n28505), .B1(n27835), 
        .B2(n27385), .Y(j202_soc_core_j22_cpu_rf_N2811) );
  sky130_fd_sc_hd__o22ai_1 U30854 ( .A1(n25981), .A2(n28505), .B1(n27836), 
        .B2(n27385), .Y(j202_soc_core_j22_cpu_rf_N3181) );
  sky130_fd_sc_hd__o22ai_1 U30855 ( .A1(n25982), .A2(n28505), .B1(n27837), 
        .B2(n27385), .Y(j202_soc_core_j22_cpu_rf_N3033) );
  sky130_fd_sc_hd__o22ai_1 U30856 ( .A1(n25983), .A2(n28505), .B1(n27838), 
        .B2(n12258), .Y(j202_soc_core_j22_cpu_rf_N3070) );
  sky130_fd_sc_hd__o22ai_1 U30857 ( .A1(n25984), .A2(n28505), .B1(n27840), 
        .B2(n27385), .Y(j202_soc_core_j22_cpu_rf_N2737) );
  sky130_fd_sc_hd__o22ai_1 U30858 ( .A1(n27841), .A2(n28505), .B1(n24712), 
        .B2(n12258), .Y(j202_soc_core_j22_cpu_rf_N3255) );
  sky130_fd_sc_hd__o22ai_1 U30859 ( .A1(n25985), .A2(n28505), .B1(n27842), 
        .B2(n12258), .Y(j202_soc_core_j22_cpu_rf_N3107) );
  sky130_fd_sc_hd__o22ai_1 U30860 ( .A1(n25986), .A2(n28505), .B1(n27843), 
        .B2(n12258), .Y(j202_soc_core_j22_cpu_rf_N2996) );
  sky130_fd_sc_hd__o22ai_1 U30861 ( .A1(n25987), .A2(n28505), .B1(n27844), 
        .B2(n27385), .Y(j202_soc_core_j22_cpu_rf_N3144) );
  sky130_fd_sc_hd__o22ai_1 U30862 ( .A1(n25988), .A2(n28505), .B1(n27845), 
        .B2(n12258), .Y(j202_soc_core_j22_cpu_rf_N2848) );
  sky130_fd_sc_hd__o22ai_1 U30863 ( .A1(n25989), .A2(n28505), .B1(n27846), 
        .B2(n12258), .Y(j202_soc_core_j22_cpu_rf_N2774) );
  sky130_fd_sc_hd__o22ai_1 U30864 ( .A1(n25964), .A2(n28505), .B1(n27847), 
        .B2(n12258), .Y(j202_soc_core_j22_cpu_rf_N2700) );
  sky130_fd_sc_hd__nand2_1 U30865 ( .A(n25662), .B(n24832), .Y(n25661) );
  sky130_fd_sc_hd__o21ai_0 U30866 ( .A1(n24832), .A2(n28505), .B1(n25661), .Y(
        j202_soc_core_j22_cpu_rf_N3292) );
  sky130_fd_sc_hd__o22ai_1 U30867 ( .A1(n28505), .A2(n27859), .B1(n27858), 
        .B2(n12258), .Y(j202_soc_core_j22_cpu_rf_N3331) );
  sky130_fd_sc_hd__a21oi_1 U30868 ( .A1(n27768), .A2(n11474), .B1(n27766), .Y(
        n25663) );
  sky130_fd_sc_hd__o21ai_1 U30869 ( .A1(n25664), .A2(n27770), .B1(n25663), .Y(
        j202_soc_core_j22_cpu_ml_maclj[20]) );
  sky130_fd_sc_hd__nand2_1 U30870 ( .A(n25665), .B(n27772), .Y(n25671) );
  sky130_fd_sc_hd__o22ai_1 U30871 ( .A1(n25672), .A2(n27775), .B1(n27774), 
        .B2(n28505), .Y(n25669) );
  sky130_fd_sc_hd__nor2_1 U30872 ( .A(n27648), .B(n25667), .Y(n25668) );
  sky130_fd_sc_hd__nor2_1 U30873 ( .A(n25669), .B(n25668), .Y(n25670) );
  sky130_fd_sc_hd__nand2_1 U30874 ( .A(n25671), .B(n25670), .Y(
        j202_soc_core_j22_cpu_rf_N3367) );
  sky130_fd_sc_hd__o22ai_1 U30875 ( .A1(n28506), .A2(n27850), .B1(n25672), 
        .B2(n27848), .Y(n25673) );
  sky130_fd_sc_hd__a21oi_1 U30876 ( .A1(n25674), .A2(n26068), .B1(n25673), .Y(
        n25675) );
  sky130_fd_sc_hd__o21ai_0 U30877 ( .A1(n27855), .A2(n28505), .B1(n25675), .Y(
        j202_soc_core_j22_cpu_rf_N318) );
  sky130_fd_sc_hd__a21oi_1 U30878 ( .A1(n25677), .A2(n27052), .B1(n26926), .Y(
        n25704) );
  sky130_fd_sc_hd__nand2_1 U30879 ( .A(n25678), .B(n25704), .Y(n25707) );
  sky130_fd_sc_hd__nand3_1 U30880 ( .A(n23485), .B(n25679), .C(n25704), .Y(
        n25706) );
  sky130_fd_sc_hd__nand3_1 U30881 ( .A(n25681), .B(n27828), .C(n25680), .Y(
        n25703) );
  sky130_fd_sc_hd__a21oi_1 U30882 ( .A1(n25697), .A2(n27785), .B1(n25682), .Y(
        n25701) );
  sky130_fd_sc_hd__o22ai_1 U30883 ( .A1(n27800), .A2(n27795), .B1(n11190), 
        .B2(n27797), .Y(n25691) );
  sky130_fd_sc_hd__o22ai_1 U30884 ( .A1(n27025), .A2(n27799), .B1(n27383), 
        .B2(n27803), .Y(n25690) );
  sky130_fd_sc_hd__a21oi_1 U30885 ( .A1(n25692), .A2(n27791), .B1(n27790), .Y(
        n25683) );
  sky130_fd_sc_hd__o22ai_1 U30886 ( .A1(n27793), .A2(n25692), .B1(n27027), 
        .B2(n25683), .Y(n25684) );
  sky130_fd_sc_hd__a21oi_1 U30887 ( .A1(n25685), .A2(n27042), .B1(n25684), .Y(
        n25687) );
  sky130_fd_sc_hd__xnor2_1 U30888 ( .A(n25692), .B(n25697), .Y(n26223) );
  sky130_fd_sc_hd__a2bb2oi_1 U30889 ( .B1(n26051), .B2(n27808), .A1_N(n25872), 
        .A2_N(n26223), .Y(n25686) );
  sky130_fd_sc_hd__o211ai_1 U30890 ( .A1(n26280), .A2(n25688), .B1(n25687), 
        .C1(n25686), .Y(n25689) );
  sky130_fd_sc_hd__nor3_1 U30891 ( .A(n25691), .B(n25690), .C(n25689), .Y(
        n25694) );
  sky130_fd_sc_hd__o22a_1 U30892 ( .A1(n28513), .A2(n27817), .B1(n26135), .B2(
        n27815), .X(n25693) );
  sky130_fd_sc_hd__nand3_1 U30893 ( .A(n25694), .B(n25693), .C(n27814), .Y(
        n25695) );
  sky130_fd_sc_hd__a21oi_1 U30894 ( .A1(n25715), .A2(n27789), .B1(n25695), .Y(
        n25700) );
  sky130_fd_sc_hd__xnor2_1 U30895 ( .A(n25697), .B(n25696), .Y(n25698) );
  sky130_fd_sc_hd__nand2_1 U30896 ( .A(n25698), .B(n27786), .Y(n25699) );
  sky130_fd_sc_hd__a21oi_2 U30897 ( .A1(n25704), .A2(n25703), .B1(n25702), .Y(
        n25705) );
  sky130_fd_sc_hd__nand3_2 U30898 ( .A(n25707), .B(n25706), .C(n25705), .Y(
        n25709) );
  sky130_fd_sc_hd__nand2_1 U30899 ( .A(n25709), .B(n24832), .Y(n25708) );
  sky130_fd_sc_hd__o21ai_0 U30900 ( .A1(n24832), .A2(n25720), .B1(n25708), .Y(
        j202_soc_core_j22_cpu_rf_N3291) );
  sky130_fd_sc_hd__o22ai_1 U30902 ( .A1(n25720), .A2(n27859), .B1(n27858), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N3330) );
  sky130_fd_sc_hd__o22ai_1 U30903 ( .A1(n27841), .A2(n25720), .B1(n24712), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N3254) );
  sky130_fd_sc_hd__o22ai_1 U30904 ( .A1(n25964), .A2(n25720), .B1(n27847), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N2699) );
  sky130_fd_sc_hd__nand2_1 U30905 ( .A(n25709), .B(n27860), .Y(n25712) );
  sky130_fd_sc_hd__o22a_1 U30906 ( .A1(n25713), .A2(n27775), .B1(n27774), .B2(
        n25720), .X(n25711) );
  sky130_fd_sc_hd__nand2_1 U30907 ( .A(n25712), .B(n25711), .Y(
        j202_soc_core_j22_cpu_rf_N3366) );
  sky130_fd_sc_hd__o22ai_1 U30908 ( .A1(n28513), .A2(n27850), .B1(n25713), 
        .B2(n27848), .Y(n25714) );
  sky130_fd_sc_hd__a21oi_1 U30909 ( .A1(n25715), .A2(n26068), .B1(n25714), .Y(
        n25716) );
  sky130_fd_sc_hd__o21ai_0 U30910 ( .A1(n27855), .A2(n25720), .B1(n25716), .Y(
        j202_soc_core_j22_cpu_rf_N317) );
  sky130_fd_sc_hd__o22ai_1 U30911 ( .A1(n25977), .A2(n25720), .B1(n28061), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N2884) );
  sky130_fd_sc_hd__o22ai_1 U30912 ( .A1(n25978), .A2(n25720), .B1(n27834), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N2958) );
  sky130_fd_sc_hd__o22ai_1 U30913 ( .A1(n25979), .A2(n25720), .B1(n28112), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N3217) );
  sky130_fd_sc_hd__o22ai_1 U30914 ( .A1(n25980), .A2(n25720), .B1(n27835), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N2810) );
  sky130_fd_sc_hd__o22ai_1 U30915 ( .A1(n25981), .A2(n25720), .B1(n27836), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N3180) );
  sky130_fd_sc_hd__o22ai_1 U30916 ( .A1(n25982), .A2(n25720), .B1(n27837), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N3032) );
  sky130_fd_sc_hd__o22ai_1 U30917 ( .A1(n25983), .A2(n25720), .B1(n27838), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N3069) );
  sky130_fd_sc_hd__o22ai_1 U30918 ( .A1(n26894), .A2(n25720), .B1(n27839), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N2921) );
  sky130_fd_sc_hd__o22ai_1 U30919 ( .A1(n25984), .A2(n25720), .B1(n27840), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N2736) );
  sky130_fd_sc_hd__o22ai_1 U30920 ( .A1(n25985), .A2(n25720), .B1(n27842), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N3106) );
  sky130_fd_sc_hd__o22ai_1 U30921 ( .A1(n25986), .A2(n25720), .B1(n27843), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N2995) );
  sky130_fd_sc_hd__o22ai_1 U30922 ( .A1(n25987), .A2(n25720), .B1(n27844), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N3143) );
  sky130_fd_sc_hd__o22ai_1 U30923 ( .A1(n25989), .A2(n25720), .B1(n27846), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N2773) );
  sky130_fd_sc_hd__nor2_1 U30924 ( .A(n29088), .B(n25717), .Y(
        j202_soc_core_wbqspiflash_00_N716) );
  sky130_fd_sc_hd__a22o_1 U30925 ( .A1(n28026), .A2(
        j202_soc_core_wbqspiflash_00_spi_out[19]), .B1(n28025), .B2(
        j202_soc_core_wbqspiflash_00_erased_sector[5]), .X(
        j202_soc_core_wbqspiflash_00_N686) );
  sky130_fd_sc_hd__o21ai_1 U30926 ( .A1(n25718), .A2(n25779), .B1(n27119), .Y(
        j202_soc_core_j22_cpu_ml_machj[19]) );
  sky130_fd_sc_hd__o22ai_1 U30927 ( .A1(n25988), .A2(n25720), .B1(n27845), 
        .B2(n25719), .Y(j202_soc_core_j22_cpu_rf_N2847) );
  sky130_fd_sc_hd__a22oi_1 U30928 ( .A1(n27862), .A2(n25725), .B1(n28525), 
        .B2(n27861), .Y(n25721) );
  sky130_fd_sc_hd__nand2_1 U30931 ( .A(n28525), .B(n25724), .Y(n25730) );
  sky130_fd_sc_hd__o22ai_1 U30932 ( .A1(n26285), .A2(n27850), .B1(n25726), 
        .B2(n27848), .Y(n25727) );
  sky130_fd_sc_hd__a21oi_1 U30933 ( .A1(n25728), .A2(n26068), .B1(n25727), .Y(
        n25729) );
  sky130_fd_sc_hd__nand2_1 U30934 ( .A(n25730), .B(n25729), .Y(
        j202_soc_core_j22_cpu_rf_N315) );
  sky130_fd_sc_hd__nand2_1 U30935 ( .A(n27624), .B(j202_soc_core_uart_div1[1]), 
        .Y(n25731) );
  sky130_fd_sc_hd__o22ai_1 U30937 ( .A1(n29149), .A2(n28064), .B1(n25741), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U30938 ( .A1(n29073), .A2(n25736), .B1(n28366), 
        .B2(n29070), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N4) );
  sky130_fd_sc_hd__nand3_1 U30939 ( .A(j202_soc_core_cmt_core_00_cmf1), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[6]), .C(n29830), .Y(
        n25737) );
  sky130_fd_sc_hd__nor3_1 U30940 ( .A(j202_soc_core_intc_core_00_rg_irqc[17]), 
        .B(n29088), .C(n25733), .Y(n25739) );
  sky130_fd_sc_hd__nand2_1 U30941 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .B(n27350), .Y(n25734) );
  sky130_fd_sc_hd__nor2_1 U30942 ( .A(n25735), .B(n25734), .Y(n27704) );
  sky130_fd_sc_hd__nand2_1 U30943 ( .A(n27704), .B(n25736), .Y(n25738) );
  sky130_fd_sc_hd__a2bb2oi_1 U30944 ( .B1(n25739), .B2(n25738), .A1_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[17]), 
        .A2_N(n25737), .Y(n25740) );
  sky130_fd_sc_hd__nor2_1 U30945 ( .A(n25741), .B(n25740), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N20) );
  sky130_fd_sc_hd__o22ai_1 U30946 ( .A1(n29149), .A2(n28310), .B1(n25742), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U30947 ( .A1(n29149), .A2(n28313), .B1(n25743), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U30948 ( .A1(n29149), .A2(n28316), .B1(n25744), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U30949 ( .A1(n29149), .A2(n26760), .B1(n25745), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U30950 ( .A1(n29149), .A2(n27575), .B1(n25746), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U30951 ( .A1(n29149), .A2(n28553), .B1(n25747), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U30952 ( .A1(n29149), .A2(n29082), .B1(n25748), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U30953 ( .A1(n29149), .A2(n29076), .B1(n25749), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__a22oi_1 U30954 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[17]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[17]), .Y(n25751) );
  sky130_fd_sc_hd__a22oi_1 U30955 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[52]), .B1(n27398), .B2(
        j202_soc_core_intc_core_00_rg_itgt[36]), .Y(n25750) );
  sky130_fd_sc_hd__nand3_1 U30956 ( .A(n25751), .B(n28238), .C(n25750), .Y(
        n25752) );
  sky130_fd_sc_hd__a21oi_1 U30957 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[113]), .B1(n25752), .Y(n25756) );
  sky130_fd_sc_hd__a22oi_1 U30958 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[60]), .B1(n28331), .B2(
        j202_soc_core_intc_core_00_rg_itgt[44]), .Y(n25755) );
  sky130_fd_sc_hd__a22oi_1 U30959 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[17]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[49]), .B2(n28330), .Y(n25754) );
  sky130_fd_sc_hd__nand2_1 U30960 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[81]), .Y(n25753) );
  sky130_fd_sc_hd__nand4_1 U30961 ( .A(n25756), .B(n25755), .C(n25754), .D(
        n25753), .Y(j202_soc_core_ahb2apb_01_N145) );
  sky130_fd_sc_hd__nor2_1 U30962 ( .A(n29088), .B(n25757), .Y(
        j202_soc_core_wbqspiflash_00_N714) );
  sky130_fd_sc_hd__a22o_1 U30963 ( .A1(n28026), .A2(
        j202_soc_core_wbqspiflash_00_spi_out[17]), .B1(n28025), .B2(
        j202_soc_core_wbqspiflash_00_erased_sector[3]), .X(
        j202_soc_core_wbqspiflash_00_N684) );
  sky130_fd_sc_hd__nand2_1 U30964 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[17]), .Y(n25758) );
  sky130_fd_sc_hd__o21ai_1 U30965 ( .A1(n25759), .A2(n28545), .B1(n25758), .Y(
        n34) );
  sky130_fd_sc_hd__a22oi_1 U30966 ( .A1(n26051), .A2(n27764), .B1(n28525), 
        .B2(n28425), .Y(n25760) );
  sky130_fd_sc_hd__nand2_1 U30967 ( .A(n24292), .B(n25760), .Y(
        j202_soc_core_j22_cpu_ml_N320) );
  sky130_fd_sc_hd__a21oi_1 U30968 ( .A1(n25761), .A2(n28056), .B1(n25776), .Y(
        n25762) );
  sky130_fd_sc_hd__o21ai_0 U30969 ( .A1(n25763), .A2(n25779), .B1(n25762), .Y(
        n29832) );
  sky130_fd_sc_hd__o22ai_1 U30970 ( .A1(n26894), .A2(n25765), .B1(n27839), 
        .B2(n12057), .Y(j202_soc_core_j22_cpu_rf_N2919) );
  sky130_fd_sc_hd__o22ai_1 U30971 ( .A1(n26894), .A2(n28477), .B1(n27839), 
        .B2(n25766), .Y(j202_soc_core_j22_cpu_rf_N2928) );
  sky130_fd_sc_hd__a22oi_1 U30972 ( .A1(n26416), .A2(n27764), .B1(n12260), 
        .B2(n28425), .Y(n25767) );
  sky130_fd_sc_hd__nand2_1 U30973 ( .A(n24292), .B(n25767), .Y(
        j202_soc_core_j22_cpu_ml_N335) );
  sky130_fd_sc_hd__a22oi_1 U30975 ( .A1(n25777), .A2(n27768), .B1(n25772), 
        .B2(n25771), .Y(n25773) );
  sky130_fd_sc_hd__o21ai_1 U30976 ( .A1(n25774), .A2(n27770), .B1(n25773), .Y(
        j202_soc_core_j22_cpu_ml_maclj[31]) );
  sky130_fd_sc_hd__a21oi_1 U30977 ( .A1(n25777), .A2(n28056), .B1(n25776), .Y(
        n25778) );
  sky130_fd_sc_hd__o21ai_1 U30978 ( .A1(n25780), .A2(n25779), .B1(n25778), .Y(
        n29834) );
  sky130_fd_sc_hd__nand2_1 U30979 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[13]), .Y(n25781) );
  sky130_fd_sc_hd__o21ai_1 U30980 ( .A1(n25782), .A2(n28545), .B1(n25781), .Y(
        n59) );
  sky130_fd_sc_hd__o22ai_1 U30981 ( .A1(n29145), .A2(n28064), .B1(n25784), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__nand2_1 U30982 ( .A(n26713), .B(n26748), .Y(n25783) );
  sky130_fd_sc_hd__nand4b_1 U30983 ( .A_N(
        j202_soc_core_intc_core_00_rg_irqc[13]), .B(n25783), .C(
        j202_soc_core_intc_core_00_in_intreq[13]), .D(n28914), .Y(n25786) );
  sky130_fd_sc_hd__nand2b_1 U30984 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[13]), 
        .B(n29566), .Y(n25785) );
  sky130_fd_sc_hd__a21oi_1 U30985 ( .A1(n25786), .A2(n25785), .B1(n25784), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N16) );
  sky130_fd_sc_hd__o22ai_1 U30986 ( .A1(n29145), .A2(n28310), .B1(n25787), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U30987 ( .A1(n29145), .A2(n28313), .B1(n25788), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U30988 ( .A1(n29145), .A2(n28316), .B1(n25789), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U30989 ( .A1(n29145), .A2(n26760), .B1(n25790), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U30990 ( .A1(n29145), .A2(n28553), .B1(n25791), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U30991 ( .A1(n29145), .A2(n29082), .B1(n25792), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U30992 ( .A1(n29145), .A2(n29076), .B1(n25793), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__a22oi_1 U30993 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[13]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[13]), .Y(n25795) );
  sky130_fd_sc_hd__a22oi_1 U30994 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[51]), .B1(n27398), .B2(
        j202_soc_core_intc_core_00_rg_itgt[35]), .Y(n25794) );
  sky130_fd_sc_hd__nand3_1 U30995 ( .A(n25795), .B(n28238), .C(n25794), .Y(
        n25796) );
  sky130_fd_sc_hd__a21oi_1 U30996 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[109]), .B1(n25796), .Y(n25800) );
  sky130_fd_sc_hd__a22oi_1 U30997 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[59]), .B1(n28331), .B2(
        j202_soc_core_intc_core_00_rg_itgt[43]), .Y(n25799) );
  sky130_fd_sc_hd__a22oi_1 U30998 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[13]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[45]), .B2(n28330), .Y(n25798) );
  sky130_fd_sc_hd__nand2_1 U30999 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[77]), .Y(n25797) );
  sky130_fd_sc_hd__nand4_1 U31000 ( .A(n25800), .B(n25799), .C(n25798), .D(
        n25797), .Y(j202_soc_core_ahb2apb_01_N141) );
  sky130_fd_sc_hd__mux2i_1 U31001 ( .A0(n26975), .A1(n26317), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N311) );
  sky130_fd_sc_hd__nand2_1 U31002 ( .A(n28055), .B(n26973), .Y(n25801) );
  sky130_fd_sc_hd__nand2_1 U31003 ( .A(n25801), .B(n12203), .Y(
        j202_soc_core_j22_cpu_ml_machj[8]) );
  sky130_fd_sc_hd__nand3_1 U31004 ( .A(n26973), .B(n27152), .C(n25812), .Y(
        n25814) );
  sky130_fd_sc_hd__nor2_1 U31005 ( .A(n26266), .B(n26341), .Y(n26256) );
  sky130_fd_sc_hd__nand2_1 U31006 ( .A(n26256), .B(n25802), .Y(n26150) );
  sky130_fd_sc_hd__xnor2_1 U31007 ( .A(j202_soc_core_j22_cpu_rfuo_sr__q_), .B(
        n26416), .Y(n25807) );
  sky130_fd_sc_hd__xor2_1 U31008 ( .A(n25807), .B(n26271), .X(n26255) );
  sky130_fd_sc_hd__a22oi_1 U31009 ( .A1(n26362), .A2(n26416), .B1(n26255), 
        .B2(n16501), .Y(n25810) );
  sky130_fd_sc_hd__nand2_1 U31010 ( .A(n28109), .B(n25808), .Y(n25815) );
  sky130_fd_sc_hd__nand3_1 U31011 ( .A(n28483), .B(n27753), .C(n25815), .Y(
        n25809) );
  sky130_fd_sc_hd__a31oi_1 U31013 ( .A1(n26978), .A2(n25812), .A3(n26150), 
        .B1(n25811), .Y(n25813) );
  sky130_fd_sc_hd__nand2_1 U31014 ( .A(n25814), .B(n25813), .Y(
        j202_soc_core_j22_cpu_rf_N2638) );
  sky130_fd_sc_hd__nand2_1 U31015 ( .A(n26865), .B(n25815), .Y(
        j202_soc_core_j22_cpu_rf_N2637) );
  sky130_fd_sc_hd__nor2_1 U31016 ( .A(n26179), .B(n12367), .Y(n25816) );
  sky130_fd_sc_hd__nand2_1 U31017 ( .A(n25817), .B(n26414), .Y(n25861) );
  sky130_fd_sc_hd__nor2_1 U31018 ( .A(n25818), .B(n25825), .Y(n25819) );
  sky130_fd_sc_hd__a21oi_1 U31019 ( .A1(n25820), .A2(n25825), .B1(n25819), .Y(
        n25844) );
  sky130_fd_sc_hd__nand2_1 U31020 ( .A(n25821), .B(n28460), .Y(n25842) );
  sky130_fd_sc_hd__nand2_1 U31021 ( .A(n27809), .B(n25825), .Y(n26305) );
  sky130_fd_sc_hd__nand2b_1 U31022 ( .A_N(n26305), .B(n25822), .Y(n25832) );
  sky130_fd_sc_hd__nor3_1 U31023 ( .A(n27026), .B(n25824), .C(n25823), .Y(
        n25828) );
  sky130_fd_sc_hd__nand2_1 U31024 ( .A(n27026), .B(n28457), .Y(n25826) );
  sky130_fd_sc_hd__nand2_1 U31025 ( .A(n25826), .B(n26305), .Y(n26234) );
  sky130_fd_sc_hd__nand2b_1 U31026 ( .A_N(n26234), .B(n25827), .Y(n25839) );
  sky130_fd_sc_hd__nand4_1 U31027 ( .A(n25829), .B(n25842), .C(n25828), .D(
        n25839), .Y(n25837) );
  sky130_fd_sc_hd__a21oi_1 U31028 ( .A1(n27809), .A2(n25831), .B1(n25830), .Y(
        n25833) );
  sky130_fd_sc_hd__nand3_1 U31029 ( .A(n25839), .B(n25833), .C(n25832), .Y(
        n25834) );
  sky130_fd_sc_hd__nor2_1 U31030 ( .A(n25834), .B(n25840), .Y(n25835) );
  sky130_fd_sc_hd__a31oi_1 U31031 ( .A1(n25835), .A2(n25844), .A3(n25842), 
        .B1(n26048), .Y(n25836) );
  sky130_fd_sc_hd__nand2_1 U31032 ( .A(n25839), .B(n27026), .Y(n25841) );
  sky130_fd_sc_hd__nor2_1 U31033 ( .A(n25841), .B(n25840), .Y(n25843) );
  sky130_fd_sc_hd__nand4_1 U31034 ( .A(n25845), .B(n25844), .C(n25843), .D(
        n25842), .Y(n25853) );
  sky130_fd_sc_hd__nand2_1 U31035 ( .A(n27809), .B(n27785), .Y(n25846) );
  sky130_fd_sc_hd__nand2_1 U31036 ( .A(n25846), .B(n27787), .Y(n25847) );
  sky130_fd_sc_hd__a22oi_1 U31037 ( .A1(n27810), .A2(n26330), .B1(n27808), 
        .B2(n27788), .Y(n25852) );
  sky130_fd_sc_hd__o22ai_1 U31038 ( .A1(n27804), .A2(n27795), .B1(n26318), 
        .B2(n27797), .Y(n25849) );
  sky130_fd_sc_hd__o22ai_1 U31039 ( .A1(n27383), .A2(n27799), .B1(n26296), 
        .B2(n27803), .Y(n25848) );
  sky130_fd_sc_hd__nor2_1 U31040 ( .A(n25849), .B(n25848), .Y(n25851) );
  sky130_fd_sc_hd__nand2_1 U31041 ( .A(n25864), .B(n27789), .Y(n25850) );
  sky130_fd_sc_hd__nand2_1 U31042 ( .A(n25856), .B(n24832), .Y(n25854) );
  sky130_fd_sc_hd__o21ai_0 U31043 ( .A1(n24832), .A2(n27389), .B1(n25854), .Y(
        j202_soc_core_j22_cpu_rf_N3302) );
  sky130_fd_sc_hd__o22ai_1 U31044 ( .A1(n27389), .A2(n27859), .B1(n27858), 
        .B2(n27386), .Y(j202_soc_core_j22_cpu_rf_N3340) );
  sky130_fd_sc_hd__o22ai_1 U31045 ( .A1(n27389), .A2(n27841), .B1(n24712), 
        .B2(n12246), .Y(j202_soc_core_j22_cpu_rf_N3265) );
  sky130_fd_sc_hd__o22ai_1 U31046 ( .A1(n27389), .A2(n25964), .B1(n27847), 
        .B2(n12246), .Y(j202_soc_core_j22_cpu_rf_N2710) );
  sky130_fd_sc_hd__o22ai_1 U31047 ( .A1(n25862), .A2(n27775), .B1(n27774), 
        .B2(n27389), .Y(n25859) );
  sky130_fd_sc_hd__nor2_1 U31048 ( .A(n27648), .B(n25857), .Y(n25858) );
  sky130_fd_sc_hd__nor2_1 U31049 ( .A(n25859), .B(n25858), .Y(n25860) );
  sky130_fd_sc_hd__o21ai_0 U31050 ( .A1(n27648), .A2(n25861), .B1(n25860), .Y(
        j202_soc_core_j22_cpu_rf_N3376) );
  sky130_fd_sc_hd__o22ai_1 U31051 ( .A1(n28457), .A2(n27850), .B1(n25862), 
        .B2(n27848), .Y(n25863) );
  sky130_fd_sc_hd__a21oi_1 U31052 ( .A1(n25864), .A2(n26068), .B1(n25863), .Y(
        n25865) );
  sky130_fd_sc_hd__o21ai_0 U31053 ( .A1(n27855), .A2(n27389), .B1(n25865), .Y(
        j202_soc_core_j22_cpu_rf_N326) );
  sky130_fd_sc_hd__o22ai_1 U31054 ( .A1(n27389), .A2(n25977), .B1(n28061), 
        .B2(n27386), .Y(j202_soc_core_j22_cpu_rf_N2895) );
  sky130_fd_sc_hd__o22ai_1 U31055 ( .A1(n27389), .A2(n25978), .B1(n27834), 
        .B2(n27386), .Y(j202_soc_core_j22_cpu_rf_N2969) );
  sky130_fd_sc_hd__o22ai_1 U31056 ( .A1(n27389), .A2(n25979), .B1(n28112), 
        .B2(n27386), .Y(j202_soc_core_j22_cpu_rf_N3228) );
  sky130_fd_sc_hd__o22ai_1 U31057 ( .A1(n27389), .A2(n25980), .B1(n27835), 
        .B2(n27386), .Y(j202_soc_core_j22_cpu_rf_N2821) );
  sky130_fd_sc_hd__o22ai_1 U31058 ( .A1(n27389), .A2(n25981), .B1(n27836), 
        .B2(n12246), .Y(j202_soc_core_j22_cpu_rf_N3191) );
  sky130_fd_sc_hd__o22ai_1 U31059 ( .A1(n27389), .A2(n25982), .B1(n27837), 
        .B2(n27386), .Y(j202_soc_core_j22_cpu_rf_N3043) );
  sky130_fd_sc_hd__o22ai_1 U31060 ( .A1(n27389), .A2(n25983), .B1(n27838), 
        .B2(n27386), .Y(j202_soc_core_j22_cpu_rf_N3080) );
  sky130_fd_sc_hd__o22ai_1 U31061 ( .A1(n27389), .A2(n25984), .B1(n27840), 
        .B2(n12246), .Y(j202_soc_core_j22_cpu_rf_N2747) );
  sky130_fd_sc_hd__o22ai_1 U31062 ( .A1(n27389), .A2(n25985), .B1(n27842), 
        .B2(n12246), .Y(j202_soc_core_j22_cpu_rf_N3117) );
  sky130_fd_sc_hd__o22ai_1 U31063 ( .A1(n27389), .A2(n25986), .B1(n27843), 
        .B2(n12246), .Y(j202_soc_core_j22_cpu_rf_N3006) );
  sky130_fd_sc_hd__o22ai_1 U31064 ( .A1(n27389), .A2(n25987), .B1(n27844), 
        .B2(n12246), .Y(j202_soc_core_j22_cpu_rf_N3154) );
  sky130_fd_sc_hd__o22ai_1 U31065 ( .A1(n27389), .A2(n25988), .B1(n27845), 
        .B2(n27386), .Y(j202_soc_core_j22_cpu_rf_N2858) );
  sky130_fd_sc_hd__o22ai_1 U31066 ( .A1(n27389), .A2(n25989), .B1(n27846), 
        .B2(n12246), .Y(j202_soc_core_j22_cpu_rf_N2784) );
  sky130_fd_sc_hd__a21oi_1 U31067 ( .A1(n28519), .A2(n27791), .B1(n27790), .Y(
        n25867) );
  sky130_fd_sc_hd__nand2b_1 U31069 ( .A_N(n25869), .B(n25868), .Y(n25886) );
  sky130_fd_sc_hd__o22ai_1 U31070 ( .A1(n27798), .A2(n27799), .B1(n26320), 
        .B2(n27795), .Y(n25871) );
  sky130_fd_sc_hd__o22ai_1 U31071 ( .A1(n27027), .A2(n27803), .B1(n27825), 
        .B2(n26943), .Y(n25870) );
  sky130_fd_sc_hd__nor2_1 U31072 ( .A(n25871), .B(n25870), .Y(n25878) );
  sky130_fd_sc_hd__xnor2_1 U31073 ( .A(n28519), .B(n27115), .Y(n26224) );
  sky130_fd_sc_hd__a2bb2oi_1 U31074 ( .B1(n27810), .B2(n26331), .A1_N(n25872), 
        .A2_N(n26224), .Y(n25877) );
  sky130_fd_sc_hd__o22ai_1 U31075 ( .A1(n26926), .A2(n25873), .B1(n27793), 
        .B2(n28519), .Y(n25875) );
  sky130_fd_sc_hd__nor2_1 U31076 ( .A(n27147), .B(n27797), .Y(n25874) );
  sky130_fd_sc_hd__a211oi_1 U31077 ( .A1(n27808), .A2(n27111), .B1(n25875), 
        .C1(n25874), .Y(n25876) );
  sky130_fd_sc_hd__nand4_1 U31078 ( .A(n27814), .B(n25878), .C(n25877), .D(
        n25876), .Y(n25880) );
  sky130_fd_sc_hd__o22ai_1 U31079 ( .A1(n26272), .A2(n27817), .B1(n26937), 
        .B2(n27815), .Y(n25879) );
  sky130_fd_sc_hd__nor2_1 U31080 ( .A(n25880), .B(n25879), .Y(n25885) );
  sky130_fd_sc_hd__nand2_1 U31081 ( .A(n27115), .B(n27785), .Y(n25881) );
  sky130_fd_sc_hd__o211ai_1 U31082 ( .A1(n11123), .A2(n27115), .B1(n26922), 
        .C1(n25881), .Y(n25882) );
  sky130_fd_sc_hd__nand2_1 U31083 ( .A(n28518), .B(n25882), .Y(n25884) );
  sky130_fd_sc_hd__nand2_1 U31084 ( .A(n25899), .B(n27789), .Y(n25883) );
  sky130_fd_sc_hd__nand4_1 U31085 ( .A(n25886), .B(n25885), .C(n25884), .D(
        n25883), .Y(n25887) );
  sky130_fd_sc_hd__nand2_1 U31086 ( .A(n25890), .B(n25889), .Y(n25891) );
  sky130_fd_sc_hd__nand2_1 U31087 ( .A(n25893), .B(n24832), .Y(n25892) );
  sky130_fd_sc_hd__o21ai_0 U31088 ( .A1(n24832), .A2(n27114), .B1(n25892), .Y(
        j202_soc_core_j22_cpu_rf_N3290) );
  sky130_fd_sc_hd__o22ai_1 U31089 ( .A1(n27859), .A2(n27114), .B1(n27858), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N3329) );
  sky130_fd_sc_hd__o22ai_1 U31090 ( .A1(n27841), .A2(n27114), .B1(n24712), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N3253) );
  sky130_fd_sc_hd__o22ai_1 U31091 ( .A1(n25964), .A2(n27114), .B1(n27847), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N2698) );
  sky130_fd_sc_hd__nand2_1 U31092 ( .A(n25893), .B(n27860), .Y(n25895) );
  sky130_fd_sc_hd__a22oi_1 U31093 ( .A1(n25896), .A2(n27862), .B1(n28518), 
        .B2(n27861), .Y(n25894) );
  sky130_fd_sc_hd__nand2_1 U31094 ( .A(n25895), .B(n25894), .Y(
        j202_soc_core_j22_cpu_rf_N3365) );
  sky130_fd_sc_hd__o22ai_1 U31095 ( .A1(n26272), .A2(n27850), .B1(n25897), 
        .B2(n27848), .Y(n25898) );
  sky130_fd_sc_hd__a21oi_1 U31096 ( .A1(n25899), .A2(n26068), .B1(n25898), .Y(
        n25900) );
  sky130_fd_sc_hd__o21ai_0 U31097 ( .A1(n27855), .A2(n27114), .B1(n25900), .Y(
        j202_soc_core_j22_cpu_rf_N316) );
  sky130_fd_sc_hd__o22ai_1 U31098 ( .A1(n25977), .A2(n27114), .B1(n28061), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N2883) );
  sky130_fd_sc_hd__o22ai_1 U31099 ( .A1(n25978), .A2(n27114), .B1(n27834), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N2957) );
  sky130_fd_sc_hd__o22ai_1 U31100 ( .A1(n25979), .A2(n27114), .B1(n28112), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N3216) );
  sky130_fd_sc_hd__o22ai_1 U31101 ( .A1(n25980), .A2(n27114), .B1(n27835), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N2809) );
  sky130_fd_sc_hd__o22ai_1 U31102 ( .A1(n25981), .A2(n27114), .B1(n27836), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N3179) );
  sky130_fd_sc_hd__o22ai_1 U31103 ( .A1(n25982), .A2(n27114), .B1(n27837), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N3031) );
  sky130_fd_sc_hd__o22ai_1 U31104 ( .A1(n25983), .A2(n27114), .B1(n27838), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N3068) );
  sky130_fd_sc_hd__o22ai_1 U31105 ( .A1(n25984), .A2(n27114), .B1(n27840), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N2735) );
  sky130_fd_sc_hd__o22ai_1 U31106 ( .A1(n25985), .A2(n27114), .B1(n27842), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N3105) );
  sky130_fd_sc_hd__o22ai_1 U31107 ( .A1(n25986), .A2(n27114), .B1(n27843), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N2994) );
  sky130_fd_sc_hd__o22ai_1 U31108 ( .A1(n25987), .A2(n27114), .B1(n27844), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N3142) );
  sky130_fd_sc_hd__o22ai_1 U31109 ( .A1(n25988), .A2(n27114), .B1(n27845), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N2846) );
  sky130_fd_sc_hd__o22ai_1 U31110 ( .A1(n25989), .A2(n27114), .B1(n27846), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N2772) );
  sky130_fd_sc_hd__nor2_1 U31111 ( .A(n28379), .B(n25904), .Y(n28079) );
  sky130_fd_sc_hd__nand2_1 U31112 ( .A(n28079), .B(n29587), .Y(n25905) );
  sky130_fd_sc_hd__nand2_1 U31113 ( .A(n28081), .B(n25905), .Y(n10530) );
  sky130_fd_sc_hd__nand2_1 U31114 ( .A(n26941), .B(n27785), .Y(n25909) );
  sky130_fd_sc_hd__o211ai_1 U31115 ( .A1(n11123), .A2(n26941), .B1(n26922), 
        .C1(n25909), .Y(n25930) );
  sky130_fd_sc_hd__o2bb2ai_1 U31116 ( .B1(n26135), .B2(n26936), .A1_N(n27042), 
        .A2_N(n26935), .Y(n25924) );
  sky130_fd_sc_hd__o21ai_1 U31117 ( .A1(n27023), .A2(n26934), .B1(n26933), .Y(
        n25923) );
  sky130_fd_sc_hd__nand2_1 U31118 ( .A(n25911), .B(n25910), .Y(n25912) );
  sky130_fd_sc_hd__nand2_1 U31119 ( .A(n25912), .B(n26414), .Y(n25914) );
  sky130_fd_sc_hd__nand3_1 U31122 ( .A(n26301), .B(n27806), .C(n26218), .Y(
        n25913) );
  sky130_fd_sc_hd__o211a_2 U31123 ( .A1(n27798), .A2(n27795), .B1(n25914), 
        .C1(n25913), .X(n25915) );
  sky130_fd_sc_hd__o21ai_0 U31124 ( .A1(n27065), .A2(n26932), .B1(n25915), .Y(
        n25922) );
  sky130_fd_sc_hd__nor2_1 U31125 ( .A(n26318), .B(n27803), .Y(n25920) );
  sky130_fd_sc_hd__o22ai_1 U31126 ( .A1(n27793), .A2(n28467), .B1(n26939), 
        .B2(n26301), .Y(n25919) );
  sky130_fd_sc_hd__o22ai_1 U31127 ( .A1(n11190), .A2(n27799), .B1(n27027), 
        .B2(n26943), .Y(n25918) );
  sky130_fd_sc_hd__a22o_1 U31128 ( .A1(n27810), .A2(n26050), .B1(n27808), .B2(
        n25916), .X(n25917) );
  sky130_fd_sc_hd__or4_1 U31129 ( .A(n25920), .B(n25919), .C(n25918), .D(
        n25917), .X(n25921) );
  sky130_fd_sc_hd__or4_1 U31130 ( .A(n25924), .B(n25923), .C(n25922), .D(
        n25921), .X(n25925) );
  sky130_fd_sc_hd__a21oi_1 U31131 ( .A1(n25926), .A2(n27789), .B1(n25925), .Y(
        n25927) );
  sky130_fd_sc_hd__a21oi_1 U31133 ( .A1(n28466), .A2(n25930), .B1(n25929), .Y(
        n25931) );
  sky130_fd_sc_hd__mux2i_1 U31134 ( .A0(n28111), .A1(n28113), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3282) );
  sky130_fd_sc_hd__nor2_1 U31135 ( .A(n27644), .B(n28111), .Y(
        j202_soc_core_j22_cpu_rf_N2654) );
  sky130_fd_sc_hd__o22ai_1 U31136 ( .A1(n28113), .A2(n27841), .B1(n24712), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N3245) );
  sky130_fd_sc_hd__o22ai_1 U31137 ( .A1(n28113), .A2(n25964), .B1(n27847), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N2690) );
  sky130_fd_sc_hd__o22ai_1 U31138 ( .A1(n25933), .A2(n27775), .B1(n27774), 
        .B2(n28113), .Y(n25934) );
  sky130_fd_sc_hd__a21oi_1 U31139 ( .A1(n25935), .A2(n27860), .B1(n25934), .Y(
        n25936) );
  sky130_fd_sc_hd__o22ai_1 U31141 ( .A1(n28113), .A2(n25977), .B1(n28061), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N2875) );
  sky130_fd_sc_hd__o22ai_1 U31142 ( .A1(n28113), .A2(n25978), .B1(n27834), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N2949) );
  sky130_fd_sc_hd__o22ai_1 U31143 ( .A1(n28113), .A2(n25980), .B1(n27835), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N2801) );
  sky130_fd_sc_hd__o22ai_1 U31144 ( .A1(n28113), .A2(n25981), .B1(n27836), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N3171) );
  sky130_fd_sc_hd__o22ai_1 U31145 ( .A1(n28113), .A2(n25982), .B1(n27837), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N3023) );
  sky130_fd_sc_hd__o22ai_1 U31146 ( .A1(n28113), .A2(n25983), .B1(n27838), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N3060) );
  sky130_fd_sc_hd__o22ai_1 U31147 ( .A1(n28113), .A2(n26894), .B1(n27839), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N2912) );
  sky130_fd_sc_hd__o22ai_1 U31148 ( .A1(n28113), .A2(n25984), .B1(n27840), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N2727) );
  sky130_fd_sc_hd__o22ai_1 U31149 ( .A1(n28113), .A2(n25985), .B1(n27842), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N3097) );
  sky130_fd_sc_hd__o22ai_1 U31150 ( .A1(n28113), .A2(n25986), .B1(n27843), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N2986) );
  sky130_fd_sc_hd__o22ai_1 U31151 ( .A1(n28113), .A2(n25987), .B1(n27844), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N3134) );
  sky130_fd_sc_hd__o22ai_1 U31152 ( .A1(n28113), .A2(n25988), .B1(n27845), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N2838) );
  sky130_fd_sc_hd__o22ai_1 U31153 ( .A1(n28113), .A2(n25989), .B1(n27846), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N2764) );
  sky130_fd_sc_hd__nand2b_1 U31155 ( .A_N(n25962), .B(n27785), .Y(n25943) );
  sky130_fd_sc_hd__nand2_1 U31156 ( .A(n25962), .B(n26916), .Y(n25942) );
  sky130_fd_sc_hd__o2bb2ai_1 U31157 ( .B1(n25944), .B2(n26936), .A1_N(n26330), 
        .A2_N(n26935), .Y(n25956) );
  sky130_fd_sc_hd__nand2_1 U31158 ( .A(n25945), .B(n26414), .Y(n25947) );
  sky130_fd_sc_hd__nand2b_1 U31159 ( .A_N(n25973), .B(n26009), .Y(n26294) );
  sky130_fd_sc_hd__nand2_1 U31160 ( .A(n26319), .B(n25973), .Y(n26216) );
  sky130_fd_sc_hd__nand3_1 U31161 ( .A(n26294), .B(n26216), .C(n27806), .Y(
        n25946) );
  sky130_fd_sc_hd__o211a_2 U31162 ( .A1(n26321), .A2(n27795), .B1(n25947), 
        .C1(n25946), .X(n25948) );
  sky130_fd_sc_hd__o21ai_0 U31163 ( .A1(n26275), .A2(n26932), .B1(n25948), .Y(
        n25955) );
  sky130_fd_sc_hd__o21ai_1 U31164 ( .A1(n25973), .A2(n26934), .B1(n26933), .Y(
        n25954) );
  sky130_fd_sc_hd__nor2_1 U31165 ( .A(n26430), .B(n27803), .Y(n25952) );
  sky130_fd_sc_hd__o22ai_1 U31166 ( .A1(n27793), .A2(n28449), .B1(n26939), 
        .B2(n26294), .Y(n25951) );
  sky130_fd_sc_hd__o22ai_1 U31167 ( .A1(n11191), .A2(n27799), .B1(n26324), 
        .B2(n26943), .Y(n25950) );
  sky130_fd_sc_hd__a22o_1 U31168 ( .A1(n27810), .A2(n27111), .B1(n27808), .B2(
        n26946), .X(n25949) );
  sky130_fd_sc_hd__or4_1 U31169 ( .A(n25952), .B(n25951), .C(n25950), .D(
        n25949), .X(n25953) );
  sky130_fd_sc_hd__or4_1 U31170 ( .A(n25956), .B(n25955), .C(n25954), .D(
        n25953), .X(n25957) );
  sky130_fd_sc_hd__a21oi_1 U31171 ( .A1(n25975), .A2(n27789), .B1(n25957), .Y(
        n25960) );
  sky130_fd_sc_hd__nand2_1 U31173 ( .A(n11181), .B(n25958), .Y(n25959) );
  sky130_fd_sc_hd__mux2i_1 U31174 ( .A0(n12262), .A1(n26896), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3286) );
  sky130_fd_sc_hd__nor2_1 U31175 ( .A(n27644), .B(n12262), .Y(
        j202_soc_core_j22_cpu_rf_N2657) );
  sky130_fd_sc_hd__mux2i_1 U31176 ( .A0(n26896), .A1(n26319), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N317) );
  sky130_fd_sc_hd__nand2_1 U31177 ( .A(n28055), .B(n25965), .Y(n25966) );
  sky130_fd_sc_hd__nand2_1 U31178 ( .A(n25966), .B(n12203), .Y(
        j202_soc_core_j22_cpu_ml_machj[14]) );
  sky130_fd_sc_hd__a2bb2oi_1 U31179 ( .B1(n25971), .B2(n27862), .A1_N(n27774), 
        .A2_N(n26896), .Y(n25967) );
  sky130_fd_sc_hd__o22ai_1 U31181 ( .A1(n25973), .A2(n27850), .B1(n25972), 
        .B2(n27848), .Y(n25974) );
  sky130_fd_sc_hd__a21oi_1 U31182 ( .A1(n25975), .A2(n26068), .B1(n25974), .Y(
        n25976) );
  sky130_fd_sc_hd__o21ai_0 U31183 ( .A1(n27855), .A2(n26896), .B1(n25976), .Y(
        j202_soc_core_j22_cpu_rf_N312) );
  sky130_fd_sc_hd__a21oi_1 U31184 ( .A1(j202_soc_core_j22_cpu_ml_bufa[12]), 
        .A2(n28056), .B1(n25990), .Y(n25992) );
  sky130_fd_sc_hd__a21oi_1 U31186 ( .A1(n28460), .A2(n27791), .B1(n27790), .Y(
        n25994) );
  sky130_fd_sc_hd__nand2_1 U31187 ( .A(n25995), .B(n26946), .Y(n26022) );
  sky130_fd_sc_hd__o21ai_1 U31188 ( .A1(n11123), .A2(n26946), .B1(n26922), .Y(
        n26020) );
  sky130_fd_sc_hd__o22ai_1 U31189 ( .A1(n26240), .A2(n26936), .B1(n28457), 
        .B2(n26932), .Y(n26014) );
  sky130_fd_sc_hd__o22ai_1 U31190 ( .A1(n27025), .A2(n27795), .B1(n27026), 
        .B2(n25996), .Y(n25998) );
  sky130_fd_sc_hd__o22ai_1 U31191 ( .A1(n27383), .A2(n26943), .B1(n26321), 
        .B2(n27803), .Y(n25997) );
  sky130_fd_sc_hd__nor2_1 U31192 ( .A(n25998), .B(n25997), .Y(n26012) );
  sky130_fd_sc_hd__xor2_1 U31193 ( .A(n28460), .B(n26946), .X(n26214) );
  sky130_fd_sc_hd__nand2b_1 U31194 ( .A_N(n26299), .B(n25999), .Y(n26007) );
  sky130_fd_sc_hd__nand2_1 U31195 ( .A(n26414), .B(
        j202_soc_core_j22_cpu_ml_bufa[12]), .Y(n26000) );
  sky130_fd_sc_hd__o22ai_1 U31196 ( .A1(n26001), .A2(n26000), .B1(n27793), 
        .B2(n28460), .Y(n26002) );
  sky130_fd_sc_hd__a21oi_1 U31197 ( .A1(n26003), .A2(n27809), .B1(n26002), .Y(
        n26006) );
  sky130_fd_sc_hd__nand2_1 U31198 ( .A(n26004), .B(n26414), .Y(n26005) );
  sky130_fd_sc_hd__nand3_1 U31199 ( .A(n26007), .B(n26006), .C(n26005), .Y(
        n26008) );
  sky130_fd_sc_hd__a21oi_1 U31200 ( .A1(n27806), .A2(n26214), .B1(n26008), .Y(
        n26011) );
  sky130_fd_sc_hd__a22oi_1 U31201 ( .A1(n27810), .A2(n26009), .B1(n27808), 
        .B2(n26923), .Y(n26010) );
  sky130_fd_sc_hd__nand4_1 U31202 ( .A(n26012), .B(n26011), .C(n26010), .D(
        n26933), .Y(n26013) );
  sky130_fd_sc_hd__a211o_1 U31203 ( .A1(n26046), .A2(n28460), .B1(n26014), 
        .C1(n26013), .X(n26015) );
  sky130_fd_sc_hd__a21oi_1 U31204 ( .A1(n26016), .A2(n27789), .B1(n26015), .Y(
        n26017) );
  sky130_fd_sc_hd__o21ai_1 U31205 ( .A1(n26926), .A2(n26018), .B1(n26017), .Y(
        n26019) );
  sky130_fd_sc_hd__a21oi_1 U31206 ( .A1(n28459), .A2(n26020), .B1(n26019), .Y(
        n26021) );
  sky130_fd_sc_hd__nor2_1 U31207 ( .A(n27644), .B(n12343), .Y(
        j202_soc_core_j22_cpu_rf_N2655) );
  sky130_fd_sc_hd__o22ai_1 U31208 ( .A1(n26670), .A2(n27841), .B1(n24712), 
        .B2(n12343), .Y(j202_soc_core_j22_cpu_rf_N3246) );
  sky130_fd_sc_hd__o22ai_1 U31209 ( .A1(n26670), .A2(n25964), .B1(n27847), 
        .B2(n12343), .Y(j202_soc_core_j22_cpu_rf_N2691) );
  sky130_fd_sc_hd__mux2i_1 U31210 ( .A0(n26670), .A1(n26318), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N315) );
  sky130_fd_sc_hd__nand2_1 U31211 ( .A(n28055), .B(n26025), .Y(n26024) );
  sky130_fd_sc_hd__nand2_1 U31212 ( .A(n26024), .B(n12203), .Y(
        j202_soc_core_j22_cpu_ml_machj[12]) );
  sky130_fd_sc_hd__nand2_1 U31213 ( .A(n26025), .B(n27772), .Y(n26030) );
  sky130_fd_sc_hd__a22oi_1 U31214 ( .A1(n26026), .A2(n27862), .B1(n28459), 
        .B2(n27861), .Y(n26029) );
  sky130_fd_sc_hd__nand2_1 U31215 ( .A(n26027), .B(n27860), .Y(n26028) );
  sky130_fd_sc_hd__nand3_1 U31216 ( .A(n26030), .B(n26029), .C(n26028), .Y(
        j202_soc_core_j22_cpu_rf_N3358) );
  sky130_fd_sc_hd__o22ai_1 U31217 ( .A1(n26670), .A2(n25977), .B1(n28061), 
        .B2(n26669), .Y(j202_soc_core_j22_cpu_rf_N2876) );
  sky130_fd_sc_hd__o22ai_1 U31218 ( .A1(n26670), .A2(n25978), .B1(n27834), 
        .B2(n26669), .Y(j202_soc_core_j22_cpu_rf_N2950) );
  sky130_fd_sc_hd__o22ai_1 U31219 ( .A1(n26670), .A2(n25979), .B1(n28112), 
        .B2(n26669), .Y(j202_soc_core_j22_cpu_rf_N3209) );
  sky130_fd_sc_hd__o22ai_1 U31220 ( .A1(n26670), .A2(n25980), .B1(n27835), 
        .B2(n26669), .Y(j202_soc_core_j22_cpu_rf_N2802) );
  sky130_fd_sc_hd__o22ai_1 U31221 ( .A1(n26670), .A2(n25981), .B1(n27836), 
        .B2(n12343), .Y(j202_soc_core_j22_cpu_rf_N3172) );
  sky130_fd_sc_hd__o22ai_1 U31222 ( .A1(n26670), .A2(n25982), .B1(n27837), 
        .B2(n26669), .Y(j202_soc_core_j22_cpu_rf_N3024) );
  sky130_fd_sc_hd__o22ai_1 U31223 ( .A1(n26670), .A2(n25983), .B1(n27838), 
        .B2(n26669), .Y(j202_soc_core_j22_cpu_rf_N3061) );
  sky130_fd_sc_hd__o22ai_1 U31224 ( .A1(n26670), .A2(n25984), .B1(n27840), 
        .B2(n12343), .Y(j202_soc_core_j22_cpu_rf_N2728) );
  sky130_fd_sc_hd__o22ai_1 U31225 ( .A1(n26670), .A2(n25985), .B1(n27842), 
        .B2(n12343), .Y(j202_soc_core_j22_cpu_rf_N3098) );
  sky130_fd_sc_hd__o22ai_1 U31226 ( .A1(n26670), .A2(n25986), .B1(n27843), 
        .B2(n12343), .Y(j202_soc_core_j22_cpu_rf_N2987) );
  sky130_fd_sc_hd__o22ai_1 U31227 ( .A1(n26670), .A2(n25987), .B1(n27844), 
        .B2(n12343), .Y(j202_soc_core_j22_cpu_rf_N3135) );
  sky130_fd_sc_hd__o22ai_1 U31228 ( .A1(n26670), .A2(n25988), .B1(n27845), 
        .B2(n12343), .Y(j202_soc_core_j22_cpu_rf_N2839) );
  sky130_fd_sc_hd__o22ai_1 U31229 ( .A1(n26670), .A2(n25989), .B1(n27846), 
        .B2(n12343), .Y(j202_soc_core_j22_cpu_rf_N2765) );
  sky130_fd_sc_hd__nand3_1 U31230 ( .A(n26032), .B(n26414), .C(n26031), .Y(
        n26067) );
  sky130_fd_sc_hd__nand2_1 U31231 ( .A(n26064), .B(n27785), .Y(n26033) );
  sky130_fd_sc_hd__o211ai_1 U31232 ( .A1(n11123), .A2(n26064), .B1(n26922), 
        .C1(n26033), .Y(n26063) );
  sky130_fd_sc_hd__o21ai_0 U31233 ( .A1(n26939), .A2(n26311), .B1(n26919), .Y(
        n26041) );
  sky130_fd_sc_hd__nand2_1 U31234 ( .A(n26311), .B(n26034), .Y(n26039) );
  sky130_fd_sc_hd__nand2_1 U31235 ( .A(n28045), .B(n26035), .Y(n26036) );
  sky130_fd_sc_hd__o211ai_1 U31236 ( .A1(j202_soc_core_j22_cpu_ml_mach[15]), 
        .A2(n26037), .B1(n27152), .C1(n26036), .Y(n26038) );
  sky130_fd_sc_hd__nand2_1 U31237 ( .A(n26039), .B(n26038), .Y(n26040) );
  sky130_fd_sc_hd__a21oi_1 U31238 ( .A1(n26041), .A2(n26064), .B1(n26040), .Y(
        n26043) );
  sky130_fd_sc_hd__o22a_1 U31239 ( .A1(n26431), .A2(n26943), .B1(n26322), .B2(
        n27803), .X(n26042) );
  sky130_fd_sc_hd__o211ai_1 U31240 ( .A1(n26044), .A2(n26926), .B1(n26043), 
        .C1(n26042), .Y(n26045) );
  sky130_fd_sc_hd__a21oi_1 U31241 ( .A1(n26046), .A2(n28443), .B1(n26045), .Y(
        n26058) );
  sky130_fd_sc_hd__xnor2_1 U31242 ( .A(n26064), .B(n26311), .Y(n26213) );
  sky130_fd_sc_hd__nand2_1 U31243 ( .A(n26213), .B(n27806), .Y(n26047) );
  sky130_fd_sc_hd__a22o_1 U31245 ( .A1(n27810), .A2(n26051), .B1(n27808), .B2(
        n26050), .X(n26052) );
  sky130_fd_sc_hd__nor2_1 U31246 ( .A(n26053), .B(n26052), .Y(n26057) );
  sky130_fd_sc_hd__o22ai_1 U31247 ( .A1(n27616), .A2(n27799), .B1(n26319), 
        .B2(n27795), .Y(n26054) );
  sky130_fd_sc_hd__a21oi_1 U31248 ( .A1(n26416), .A2(n26935), .B1(n26054), .Y(
        n26056) );
  sky130_fd_sc_hd__o22a_1 U31249 ( .A1(n26309), .A2(n26936), .B1(n26408), .B2(
        n26932), .X(n26055) );
  sky130_fd_sc_hd__nand4_1 U31250 ( .A(n26058), .B(n26057), .C(n26056), .D(
        n26055), .Y(n26059) );
  sky130_fd_sc_hd__a21oi_1 U31251 ( .A1(n26069), .A2(n27789), .B1(n26059), .Y(
        n26060) );
  sky130_fd_sc_hd__a21oi_1 U31253 ( .A1(n28442), .A2(n26063), .B1(n26062), .Y(
        n26066) );
  sky130_fd_sc_hd__o22ai_1 U31254 ( .A1(n27859), .A2(n12264), .B1(n27858), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N3326) );
  sky130_fd_sc_hd__a22oi_1 U31255 ( .A1(n26070), .A2(n28443), .B1(n26069), 
        .B2(n26068), .Y(n26073) );
  sky130_fd_sc_hd__nand2_1 U31256 ( .A(n26071), .B(n26074), .Y(n26072) );
  sky130_fd_sc_hd__o211ai_1 U31257 ( .A1(n27855), .A2(n12264), .B1(n26073), 
        .C1(n26072), .Y(j202_soc_core_j22_cpu_rf_N313) );
  sky130_fd_sc_hd__nor2_1 U31258 ( .A(n27644), .B(n11115), .Y(
        j202_soc_core_j22_cpu_rf_N2658) );
  sky130_fd_sc_hd__o22ai_1 U31259 ( .A1(n27841), .A2(n12264), .B1(n24712), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N3250) );
  sky130_fd_sc_hd__o22ai_1 U31260 ( .A1(n25977), .A2(n12264), .B1(n28061), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N2880) );
  sky130_fd_sc_hd__o22ai_1 U31261 ( .A1(n25978), .A2(n12264), .B1(n27834), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N2954) );
  sky130_fd_sc_hd__o22ai_1 U31262 ( .A1(n25979), .A2(n12264), .B1(n28112), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N3213) );
  sky130_fd_sc_hd__o22ai_1 U31263 ( .A1(n25980), .A2(n12264), .B1(n27835), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N2806) );
  sky130_fd_sc_hd__o22ai_1 U31264 ( .A1(n25981), .A2(n12264), .B1(n27836), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N3176) );
  sky130_fd_sc_hd__o22ai_1 U31265 ( .A1(n25982), .A2(n12264), .B1(n27837), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N3028) );
  sky130_fd_sc_hd__o22ai_1 U31266 ( .A1(n25983), .A2(n12264), .B1(n27838), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N3065) );
  sky130_fd_sc_hd__o22ai_1 U31267 ( .A1(n25984), .A2(n12264), .B1(n27840), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N2732) );
  sky130_fd_sc_hd__o22ai_1 U31268 ( .A1(n25985), .A2(n12264), .B1(n27842), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N3102) );
  sky130_fd_sc_hd__o22ai_1 U31269 ( .A1(n25986), .A2(n12264), .B1(n27843), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N2991) );
  sky130_fd_sc_hd__o22ai_1 U31270 ( .A1(n25987), .A2(n12264), .B1(n27844), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N3139) );
  sky130_fd_sc_hd__o22ai_1 U31271 ( .A1(n25988), .A2(n12264), .B1(n27845), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N2843) );
  sky130_fd_sc_hd__o22ai_1 U31272 ( .A1(n25989), .A2(n12264), .B1(n27846), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N2769) );
  sky130_fd_sc_hd__o22ai_1 U31273 ( .A1(n25964), .A2(n12264), .B1(n27847), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N2695) );
  sky130_fd_sc_hd__a22oi_1 U31274 ( .A1(n27862), .A2(n26074), .B1(n28442), 
        .B2(n27861), .Y(n26075) );
  sky130_fd_sc_hd__o21ai_0 U31275 ( .A1(n27648), .A2(n11115), .B1(n26075), .Y(
        j202_soc_core_j22_cpu_rf_N3361) );
  sky130_fd_sc_hd__mux2i_1 U31276 ( .A0(n12264), .A1(n26430), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N318) );
  sky130_fd_sc_hd__nand2_1 U31277 ( .A(n26077), .B(n26076), .Y(n26078) );
  sky130_fd_sc_hd__nand2_1 U31278 ( .A(n26078), .B(n27119), .Y(
        j202_soc_core_j22_cpu_ml_machj[15]) );
  sky130_fd_sc_hd__nand2_1 U31279 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[15]), .Y(n26079) );
  sky130_fd_sc_hd__o21ai_1 U31280 ( .A1(n26093), .A2(n28289), .B1(n26079), .Y(
        n122) );
  sky130_fd_sc_hd__nand2_1 U31281 ( .A(n26080), .B(n26990), .Y(n26081) );
  sky130_fd_sc_hd__nand2_1 U31282 ( .A(n26082), .B(n26081), .Y(n26089) );
  sky130_fd_sc_hd__o21ai_1 U31284 ( .A1(n27723), .A2(n27530), .B1(n26083), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[13]) );
  sky130_fd_sc_hd__nor3_1 U31285 ( .A(n27540), .B(
        j202_soc_core_cmt_core_00_cnt1[14]), .C(n26089), .Y(n26084) );
  sky130_fd_sc_hd__a21oi_1 U31286 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[14]), .A2(n27544), .B1(n26084), 
        .Y(n26085) );
  sky130_fd_sc_hd__o21ai_1 U31288 ( .A1(j202_soc_core_cmt_core_00_cnt1[15]), 
        .A2(n26089), .B1(j202_soc_core_cmt_core_00_cnt1[14]), .Y(n26088) );
  sky130_fd_sc_hd__o211ai_1 U31289 ( .A1(j202_soc_core_cmt_core_00_cnt1[14]), 
        .A2(j202_soc_core_cmt_core_00_cnt1[15]), .B1(n26990), .C1(n26088), .Y(
        n26091) );
  sky130_fd_sc_hd__a22oi_1 U31290 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[15]), .A2(n27544), .B1(n26089), 
        .B2(j202_soc_core_cmt_core_00_cnt1[15]), .Y(n26090) );
  sky130_fd_sc_hd__nand2_1 U31291 ( .A(n26091), .B(n26090), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[15]) );
  sky130_fd_sc_hd__nand2_1 U31292 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[15]), .Y(n26092) );
  sky130_fd_sc_hd__o21ai_1 U31293 ( .A1(n26093), .A2(n28291), .B1(n26092), .Y(
        n128) );
  sky130_fd_sc_hd__a31oi_1 U31294 ( .A1(n26095), .A2(n26096), .A3(
        j202_soc_core_cmt_core_00_cnt0[12]), .B1(
        j202_soc_core_cmt_core_00_cnt0[13]), .Y(n26098) );
  sky130_fd_sc_hd__and3_1 U31295 ( .A(n26096), .B(
        j202_soc_core_cmt_core_00_cnt0[12]), .C(
        j202_soc_core_cmt_core_00_cnt0[13]), .X(n26099) );
  sky130_fd_sc_hd__o22ai_1 U31297 ( .A1(n27482), .A2(n27723), .B1(n26098), 
        .B2(n26101), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[13])
         );
  sky130_fd_sc_hd__nor3_1 U31298 ( .A(j202_soc_core_cmt_core_00_cnt0[14]), .B(
        n26106), .C(n26104), .Y(n26103) );
  sky130_fd_sc_hd__a21oi_1 U31299 ( .A1(n27486), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[14]), .B1(n26103), .Y(n26100) );
  sky130_fd_sc_hd__nor4_1 U31302 ( .A(j202_soc_core_cmt_core_00_cnt0[15]), .B(
        n26106), .C(n26105), .D(n26104), .Y(n26107) );
  sky130_fd_sc_hd__a21oi_1 U31303 ( .A1(n27486), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[15]), .B1(n26107), .Y(n26108) );
  sky130_fd_sc_hd__nand2_1 U31304 ( .A(n26109), .B(n26108), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[15]) );
  sky130_fd_sc_hd__a22oi_1 U31305 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[15]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[15]), 
        .Y(n26111) );
  sky130_fd_sc_hd__a22oi_1 U31306 ( .A1(n28297), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[15]), 
        .B1(n28301), .B2(j202_soc_core_cmt_core_00_const0[15]), .Y(n26110) );
  sky130_fd_sc_hd__nand2_1 U31307 ( .A(n26111), .B(n26110), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[15]) );
  sky130_fd_sc_hd__nand2_1 U31308 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[15]), .Y(n26112) );
  sky130_fd_sc_hd__o21ai_1 U31309 ( .A1(n26113), .A2(n28545), .B1(n26112), .Y(
        n61) );
  sky130_fd_sc_hd__o22ai_1 U31310 ( .A1(n29154), .A2(n28064), .B1(n26116), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__nor2_1 U31311 ( .A(n26114), .B(n27349), .Y(n28066) );
  sky130_fd_sc_hd__nand2_1 U31312 ( .A(n28066), .B(n26748), .Y(n26115) );
  sky130_fd_sc_hd__nand4b_1 U31313 ( .A_N(
        j202_soc_core_intc_core_00_rg_irqc[15]), .B(n26115), .C(
        j202_soc_core_intc_core_00_in_intreq[15]), .D(n12069), .Y(n26118) );
  sky130_fd_sc_hd__nand2b_1 U31314 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[15]), 
        .B(n29567), .Y(n26117) );
  sky130_fd_sc_hd__a21oi_1 U31315 ( .A1(n26118), .A2(n26117), .B1(n26116), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N18) );
  sky130_fd_sc_hd__o22ai_1 U31316 ( .A1(n29154), .A2(n28310), .B1(n26119), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U31317 ( .A1(n29154), .A2(n28313), .B1(n26120), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U31318 ( .A1(n29154), .A2(n28316), .B1(n26121), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U31319 ( .A1(n29154), .A2(n26760), .B1(n26122), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U31320 ( .A1(n29154), .A2(n27575), .B1(n26123), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U31321 ( .A1(n29154), .A2(n28553), .B1(n26124), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U31322 ( .A1(n29154), .A2(n29082), .B1(n26125), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U31323 ( .A1(n29154), .A2(n29076), .B1(n26126), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__a22oi_1 U31324 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[15]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[15]), .Y(n26128) );
  sky130_fd_sc_hd__a22oi_1 U31325 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[115]), .B1(n27398), .B2(
        j202_soc_core_intc_core_00_rg_itgt[99]), .Y(n26127) );
  sky130_fd_sc_hd__nand3_1 U31326 ( .A(n26128), .B(n28238), .C(n26127), .Y(
        n26129) );
  sky130_fd_sc_hd__a21oi_1 U31327 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[111]), .B1(n26129), .Y(n26133) );
  sky130_fd_sc_hd__a22oi_1 U31328 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[123]), .B1(n28331), .B2(
        j202_soc_core_intc_core_00_rg_itgt[107]), .Y(n26132) );
  sky130_fd_sc_hd__a22oi_1 U31329 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[15]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[47]), .B2(n28330), .Y(n26131) );
  sky130_fd_sc_hd__nand2_1 U31330 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[79]), .Y(n26130) );
  sky130_fd_sc_hd__nand4_1 U31331 ( .A(n26133), .B(n26132), .C(n26131), .D(
        n26130), .Y(j202_soc_core_ahb2apb_01_N143) );
  sky130_fd_sc_hd__nor2_1 U31332 ( .A(n29088), .B(n26134), .Y(
        j202_soc_core_wbqspiflash_00_N712) );
  sky130_fd_sc_hd__a22o_1 U31333 ( .A1(n28026), .A2(
        j202_soc_core_wbqspiflash_00_spi_out[15]), .B1(n28025), .B2(
        j202_soc_core_wbqspiflash_00_erased_sector[1]), .X(
        j202_soc_core_wbqspiflash_00_N682) );
  sky130_fd_sc_hd__nor2_1 U31334 ( .A(n28489), .B(n28495), .Y(n26136) );
  sky130_fd_sc_hd__nand4_1 U31335 ( .A(n26136), .B(n26135), .C(n26240), .D(
        n11144), .Y(n26137) );
  sky130_fd_sc_hd__nand2_1 U31336 ( .A(n26137), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[3]), .Y(n26138) );
  sky130_fd_sc_hd__nand2_1 U31337 ( .A(n26138), .B(n26362), .Y(n26155) );
  sky130_fd_sc_hd__nand3_1 U31338 ( .A(n26205), .B(n26208), .C(n26345), .Y(
        n26365) );
  sky130_fd_sc_hd__nand2_1 U31339 ( .A(n26140), .B(n26139), .Y(n26141) );
  sky130_fd_sc_hd__nand2_1 U31340 ( .A(n26365), .B(n26141), .Y(n26147) );
  sky130_fd_sc_hd__nor2_1 U31341 ( .A(n26142), .B(n26341), .Y(n26347) );
  sky130_fd_sc_hd__o22ai_1 U31342 ( .A1(n26145), .A2(n26144), .B1(n26424), 
        .B2(n26143), .Y(n26146) );
  sky130_fd_sc_hd__nor2_1 U31343 ( .A(n26147), .B(n26146), .Y(n26154) );
  sky130_fd_sc_hd__nand2_1 U31344 ( .A(n26149), .B(n26148), .Y(n26339) );
  sky130_fd_sc_hd__o21ai_1 U31345 ( .A1(n26345), .A2(n26373), .B1(n26339), .Y(
        n26152) );
  sky130_fd_sc_hd__o21ai_1 U31346 ( .A1(n26210), .A2(n26374), .B1(n26150), .Y(
        n26151) );
  sky130_fd_sc_hd__nor2_1 U31347 ( .A(n26152), .B(n26151), .Y(n26153) );
  sky130_fd_sc_hd__nand3_1 U31348 ( .A(n26155), .B(n26154), .C(n26153), .Y(
        n26392) );
  sky130_fd_sc_hd__nand3_1 U31349 ( .A(n28109), .B(n26157), .C(n26156), .Y(
        n26396) );
  sky130_fd_sc_hd__nor2_1 U31351 ( .A(n12222), .B(n28470), .Y(n26204) );
  sky130_fd_sc_hd__nor2_1 U31352 ( .A(n28508), .B(n28501), .Y(n26161) );
  sky130_fd_sc_hd__nor2_1 U31353 ( .A(n26163), .B(n12260), .Y(n26203) );
  sky130_fd_sc_hd__nand2_1 U31354 ( .A(n12367), .B(n12423), .Y(n26167) );
  sky130_fd_sc_hd__nor2_1 U31355 ( .A(n26168), .B(n26167), .Y(n26170) );
  sky130_fd_sc_hd__nand4_1 U31356 ( .A(n26172), .B(n26171), .C(n26170), .D(
        n26169), .Y(n26173) );
  sky130_fd_sc_hd__nand2_1 U31357 ( .A(n26173), .B(n26189), .Y(n26176) );
  sky130_fd_sc_hd__nand4_1 U31358 ( .A(n26176), .B(n26175), .C(n26174), .D(
        n27668), .Y(n26184) );
  sky130_fd_sc_hd__a31oi_1 U31359 ( .A1(n26182), .A2(n26181), .A3(n26180), 
        .B1(n26179), .Y(n26183) );
  sky130_fd_sc_hd__nor2_1 U31360 ( .A(n26184), .B(n26183), .Y(n26202) );
  sky130_fd_sc_hd__nand3_1 U31361 ( .A(n26187), .B(n26186), .C(n26185), .Y(
        n26188) );
  sky130_fd_sc_hd__o31a_1 U31362 ( .A1(n26191), .A2(n26190), .A3(n10971), .B1(
        n26189), .X(n26193) );
  sky130_fd_sc_hd__nor2_1 U31363 ( .A(n26193), .B(n26192), .Y(n26198) );
  sky130_fd_sc_hd__nor3_1 U31364 ( .A(n26196), .B(n26195), .C(n26194), .Y(
        n26197) );
  sky130_fd_sc_hd__nand4_1 U31365 ( .A(n26199), .B(n27461), .C(n26198), .D(
        n26197), .Y(n26200) );
  sky130_fd_sc_hd__nor2_1 U31366 ( .A(n26200), .B(n28453), .Y(n26201) );
  sky130_fd_sc_hd__nand4_1 U31367 ( .A(n26204), .B(n26203), .C(n26202), .D(
        n26201), .Y(n26391) );
  sky130_fd_sc_hd__xor2_1 U31368 ( .A(n26206), .B(n26271), .X(n26261) );
  sky130_fd_sc_hd__xor2_1 U31369 ( .A(n26417), .B(n26261), .X(n26364) );
  sky130_fd_sc_hd__o22ai_1 U31370 ( .A1(n26271), .A2(n26207), .B1(n26341), 
        .B2(n26364), .Y(n26209) );
  sky130_fd_sc_hd__nand2_1 U31371 ( .A(n26209), .B(n26208), .Y(n26260) );
  sky130_fd_sc_hd__a21oi_1 U31372 ( .A1(n26300), .A2(n26212), .B1(n26211), .Y(
        n26222) );
  sky130_fd_sc_hd__nor2_1 U31373 ( .A(n26214), .B(n26213), .Y(n26221) );
  sky130_fd_sc_hd__nand2_1 U31374 ( .A(n26944), .B(n26215), .Y(n26217) );
  sky130_fd_sc_hd__a22oi_1 U31375 ( .A1(n26217), .A2(n26292), .B1(n26294), 
        .B2(n26216), .Y(n26220) );
  sky130_fd_sc_hd__nand2b_1 U31376 ( .A_N(n27816), .B(n26923), .Y(n26938) );
  sky130_fd_sc_hd__nand2_1 U31377 ( .A(n27798), .B(n27816), .Y(n26924) );
  sky130_fd_sc_hd__a22oi_1 U31378 ( .A1(n26301), .A2(n26218), .B1(n26938), 
        .B2(n26924), .Y(n26219) );
  sky130_fd_sc_hd__nand4_1 U31379 ( .A(n26222), .B(n26221), .C(n26220), .D(
        n26219), .Y(n26348) );
  sky130_fd_sc_hd__nand4_1 U31380 ( .A(n26226), .B(n26225), .C(n26224), .D(
        n26223), .Y(n26232) );
  sky130_fd_sc_hd__nor2_1 U31381 ( .A(n26228), .B(n26227), .Y(n26231) );
  sky130_fd_sc_hd__nand4b_1 U31382 ( .A_N(n26232), .B(n26231), .C(n26230), .D(
        n26229), .Y(n26350) );
  sky130_fd_sc_hd__nand4_1 U31383 ( .A(n26236), .B(n26235), .C(n26234), .D(
        n26233), .Y(n26239) );
  sky130_fd_sc_hd__xor2_1 U31384 ( .A(n28471), .B(n27788), .X(n27805) );
  sky130_fd_sc_hd__xor2_1 U31385 ( .A(n28463), .B(n27042), .X(n27031) );
  sky130_fd_sc_hd__nor2_1 U31386 ( .A(n27805), .B(n27031), .Y(n26238) );
  sky130_fd_sc_hd__xor2_1 U31387 ( .A(n26416), .B(n26408), .X(n26434) );
  sky130_fd_sc_hd__nand4b_1 U31388 ( .A_N(n26239), .B(n26238), .C(n26434), .D(
        n26237), .Y(n26351) );
  sky130_fd_sc_hd__nand2_1 U31389 ( .A(n27365), .B(n26240), .Y(n26241) );
  sky130_fd_sc_hd__nand2_1 U31390 ( .A(n26299), .B(n26241), .Y(n26244) );
  sky130_fd_sc_hd__nand2_1 U31391 ( .A(n26242), .B(n26293), .Y(n26243) );
  sky130_fd_sc_hd__nand2_1 U31392 ( .A(n26244), .B(n26243), .Y(n26246) );
  sky130_fd_sc_hd__nor2_1 U31393 ( .A(n26246), .B(n26245), .Y(n26254) );
  sky130_fd_sc_hd__a21oi_1 U31394 ( .A1(n26307), .A2(n26248), .B1(n26247), .Y(
        n26253) );
  sky130_fd_sc_hd__nor2b_1 U31395 ( .B_N(n26250), .A(n26249), .Y(n26251) );
  sky130_fd_sc_hd__nand4_1 U31396 ( .A(n26254), .B(n26253), .C(n26252), .D(
        n26251), .Y(n26352) );
  sky130_fd_sc_hd__nand4_1 U31397 ( .A(n26348), .B(n26350), .C(n26351), .D(
        n26352), .Y(n26258) );
  sky130_fd_sc_hd__xnor2_1 U31398 ( .A(j202_soc_core_j22_cpu_rfuo_sr__m_), .B(
        n26255), .Y(n26257) );
  sky130_fd_sc_hd__a22oi_1 U31399 ( .A1(n26346), .A2(n26258), .B1(n26257), 
        .B2(n26256), .Y(n26259) );
  sky130_fd_sc_hd__nand2_1 U31400 ( .A(n26260), .B(n26259), .Y(n26372) );
  sky130_fd_sc_hd__nand3_1 U31401 ( .A(n26271), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[4]), .C(n28104), .Y(n26262) );
  sky130_fd_sc_hd__o21a_1 U31402 ( .A1(n26264), .A2(n26263), .B1(n26262), .X(
        n26370) );
  sky130_fd_sc_hd__a21oi_1 U31403 ( .A1(n26265), .A2(n26416), .B1(n26420), .Y(
        n26267) );
  sky130_fd_sc_hd__o22ai_1 U31404 ( .A1(n26268), .A2(n26267), .B1(n26266), 
        .B2(n26434), .Y(n26269) );
  sky130_fd_sc_hd__a21o_1 U31405 ( .A1(n26271), .A2(n26270), .B1(n26269), .X(
        n26363) );
  sky130_fd_sc_hd__o22ai_1 U31406 ( .A1(n26408), .A2(n28429), .B1(n27800), 
        .B2(n26272), .Y(n26274) );
  sky130_fd_sc_hd__o22ai_1 U31407 ( .A1(n27065), .A2(n27804), .B1(n27027), 
        .B2(n28513), .Y(n26273) );
  sky130_fd_sc_hd__nor2_1 U31408 ( .A(n26274), .B(n26273), .Y(n26291) );
  sky130_fd_sc_hd__o22ai_1 U31409 ( .A1(n26276), .A2(n27796), .B1(n26275), 
        .B2(n26435), .Y(n26279) );
  sky130_fd_sc_hd__o22ai_1 U31410 ( .A1(n27851), .A2(n27825), .B1(n26324), 
        .B2(n26277), .Y(n26278) );
  sky130_fd_sc_hd__nor2_1 U31411 ( .A(n26279), .B(n26278), .Y(n26290) );
  sky130_fd_sc_hd__o22ai_1 U31412 ( .A1(n28506), .A2(n27383), .B1(n27147), 
        .B2(n26937), .Y(n26283) );
  sky130_fd_sc_hd__o22ai_1 U31413 ( .A1(n26281), .A2(n26280), .B1(n26323), 
        .B2(n28481), .Y(n26282) );
  sky130_fd_sc_hd__nor2_1 U31414 ( .A(n26283), .B(n26282), .Y(n26289) );
  sky130_fd_sc_hd__o22ai_1 U31415 ( .A1(n26421), .A2(n11189), .B1(n26284), 
        .B2(n11144), .Y(n26287) );
  sky130_fd_sc_hd__o22ai_1 U31416 ( .A1(n26285), .A2(n26320), .B1(n26322), 
        .B2(n28532), .Y(n26286) );
  sky130_fd_sc_hd__nor2_1 U31417 ( .A(n26287), .B(n26286), .Y(n26288) );
  sky130_fd_sc_hd__nand4_1 U31418 ( .A(n26291), .B(n26290), .C(n26289), .D(
        n26288), .Y(n26360) );
  sky130_fd_sc_hd__nand4_1 U31419 ( .A(n26294), .B(n26938), .C(n26293), .D(
        n26292), .Y(n26304) );
  sky130_fd_sc_hd__nor2_1 U31420 ( .A(n28451), .B(n26296), .Y(n26297) );
  sky130_fd_sc_hd__nor3_1 U31421 ( .A(n26298), .B(n26373), .C(n26297), .Y(
        n26302) );
  sky130_fd_sc_hd__nand4_1 U31422 ( .A(n26302), .B(n26301), .C(n26300), .D(
        n26299), .Y(n26303) );
  sky130_fd_sc_hd__nor2_1 U31423 ( .A(n26304), .B(n26303), .Y(n26316) );
  sky130_fd_sc_hd__nand4_1 U31424 ( .A(n26308), .B(n26307), .C(n26306), .D(
        n26305), .Y(n26314) );
  sky130_fd_sc_hd__o22ai_1 U31425 ( .A1(n26309), .A2(n27616), .B1(n26431), 
        .B2(n28487), .Y(n26313) );
  sky130_fd_sc_hd__o22ai_1 U31426 ( .A1(n26311), .A2(n26430), .B1(n26318), 
        .B2(n26310), .Y(n26312) );
  sky130_fd_sc_hd__nor3_1 U31427 ( .A(n26314), .B(n26313), .C(n26312), .Y(
        n26315) );
  sky130_fd_sc_hd__nand2_1 U31428 ( .A(n26316), .B(n26315), .Y(n26359) );
  sky130_fd_sc_hd__nand4_1 U31429 ( .A(n26430), .B(n26317), .C(
        j202_soc_core_j22_cpu_exuop_EXU_[0]), .D(n27798), .Y(n26328) );
  sky130_fd_sc_hd__nand4_1 U31430 ( .A(n27025), .B(n26319), .C(n26944), .D(
        n26318), .Y(n26327) );
  sky130_fd_sc_hd__nand4_1 U31431 ( .A(n27800), .B(n26322), .C(n26321), .D(
        n26320), .Y(n26326) );
  sky130_fd_sc_hd__nand4_1 U31432 ( .A(n26324), .B(n27027), .C(n26431), .D(
        n26323), .Y(n26325) );
  sky130_fd_sc_hd__nor4_1 U31433 ( .A(n26328), .B(n26327), .C(n26326), .D(
        n26325), .Y(n26338) );
  sky130_fd_sc_hd__nor4_1 U31434 ( .A(n27032), .B(n27042), .C(n27033), .D(
        n26329), .Y(n26337) );
  sky130_fd_sc_hd__nor4_1 U31435 ( .A(n27788), .B(n27809), .C(n26331), .D(
        n26330), .Y(n26336) );
  sky130_fd_sc_hd__nand4_1 U31436 ( .A(n27365), .B(n11189), .C(n11191), .D(
        n27616), .Y(n26333) );
  sky130_fd_sc_hd__nor4_1 U31437 ( .A(n26334), .B(n26377), .C(n26333), .D(
        n26332), .Y(n26335) );
  sky130_fd_sc_hd__nand4_1 U31438 ( .A(n26338), .B(n26337), .C(n26336), .D(
        n26335), .Y(n26344) );
  sky130_fd_sc_hd__nor2_1 U31439 ( .A(n26339), .B(n26416), .Y(n26343) );
  sky130_fd_sc_hd__nor3_1 U31440 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[3]), 
        .B(n26341), .C(n26340), .Y(n26342) );
  sky130_fd_sc_hd__a21oi_1 U31441 ( .A1(n26344), .A2(n26343), .B1(n26342), .Y(
        n26358) );
  sky130_fd_sc_hd__nor2_1 U31443 ( .A(n26349), .B(n26348), .Y(n26356) );
  sky130_fd_sc_hd__clkinv_1 U31444 ( .A(n26350), .Y(n26355) );
  sky130_fd_sc_hd__clkinv_1 U31445 ( .A(n26351), .Y(n26354) );
  sky130_fd_sc_hd__clkinv_1 U31446 ( .A(n26352), .Y(n26353) );
  sky130_fd_sc_hd__nand4_1 U31447 ( .A(n26356), .B(n26355), .C(n26354), .D(
        n26353), .Y(n26357) );
  sky130_fd_sc_hd__o211ai_1 U31448 ( .A1(n26360), .A2(n26359), .B1(n26358), 
        .C1(n26357), .Y(n26361) );
  sky130_fd_sc_hd__a21oi_1 U31449 ( .A1(n26363), .A2(n26362), .B1(n26361), .Y(
        n26369) );
  sky130_fd_sc_hd__nand2_1 U31450 ( .A(n26367), .B(n26366), .Y(n26368) );
  sky130_fd_sc_hd__o211ai_1 U31451 ( .A1(j202_soc_core_j22_cpu_exuop_EXU_[2]), 
        .A2(n26370), .B1(n26369), .C1(n26368), .Y(n26371) );
  sky130_fd_sc_hd__a31oi_1 U31452 ( .A1(n26372), .A2(
        j202_soc_core_j22_cpu_exuop_EXU_[1]), .A3(n28104), .B1(n26371), .Y(
        n26390) );
  sky130_fd_sc_hd__nor2_1 U31453 ( .A(n26374), .B(n26373), .Y(n26380) );
  sky130_fd_sc_hd__nand2_1 U31454 ( .A(n12431), .B(n26375), .Y(n26385) );
  sky130_fd_sc_hd__inv_2 U31455 ( .A(n28508), .Y(n28059) );
  sky130_fd_sc_hd__o21a_1 U31456 ( .A1(n27365), .A2(n28059), .B1(n26376), .X(
        n26387) );
  sky130_fd_sc_hd__nand2_1 U31457 ( .A(n12402), .B(n26378), .Y(n26382) );
  sky130_fd_sc_hd__nand4_1 U31458 ( .A(n13057), .B(n26387), .C(n26379), .D(
        n26382), .Y(n26389) );
  sky130_fd_sc_hd__nand4_1 U31459 ( .A(n26382), .B(n27616), .C(n26381), .D(
        n26380), .Y(n26383) );
  sky130_fd_sc_hd__nor2_1 U31460 ( .A(n26384), .B(n26383), .Y(n26386) );
  sky130_fd_sc_hd__nand3_1 U31461 ( .A(n26387), .B(n26386), .C(n26385), .Y(
        n26388) );
  sky130_fd_sc_hd__nand4_1 U31462 ( .A(n26391), .B(n26390), .C(n26389), .D(
        n26388), .Y(n26394) );
  sky130_fd_sc_hd__nand2_1 U31463 ( .A(n28109), .B(n26392), .Y(n26397) );
  sky130_fd_sc_hd__nand2_1 U31464 ( .A(n26865), .B(n26397), .Y(
        j202_soc_core_j22_cpu_rf_N2625) );
  sky130_fd_sc_hd__nand4_1 U31465 ( .A(n26399), .B(n27828), .C(n26398), .D(
        n26400), .Y(n26407) );
  sky130_fd_sc_hd__and3_1 U31466 ( .A(n26401), .B(n27052), .C(n26400), .X(
        n26402) );
  sky130_fd_sc_hd__nand2_1 U31467 ( .A(n26403), .B(n26402), .Y(n26415) );
  sky130_fd_sc_hd__nand2_1 U31468 ( .A(n26405), .B(n26404), .Y(n26406) );
  sky130_fd_sc_hd__nand3_1 U31469 ( .A(n26407), .B(n26414), .C(n26406), .Y(
        n26413) );
  sky130_fd_sc_hd__o21a_1 U31470 ( .A1(n26408), .A2(n26939), .B1(n26919), .X(
        n26410) );
  sky130_fd_sc_hd__nand2_1 U31471 ( .A(n26415), .B(n26414), .Y(n26449) );
  sky130_fd_sc_hd__nand2_1 U31473 ( .A(n26417), .B(n27789), .Y(n26444) );
  sky130_fd_sc_hd__nand2_1 U31474 ( .A(n28429), .B(n26937), .Y(n26418) );
  sky130_fd_sc_hd__o211ai_1 U31475 ( .A1(j202_soc_core_j22_cpu_rfuo_sr__t_), 
        .A2(n26937), .B1(n26418), .C1(n26942), .Y(n26423) );
  sky130_fd_sc_hd__nand3_1 U31476 ( .A(n26420), .B(n26419), .C(n28521), .Y(
        n26422) );
  sky130_fd_sc_hd__mux2i_1 U31477 ( .A0(n26423), .A1(n26422), .S(n26421), .Y(
        n26442) );
  sky130_fd_sc_hd__nand2_1 U31478 ( .A(n27808), .B(n27033), .Y(n26429) );
  sky130_fd_sc_hd__o21ai_1 U31479 ( .A1(n26929), .A2(n26425), .B1(n26424), .Y(
        n26427) );
  sky130_fd_sc_hd__nand3_1 U31480 ( .A(n26427), .B(n26426), .C(n28443), .Y(
        n26428) );
  sky130_fd_sc_hd__nand2_1 U31481 ( .A(n26429), .B(n26428), .Y(n26433) );
  sky130_fd_sc_hd__o22ai_1 U31482 ( .A1(n26431), .A2(n27799), .B1(n26430), 
        .B2(n27797), .Y(n26432) );
  sky130_fd_sc_hd__nor2_1 U31483 ( .A(n26433), .B(n26432), .Y(n26440) );
  sky130_fd_sc_hd__o22ai_1 U31484 ( .A1(n28431), .A2(n27793), .B1(n26435), 
        .B2(n27795), .Y(n26436) );
  sky130_fd_sc_hd__a21oi_1 U31485 ( .A1(n26437), .A2(n27806), .B1(n26436), .Y(
        n26439) );
  sky130_fd_sc_hd__nand2_1 U31486 ( .A(n27039), .B(n28431), .Y(n26438) );
  sky130_fd_sc_hd__nand4_1 U31487 ( .A(n27814), .B(n26440), .C(n26439), .D(
        n26438), .Y(n26441) );
  sky130_fd_sc_hd__nor2_1 U31488 ( .A(n26442), .B(n26441), .Y(n26443) );
  sky130_fd_sc_hd__nand2_1 U31489 ( .A(n26444), .B(n26443), .Y(n26445) );
  sky130_fd_sc_hd__o22ai_1 U31491 ( .A1(n25977), .A2(n27586), .B1(n28061), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N2898) );
  sky130_fd_sc_hd__o22ai_1 U31492 ( .A1(n25981), .A2(n27586), .B1(n27836), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N3194) );
  sky130_fd_sc_hd__o22ai_1 U31493 ( .A1(n25982), .A2(n27586), .B1(n27837), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N3046) );
  sky130_fd_sc_hd__o22ai_1 U31494 ( .A1(n25987), .A2(n27586), .B1(n27844), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N3157) );
  sky130_fd_sc_hd__o22ai_1 U31495 ( .A1(n25989), .A2(n27586), .B1(n27846), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N2787) );
  sky130_fd_sc_hd__o22ai_1 U31496 ( .A1(n25984), .A2(n27586), .B1(n27840), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N2750) );
  sky130_fd_sc_hd__o22ai_1 U31497 ( .A1(n25988), .A2(n27586), .B1(n27845), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N2861) );
  sky130_fd_sc_hd__o22ai_1 U31498 ( .A1(n25978), .A2(n27586), .B1(n27834), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N2972) );
  sky130_fd_sc_hd__o22ai_1 U31499 ( .A1(n26894), .A2(n27586), .B1(n27839), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N2935) );
  sky130_fd_sc_hd__o22ai_1 U31500 ( .A1(n25980), .A2(n27586), .B1(n27835), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N2824) );
  sky130_fd_sc_hd__o22ai_1 U31501 ( .A1(n25983), .A2(n27586), .B1(n27838), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N3083) );
  sky130_fd_sc_hd__o22ai_1 U31502 ( .A1(n25979), .A2(n27586), .B1(n28112), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N3231) );
  sky130_fd_sc_hd__o22ai_1 U31503 ( .A1(n25986), .A2(n27586), .B1(n27843), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N3009) );
  sky130_fd_sc_hd__o22ai_1 U31504 ( .A1(n25964), .A2(n27586), .B1(n27847), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N2713) );
  sky130_fd_sc_hd__o22ai_1 U31505 ( .A1(n25985), .A2(n27586), .B1(n27842), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N3120) );
  sky130_fd_sc_hd__nor2_1 U31506 ( .A(n27644), .B(n27583), .Y(
        j202_soc_core_j22_cpu_rf_N2676) );
  sky130_fd_sc_hd__o22ai_1 U31507 ( .A1(n27841), .A2(n27586), .B1(n24712), 
        .B2(n27583), .Y(j202_soc_core_j22_cpu_rf_N3268) );
  sky130_fd_sc_hd__o22ai_1 U31508 ( .A1(n25983), .A2(n25245), .B1(n27838), 
        .B2(n26451), .Y(j202_soc_core_j22_cpu_rf_N3074) );
  sky130_fd_sc_hd__nand2_1 U31509 ( .A(n26454), .B(n24832), .Y(n26452) );
  sky130_fd_sc_hd__o21ai_0 U31510 ( .A1(n24832), .A2(n26456), .B1(n26452), .Y(
        j202_soc_core_j22_cpu_rf_N3297) );
  sky130_fd_sc_hd__o22ai_1 U31511 ( .A1(n26456), .A2(n27859), .B1(n27858), 
        .B2(n26453), .Y(j202_soc_core_j22_cpu_rf_N3336) );
  sky130_fd_sc_hd__nand2_1 U31512 ( .A(n26454), .B(n27860), .Y(n26458) );
  sky130_fd_sc_hd__o22a_1 U31513 ( .A1(n26459), .A2(n27775), .B1(n27774), .B2(
        n26456), .X(n26457) );
  sky130_fd_sc_hd__nand2_1 U31514 ( .A(n26458), .B(n26457), .Y(
        j202_soc_core_j22_cpu_rf_N3372) );
  sky130_fd_sc_hd__o22ai_1 U31515 ( .A1(n28481), .A2(n27850), .B1(n26459), 
        .B2(n27848), .Y(n26460) );
  sky130_fd_sc_hd__a21oi_1 U31516 ( .A1(n26461), .A2(n26068), .B1(n26460), .Y(
        n26462) );
  sky130_fd_sc_hd__o21ai_0 U31517 ( .A1(n27855), .A2(n26456), .B1(n26462), .Y(
        j202_soc_core_j22_cpu_rf_N322) );
  sky130_fd_sc_hd__nor2_1 U31519 ( .A(n26465), .B(n26464), .Y(n29167) );
  sky130_fd_sc_hd__nand2_1 U31520 ( .A(n26466), .B(n29167), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N313) );
  sky130_fd_sc_hd__a211oi_1 U31521 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[7]), .A2(n28653), .B1(
        n28647), .C1(n26469), .Y(n26468) );
  sky130_fd_sc_hd__nor2_1 U31522 ( .A(n26468), .B(n28651), .Y(
        j202_soc_core_wbqspiflash_00_N621) );
  sky130_fd_sc_hd__xnor2_1 U31523 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[8]), .B(n26469), .Y(n26470)
         );
  sky130_fd_sc_hd__a21oi_1 U31524 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), 
        .A2(n26470), .B1(n28651), .Y(j202_soc_core_wbqspiflash_00_N622) );
  sky130_fd_sc_hd__a21oi_1 U31525 ( .A1(n26471), .A2(
        j202_soc_core_wbqspiflash_00_reset_counter[9]), .B1(n28647), .Y(n26472) );
  sky130_fd_sc_hd__a21oi_1 U31526 ( .A1(n26472), .A2(n26651), .B1(n28651), .Y(
        j202_soc_core_wbqspiflash_00_N623) );
  sky130_fd_sc_hd__nor2_1 U31527 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[0]), .B(n29276), .Y(
        j202_soc_core_wbqspiflash_00_N614) );
  sky130_fd_sc_hd__xor2_1 U31528 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[2]), .B(n26474), .X(n26473)
         );
  sky130_fd_sc_hd__a21oi_1 U31529 ( .A1(n26473), .A2(
        j202_soc_core_wbqspiflash_00_state[0]), .B1(n28651), .Y(
        j202_soc_core_wbqspiflash_00_N616) );
  sky130_fd_sc_hd__a21oi_1 U31530 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[2]), .A2(
        j202_soc_core_wbqspiflash_00_reset_counter[3]), .B1(n28647), .Y(n26476) );
  sky130_fd_sc_hd__nand2_1 U31531 ( .A(n26474), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[3]), .Y(n26475) );
  sky130_fd_sc_hd__a31oi_1 U31532 ( .A1(n28645), .A2(n26476), .A3(n26475), 
        .B1(n28651), .Y(j202_soc_core_wbqspiflash_00_N617) );
  sky130_fd_sc_hd__nor2_1 U31533 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[8]), .B(n26477), .Y(n28682)
         );
  sky130_fd_sc_hd__nand2_1 U31534 ( .A(n28682), .B(n26478), .Y(
        j202_soc_core_wbqspiflash_00_N85) );
  sky130_fd_sc_hd__o21ai_1 U31535 ( .A1(n28651), .A2(n26480), .B1(n29827), .Y(
        j202_soc_core_wbqspiflash_00_N742) );
  sky130_fd_sc_hd__nor2_1 U31536 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .B(n26481), .Y(n28858)
         );
  sky130_fd_sc_hd__nand2_1 U31537 ( .A(n28858), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .Y(n27272) );
  sky130_fd_sc_hd__nand2_1 U31538 ( .A(n28729), .B(n27296), .Y(n26503) );
  sky130_fd_sc_hd__o21ai_1 U31539 ( .A1(j202_soc_core_wbqspiflash_00_spif_cmd), 
        .A2(n27272), .B1(n26503), .Y(n27265) );
  sky130_fd_sc_hd__a21oi_1 U31540 ( .A1(n26482), .A2(n27265), .B1(n26635), .Y(
        n26494) );
  sky130_fd_sc_hd__nand2_1 U31541 ( .A(n27228), .B(n26484), .Y(n28863) );
  sky130_fd_sc_hd__nand2_1 U31542 ( .A(n26486), .B(n27287), .Y(n26495) );
  sky130_fd_sc_hd__a31oi_1 U31543 ( .A1(n26487), .A2(n28864), .A3(n27430), 
        .B1(n26630), .Y(n26488) );
  sky130_fd_sc_hd__nand2_1 U31544 ( .A(n26519), .B(n28688), .Y(n28671) );
  sky130_fd_sc_hd__nand3_1 U31545 ( .A(n26488), .B(n27240), .C(n28671), .Y(
        n27256) );
  sky130_fd_sc_hd__nand2_1 U31546 ( .A(n27228), .B(n28647), .Y(n27187) );
  sky130_fd_sc_hd__nand2b_1 U31547 ( .A_N(n27187), .B(n27219), .Y(n28844) );
  sky130_fd_sc_hd__nor2_1 U31548 ( .A(j202_soc_core_wbqspiflash_00_state[3]), 
        .B(n27279), .Y(n27274) );
  sky130_fd_sc_hd__nand2_1 U31549 ( .A(n27274), .B(
        j202_soc_core_wbqspiflash_00_state[4]), .Y(n27259) );
  sky130_fd_sc_hd__nand2_1 U31550 ( .A(n28844), .B(n27259), .Y(n26562) );
  sky130_fd_sc_hd__nor3_1 U31551 ( .A(n28687), .B(n27256), .C(n26562), .Y(
        n26493) );
  sky130_fd_sc_hd__nand2_1 U31552 ( .A(n27296), .B(n26489), .Y(n27194) );
  sky130_fd_sc_hd__o21ai_1 U31554 ( .A1(n26491), .A2(n27250), .B1(n28843), .Y(
        n26492) );
  sky130_fd_sc_hd__a31oi_1 U31555 ( .A1(n26494), .A2(n26493), .A3(n26492), 
        .B1(j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N736) );
  sky130_fd_sc_hd__nand2_1 U31556 ( .A(n28685), .B(n26495), .Y(n26520) );
  sky130_fd_sc_hd__a31oi_1 U31557 ( .A1(n27285), .A2(n28647), .A3(n27264), 
        .B1(n29088), .Y(n26496) );
  sky130_fd_sc_hd__nand3_1 U31558 ( .A(n27248), .B(n27186), .C(n26496), .Y(
        n26501) );
  sky130_fd_sc_hd__a21oi_1 U31559 ( .A1(n28840), .A2(n26499), .B1(n26498), .Y(
        n26500) );
  sky130_fd_sc_hd__or3_1 U31560 ( .A(n26502), .B(n26501), .C(n26500), .X(
        j202_soc_core_wbqspiflash_00_N735) );
  sky130_fd_sc_hd__o22a_1 U31561 ( .A1(n27183), .A2(n27194), .B1(n26504), .B2(
        n26503), .X(n26505) );
  sky130_fd_sc_hd__nand3_1 U31562 ( .A(n26507), .B(n26506), .C(n26505), .Y(
        n26508) );
  sky130_fd_sc_hd__nor4_1 U31563 ( .A(n28744), .B(n28861), .C(n26508), .D(
        n28878), .Y(n26509) );
  sky130_fd_sc_hd__nor2_1 U31564 ( .A(n29088), .B(n26509), .Y(
        j202_soc_core_wbqspiflash_00_N737) );
  sky130_fd_sc_hd__a21oi_1 U31565 ( .A1(n28708), .A2(
        j202_soc_core_wbqspiflash_00_spi_valid), .B1(n26511), .Y(n26617) );
  sky130_fd_sc_hd__o31ai_1 U31566 ( .A1(n26580), .A2(n27279), .A3(n27278), 
        .B1(n26512), .Y(n26610) );
  sky130_fd_sc_hd__a21oi_1 U31567 ( .A1(n26514), .A2(n26513), .B1(n26610), .Y(
        n26515) );
  sky130_fd_sc_hd__nand2_1 U31568 ( .A(n28731), .B(n26515), .Y(n26518) );
  sky130_fd_sc_hd__nor2_1 U31569 ( .A(j202_soc_core_wbqspiflash_00_spi_valid), 
        .B(n26516), .Y(n26517) );
  sky130_fd_sc_hd__nor4_1 U31570 ( .A(n26617), .B(n28886), .C(n26518), .D(
        n26517), .Y(n26524) );
  sky130_fd_sc_hd__nor2_1 U31571 ( .A(j202_soc_core_wbqspiflash_00_state[3]), 
        .B(n26519), .Y(n28852) );
  sky130_fd_sc_hd__nor3_1 U31572 ( .A(n26520), .B(n26594), .C(n28852), .Y(
        n26523) );
  sky130_fd_sc_hd__a21oi_1 U31573 ( .A1(n27429), .A2(n26612), .B1(n28828), .Y(
        n26522) );
  sky130_fd_sc_hd__nand2b_1 U31574 ( .A_N(n27280), .B(n26521), .Y(n28656) );
  sky130_fd_sc_hd__nor2_1 U31575 ( .A(n27220), .B(n28878), .Y(n28679) );
  sky130_fd_sc_hd__nand4_1 U31576 ( .A(n26524), .B(n26523), .C(n26522), .D(
        n28679), .Y(n26526) );
  sky130_fd_sc_hd__o22ai_1 U31577 ( .A1(n28866), .A2(n27613), .B1(n27246), 
        .B2(n26597), .Y(n26525) );
  sky130_fd_sc_hd__a31oi_1 U31578 ( .A1(n26526), .A2(j202_soc_core_qspi_wb_cyc), .A3(j202_soc_core_wbqspiflash_00_spif_req), .B1(n26525), .Y(n26527) );
  sky130_fd_sc_hd__nor2_1 U31580 ( .A(n29088), .B(n28843), .Y(n27308) );
  sky130_fd_sc_hd__o22ai_1 U31581 ( .A1(
        j202_soc_core_wbqspiflash_00_spif_data[28]), .A2(n26529), .B1(n29568), 
        .B2(n27308), .Y(j202_soc_core_wbqspiflash_00_N722) );
  sky130_fd_sc_hd__nand3_1 U31582 ( .A(n28836), .B(n26647), .C(io_out[8]), .Y(
        n26536) );
  sky130_fd_sc_hd__nand3_1 U31583 ( .A(n28843), .B(n27193), .C(n28739), .Y(
        n26593) );
  sky130_fd_sc_hd__a21oi_1 U31584 ( .A1(n26603), .A2(n26530), .B1(n29088), .Y(
        n26531) );
  sky130_fd_sc_hd__o31ai_1 U31585 ( .A1(n26532), .A2(n27430), .A3(n26536), 
        .B1(n26531), .Y(j202_soc_core_wbqspiflash_00_N721) );
  sky130_fd_sc_hd__nand2_1 U31586 ( .A(n28730), .B(n28859), .Y(n26581) );
  sky130_fd_sc_hd__nor2_1 U31587 ( .A(n26612), .B(n26533), .Y(n26599) );
  sky130_fd_sc_hd__nor3_1 U31589 ( .A(n26538), .B(n26537), .C(n26536), .Y(
        n26541) );
  sky130_fd_sc_hd__nor2_1 U31590 ( .A(n27257), .B(n26634), .Y(n26540) );
  sky130_fd_sc_hd__nor4_1 U31591 ( .A(n26599), .B(n26541), .C(n26540), .D(
        n26539), .Y(n26542) );
  sky130_fd_sc_hd__o31ai_1 U31592 ( .A1(n26633), .A2(
        j202_soc_core_wbqspiflash_00_spi_busy), .A3(n26581), .B1(n26542), .Y(
        n26551) );
  sky130_fd_sc_hd__a21oi_1 U31593 ( .A1(n26544), .A2(n26543), .B1(n27193), .Y(
        n26545) );
  sky130_fd_sc_hd__a21oi_1 U31594 ( .A1(j202_soc_core_qspi_wb_ack), .A2(n26546), .B1(n26545), .Y(n26547) );
  sky130_fd_sc_hd__a21oi_1 U31595 ( .A1(n27197), .A2(
        j202_soc_core_wbqspiflash_00_write_protect), .B1(n26547), .Y(n26549)
         );
  sky130_fd_sc_hd__a21oi_1 U31597 ( .A1(n26551), .A2(
        j202_soc_core_wbqspiflash_00_spif_req), .B1(n26550), .Y(n26553) );
  sky130_fd_sc_hd__nand3_1 U31598 ( .A(n28843), .B(n27193), .C(n29569), .Y(
        n26552) );
  sky130_fd_sc_hd__o21ai_1 U31599 ( .A1(n29088), .A2(n26553), .B1(n26552), .Y(
        j202_soc_core_wbqspiflash_00_N730) );
  sky130_fd_sc_hd__o21ai_1 U31600 ( .A1(n28861), .A2(n27220), .B1(n12069), .Y(
        j202_soc_core_wbqspiflash_00_N729) );
  sky130_fd_sc_hd__a31oi_1 U31601 ( .A1(n26556), .A2(n26555), .A3(n26558), 
        .B1(n27226), .Y(n27191) );
  sky130_fd_sc_hd__nand2_1 U31602 ( .A(n28688), .B(n26557), .Y(n26638) );
  sky130_fd_sc_hd__nor2_1 U31603 ( .A(n27226), .B(n26559), .Y(n27245) );
  sky130_fd_sc_hd__a21oi_1 U31604 ( .A1(n26559), .A2(n26558), .B1(n27245), .Y(
        n26560) );
  sky130_fd_sc_hd__o22ai_1 U31605 ( .A1(n26580), .A2(n26638), .B1(n26597), 
        .B2(n26560), .Y(n26561) );
  sky130_fd_sc_hd__a211o_1 U31606 ( .A1(n27191), .A2(n26594), .B1(n26562), 
        .C1(n26561), .X(j202_soc_core_wbqspiflash_00_N590) );
  sky130_fd_sc_hd__nand2_1 U31607 ( .A(n27219), .B(
        j202_soc_core_wbqspiflash_00_spi_busy), .Y(n27185) );
  sky130_fd_sc_hd__a21oi_1 U31608 ( .A1(n28840), .A2(
        j202_soc_core_wbqspiflash_00_state[0]), .B1(
        j202_soc_core_wbqspiflash_00_state[1]), .Y(n26563) );
  sky130_fd_sc_hd__o21ai_1 U31609 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), 
        .A2(n27185), .B1(n26563), .Y(n26566) );
  sky130_fd_sc_hd__a21oi_1 U31610 ( .A1(n26566), .A2(n26565), .B1(n29088), .Y(
        j202_soc_core_wbqspiflash_00_N745) );
  sky130_fd_sc_hd__a31oi_1 U31611 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_state[0]), .A2(
        j202_soc_core_wbqspiflash_00_spi_wr), .A3(n26568), .B1(n26567), .Y(
        n26573) );
  sky130_fd_sc_hd__nand2_1 U31613 ( .A(n29257), .B(n26570), .Y(n28693) );
  sky130_fd_sc_hd__nand2_1 U31614 ( .A(n28693), .B(n26571), .Y(n26656) );
  sky130_fd_sc_hd__or4_1 U31615 ( .A(n26573), .B(n26662), .C(n26572), .D(
        n26656), .X(j202_soc_core_wbqspiflash_00_lldriver_N321) );
  sky130_fd_sc_hd__nor3_1 U31616 ( .A(n26612), .B(n26575), .C(n27278), .Y(
        n26577) );
  sky130_fd_sc_hd__nor4_1 U31617 ( .A(n26594), .B(n26577), .C(n26576), .D(
        j202_soc_core_wbqspiflash_00_N710), .Y(n26578) );
  sky130_fd_sc_hd__nand2_1 U31619 ( .A(n28688), .B(n26580), .Y(n26582) );
  sky130_fd_sc_hd__nand4_1 U31620 ( .A(n26583), .B(n26582), .C(n26581), .D(
        n26640), .Y(n26591) );
  sky130_fd_sc_hd__nand2_1 U31621 ( .A(n28837), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .Y(n27202) );
  sky130_fd_sc_hd__nand2_1 U31622 ( .A(n27202), .B(n27251), .Y(n26584) );
  sky130_fd_sc_hd__a21oi_1 U31623 ( .A1(n28730), .A2(n26584), .B1(n28836), .Y(
        n28882) );
  sky130_fd_sc_hd__nor3_1 U31626 ( .A(n26588), .B(n27254), .C(n27191), .Y(
        n26589) );
  sky130_fd_sc_hd__o31ai_1 U31627 ( .A1(n26591), .A2(n26590), .A3(n26589), 
        .B1(n29830), .Y(n26592) );
  sky130_fd_sc_hd__o31ai_1 U31628 ( .A1(
        j202_soc_core_wbqspiflash_00_write_in_progress), .A2(n26593), .A3(
        n27601), .B1(n26592), .Y(j202_soc_core_wbqspiflash_00_N727) );
  sky130_fd_sc_hd__o21ai_1 U31629 ( .A1(n26596), .A2(n26595), .B1(n26594), .Y(
        n26628) );
  sky130_fd_sc_hd__nand2_1 U31630 ( .A(j202_soc_core_wbqspiflash_00_spi_len[1]), .B(j202_soc_core_wbqspiflash_00_spi_len[0]), .Y(n28722) );
  sky130_fd_sc_hd__o22ai_1 U31631 ( .A1(n28651), .A2(n26651), .B1(n27245), 
        .B2(n26597), .Y(n26598) );
  sky130_fd_sc_hd__a31oi_1 U31632 ( .A1(n28717), .A2(
        j202_soc_core_wbqspiflash_00_spi_valid), .A3(n28878), .B1(n26598), .Y(
        n26607) );
  sky130_fd_sc_hd__nor2_1 U31633 ( .A(n26599), .B(n26635), .Y(n26606) );
  sky130_fd_sc_hd__nor2_1 U31634 ( .A(n28656), .B(n26600), .Y(n26602) );
  sky130_fd_sc_hd__nor2_1 U31635 ( .A(n26623), .B(n28731), .Y(n26601) );
  sky130_fd_sc_hd__nor4_1 U31636 ( .A(n29088), .B(n26602), .C(n26601), .D(
        n28888), .Y(n26605) );
  sky130_fd_sc_hd__nand3_1 U31637 ( .A(n26603), .B(
        j202_soc_core_qspi_wb_wdat[31]), .C(
        j202_soc_core_wbqspiflash_00_write_in_progress), .Y(n26604) );
  sky130_fd_sc_hd__nand4_1 U31638 ( .A(n26607), .B(n26606), .C(n26605), .D(
        n26604), .Y(n26615) );
  sky130_fd_sc_hd__a22oi_1 U31639 ( .A1(n27287), .A2(n27286), .B1(n26608), 
        .B2(j202_soc_core_wbqspiflash_00_state[1]), .Y(n26609) );
  sky130_fd_sc_hd__o21ai_1 U31640 ( .A1(j202_soc_core_wbqspiflash_00_state[4]), 
        .A2(n27187), .B1(n26609), .Y(n26611) );
  sky130_fd_sc_hd__a211oi_1 U31641 ( .A1(io_out[8]), .A2(n26611), .B1(n27431), 
        .C1(n26610), .Y(n26613) );
  sky130_fd_sc_hd__a211oi_1 U31643 ( .A1(n28843), .A2(n26616), .B1(n26615), 
        .C1(n26614), .Y(n26627) );
  sky130_fd_sc_hd__nand3_1 U31644 ( .A(n28840), .B(n27287), .C(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n28686) );
  sky130_fd_sc_hd__o31ai_1 U31646 ( .A1(n28686), .A2(n28722), .A3(io_out[8]), 
        .B1(n26618), .Y(n26625) );
  sky130_fd_sc_hd__nand2_1 U31647 ( .A(n27268), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n26619) );
  sky130_fd_sc_hd__o21ai_1 U31648 ( .A1(io_out[8]), .A2(n26619), .B1(n27181), 
        .Y(n26621) );
  sky130_fd_sc_hd__nor4_1 U31649 ( .A(j202_soc_core_wbqspiflash_00_spi_in[28]), 
        .B(j202_soc_core_wbqspiflash_00_spi_in[30]), .C(n29133), .D(n26640), 
        .Y(n26620) );
  sky130_fd_sc_hd__a22oi_1 U31650 ( .A1(n27228), .A2(n26621), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[29]), .B2(n26620), .Y(n26622) );
  sky130_fd_sc_hd__o211ai_1 U31651 ( .A1(n28727), .A2(n28734), .B1(n26622), 
        .C1(n28724), .Y(n26624) );
  sky130_fd_sc_hd__nand3_1 U31653 ( .A(n26628), .B(n26627), .C(n26626), .Y(
        j202_soc_core_wbqspiflash_00_N723) );
  sky130_fd_sc_hd__nand3_1 U31654 ( .A(n26629), .B(n28687), .C(n28841), .Y(
        n26650) );
  sky130_fd_sc_hd__a21oi_1 U31655 ( .A1(n26631), .A2(n27274), .B1(n26630), .Y(
        n26632) );
  sky130_fd_sc_hd__nand2_1 U31656 ( .A(n27221), .B(
        j202_soc_core_wbqspiflash_00_state[4]), .Y(n27253) );
  sky130_fd_sc_hd__o21ai_1 U31657 ( .A1(n26633), .A2(n26632), .B1(n27253), .Y(
        n26646) );
  sky130_fd_sc_hd__o21ai_1 U31658 ( .A1(n26634), .A2(n27187), .B1(n28686), .Y(
        n26636) );
  sky130_fd_sc_hd__nor3_1 U31659 ( .A(n28888), .B(n26636), .C(n26635), .Y(
        n26644) );
  sky130_fd_sc_hd__o211ai_1 U31660 ( .A1(n28866), .A2(n27226), .B1(
        j202_soc_core_wbqspiflash_00_write_in_progress), .C1(n26637), .Y(
        n26639) );
  sky130_fd_sc_hd__nand4_1 U31661 ( .A(n26640), .B(n26639), .C(n27259), .D(
        n26638), .Y(n26642) );
  sky130_fd_sc_hd__nor2_1 U31662 ( .A(n26642), .B(n26641), .Y(n26643) );
  sky130_fd_sc_hd__nand3_1 U31663 ( .A(n26644), .B(n28679), .C(n26643), .Y(
        n26645) );
  sky130_fd_sc_hd__a21oi_1 U31664 ( .A1(n26647), .A2(n26646), .B1(n26645), .Y(
        n26648) );
  sky130_fd_sc_hd__a31oi_1 U31665 ( .A1(n26650), .A2(n26649), .A3(n26648), 
        .B1(j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N734) );
  sky130_fd_sc_hd__nand3_1 U31666 ( .A(n26652), .B(n29745), .C(n26651), .Y(
        j202_soc_core_wbqspiflash_00_N733) );
  sky130_fd_sc_hd__nor4_1 U31667 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[3]), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[1]), .C(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[4]), .D(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[5]), .Y(n26658) );
  sky130_fd_sc_hd__nor2_1 U31668 ( .A(n28726), .B(n26667), .Y(n28694) );
  sky130_fd_sc_hd__nand2_1 U31669 ( .A(n28694), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[2]), .Y(n26655) );
  sky130_fd_sc_hd__nand2_1 U31670 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[0]), .B(n26653), .Y(
        n26654) );
  sky130_fd_sc_hd__o22ai_1 U31671 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[0]), .A2(n26655), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[2]), .B2(n26654), .Y(
        n26657) );
  sky130_fd_sc_hd__a21oi_1 U31672 ( .A1(n26658), .A2(n26657), .B1(n26656), .Y(
        n26659) );
  sky130_fd_sc_hd__o211ai_1 U31673 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_sck), .A2(n26661), .B1(n26660), 
        .C1(n26659), .Y(j202_soc_core_wbqspiflash_00_lldriver_N307) );
  sky130_fd_sc_hd__o21ai_1 U31674 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .A2(n26664), .B1(
        n26663), .Y(j202_soc_core_wbqspiflash_00_lldriver_N309) );
  sky130_fd_sc_hd__nor2_1 U31675 ( .A(j202_soc_core_wbqspiflash_00_spi_hold), 
        .B(n26665), .Y(n26668) );
  sky130_fd_sc_hd__nand4b_1 U31676 ( .A_N(n26668), .B(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .C(n26667), .D(n26666), 
        .Y(j202_soc_core_wbqspiflash_00_lldriver_N308) );
  sky130_fd_sc_hd__o22ai_1 U31677 ( .A1(n26670), .A2(n26894), .B1(n27839), 
        .B2(n12343), .Y(j202_soc_core_j22_cpu_rf_N2913) );
  sky130_fd_sc_hd__o22ai_1 U31678 ( .A1(n26670), .A2(n27859), .B1(n27858), 
        .B2(n12343), .Y(j202_soc_core_j22_cpu_rf_N3323) );
  sky130_fd_sc_hd__o22ai_1 U31679 ( .A1(n29147), .A2(n27575), .B1(n26671), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U31680 ( .A1(n29155), .A2(n27575), .B1(n26672), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U31681 ( .A1(n29153), .A2(n27575), .B1(n30173), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U31682 ( .A1(n29159), .A2(n28064), .B1(n26676), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__nor2_1 U31683 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[3]), .B(n26674), .Y(n26696) );
  sky130_fd_sc_hd__nand2_1 U31684 ( .A(n26713), .B(n26696), .Y(n26675) );
  sky130_fd_sc_hd__nand4b_1 U31685 ( .A_N(
        j202_soc_core_intc_core_00_rg_irqc[5]), .B(n26675), .C(
        j202_soc_core_intc_core_00_in_intreq[5]), .D(n29827), .Y(n26678) );
  sky130_fd_sc_hd__nand2b_1 U31686 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[5]), 
        .B(n29570), .Y(n26677) );
  sky130_fd_sc_hd__a21oi_1 U31687 ( .A1(n26678), .A2(n26677), .B1(n26676), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N8) );
  sky130_fd_sc_hd__nor2_1 U31688 ( .A(n29088), .B(
        j202_soc_core_qspi_wb_wdat[20]), .Y(n29047) );
  sky130_fd_sc_hd__o22ai_1 U31689 ( .A1(n26704), .A2(n26679), .B1(n29047), 
        .B2(n26702), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U31690 ( .A1(n29160), .A2(n28064), .B1(n26684), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__a21oi_1 U31691 ( .A1(n26696), .A2(n26719), .B1(
        j202_soc_core_intc_core_00_rg_irqc[4]), .Y(n26682) );
  sky130_fd_sc_hd__nor2_1 U31692 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[4]), 
        .B(n26680), .Y(n26681) );
  sky130_fd_sc_hd__a31oi_1 U31693 ( .A1(n26682), .A2(
        j202_soc_core_intc_core_00_in_intreq[4]), .A3(n29830), .B1(n26681), 
        .Y(n26683) );
  sky130_fd_sc_hd__nor2_1 U31694 ( .A(n26684), .B(n26683), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N7) );
  sky130_fd_sc_hd__nor2_1 U31695 ( .A(n29088), .B(
        j202_soc_core_qspi_wb_wdat[16]), .Y(n29016) );
  sky130_fd_sc_hd__o22ai_1 U31696 ( .A1(n26704), .A2(n26685), .B1(n29016), 
        .B2(n26702), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U31697 ( .A1(n29151), .A2(n27575), .B1(n26686), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U31698 ( .A1(n29152), .A2(n27575), .B1(n26687), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U31699 ( .A1(n27633), .A2(n27575), .B1(n26688), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U31700 ( .A1(n28002), .A2(n27575), .B1(n26689), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U31701 ( .A1(n27875), .A2(n27575), .B1(n26690), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U31702 ( .A1(n29157), .A2(n28064), .B1(n26692), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__nand2_1 U31703 ( .A(n28066), .B(n26696), .Y(n26691) );
  sky130_fd_sc_hd__nand4b_1 U31704 ( .A_N(
        j202_soc_core_intc_core_00_rg_irqc[7]), .B(n26691), .C(
        j202_soc_core_intc_core_00_in_intreq[7]), .D(n12069), .Y(n26694) );
  sky130_fd_sc_hd__nand2b_1 U31705 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[7]), 
        .B(n29572), .Y(n26693) );
  sky130_fd_sc_hd__a21oi_1 U31706 ( .A1(n26694), .A2(n26693), .B1(n26692), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N10) );
  sky130_fd_sc_hd__nor2_1 U31707 ( .A(n29088), .B(
        j202_soc_core_qspi_wb_wdat[28]), .Y(n29062) );
  sky130_fd_sc_hd__o22ai_1 U31708 ( .A1(n26704), .A2(n26695), .B1(n29062), 
        .B2(n26702), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U31709 ( .A1(n29158), .A2(n28064), .B1(n26701), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__a21oi_1 U31710 ( .A1(n26696), .A2(n26747), .B1(
        j202_soc_core_intc_core_00_rg_irqc[6]), .Y(n26699) );
  sky130_fd_sc_hd__nor2_1 U31711 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[6]), 
        .B(n26697), .Y(n26698) );
  sky130_fd_sc_hd__a31oi_1 U31712 ( .A1(n26699), .A2(
        j202_soc_core_intc_core_00_in_intreq[6]), .A3(n29827), .B1(n26698), 
        .Y(n26700) );
  sky130_fd_sc_hd__nor2_1 U31713 ( .A(n26701), .B(n26700), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N9) );
  sky130_fd_sc_hd__nor2_1 U31714 ( .A(n29088), .B(
        j202_soc_core_qspi_wb_wdat[24]), .Y(n29054) );
  sky130_fd_sc_hd__o22ai_1 U31715 ( .A1(n26704), .A2(n26703), .B1(n29054), 
        .B2(n26702), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U31716 ( .A1(n27172), .A2(n27575), .B1(n26705), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U31717 ( .A1(n27655), .A2(n27575), .B1(n26706), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U31718 ( .A1(n27395), .A2(n27575), .B1(n26707), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U31719 ( .A1(n27078), .A2(n27575), .B1(n26708), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U31720 ( .A1(n27601), .A2(n27575), .B1(n26709), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U31721 ( .A1(n29158), .A2(n26760), .B1(n26710), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U31722 ( .A1(n29162), .A2(n26760), .B1(n26711), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U31723 ( .A1(n26746), .A2(n26712), .B1(n28931), 
        .B2(n26744), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U31724 ( .A1(n29148), .A2(n28064), .B1(n26715), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__nand2_1 U31725 ( .A(n26713), .B(n28065), .Y(n26714) );
  sky130_fd_sc_hd__nand4b_1 U31726 ( .A_N(
        j202_soc_core_intc_core_00_rg_irqc[9]), .B(n26714), .C(
        j202_soc_core_intc_core_00_in_intreq[9]), .D(n29830), .Y(n26717) );
  sky130_fd_sc_hd__nand2b_1 U31727 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[9]), 
        .B(n29574), .Y(n26716) );
  sky130_fd_sc_hd__a21oi_1 U31728 ( .A1(n26717), .A2(n26716), .B1(n26715), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N12) );
  sky130_fd_sc_hd__o22ai_1 U31729 ( .A1(n26746), .A2(n26718), .B1(n28246), 
        .B2(n26744), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U31730 ( .A1(n29146), .A2(n28064), .B1(n26724), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__a21oi_1 U31731 ( .A1(n28065), .A2(n26719), .B1(
        j202_soc_core_intc_core_00_rg_irqc[8]), .Y(n26722) );
  sky130_fd_sc_hd__nor2_1 U31732 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[8]), 
        .B(n26720), .Y(n26721) );
  sky130_fd_sc_hd__a31oi_1 U31733 ( .A1(n26722), .A2(
        j202_soc_core_intc_core_00_in_intreq[8]), .A3(n12069), .B1(n26721), 
        .Y(n26723) );
  sky130_fd_sc_hd__nor2_1 U31734 ( .A(n26724), .B(n26723), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N11) );
  sky130_fd_sc_hd__o22ai_1 U31735 ( .A1(n29163), .A2(n26760), .B1(n26725), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U31736 ( .A1(n29159), .A2(n26760), .B1(n26726), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U31737 ( .A1(n29165), .A2(n26760), .B1(n26727), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U31738 ( .A1(n29160), .A2(n26760), .B1(n26728), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U31739 ( .A1(n29161), .A2(n26760), .B1(n26729), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U31740 ( .A1(n29157), .A2(n26760), .B1(n26730), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U31741 ( .A1(n29144), .A2(n26760), .B1(n26731), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U31742 ( .A1(n26746), .A2(n26732), .B1(n28959), 
        .B2(n26744), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U31743 ( .A1(n29148), .A2(n26760), .B1(n26733), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U31744 ( .A1(n29146), .A2(n26760), .B1(n26734), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U31745 ( .A1(n29155), .A2(n26760), .B1(n26735), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U31746 ( .A1(n29153), .A2(n26760), .B1(n26736), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U31747 ( .A1(n26746), .A2(n26737), .B1(n29047), 
        .B2(n26744), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U31748 ( .A1(n26746), .A2(n26738), .B1(n29016), 
        .B2(n26744), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U31749 ( .A1(n29151), .A2(n26760), .B1(n26739), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U31750 ( .A1(n29152), .A2(n26760), .B1(n12695), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U31751 ( .A1(n27633), .A2(n26760), .B1(n26740), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U31752 ( .A1(n28002), .A2(n26760), .B1(n26741), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U31753 ( .A1(n27875), .A2(n26760), .B1(n26742), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U31754 ( .A1(n26746), .A2(n26743), .B1(n29062), 
        .B2(n26744), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U31755 ( .A1(n26746), .A2(n26745), .B1(n29054), 
        .B2(n26744), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U31756 ( .A1(n29144), .A2(n28064), .B1(n26753), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__a21oi_1 U31757 ( .A1(n26748), .A2(n26747), .B1(
        j202_soc_core_intc_core_00_rg_irqc[14]), .Y(n26751) );
  sky130_fd_sc_hd__nor2_1 U31758 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[14]), 
        .B(n26749), .Y(n26750) );
  sky130_fd_sc_hd__a31oi_1 U31759 ( .A1(n26751), .A2(
        j202_soc_core_intc_core_00_in_intreq[14]), .A3(n12069), .B1(n26750), 
        .Y(n26752) );
  sky130_fd_sc_hd__nor2_1 U31760 ( .A(n26753), .B(n26752), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N17) );
  sky130_fd_sc_hd__o22ai_1 U31761 ( .A1(n27172), .A2(n26760), .B1(n26754), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U31762 ( .A1(n27655), .A2(n26760), .B1(n26755), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U31763 ( .A1(n27395), .A2(n26760), .B1(n26756), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U31764 ( .A1(n27078), .A2(n26760), .B1(n26757), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U31765 ( .A1(n27601), .A2(n26760), .B1(n26759), 
        .B2(n26758), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U31766 ( .A1(n29158), .A2(n28553), .B1(n26761), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U31767 ( .A1(n27658), .A2(n26762), .B1(n28931), 
        .B2(n27656), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U31768 ( .A1(n29151), .A2(n28064), .B1(n26763), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U31769 ( .A1(n27658), .A2(n26765), .B1(n28246), 
        .B2(n27656), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U31770 ( .A1(n29157), .A2(n28553), .B1(n26766), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U31771 ( .A1(n29155), .A2(n28553), .B1(n26767), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U31772 ( .A1(n29153), .A2(n28064), .B1(n26855), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__nand2_1 U31773 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[0]), 
        .B(j202_soc_core_ahb2apb_02_hsize_buf[1]), .Y(
        j202_soc_core_ahb2apb_02_N123) );
  sky130_fd_sc_hd__clkinv_1 U31774 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[0]), 
        .Y(n26771) );
  sky130_fd_sc_hd__nand2_1 U31775 ( .A(n26773), .B(n26771), .Y(n26770) );
  sky130_fd_sc_hd__nor2_1 U31776 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[1]), 
        .B(n26771), .Y(n26774) );
  sky130_fd_sc_hd__clkinv_1 U31777 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[1]), 
        .Y(n26768) );
  sky130_fd_sc_hd__nor2_1 U31778 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[0]), 
        .B(n26768), .Y(n26772) );
  sky130_fd_sc_hd__a21oi_1 U31779 ( .A1(j202_soc_core_gpio_core_00_reg_addr[1]), .A2(n26774), .B1(n26772), .Y(n26769) );
  sky130_fd_sc_hd__o21ai_0 U31780 ( .A1(j202_soc_core_gpio_core_00_reg_addr[0]), .A2(n26770), .B1(n26769), .Y(n10945) );
  sky130_fd_sc_hd__o21ai_0 U31781 ( .A1(n26770), .A2(n26777), .B1(n26769), .Y(
        n10944) );
  sky130_fd_sc_hd__nand2_1 U31782 ( .A(j202_soc_core_gpio_core_00_reg_addr[1]), 
        .B(n26771), .Y(n26776) );
  sky130_fd_sc_hd__a21oi_1 U31783 ( .A1(n26774), .A2(n26773), .B1(n26772), .Y(
        n26775) );
  sky130_fd_sc_hd__o21ai_0 U31784 ( .A1(j202_soc_core_gpio_core_00_reg_addr[0]), .A2(n26776), .B1(n26775), .Y(n10943) );
  sky130_fd_sc_hd__o21ai_0 U31785 ( .A1(n26777), .A2(n26776), .B1(n26775), .Y(
        n10942) );
  sky130_fd_sc_hd__nand2_1 U31786 ( .A(n12069), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[31]), .Y(n26781) );
  sky130_fd_sc_hd__a21oi_1 U31787 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[31]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[31]), .B1(gpio_en_o[31]), 
        .Y(n26778) );
  sky130_fd_sc_hd__nand2_1 U31788 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[31]), .B(n26778), .Y(
        n26779) );
  sky130_fd_sc_hd__a21oi_1 U31789 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[31]), .A2(n26780), 
        .B1(n26779), .Y(n26786) );
  sky130_fd_sc_hd__o21ai_1 U31790 ( .A1(j202_soc_core_rst), .A2(n26782), .B1(
        n26781), .Y(n26785) );
  sky130_fd_sc_hd__o21ai_1 U31791 ( .A1(n29088), .A2(
        j202_soc_core_qspi_wb_wdat[31]), .B1(n29039), .Y(n26784) );
  sky130_fd_sc_hd__a22o_1 U31792 ( .A1(n26786), .A2(n26785), .B1(n26784), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[31]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N71) );
  sky130_fd_sc_hd__nand2_1 U31793 ( .A(n29827), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[30]), .Y(n26790) );
  sky130_fd_sc_hd__a21oi_1 U31794 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[30]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[30]), .B1(gpio_en_o[30]), 
        .Y(n26787) );
  sky130_fd_sc_hd__nand2_1 U31795 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[30]), .B(n26787), .Y(
        n26788) );
  sky130_fd_sc_hd__a21oi_1 U31796 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[30]), .A2(n26789), 
        .B1(n26788), .Y(n26794) );
  sky130_fd_sc_hd__o21ai_1 U31797 ( .A1(n29088), .A2(n26791), .B1(n26790), .Y(
        n26793) );
  sky130_fd_sc_hd__a22o_1 U31799 ( .A1(n26794), .A2(n26793), .B1(n26792), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[30]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N70) );
  sky130_fd_sc_hd__nand2_1 U31800 ( .A(n29745), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[29]), .Y(n26798) );
  sky130_fd_sc_hd__clkinv_1 U31801 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[29]), .Y(n26795) );
  sky130_fd_sc_hd__a21oi_1 U31802 ( .A1(n26795), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[29]), .B1(
        gpio_en_o[29]), .Y(n26796) );
  sky130_fd_sc_hd__nand2_1 U31803 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[29]), .B(n26796), .Y(
        n26797) );
  sky130_fd_sc_hd__a21oi_1 U31804 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[29]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[29]), .B1(n26797), .Y(
        n26802) );
  sky130_fd_sc_hd__o21ai_1 U31805 ( .A1(n29088), .A2(n26799), .B1(n26798), .Y(
        n26801) );
  sky130_fd_sc_hd__o21ai_1 U31806 ( .A1(n29088), .A2(
        j202_soc_core_qspi_wb_wdat[29]), .B1(n29039), .Y(n26800) );
  sky130_fd_sc_hd__a22o_1 U31807 ( .A1(n26802), .A2(n26801), .B1(n26800), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[29]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N69) );
  sky130_fd_sc_hd__clkinv_1 U31808 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[27]), .Y(n26803) );
  sky130_fd_sc_hd__o21ai_1 U31809 ( .A1(n26803), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[27]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[27]), .Y(n26804) );
  sky130_fd_sc_hd__a21oi_1 U31810 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[27]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[27]), .B1(n26804), 
        .Y(n26808) );
  sky130_fd_sc_hd__a21oi_1 U31811 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[27]), .A2(n12069), 
        .B1(n29577), .Y(n26805) );
  sky130_fd_sc_hd__nor2_1 U31812 ( .A(gpio_en_o[27]), .B(n26805), .Y(n26807)
         );
  sky130_fd_sc_hd__a22o_1 U31814 ( .A1(n26808), .A2(n26807), .B1(n26806), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[27]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N67) );
  sky130_fd_sc_hd__a21oi_1 U31815 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[26]), .A2(n29830), 
        .B1(n29578), .Y(n26815) );
  sky130_fd_sc_hd__o2bb2ai_1 U31816 ( .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[26]), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[26]), .A1_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[26]), .A2_N(n26809), .Y(
        n26811) );
  sky130_fd_sc_hd__clkinv_1 U31817 ( .A(gpio_en_o[26]), .Y(n26810) );
  sky130_fd_sc_hd__nand3_1 U31818 ( .A(n26811), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[26]), .C(n26810), .Y(
        n26814) );
  sky130_fd_sc_hd__a21oi_1 U31819 ( .A1(n29827), .A2(n27867), .B1(n29061), .Y(
        n26812) );
  sky130_fd_sc_hd__o22ai_1 U31820 ( .A1(n26815), .A2(n26814), .B1(n26813), 
        .B2(n26812), .Y(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N66)
         );
  sky130_fd_sc_hd__nand2_1 U31821 ( .A(n29827), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[25]), .Y(n26819) );
  sky130_fd_sc_hd__clkinv_1 U31822 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[25]), .Y(n26816) );
  sky130_fd_sc_hd__a21oi_1 U31823 ( .A1(n26816), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[25]), .B1(
        gpio_en_o[25]), .Y(n26817) );
  sky130_fd_sc_hd__nand2_1 U31824 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[25]), .B(n26817), .Y(
        n26818) );
  sky130_fd_sc_hd__a21oi_1 U31825 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[25]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[25]), .B1(n26818), .Y(
        n26823) );
  sky130_fd_sc_hd__clkinv_1 U31826 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[25]), .Y(n26820) );
  sky130_fd_sc_hd__o21ai_1 U31827 ( .A1(j202_soc_core_rst), .A2(n26820), .B1(
        n26819), .Y(n26822) );
  sky130_fd_sc_hd__o21ai_1 U31828 ( .A1(j202_soc_core_rst), .A2(
        j202_soc_core_qspi_wb_wdat[25]), .B1(n29039), .Y(n26821) );
  sky130_fd_sc_hd__a22o_1 U31829 ( .A1(n26823), .A2(n26822), .B1(n26821), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[25]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N65) );
  sky130_fd_sc_hd__nor2_1 U31830 ( .A(j202_soc_core_rst), .B(n26824), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N26) );
  sky130_fd_sc_hd__a21oi_1 U31831 ( .A1(n29827), .A2(n27625), .B1(n29061), .Y(
        n26829) );
  sky130_fd_sc_hd__a21oi_1 U31832 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[23]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[23]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[23]), .Y(n26827) );
  sky130_fd_sc_hd__nor2_1 U31833 ( .A(j202_soc_core_rst), .B(gpio_en_o[23]), 
        .Y(n26826) );
  sky130_fd_sc_hd__nand4b_1 U31835 ( .A_N(n26827), .B(n26826), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[23]), .D(n26825), .Y(
        n26828) );
  sky130_fd_sc_hd__o21ai_1 U31836 ( .A1(n26830), .A2(n26829), .B1(n26828), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N63) );
  sky130_fd_sc_hd__a21oi_1 U31837 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[22]), .A2(n29745), 
        .B1(n29579), .Y(n26838) );
  sky130_fd_sc_hd__o2bb2ai_1 U31838 ( .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[22]), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[22]), .A1_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[22]), .A2_N(n26831), .Y(
        n26833) );
  sky130_fd_sc_hd__clkinv_1 U31839 ( .A(gpio_en_o[22]), .Y(n26832) );
  sky130_fd_sc_hd__nand3_1 U31840 ( .A(n26833), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[22]), .C(n26832), .Y(
        n26837) );
  sky130_fd_sc_hd__a21oi_1 U31841 ( .A1(n29745), .A2(n26834), .B1(n29061), .Y(
        n26835) );
  sky130_fd_sc_hd__o22ai_1 U31842 ( .A1(n26838), .A2(n26837), .B1(n26836), 
        .B2(n26835), .Y(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N62)
         );
  sky130_fd_sc_hd__nand2_1 U31843 ( .A(n29745), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[21]), .Y(n26842) );
  sky130_fd_sc_hd__a21oi_1 U31844 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[21]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[21]), .B1(gpio_en_o[21]), 
        .Y(n26839) );
  sky130_fd_sc_hd__nand2_1 U31845 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[21]), .B(n26839), .Y(
        n26840) );
  sky130_fd_sc_hd__a21oi_1 U31846 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[21]), .A2(n26841), 
        .B1(n26840), .Y(n26846) );
  sky130_fd_sc_hd__o21ai_1 U31847 ( .A1(n29088), .A2(n26843), .B1(n26842), .Y(
        n26845) );
  sky130_fd_sc_hd__a22o_1 U31849 ( .A1(n26846), .A2(n26845), .B1(n26844), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[21]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N61) );
  sky130_fd_sc_hd__a21oi_1 U31850 ( .A1(n29745), .A2(n28902), .B1(n29061), .Y(
        n26851) );
  sky130_fd_sc_hd__clkinv_1 U31851 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[1]), .Y(n26847) );
  sky130_fd_sc_hd__o22ai_1 U31852 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[1]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]), .B1(n26847), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[1]), .Y(n26848)
         );
  sky130_fd_sc_hd__a21oi_1 U31853 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[1]), .B1(n26848), 
        .Y(n26849) );
  sky130_fd_sc_hd__nand4_1 U31854 ( .A(n26849), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[1]), .C(n29745), .D(
        io_oeb[1]), .Y(n26850) );
  sky130_fd_sc_hd__o21ai_1 U31855 ( .A1(n26852), .A2(n26851), .B1(n26850), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N41) );
  sky130_fd_sc_hd__nand2b_1 U31856 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[18]), 
        .B(n29580), .Y(n26857) );
  sky130_fd_sc_hd__nand3_1 U31857 ( .A(n26853), .B(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[1]), .C(n27350), .Y(n26854) );
  sky130_fd_sc_hd__nand4b_1 U31858 ( .A_N(
        j202_soc_core_intc_core_00_rg_irqc[18]), .B(n26854), .C(
        j202_soc_core_intc_core_00_in_intreq[18]), .D(n12069), .Y(n26856) );
  sky130_fd_sc_hd__a21oi_1 U31859 ( .A1(n26857), .A2(n26856), .B1(n26855), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N21) );
  sky130_fd_sc_hd__o22ai_1 U31860 ( .A1(n27658), .A2(n26858), .B1(n28959), 
        .B2(n27656), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U31861 ( .A1(n29153), .A2(n28553), .B1(n26859), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__nand2_1 U31862 ( .A(n27753), .B(n26860), .Y(n27580) );
  sky130_fd_sc_hd__nand2_1 U31863 ( .A(n27578), .B(
        j202_soc_core_intr_level__4_), .Y(n26861) );
  sky130_fd_sc_hd__o21ai_1 U31864 ( .A1(n27578), .A2(
        j202_soc_core_j22_cpu_rf_N2627), .B1(n26861), .Y(n27577) );
  sky130_fd_sc_hd__a21oi_1 U31865 ( .A1(j202_soc_core_intr_level__2_), .A2(
        n27578), .B1(n27577), .Y(n26863) );
  sky130_fd_sc_hd__nor2_1 U31866 ( .A(j202_soc_core_j22_cpu_intack), .B(n27753), .Y(n27576) );
  sky130_fd_sc_hd__o211ai_1 U31867 ( .A1(n27461), .A2(n27580), .B1(n26863), 
        .C1(n26862), .Y(j202_soc_core_j22_cpu_rf_N3390) );
  sky130_fd_sc_hd__nand2_1 U31868 ( .A(n26865), .B(n26864), .Y(
        j202_soc_core_j22_cpu_rf_N3391) );
  sky130_fd_sc_hd__o22ai_1 U31869 ( .A1(n27461), .A2(n25977), .B1(n28061), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N2869) );
  sky130_fd_sc_hd__o22ai_1 U31870 ( .A1(n27461), .A2(n25978), .B1(n27834), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N2943) );
  sky130_fd_sc_hd__o22ai_1 U31871 ( .A1(n27461), .A2(n25979), .B1(n28112), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N3202) );
  sky130_fd_sc_hd__o22ai_1 U31872 ( .A1(n27461), .A2(n25980), .B1(n27835), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N2795) );
  sky130_fd_sc_hd__o22ai_1 U31873 ( .A1(n27461), .A2(n25981), .B1(n27836), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N3165) );
  sky130_fd_sc_hd__o22ai_1 U31874 ( .A1(n27461), .A2(n25982), .B1(n27837), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N3017) );
  sky130_fd_sc_hd__o22ai_1 U31875 ( .A1(n27461), .A2(n26894), .B1(n27839), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N2906) );
  sky130_fd_sc_hd__o22ai_1 U31876 ( .A1(n27461), .A2(n25984), .B1(n27840), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N2721) );
  sky130_fd_sc_hd__o22ai_1 U31877 ( .A1(n27461), .A2(n25985), .B1(n27842), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N3091) );
  sky130_fd_sc_hd__o22ai_1 U31878 ( .A1(n27461), .A2(n25986), .B1(n27843), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N2980) );
  sky130_fd_sc_hd__o22ai_1 U31879 ( .A1(n27461), .A2(n25987), .B1(n27844), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N3128) );
  sky130_fd_sc_hd__o22ai_1 U31880 ( .A1(n27461), .A2(n25988), .B1(n27845), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N2832) );
  sky130_fd_sc_hd__o22ai_1 U31881 ( .A1(n27461), .A2(n25989), .B1(n27846), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N2758) );
  sky130_fd_sc_hd__nand3_1 U31882 ( .A(n26868), .B(n26867), .C(n26866), .Y(
        n26869) );
  sky130_fd_sc_hd__nand2_1 U31883 ( .A(n26869), .B(n27717), .Y(n26870) );
  sky130_fd_sc_hd__nand3_1 U31884 ( .A(n26872), .B(n26871), .C(n26870), .Y(
        n10651) );
  sky130_fd_sc_hd__nand2_1 U31885 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[14]), .Y(n26873) );
  sky130_fd_sc_hd__o21ai_1 U31886 ( .A1(n26875), .A2(n28289), .B1(n26873), .Y(
        n127) );
  sky130_fd_sc_hd__nand2_1 U31887 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[14]), .Y(n26874) );
  sky130_fd_sc_hd__a22oi_1 U31889 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[14]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[14]), 
        .Y(n26877) );
  sky130_fd_sc_hd__a22oi_1 U31890 ( .A1(n28297), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[14]), 
        .B1(n28301), .B2(j202_soc_core_cmt_core_00_const0[14]), .Y(n26876) );
  sky130_fd_sc_hd__nand2_1 U31891 ( .A(n26877), .B(n26876), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[14]) );
  sky130_fd_sc_hd__nand2_1 U31892 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[14]), .Y(n26878) );
  sky130_fd_sc_hd__o22ai_1 U31894 ( .A1(n29144), .A2(n28310), .B1(n26880), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U31895 ( .A1(n29144), .A2(n28313), .B1(n26881), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U31896 ( .A1(n29144), .A2(n28316), .B1(n26882), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U31897 ( .A1(n29144), .A2(n28553), .B1(n26883), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U31898 ( .A1(n29144), .A2(n29082), .B1(n26884), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U31899 ( .A1(n29144), .A2(n29076), .B1(n26885), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__a22oi_1 U31900 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[14]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[14]), .Y(n26887) );
  sky130_fd_sc_hd__a22oi_1 U31901 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[83]), .B1(n27398), .B2(
        j202_soc_core_intc_core_00_rg_itgt[67]), .Y(n26886) );
  sky130_fd_sc_hd__nand3_1 U31902 ( .A(n26887), .B(n28238), .C(n26886), .Y(
        n26888) );
  sky130_fd_sc_hd__a21oi_1 U31903 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[110]), .B1(n26888), .Y(n26892) );
  sky130_fd_sc_hd__a22oi_1 U31904 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[91]), .B1(n28331), .B2(
        j202_soc_core_intc_core_00_rg_itgt[75]), .Y(n26891) );
  sky130_fd_sc_hd__a22oi_1 U31905 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[14]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[46]), .B2(n28330), .Y(n26890) );
  sky130_fd_sc_hd__nand2_1 U31906 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[78]), .Y(n26889) );
  sky130_fd_sc_hd__nand4_1 U31907 ( .A(n26892), .B(n26891), .C(n26890), .D(
        n26889), .Y(j202_soc_core_ahb2apb_01_N142) );
  sky130_fd_sc_hd__nor2_1 U31908 ( .A(n29088), .B(n26893), .Y(
        j202_soc_core_wbqspiflash_00_N711) );
  sky130_fd_sc_hd__a22o_1 U31909 ( .A1(n28026), .A2(
        j202_soc_core_wbqspiflash_00_spi_out[14]), .B1(n28025), .B2(
        j202_soc_core_wbqspiflash_00_erased_sector[0]), .X(
        j202_soc_core_wbqspiflash_00_N681) );
  sky130_fd_sc_hd__o22ai_1 U31910 ( .A1(n25977), .A2(n28448), .B1(n28061), 
        .B2(n26897), .Y(j202_soc_core_j22_cpu_rf_N2897) );
  sky130_fd_sc_hd__nand3_1 U31911 ( .A(n26900), .B(n26899), .C(n26898), .Y(
        n26906) );
  sky130_fd_sc_hd__nand2b_1 U31912 ( .A_N(n26906), .B(n26902), .Y(n29311) );
  sky130_fd_sc_hd__nor2_1 U31913 ( .A(n26906), .B(n26903), .Y(n26911) );
  sky130_fd_sc_hd__a22oi_1 U31914 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[10]), .A2(n29390), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[10]), .B2(n29391), .Y(
        n26914) );
  sky130_fd_sc_hd__nand3_1 U31915 ( .A(n26911), .B(n26909), .C(n26908), .Y(
        n28257) );
  sky130_fd_sc_hd__nand2_1 U31916 ( .A(n26911), .B(n26910), .Y(n29310) );
  sky130_fd_sc_hd__o22ai_1 U31917 ( .A1(n28912), .A2(n28257), .B1(io_oeb[30]), 
        .B2(n29310), .Y(n26912) );
  sky130_fd_sc_hd__a21oi_1 U31918 ( .A1(n29389), .A2(la_data_out[10]), .B1(
        n26912), .Y(n26913) );
  sky130_fd_sc_hd__o211ai_1 U31919 ( .A1(n29311), .A2(n28971), .B1(n26914), 
        .C1(n26913), .Y(j202_soc_core_ahb2apb_02_N138) );
  sky130_fd_sc_hd__mux2i_1 U31920 ( .A0(n26965), .A1(n27798), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N313) );
  sky130_fd_sc_hd__nand2_1 U31921 ( .A(n28055), .B(n27773), .Y(n26915) );
  sky130_fd_sc_hd__nand2_1 U31922 ( .A(n26915), .B(n12203), .Y(
        j202_soc_core_j22_cpu_ml_machj[10]) );
  sky130_fd_sc_hd__nand2_1 U31923 ( .A(n26917), .B(n26916), .Y(n26918) );
  sky130_fd_sc_hd__nand2_1 U31924 ( .A(n26921), .B(n26923), .Y(n26963) );
  sky130_fd_sc_hd__o21ai_1 U31925 ( .A1(n11123), .A2(n26923), .B1(n26922), .Y(
        n26960) );
  sky130_fd_sc_hd__nand3_1 U31926 ( .A(n26938), .B(n26924), .C(n27806), .Y(
        n26925) );
  sky130_fd_sc_hd__o21ai_0 U31927 ( .A1(n26927), .A2(n26926), .B1(n26925), .Y(
        n26928) );
  sky130_fd_sc_hd__a21oi_1 U31928 ( .A1(n26930), .A2(n26929), .B1(n26928), .Y(
        n26931) );
  sky130_fd_sc_hd__o21ai_0 U31929 ( .A1(n27851), .A2(n26932), .B1(n26931), .Y(
        n26954) );
  sky130_fd_sc_hd__o21ai_0 U31930 ( .A1(n27816), .A2(n26934), .B1(n26933), .Y(
        n26953) );
  sky130_fd_sc_hd__o2bb2ai_1 U31931 ( .B1(n26937), .B2(n26936), .A1_N(n27788), 
        .A2_N(n26935), .Y(n26952) );
  sky130_fd_sc_hd__o22ai_1 U31932 ( .A1(n27793), .A2(n28473), .B1(n26939), 
        .B2(n26938), .Y(n26940) );
  sky130_fd_sc_hd__a21oi_1 U31933 ( .A1(n26942), .A2(n26941), .B1(n26940), .Y(
        n26950) );
  sky130_fd_sc_hd__o22a_1 U31934 ( .A1(n26944), .A2(n27795), .B1(n27800), .B2(
        n26943), .X(n26949) );
  sky130_fd_sc_hd__nand2_1 U31935 ( .A(n27808), .B(n26945), .Y(n26948) );
  sky130_fd_sc_hd__nand2_1 U31936 ( .A(n27810), .B(n26946), .Y(n26947) );
  sky130_fd_sc_hd__nand4_1 U31937 ( .A(n26950), .B(n26949), .C(n26948), .D(
        n26947), .Y(n26951) );
  sky130_fd_sc_hd__or4_1 U31938 ( .A(n26954), .B(n26953), .C(n26952), .D(
        n26951), .X(n26955) );
  sky130_fd_sc_hd__a21oi_1 U31939 ( .A1(n26956), .A2(n27789), .B1(n26955), .Y(
        n26957) );
  sky130_fd_sc_hd__o21ai_1 U31940 ( .A1(n26926), .A2(n26958), .B1(n26957), .Y(
        n26959) );
  sky130_fd_sc_hd__a21oi_1 U31941 ( .A1(n26961), .A2(n26960), .B1(n26959), .Y(
        n26962) );
  sky130_fd_sc_hd__buf_6 U31942 ( .A(n26964), .X(n27771) );
  sky130_fd_sc_hd__o22ai_1 U31943 ( .A1(n26965), .A2(n26894), .B1(n27839), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N2911) );
  sky130_fd_sc_hd__o22ai_1 U31944 ( .A1(n26965), .A2(n25983), .B1(n27838), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N3059) );
  sky130_fd_sc_hd__o22ai_1 U31945 ( .A1(n26965), .A2(n25977), .B1(n28061), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N2874) );
  sky130_fd_sc_hd__o22ai_1 U31946 ( .A1(n26965), .A2(n25981), .B1(n27836), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N3170) );
  sky130_fd_sc_hd__o22ai_1 U31947 ( .A1(n26965), .A2(n25982), .B1(n27837), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N3022) );
  sky130_fd_sc_hd__o22ai_1 U31948 ( .A1(n26965), .A2(n25964), .B1(n27847), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N2689) );
  sky130_fd_sc_hd__o22ai_1 U31949 ( .A1(n26965), .A2(n25985), .B1(n27842), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N3096) );
  sky130_fd_sc_hd__o22ai_1 U31950 ( .A1(n26965), .A2(n25989), .B1(n27846), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N2763) );
  sky130_fd_sc_hd__nor2_1 U31951 ( .A(n27644), .B(n27771), .Y(
        j202_soc_core_j22_cpu_rf_N2653) );
  sky130_fd_sc_hd__o22ai_1 U31952 ( .A1(n26965), .A2(n25988), .B1(n27845), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N2837) );
  sky130_fd_sc_hd__o22ai_1 U31953 ( .A1(n26965), .A2(n25980), .B1(n27835), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N2800) );
  sky130_fd_sc_hd__o22ai_1 U31954 ( .A1(n26965), .A2(n25979), .B1(n28112), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N3207) );
  sky130_fd_sc_hd__o22ai_1 U31955 ( .A1(n26965), .A2(n25986), .B1(n27843), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N2985) );
  sky130_fd_sc_hd__o22ai_1 U31956 ( .A1(n26965), .A2(n25987), .B1(n27844), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N3133) );
  sky130_fd_sc_hd__o22ai_1 U31957 ( .A1(n26965), .A2(n25984), .B1(n27840), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N2726) );
  sky130_fd_sc_hd__o22ai_1 U31958 ( .A1(n26965), .A2(n25978), .B1(n27834), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N2948) );
  sky130_fd_sc_hd__o22ai_1 U31959 ( .A1(n26965), .A2(n27841), .B1(n24712), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N3244) );
  sky130_fd_sc_hd__nand2_1 U31960 ( .A(n26967), .B(n26966), .Y(n26971) );
  sky130_fd_sc_hd__nand2b_1 U31961 ( .A_N(n26968), .B(
        j202_soc_core_j22_cpu_ml_macl[8]), .Y(n26970) );
  sky130_fd_sc_hd__a21oi_1 U31962 ( .A1(n27768), .A2(
        j202_soc_core_j22_cpu_ml_bufa[8]), .B1(n27766), .Y(n26969) );
  sky130_fd_sc_hd__nand3_1 U31963 ( .A(n26971), .B(n26970), .C(n26969), .Y(
        j202_soc_core_j22_cpu_ml_maclj[8]) );
  sky130_fd_sc_hd__o22ai_1 U31964 ( .A1(n26975), .A2(n25977), .B1(n28061), 
        .B2(n30071), .Y(j202_soc_core_j22_cpu_rf_N2872) );
  sky130_fd_sc_hd__o22ai_1 U31965 ( .A1(n26975), .A2(n27859), .B1(n27858), 
        .B2(n26972), .Y(j202_soc_core_j22_cpu_rf_N3318) );
  sky130_fd_sc_hd__mux2i_1 U31966 ( .A0(n26972), .A1(n26975), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3279) );
  sky130_fd_sc_hd__inv_1 U31967 ( .A(n26973), .Y(n26980) );
  sky130_fd_sc_hd__o22ai_1 U31968 ( .A1(n26976), .A2(n27775), .B1(n27774), 
        .B2(n26975), .Y(n26977) );
  sky130_fd_sc_hd__a21oi_1 U31969 ( .A1(n26978), .A2(n27860), .B1(n26977), .Y(
        n26979) );
  sky130_fd_sc_hd__a21oi_1 U31971 ( .A1(n26982), .A2(
        j202_soc_core_cmt_core_00_cnt1[7]), .B1(
        j202_soc_core_cmt_core_00_cnt1[8]), .Y(n26983) );
  sky130_fd_sc_hd__a21oi_1 U31972 ( .A1(n26990), .A2(n26984), .B1(n27545), .Y(
        n26987) );
  sky130_fd_sc_hd__o22ai_1 U31973 ( .A1(n27530), .A2(n27964), .B1(n26983), 
        .B2(n26987), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[8])
         );
  sky130_fd_sc_hd__nor3_1 U31974 ( .A(j202_soc_core_cmt_core_00_cnt1[9]), .B(
        n26984), .C(n27548), .Y(n26985) );
  sky130_fd_sc_hd__a21oi_1 U31975 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[9]), .A2(n27544), .B1(n26985), 
        .Y(n26986) );
  sky130_fd_sc_hd__nand3_1 U31977 ( .A(n26991), .B(n26990), .C(n26989), .Y(
        n26994) );
  sky130_fd_sc_hd__nand2_1 U31978 ( .A(n26992), .B(
        j202_soc_core_cmt_core_00_cnt1[11]), .Y(n26993) );
  sky130_fd_sc_hd__o211ai_1 U31979 ( .A1(n26996), .A2(n27530), .B1(n26994), 
        .C1(n26993), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[11])
         );
  sky130_fd_sc_hd__nand2_1 U31980 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[11]), .Y(n26995) );
  sky130_fd_sc_hd__o21ai_1 U31981 ( .A1(n26996), .A2(n28291), .B1(n26995), .Y(
        n131) );
  sky130_fd_sc_hd__a22oi_1 U31982 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[11]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[11]), 
        .Y(n26998) );
  sky130_fd_sc_hd__a22oi_1 U31983 ( .A1(n28297), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[11]), 
        .B1(n28301), .B2(j202_soc_core_cmt_core_00_const0[11]), .Y(n26997) );
  sky130_fd_sc_hd__nand2_1 U31984 ( .A(n26998), .B(n26997), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[11]) );
  sky130_fd_sc_hd__nand2_1 U31985 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[11]), .Y(n26999) );
  sky130_fd_sc_hd__o21ai_1 U31986 ( .A1(n27000), .A2(n28545), .B1(n26999), .Y(
        n57) );
  sky130_fd_sc_hd__o22ai_1 U31987 ( .A1(n29155), .A2(n28310), .B1(n27001), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U31988 ( .A1(n29155), .A2(n28313), .B1(n27002), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U31989 ( .A1(n29155), .A2(n28316), .B1(n27003), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U31990 ( .A1(n29155), .A2(n29082), .B1(n27004), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U31991 ( .A1(n29155), .A2(n29076), .B1(n27005), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__a22oi_1 U31992 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[11]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[11]), .Y(n27007) );
  sky130_fd_sc_hd__a22oi_1 U31993 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[114]), .B1(n27398), .B2(
        j202_soc_core_intc_core_00_rg_itgt[98]), .Y(n27006) );
  sky130_fd_sc_hd__nand3_1 U31994 ( .A(n27007), .B(n28238), .C(n27006), .Y(
        n27008) );
  sky130_fd_sc_hd__a21oi_1 U31995 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[107]), .B1(n27008), .Y(n27012) );
  sky130_fd_sc_hd__a22oi_1 U31996 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[122]), .B1(n28331), .B2(
        j202_soc_core_intc_core_00_rg_itgt[106]), .Y(n27011) );
  sky130_fd_sc_hd__a22oi_1 U31997 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[11]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[43]), .B2(n28330), .Y(n27010) );
  sky130_fd_sc_hd__nand2_1 U31998 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[75]), .Y(n27009) );
  sky130_fd_sc_hd__nand4_1 U31999 ( .A(n27012), .B(n27011), .C(n27010), .D(
        n27009), .Y(j202_soc_core_ahb2apb_01_N139) );
  sky130_fd_sc_hd__o22ai_1 U32000 ( .A1(n28913), .A2(n28257), .B1(n28978), 
        .B2(n29311), .Y(n27013) );
  sky130_fd_sc_hd__a21oi_1 U32001 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[11]), .A2(n29391), .B1(
        n27013), .Y(n27015) );
  sky130_fd_sc_hd__a22oi_1 U32002 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[11]), .A2(n29390), .B1(
        n29389), .B2(la_data_out[11]), .Y(n27014) );
  sky130_fd_sc_hd__o211ai_1 U32003 ( .A1(n29310), .A2(io_oeb[31]), .B1(n27015), 
        .C1(n27014), .Y(j202_soc_core_ahb2apb_02_N139) );
  sky130_fd_sc_hd__mux2i_1 U32004 ( .A0(n28113), .A1(n27025), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N314) );
  sky130_fd_sc_hd__nand2_1 U32005 ( .A(n28055), .B(n27016), .Y(n27018) );
  sky130_fd_sc_hd__nand2_1 U32006 ( .A(n28056), .B(n21280), .Y(n27017) );
  sky130_fd_sc_hd__nand3_1 U32007 ( .A(n27018), .B(n12203), .C(n27017), .Y(
        j202_soc_core_j22_cpu_ml_machj[11]) );
  sky130_fd_sc_hd__o22ai_1 U32008 ( .A1(n28113), .A2(n27859), .B1(n27858), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N3322) );
  sky130_fd_sc_hd__o22ai_1 U32009 ( .A1(n27064), .A2(n27775), .B1(n27774), 
        .B2(n27019), .Y(n27062) );
  sky130_fd_sc_hd__a21oi_1 U32010 ( .A1(n27021), .A2(n27052), .B1(n26926), .Y(
        n27056) );
  sky130_fd_sc_hd__nand2_1 U32011 ( .A(n27022), .B(n27056), .Y(n27060) );
  sky130_fd_sc_hd__nand2_1 U32012 ( .A(n27042), .B(n27786), .Y(n27048) );
  sky130_fd_sc_hd__nor2_1 U32013 ( .A(n27048), .B(n27044), .Y(n27050) );
  sky130_fd_sc_hd__nor2_1 U32014 ( .A(n27023), .B(n27815), .Y(n27038) );
  sky130_fd_sc_hd__a21oi_1 U32015 ( .A1(n28463), .A2(n27791), .B1(n27790), .Y(
        n27024) );
  sky130_fd_sc_hd__o22ai_1 U32016 ( .A1(n28463), .A2(n27793), .B1(n27804), 
        .B2(n27024), .Y(n27030) );
  sky130_fd_sc_hd__nor2_1 U32017 ( .A(n27025), .B(n27797), .Y(n27029) );
  sky130_fd_sc_hd__o22ai_1 U32018 ( .A1(n27027), .A2(n27799), .B1(n27026), 
        .B2(n27803), .Y(n27028) );
  sky130_fd_sc_hd__nor3_1 U32019 ( .A(n27030), .B(n27029), .C(n27028), .Y(
        n27036) );
  sky130_fd_sc_hd__a2bb2oi_1 U32020 ( .B1(n27806), .B2(n27031), .A1_N(n27825), 
        .A2_N(n27795), .Y(n27035) );
  sky130_fd_sc_hd__a22oi_1 U32021 ( .A1(n27810), .A2(n27033), .B1(n27808), 
        .B2(n27032), .Y(n27034) );
  sky130_fd_sc_hd__nand4_1 U32022 ( .A(n27814), .B(n27036), .C(n27035), .D(
        n27034), .Y(n27037) );
  sky130_fd_sc_hd__a211o_1 U32023 ( .A1(n27039), .A2(n28463), .B1(n27038), 
        .C1(n27037), .X(n27040) );
  sky130_fd_sc_hd__a21oi_1 U32024 ( .A1(n27067), .A2(n27789), .B1(n27040), .Y(
        n27046) );
  sky130_fd_sc_hd__nand2_1 U32025 ( .A(n27042), .B(n27785), .Y(n27041) );
  sky130_fd_sc_hd__o211ai_1 U32026 ( .A1(n26411), .A2(n27042), .B1(n27787), 
        .C1(n27041), .Y(n27043) );
  sky130_fd_sc_hd__nand3_1 U32027 ( .A(n27047), .B(n27044), .C(n27043), .Y(
        n27045) );
  sky130_fd_sc_hd__o211ai_1 U32028 ( .A1(n27048), .A2(n27047), .B1(n27046), 
        .C1(n27045), .Y(n27049) );
  sky130_fd_sc_hd__nor2_1 U32029 ( .A(n27050), .B(n27049), .Y(n27059) );
  sky130_fd_sc_hd__nor2_1 U32030 ( .A(n27052), .B(n27051), .Y(n27054) );
  sky130_fd_sc_hd__nand3_1 U32031 ( .A(n27055), .B(n27054), .C(n27053), .Y(
        n27057) );
  sky130_fd_sc_hd__nand2_1 U32032 ( .A(n27057), .B(n27056), .Y(n27058) );
  sky130_fd_sc_hd__nand3_2 U32033 ( .A(n27059), .B(n27060), .C(n27058), .Y(
        n27087) );
  sky130_fd_sc_hd__nand2_1 U32034 ( .A(n27087), .B(n27860), .Y(n27061) );
  sky130_fd_sc_hd__o22ai_1 U32036 ( .A1(n27841), .A2(n27019), .B1(n24712), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N3263) );
  sky130_fd_sc_hd__o22ai_1 U32037 ( .A1(n25977), .A2(n27019), .B1(n28061), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N2893) );
  sky130_fd_sc_hd__o22ai_1 U32038 ( .A1(n25978), .A2(n27019), .B1(n27834), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N2967) );
  sky130_fd_sc_hd__o22ai_1 U32039 ( .A1(n25979), .A2(n27019), .B1(n28112), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N3226) );
  sky130_fd_sc_hd__o22ai_1 U32040 ( .A1(n25981), .A2(n27019), .B1(n27836), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N3189) );
  sky130_fd_sc_hd__o22ai_1 U32041 ( .A1(n25982), .A2(n27019), .B1(n27837), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N3041) );
  sky130_fd_sc_hd__o22ai_1 U32042 ( .A1(n25983), .A2(n27019), .B1(n27838), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N3078) );
  sky130_fd_sc_hd__o22ai_1 U32043 ( .A1(n26894), .A2(n27019), .B1(n27839), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N2930) );
  sky130_fd_sc_hd__o22ai_1 U32044 ( .A1(n25984), .A2(n27019), .B1(n27840), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N2745) );
  sky130_fd_sc_hd__o22ai_1 U32045 ( .A1(n25985), .A2(n27019), .B1(n27842), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N3115) );
  sky130_fd_sc_hd__o22ai_1 U32046 ( .A1(n25986), .A2(n27019), .B1(n27843), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N3004) );
  sky130_fd_sc_hd__o22ai_1 U32047 ( .A1(n25987), .A2(n27019), .B1(n27844), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N3152) );
  sky130_fd_sc_hd__o22ai_1 U32048 ( .A1(n25988), .A2(n27019), .B1(n27845), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N2856) );
  sky130_fd_sc_hd__o22ai_1 U32049 ( .A1(n25989), .A2(n27019), .B1(n27846), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N2782) );
  sky130_fd_sc_hd__o22ai_1 U32050 ( .A1(n25964), .A2(n27019), .B1(n27847), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N2708) );
  sky130_fd_sc_hd__o22ai_1 U32051 ( .A1(n27065), .A2(n27850), .B1(n27064), 
        .B2(n27848), .Y(n27066) );
  sky130_fd_sc_hd__a21oi_1 U32052 ( .A1(n27067), .A2(n26068), .B1(n27066), .Y(
        n27068) );
  sky130_fd_sc_hd__o21ai_0 U32053 ( .A1(n27855), .A2(n27019), .B1(n27068), .Y(
        j202_soc_core_j22_cpu_rf_N325) );
  sky130_fd_sc_hd__o22ai_1 U32054 ( .A1(n27859), .A2(n27019), .B1(n27858), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N3339) );
  sky130_fd_sc_hd__nand2_1 U32055 ( .A(n27994), .B(j202_soc_core_uart_div0[3]), 
        .Y(n27069) );
  sky130_fd_sc_hd__o21ai_1 U32056 ( .A1(n27994), .A2(n27070), .B1(n27069), .Y(
        n70) );
  sky130_fd_sc_hd__o22ai_1 U32057 ( .A1(n27078), .A2(n28310), .B1(n27071), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U32058 ( .A1(n27078), .A2(n28313), .B1(n27072), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U32059 ( .A1(n27078), .A2(n28316), .B1(n27073), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U32060 ( .A1(n27078), .A2(n28064), .B1(n27074), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U32061 ( .A1(n27078), .A2(n28553), .B1(n27075), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U32062 ( .A1(n27078), .A2(n29082), .B1(n27076), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U32063 ( .A1(n27078), .A2(n29076), .B1(n27077), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__a21oi_1 U32064 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[126]), .B1(n28326), .Y(n27086) );
  sky130_fd_sc_hd__nand2_1 U32065 ( .A(n28236), .B(
        j202_soc_core_intc_core_00_rg_ie[27]), .Y(n27081) );
  sky130_fd_sc_hd__a22oi_1 U32066 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[118]), .B1(n27398), .B2(
        j202_soc_core_intc_core_00_rg_itgt[102]), .Y(n27080) );
  sky130_fd_sc_hd__nand2_1 U32067 ( .A(n28331), .B(
        j202_soc_core_intc_core_00_rg_itgt[110]), .Y(n27079) );
  sky130_fd_sc_hd__nand3_1 U32068 ( .A(n27081), .B(n27080), .C(n27079), .Y(
        n27082) );
  sky130_fd_sc_hd__a21oi_1 U32069 ( .A1(j202_soc_core_intc_core_00_rg_ipr[59]), 
        .A2(n28330), .B1(n27082), .Y(n27085) );
  sky130_fd_sc_hd__a22oi_1 U32070 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[27]), .B1(n28329), .B2(
        j202_soc_core_intc_core_00_rg_ipr[123]), .Y(n27084) );
  sky130_fd_sc_hd__nand2_1 U32071 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[91]), .Y(n27083) );
  sky130_fd_sc_hd__nand4_1 U32072 ( .A(n27086), .B(n27085), .C(n27084), .D(
        n27083), .Y(j202_soc_core_ahb2apb_01_N155) );
  sky130_fd_sc_hd__a22o_1 U32073 ( .A1(n28026), .A2(
        j202_soc_core_wbqspiflash_00_spi_out[27]), .B1(n28025), .B2(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled), .X(
        j202_soc_core_wbqspiflash_00_N694) );
  sky130_fd_sc_hd__nand2_1 U32074 ( .A(n27087), .B(n24832), .Y(n27088) );
  sky130_fd_sc_hd__o21ai_0 U32075 ( .A1(n24832), .A2(n27019), .B1(n27088), .Y(
        j202_soc_core_j22_cpu_rf_N3300) );
  sky130_fd_sc_hd__o22ai_1 U32076 ( .A1(n25980), .A2(n27019), .B1(n27835), 
        .B2(n27089), .Y(j202_soc_core_j22_cpu_rf_N2819) );
  sky130_fd_sc_hd__nand2_1 U32077 ( .A(n27091), .B(n27090), .Y(n27092) );
  sky130_fd_sc_hd__o21ai_1 U32078 ( .A1(n29581), .A2(n27918), .B1(n27094), .Y(
        j202_soc_core_ahb2aqu_00_N163) );
  sky130_fd_sc_hd__nand2_1 U32079 ( .A(n27624), .B(j202_soc_core_uart_div1[0]), 
        .Y(n27095) );
  sky130_fd_sc_hd__o22ai_1 U32081 ( .A1(n29151), .A2(n28316), .B1(n27097), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U32082 ( .A1(n29151), .A2(n28553), .B1(n27098), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U32083 ( .A1(n27658), .A2(n27099), .B1(n29016), 
        .B2(n27656), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U32084 ( .A1(n28235), .A2(n27100), .B1(n29016), 
        .B2(n28233), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__a22oi_1 U32085 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[16]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[16]), .Y(n27102) );
  sky130_fd_sc_hd__a22oi_1 U32086 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[20]), .B1(n27398), .B2(
        j202_soc_core_intc_core_00_rg_itgt[4]), .Y(n27101) );
  sky130_fd_sc_hd__nand3_1 U32087 ( .A(n27102), .B(n28238), .C(n27101), .Y(
        n27103) );
  sky130_fd_sc_hd__a21oi_1 U32088 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[112]), .B1(n27103), .Y(n27107) );
  sky130_fd_sc_hd__a22oi_1 U32089 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[28]), .B1(
        j202_soc_core_intc_core_00_rg_itgt[12]), .B2(n28331), .Y(n27106) );
  sky130_fd_sc_hd__a22oi_1 U32090 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[16]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[48]), .B2(n28330), .Y(n27105) );
  sky130_fd_sc_hd__nand2_1 U32091 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[80]), .Y(n27104) );
  sky130_fd_sc_hd__nand4_1 U32092 ( .A(n27107), .B(n27106), .C(n27105), .D(
        n27104), .Y(j202_soc_core_ahb2apb_01_N144) );
  sky130_fd_sc_hd__nor2_1 U32093 ( .A(n29088), .B(n27108), .Y(
        j202_soc_core_wbqspiflash_00_N713) );
  sky130_fd_sc_hd__a22o_1 U32094 ( .A1(n28026), .A2(
        j202_soc_core_wbqspiflash_00_spi_out[16]), .B1(n28025), .B2(
        j202_soc_core_wbqspiflash_00_erased_sector[2]), .X(
        j202_soc_core_wbqspiflash_00_N683) );
  sky130_fd_sc_hd__nand2_1 U32095 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[16]), .Y(n27109) );
  sky130_fd_sc_hd__o21ai_1 U32096 ( .A1(n27110), .A2(n28545), .B1(n27109), .Y(
        n38) );
  sky130_fd_sc_hd__nand2_1 U32097 ( .A(n27764), .B(n27111), .Y(n27112) );
  sky130_fd_sc_hd__o211ai_1 U32098 ( .A1(n27388), .A2(n28537), .B1(n27112), 
        .C1(n24292), .Y(j202_soc_core_j22_cpu_ml_N319) );
  sky130_fd_sc_hd__o22ai_1 U32099 ( .A1(n26894), .A2(n28537), .B1(n27839), 
        .B2(n12256), .Y(j202_soc_core_j22_cpu_rf_N2918) );
  sky130_fd_sc_hd__o22ai_1 U32100 ( .A1(n25980), .A2(n28537), .B1(n27835), 
        .B2(n28060), .Y(j202_soc_core_j22_cpu_rf_N2807) );
  sky130_fd_sc_hd__o22ai_1 U32101 ( .A1(n25983), .A2(n28537), .B1(n27838), 
        .B2(n28060), .Y(j202_soc_core_j22_cpu_rf_N3066) );
  sky130_fd_sc_hd__o22ai_1 U32102 ( .A1(n25979), .A2(n28537), .B1(n28112), 
        .B2(n28060), .Y(j202_soc_core_j22_cpu_rf_N3214) );
  sky130_fd_sc_hd__o22ai_1 U32103 ( .A1(n25981), .A2(n28537), .B1(n27836), 
        .B2(n12256), .Y(j202_soc_core_j22_cpu_rf_N3177) );
  sky130_fd_sc_hd__o22ai_1 U32104 ( .A1(n25986), .A2(n28537), .B1(n27843), 
        .B2(n12256), .Y(j202_soc_core_j22_cpu_rf_N2992) );
  sky130_fd_sc_hd__o22ai_1 U32105 ( .A1(n25982), .A2(n28537), .B1(n27837), 
        .B2(n28060), .Y(j202_soc_core_j22_cpu_rf_N3029) );
  sky130_fd_sc_hd__o22ai_1 U32106 ( .A1(n25985), .A2(n28537), .B1(n27842), 
        .B2(n28060), .Y(j202_soc_core_j22_cpu_rf_N3103) );
  sky130_fd_sc_hd__o22ai_1 U32107 ( .A1(n25987), .A2(n28537), .B1(n27844), 
        .B2(n28060), .Y(j202_soc_core_j22_cpu_rf_N3140) );
  sky130_fd_sc_hd__o22ai_1 U32108 ( .A1(n25989), .A2(n28537), .B1(n27846), 
        .B2(n12256), .Y(j202_soc_core_j22_cpu_rf_N2770) );
  sky130_fd_sc_hd__o22ai_1 U32109 ( .A1(n25984), .A2(n28537), .B1(n27840), 
        .B2(n28060), .Y(j202_soc_core_j22_cpu_rf_N2733) );
  sky130_fd_sc_hd__o22ai_1 U32110 ( .A1(n25988), .A2(n28537), .B1(n27845), 
        .B2(n12256), .Y(j202_soc_core_j22_cpu_rf_N2844) );
  sky130_fd_sc_hd__o22ai_1 U32111 ( .A1(n25978), .A2(n28537), .B1(n27834), 
        .B2(n28060), .Y(j202_soc_core_j22_cpu_rf_N2955) );
  sky130_fd_sc_hd__o22ai_1 U32112 ( .A1(n26894), .A2(n27114), .B1(n27839), 
        .B2(n27113), .Y(j202_soc_core_j22_cpu_rf_N2920) );
  sky130_fd_sc_hd__a22oi_1 U32113 ( .A1(n27115), .A2(n27764), .B1(n28518), 
        .B2(n28425), .Y(n27116) );
  sky130_fd_sc_hd__nand2_1 U32114 ( .A(n24292), .B(n27116), .Y(
        j202_soc_core_j22_cpu_ml_N321) );
  sky130_fd_sc_hd__nand2_1 U32115 ( .A(n28056), .B(n11392), .Y(n27118) );
  sky130_fd_sc_hd__nand3_1 U32116 ( .A(n11460), .B(n30015), .C(n30127), .Y(
        n27124) );
  sky130_fd_sc_hd__o22ai_1 U32117 ( .A1(n27148), .A2(n27859), .B1(n27858), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N3311) );
  sky130_fd_sc_hd__mux2i_1 U32118 ( .A0(n27146), .A1(n27148), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3272) );
  sky130_fd_sc_hd__nor2_1 U32119 ( .A(n27644), .B(n27146), .Y(
        j202_soc_core_j22_cpu_rf_N2644) );
  sky130_fd_sc_hd__o22ai_1 U32120 ( .A1(n27148), .A2(n27841), .B1(n24712), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N3235) );
  sky130_fd_sc_hd__o22ai_1 U32121 ( .A1(n27148), .A2(n25977), .B1(n28061), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N2865) );
  sky130_fd_sc_hd__o22ai_1 U32122 ( .A1(n27148), .A2(n25978), .B1(n27834), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N2939) );
  sky130_fd_sc_hd__o22ai_1 U32123 ( .A1(n27148), .A2(n25979), .B1(n28112), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N3198) );
  sky130_fd_sc_hd__o22ai_1 U32124 ( .A1(n27148), .A2(n25980), .B1(n27835), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N2791) );
  sky130_fd_sc_hd__o22ai_1 U32125 ( .A1(n27148), .A2(n25981), .B1(n27836), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N3161) );
  sky130_fd_sc_hd__o22ai_1 U32126 ( .A1(n27148), .A2(n25982), .B1(n27837), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N3013) );
  sky130_fd_sc_hd__o22ai_1 U32127 ( .A1(n27148), .A2(n25983), .B1(n27838), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N3050) );
  sky130_fd_sc_hd__o22ai_1 U32128 ( .A1(n27148), .A2(n25984), .B1(n27840), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N2717) );
  sky130_fd_sc_hd__o22ai_1 U32129 ( .A1(n27148), .A2(n25985), .B1(n27842), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N3087) );
  sky130_fd_sc_hd__o22ai_1 U32130 ( .A1(n27148), .A2(n25986), .B1(n27843), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N2976) );
  sky130_fd_sc_hd__o22ai_1 U32131 ( .A1(n27148), .A2(n25987), .B1(n27844), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N3124) );
  sky130_fd_sc_hd__o22ai_1 U32132 ( .A1(n27148), .A2(n25988), .B1(n27845), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N2828) );
  sky130_fd_sc_hd__o22ai_1 U32133 ( .A1(n27148), .A2(n25989), .B1(n27846), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N2754) );
  sky130_fd_sc_hd__o22ai_1 U32134 ( .A1(n27148), .A2(n25964), .B1(n27847), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N2680) );
  sky130_fd_sc_hd__o21ai_0 U32135 ( .A1(n27648), .A2(n27146), .B1(n27126), .Y(
        j202_soc_core_j22_cpu_rf_N3347) );
  sky130_fd_sc_hd__nand2_1 U32136 ( .A(n27624), .B(j202_soc_core_uart_div1[2]), 
        .Y(n27127) );
  sky130_fd_sc_hd__o22ai_1 U32138 ( .A1(n29153), .A2(n28310), .B1(n27129), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U32139 ( .A1(n29153), .A2(n28313), .B1(n27130), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U32140 ( .A1(n29153), .A2(n28316), .B1(n27131), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U32141 ( .A1(n29153), .A2(n29082), .B1(n27132), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U32142 ( .A1(n29153), .A2(n29076), .B1(n27133), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__a22oi_1 U32143 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[18]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[18]), .Y(n27135) );
  sky130_fd_sc_hd__a22oi_1 U32144 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[84]), .B1(n27398), .B2(
        j202_soc_core_intc_core_00_rg_itgt[68]), .Y(n27134) );
  sky130_fd_sc_hd__nand3_1 U32145 ( .A(n27135), .B(n28238), .C(n27134), .Y(
        n27136) );
  sky130_fd_sc_hd__a21oi_1 U32146 ( .A1(j202_soc_core_intc_core_00_rg_ipr[50]), 
        .A2(n28330), .B1(n27136), .Y(n27140) );
  sky130_fd_sc_hd__a22oi_1 U32147 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[92]), .B1(n28331), .B2(
        j202_soc_core_intc_core_00_rg_itgt[76]), .Y(n27139) );
  sky130_fd_sc_hd__a22oi_1 U32148 ( .A1(n28321), .A2(
        j202_soc_core_intc_core_00_rg_ipr[82]), .B1(n28329), .B2(
        j202_soc_core_intc_core_00_rg_ipr[114]), .Y(n27138) );
  sky130_fd_sc_hd__nand2_1 U32149 ( .A(n28323), .B(
        j202_soc_core_intc_core_00_rg_ipr[18]), .Y(n27137) );
  sky130_fd_sc_hd__nand4_1 U32150 ( .A(n27140), .B(n27139), .C(n27138), .D(
        n27137), .Y(j202_soc_core_ahb2apb_01_N146) );
  sky130_fd_sc_hd__nor2_1 U32151 ( .A(j202_soc_core_rst), .B(n27141), .Y(
        j202_soc_core_wbqspiflash_00_N715) );
  sky130_fd_sc_hd__a22o_1 U32152 ( .A1(n28026), .A2(
        j202_soc_core_wbqspiflash_00_spi_out[18]), .B1(n28025), .B2(
        j202_soc_core_wbqspiflash_00_erased_sector[4]), .X(
        j202_soc_core_wbqspiflash_00_N685) );
  sky130_fd_sc_hd__nand2_1 U32153 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[18]), .Y(n27142) );
  sky130_fd_sc_hd__o21ai_1 U32154 ( .A1(n27143), .A2(n28545), .B1(n27142), .Y(
        n62) );
  sky130_fd_sc_hd__nand2_1 U32155 ( .A(n28055), .B(n27144), .Y(n27145) );
  sky130_fd_sc_hd__nand2_1 U32156 ( .A(n27145), .B(n12203), .Y(
        j202_soc_core_j22_cpu_ml_machj[2]) );
  sky130_fd_sc_hd__o22ai_1 U32157 ( .A1(n27148), .A2(n26894), .B1(n27839), 
        .B2(n27146), .Y(j202_soc_core_j22_cpu_rf_N2902) );
  sky130_fd_sc_hd__mux2i_1 U32158 ( .A0(n27148), .A1(n27147), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N305) );
  sky130_fd_sc_hd__o22ai_1 U32159 ( .A1(n29162), .A2(n27575), .B1(n27149), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U32160 ( .A1(n29157), .A2(n27575), .B1(n27150), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U32161 ( .A1(n29159), .A2(n28553), .B1(n27151), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__nand3_1 U32162 ( .A(n27153), .B(n27152), .C(n27576), .Y(
        n27161) );
  sky130_fd_sc_hd__nand2_1 U32163 ( .A(n28501), .B(n27154), .Y(n27157) );
  sky130_fd_sc_hd__nand2_1 U32164 ( .A(n27578), .B(
        j202_soc_core_intr_level__1_), .Y(n27155) );
  sky130_fd_sc_hd__nand3_1 U32165 ( .A(n27157), .B(n27156), .C(n27155), .Y(
        n27158) );
  sky130_fd_sc_hd__a21oi_1 U32166 ( .A1(n27159), .A2(n27576), .B1(n27158), .Y(
        n27160) );
  sky130_fd_sc_hd__nand2_1 U32167 ( .A(n27161), .B(n27160), .Y(
        j202_soc_core_j22_cpu_rf_N3388) );
  sky130_fd_sc_hd__o22ai_1 U32168 ( .A1(n28480), .A2(n25983), .B1(n27838), 
        .B2(n27162), .Y(j202_soc_core_j22_cpu_rf_N3058) );
  sky130_fd_sc_hd__nand2_1 U32169 ( .A(n27994), .B(j202_soc_core_uart_div0[1]), 
        .Y(n27163) );
  sky130_fd_sc_hd__o21ai_1 U32170 ( .A1(n27994), .A2(n27164), .B1(n27163), .Y(
        n135) );
  sky130_fd_sc_hd__o22ai_1 U32171 ( .A1(n27172), .A2(n28310), .B1(n27165), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U32172 ( .A1(n27172), .A2(n28313), .B1(n27166), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U32173 ( .A1(n27172), .A2(n28316), .B1(n27167), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U32174 ( .A1(n27172), .A2(n28064), .B1(n27168), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U32175 ( .A1(n27172), .A2(n28553), .B1(n27169), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U32176 ( .A1(n27172), .A2(n29082), .B1(n27170), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U32177 ( .A1(n27172), .A2(n29076), .B1(n27171), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__a21oi_1 U32178 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[62]), .B1(n28326), .Y(n27180) );
  sky130_fd_sc_hd__nand2_1 U32179 ( .A(n28236), .B(
        j202_soc_core_intc_core_00_rg_ie[25]), .Y(n27175) );
  sky130_fd_sc_hd__a22oi_1 U32180 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[54]), .B1(n27398), .B2(
        j202_soc_core_intc_core_00_rg_itgt[38]), .Y(n27174) );
  sky130_fd_sc_hd__nand2_1 U32181 ( .A(n28331), .B(
        j202_soc_core_intc_core_00_rg_itgt[46]), .Y(n27173) );
  sky130_fd_sc_hd__nand3_1 U32182 ( .A(n27175), .B(n27174), .C(n27173), .Y(
        n27176) );
  sky130_fd_sc_hd__a21oi_1 U32183 ( .A1(j202_soc_core_intc_core_00_rg_ipr[57]), 
        .A2(n28330), .B1(n27176), .Y(n27179) );
  sky130_fd_sc_hd__a22oi_1 U32184 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[25]), .B1(n28329), .B2(
        j202_soc_core_intc_core_00_rg_ipr[121]), .Y(n27178) );
  sky130_fd_sc_hd__nand2_1 U32185 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[89]), .Y(n27177) );
  sky130_fd_sc_hd__nand4_1 U32186 ( .A(n27180), .B(n27179), .C(n27178), .D(
        n27177), .Y(j202_soc_core_ahb2apb_01_N153) );
  sky130_fd_sc_hd__nand3_1 U32187 ( .A(n28861), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .C(
        j202_soc_core_wbqspiflash_00_spi_busy), .Y(n27182) );
  sky130_fd_sc_hd__nor4_1 U32190 ( .A(n28669), .B(n27189), .C(n28730), .D(
        n27220), .Y(n28690) );
  sky130_fd_sc_hd__a21oi_1 U32191 ( .A1(n28690), .A2(n27190), .B1(
        j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N746) );
  sky130_fd_sc_hd__o22ai_1 U32192 ( .A1(n27231), .A2(n27296), .B1(n27264), 
        .B2(n27191), .Y(n27192) );
  sky130_fd_sc_hd__nand2_1 U32193 ( .A(n27192), .B(n28870), .Y(n27218) );
  sky130_fd_sc_hd__nor2_1 U32194 ( .A(j202_soc_core_qspi_wb_addr[3]), .B(
        n28739), .Y(n28676) );
  sky130_fd_sc_hd__nor3_1 U32196 ( .A(
        j202_soc_core_wbqspiflash_00_write_in_progress), .B(
        j202_soc_core_qspi_wb_addr[3]), .C(n27294), .Y(n27199) );
  sky130_fd_sc_hd__nand3_1 U32197 ( .A(n27197), .B(n27407), .C(n27614), .Y(
        n27295) );
  sky130_fd_sc_hd__o21ai_1 U32198 ( .A1(n27288), .A2(n28676), .B1(n27295), .Y(
        n27198) );
  sky130_fd_sc_hd__nor3_1 U32199 ( .A(n27200), .B(n27199), .C(n27198), .Y(
        n27207) );
  sky130_fd_sc_hd__nand2_1 U32200 ( .A(n28729), .B(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled), .Y(n27205) );
  sky130_fd_sc_hd__a31oi_1 U32201 ( .A1(n27203), .A2(n27233), .A3(n27202), 
        .B1(n27201), .Y(n27204) );
  sky130_fd_sc_hd__a31oi_1 U32202 ( .A1(n27219), .A2(n28647), .A3(n27205), 
        .B1(n27204), .Y(n27206) );
  sky130_fd_sc_hd__o21ai_1 U32204 ( .A1(j202_soc_core_wbqspiflash_00_spi_spd), 
        .A2(n27245), .B1(n27246), .Y(n27209) );
  sky130_fd_sc_hd__nand2_1 U32205 ( .A(n27209), .B(n27208), .Y(n27214) );
  sky130_fd_sc_hd__a211oi_1 U32206 ( .A1(n27212), .A2(n27287), .B1(n27211), 
        .C1(n28744), .Y(n27213) );
  sky130_fd_sc_hd__nand4_1 U32207 ( .A(n27214), .B(n27213), .C(n28817), .D(
        n27253), .Y(n27215) );
  sky130_fd_sc_hd__a21oi_1 U32208 ( .A1(n27216), .A2(n27224), .B1(n27215), .Y(
        n27217) );
  sky130_fd_sc_hd__a21oi_1 U32209 ( .A1(n27218), .A2(n27217), .B1(
        j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N724) );
  sky130_fd_sc_hd__a21oi_1 U32210 ( .A1(n27219), .A2(n28688), .B1(n27431), .Y(
        n29087) );
  sky130_fd_sc_hd__nand2_1 U32211 ( .A(n28828), .B(
        j202_soc_core_wbqspiflash_00_spif_data[6]), .Y(n28825) );
  sky130_fd_sc_hd__o21ai_1 U32212 ( .A1(n29087), .A2(n27459), .B1(n28825), .Y(
        j202_soc_core_wbqspiflash_00_N612) );
  sky130_fd_sc_hd__a31oi_1 U32213 ( .A1(j202_soc_core_wbqspiflash_00_state[2]), 
        .A2(j202_soc_core_wbqspiflash_00_spi_valid), .A3(n27221), .B1(n27220), 
        .Y(n27222) );
  sky130_fd_sc_hd__a21oi_1 U32214 ( .A1(n27223), .A2(n27222), .B1(n29088), .Y(
        j202_soc_core_wbqspiflash_00_N750) );
  sky130_fd_sc_hd__nand2_1 U32215 ( .A(n28828), .B(
        j202_soc_core_wbqspiflash_00_spif_data[5]), .Y(n28820) );
  sky130_fd_sc_hd__o21ai_1 U32216 ( .A1(n29087), .A2(n27432), .B1(n28820), .Y(
        j202_soc_core_wbqspiflash_00_N611) );
  sky130_fd_sc_hd__nand2_1 U32217 ( .A(n27224), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n28838) );
  sky130_fd_sc_hd__nor3_1 U32218 ( .A(n27226), .B(n28838), .C(n27225), .Y(
        n27227) );
  sky130_fd_sc_hd__o21ai_1 U32220 ( .A1(n27614), .A2(n27229), .B1(n27289), .Y(
        n27237) );
  sky130_fd_sc_hd__nand2_1 U32221 ( .A(n28647), .B(
        j202_soc_core_wbqspiflash_00_state[4]), .Y(n27266) );
  sky130_fd_sc_hd__or3_1 U32222 ( .A(j202_soc_core_wbqspiflash_00_state[3]), 
        .B(n27266), .C(n27251), .X(n27230) );
  sky130_fd_sc_hd__o21ai_1 U32223 ( .A1(n27232), .A2(n27231), .B1(n27230), .Y(
        n27236) );
  sky130_fd_sc_hd__a31oi_1 U32224 ( .A1(n27234), .A2(n27233), .A3(n27275), 
        .B1(n28863), .Y(n27235) );
  sky130_fd_sc_hd__a211oi_1 U32225 ( .A1(n28843), .A2(n27237), .B1(n27236), 
        .C1(n27235), .Y(n27243) );
  sky130_fd_sc_hd__nor3_1 U32226 ( .A(n28866), .B(n27238), .C(n28865), .Y(
        n28879) );
  sky130_fd_sc_hd__nor2_1 U32227 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[5]), .B(
        j202_soc_core_wbqspiflash_00_spif_data[6]), .Y(n27239) );
  sky130_fd_sc_hd__nor2_1 U32229 ( .A(n27283), .B(n27240), .Y(n27241) );
  sky130_fd_sc_hd__nor4_1 U32230 ( .A(n28814), .B(n28869), .C(n28879), .D(
        n27241), .Y(n27242) );
  sky130_fd_sc_hd__a31oi_1 U32231 ( .A1(n27244), .A2(n27243), .A3(n27242), 
        .B1(j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N728) );
  sky130_fd_sc_hd__nand2_1 U32232 ( .A(n27247), .B(n27246), .Y(n27281) );
  sky130_fd_sc_hd__nor3_1 U32233 ( .A(j202_soc_core_wbqspiflash_00_spi_spd), 
        .B(n27248), .C(n27281), .Y(n27249) );
  sky130_fd_sc_hd__a21oi_1 U32234 ( .A1(n27298), .A2(n27250), .B1(n27249), .Y(
        n27263) );
  sky130_fd_sc_hd__nor2_1 U32235 ( .A(n27266), .B(n27252), .Y(n28851) );
  sky130_fd_sc_hd__a21oi_1 U32236 ( .A1(n27254), .A2(n27253), .B1(n27268), .Y(
        n27255) );
  sky130_fd_sc_hd__nor2_1 U32237 ( .A(n27256), .B(n27255), .Y(n27258) );
  sky130_fd_sc_hd__nand3_1 U32238 ( .A(n27259), .B(n27258), .C(n27257), .Y(
        n27260) );
  sky130_fd_sc_hd__a31oi_1 U32239 ( .A1(n27261), .A2(n28870), .A3(n28851), 
        .B1(n27260), .Y(n27262) );
  sky130_fd_sc_hd__a31oi_1 U32240 ( .A1(n27263), .A2(n27262), .A3(n28747), 
        .B1(n29088), .Y(j202_soc_core_wbqspiflash_00_N726) );
  sky130_fd_sc_hd__o211ai_1 U32241 ( .A1(n27266), .A2(n27265), .B1(n27279), 
        .C1(n27264), .Y(n27270) );
  sky130_fd_sc_hd__o21bai_1 U32242 ( .A1(n27268), .A2(n27267), .B1_N(n28869), 
        .Y(n27269) );
  sky130_fd_sc_hd__a21oi_1 U32243 ( .A1(n28870), .A2(n27270), .B1(n27269), .Y(
        n27277) );
  sky130_fd_sc_hd__nand2_1 U32244 ( .A(n27271), .B(
        j202_soc_core_wbqspiflash_00_write_in_progress), .Y(n27273) );
  sky130_fd_sc_hd__nand4_1 U32245 ( .A(n27275), .B(n27274), .C(n27273), .D(
        n27272), .Y(n27276) );
  sky130_fd_sc_hd__o211ai_1 U32246 ( .A1(n27279), .A2(n27278), .B1(n27277), 
        .C1(n27276), .Y(n27305) );
  sky130_fd_sc_hd__a21oi_1 U32247 ( .A1(n28840), .A2(n27281), .B1(n27280), .Y(
        n27282) );
  sky130_fd_sc_hd__a31oi_1 U32248 ( .A1(n27285), .A2(n27284), .A3(n27283), 
        .B1(n27282), .Y(n27303) );
  sky130_fd_sc_hd__nand2_1 U32249 ( .A(n27287), .B(n27286), .Y(n27302) );
  sky130_fd_sc_hd__a21oi_1 U32250 ( .A1(n27291), .A2(
        j202_soc_core_qspi_wb_addr[2]), .B1(n27290), .Y(n27292) );
  sky130_fd_sc_hd__o21ai_1 U32251 ( .A1(n27294), .A2(n27293), .B1(n27292), .Y(
        n27300) );
  sky130_fd_sc_hd__o21ai_1 U32252 ( .A1(n27297), .A2(n27296), .B1(n27295), .Y(
        n27299) );
  sky130_fd_sc_hd__o21ai_1 U32253 ( .A1(n27300), .A2(n27299), .B1(n27298), .Y(
        n27301) );
  sky130_fd_sc_hd__nand4_1 U32254 ( .A(n27303), .B(n28817), .C(n27302), .D(
        n27301), .Y(n27304) );
  sky130_fd_sc_hd__o21a_1 U32255 ( .A1(n27305), .A2(n27304), .B1(n29830), .X(
        j202_soc_core_wbqspiflash_00_N725) );
  sky130_fd_sc_hd__nor2_1 U32256 ( .A(n27306), .B(n28685), .Y(
        j202_soc_core_wbqspiflash_00_N741) );
  sky130_fd_sc_hd__a21oi_1 U32257 ( .A1(n28780), .A2(
        j202_soc_core_wbqspiflash_00_write_in_progress), .B1(n27307), .Y(
        n27309) );
  sky130_fd_sc_hd__nand2b_1 U32259 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[20]), 
        .B(n29582), .Y(n27314) );
  sky130_fd_sc_hd__nand2_1 U32260 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]), .B(n27310), .Y(n27311) );
  sky130_fd_sc_hd__nand4b_1 U32261 ( .A_N(
        j202_soc_core_intc_core_00_rg_irqc[20]), .B(n27311), .C(
        j202_soc_core_intc_core_00_in_intreq[20]), .D(n12069), .Y(n27313) );
  sky130_fd_sc_hd__a21oi_1 U32262 ( .A1(n27314), .A2(n27313), .B1(n27312), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N23) );
  sky130_fd_sc_hd__mux2i_1 U32263 ( .A0(n27317), .A1(n27316), .S(n23228), .Y(
        n27324) );
  sky130_fd_sc_hd__a22oi_1 U32264 ( .A1(n27321), .A2(n27320), .B1(n30169), 
        .B2(n27318), .Y(n27323) );
  sky130_fd_sc_hd__mux2i_1 U32265 ( .A0(n27324), .A1(n27323), .S(n27322), .Y(
        n27338) );
  sky130_fd_sc_hd__a22oi_1 U32266 ( .A1(n27328), .A2(n27327), .B1(n27326), 
        .B2(n27325), .Y(n27335) );
  sky130_fd_sc_hd__a22oi_1 U32267 ( .A1(n27332), .A2(n27331), .B1(n27330), 
        .B2(n27329), .Y(n27334) );
  sky130_fd_sc_hd__mux2i_1 U32268 ( .A0(n27335), .A1(n27334), .S(n27333), .Y(
        n27337) );
  sky130_fd_sc_hd__mux2i_1 U32269 ( .A0(n27338), .A1(n27337), .S(n27336), .Y(
        n27347) );
  sky130_fd_sc_hd__a21oi_1 U32271 ( .A1(n27342), .A2(n27341), .B1(n27340), .Y(
        n27343) );
  sky130_fd_sc_hd__o21ai_1 U32273 ( .A1(n27347), .A2(n27712), .B1(n27346), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N3) );
  sky130_fd_sc_hd__o22ai_1 U32274 ( .A1(n29073), .A2(n27349), .B1(n27348), 
        .B2(n29070), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N3) );
  sky130_fd_sc_hd__nand2_1 U32275 ( .A(n28066), .B(n27350), .Y(n27351) );
  sky130_fd_sc_hd__nand4b_1 U32276 ( .A_N(
        j202_soc_core_intc_core_00_rg_irqc[3]), .B(n27351), .C(
        j202_soc_core_intc_core_00_in_intreq[3]), .D(n12069), .Y(n27354) );
  sky130_fd_sc_hd__nand2b_1 U32277 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[3]), 
        .B(n29584), .Y(n27353) );
  sky130_fd_sc_hd__a21oi_1 U32278 ( .A1(n27354), .A2(n27353), .B1(n27352), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N6) );
  sky130_fd_sc_hd__a21oi_1 U32279 ( .A1(n27357), .A2(n27356), .B1(n27355), .Y(
        n27358) );
  sky130_fd_sc_hd__nor2_1 U32280 ( .A(n27358), .B(n12352), .Y(n27360) );
  sky130_fd_sc_hd__o22ai_1 U32281 ( .A1(n28059), .A2(n26894), .B1(n27839), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N2904) );
  sky130_fd_sc_hd__o22ai_1 U32282 ( .A1(n28059), .A2(n25980), .B1(n27835), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N2793) );
  sky130_fd_sc_hd__o22ai_1 U32283 ( .A1(n28059), .A2(n25983), .B1(n27838), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N3052) );
  sky130_fd_sc_hd__o22ai_1 U32284 ( .A1(n28059), .A2(n25979), .B1(n28112), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N3200) );
  sky130_fd_sc_hd__o22ai_1 U32285 ( .A1(n28059), .A2(n25986), .B1(n27843), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N2978) );
  sky130_fd_sc_hd__o22ai_1 U32286 ( .A1(n28059), .A2(n25982), .B1(n27837), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N3015) );
  sky130_fd_sc_hd__o22ai_1 U32287 ( .A1(n28059), .A2(n25964), .B1(n27847), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N2682) );
  sky130_fd_sc_hd__o22ai_1 U32288 ( .A1(n28059), .A2(n25989), .B1(n27846), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N2756) );
  sky130_fd_sc_hd__o21ai_0 U32289 ( .A1(n27644), .A2(n12344), .B1(n27364), .Y(
        j202_soc_core_j22_cpu_rf_N2646) );
  sky130_fd_sc_hd__o22ai_1 U32290 ( .A1(n28059), .A2(n27841), .B1(n24712), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N3237) );
  sky130_fd_sc_hd__o22ai_1 U32291 ( .A1(n28059), .A2(n25981), .B1(n27836), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N3163) );
  sky130_fd_sc_hd__o22ai_1 U32292 ( .A1(n28059), .A2(n25985), .B1(n27842), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N3089) );
  sky130_fd_sc_hd__o22ai_1 U32293 ( .A1(n28059), .A2(n25987), .B1(n27844), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N3126) );
  sky130_fd_sc_hd__o22ai_1 U32294 ( .A1(n28059), .A2(n25984), .B1(n27840), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N2719) );
  sky130_fd_sc_hd__o22ai_1 U32295 ( .A1(n28059), .A2(n25988), .B1(n27845), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N2830) );
  sky130_fd_sc_hd__o22ai_1 U32296 ( .A1(n28059), .A2(n25978), .B1(n27834), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N2941) );
  sky130_fd_sc_hd__mux2i_1 U32297 ( .A0(n28059), .A1(n27365), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N307) );
  sky130_fd_sc_hd__nand2_1 U32298 ( .A(n27624), .B(j202_soc_core_uart_div1[4]), 
        .Y(n27366) );
  sky130_fd_sc_hd__o22ai_1 U32300 ( .A1(n29152), .A2(n28316), .B1(n27368), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U32301 ( .A1(n29152), .A2(n28553), .B1(n27369), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U32302 ( .A1(n27658), .A2(n27370), .B1(n29047), 
        .B2(n27656), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U32303 ( .A1(n28235), .A2(n27371), .B1(n29047), 
        .B2(n28233), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__a22oi_1 U32304 ( .A1(n28318), .A2(
        j202_soc_core_intc_core_00_rg_ie[20]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[20]), .Y(n27373) );
  sky130_fd_sc_hd__a22oi_1 U32305 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[21]), .B1(n27398), .B2(
        j202_soc_core_intc_core_00_rg_itgt[5]), .Y(n27372) );
  sky130_fd_sc_hd__nand3_1 U32306 ( .A(n27373), .B(n28238), .C(n27372), .Y(
        n27374) );
  sky130_fd_sc_hd__a21oi_1 U32307 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[116]), .B1(n27374), .Y(n27378) );
  sky130_fd_sc_hd__a22oi_1 U32308 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[29]), .B1(
        j202_soc_core_intc_core_00_rg_itgt[13]), .B2(n28331), .Y(n27377) );
  sky130_fd_sc_hd__a22oi_1 U32309 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[20]), .B1(n28330), .B2(
        j202_soc_core_intc_core_00_rg_ipr[52]), .Y(n27376) );
  sky130_fd_sc_hd__nand2_1 U32310 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[84]), .Y(n27375) );
  sky130_fd_sc_hd__nand4_1 U32311 ( .A(n27378), .B(n27377), .C(n27376), .D(
        n27375), .Y(j202_soc_core_ahb2apb_01_N148) );
  sky130_fd_sc_hd__nor2_1 U32312 ( .A(n29088), .B(n27379), .Y(
        j202_soc_core_wbqspiflash_00_N717) );
  sky130_fd_sc_hd__a22o_1 U32313 ( .A1(n28026), .A2(
        j202_soc_core_wbqspiflash_00_spi_out[20]), .B1(n28025), .B2(
        j202_soc_core_wbqspiflash_00_erased_sector[6]), .X(
        j202_soc_core_wbqspiflash_00_N687) );
  sky130_fd_sc_hd__nand2_1 U32314 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[20]), .Y(n27380) );
  sky130_fd_sc_hd__o21ai_1 U32315 ( .A1(n27381), .A2(n28545), .B1(n27380), .Y(
        n63) );
  sky130_fd_sc_hd__o22a_1 U32316 ( .A1(n27383), .A2(n27382), .B1(n27388), .B2(
        n28505), .X(n27384) );
  sky130_fd_sc_hd__nand2_1 U32317 ( .A(n24292), .B(n27384), .Y(
        j202_soc_core_j22_cpu_ml_N324) );
  sky130_fd_sc_hd__o22ai_1 U32318 ( .A1(n26894), .A2(n28505), .B1(n27839), 
        .B2(n27385), .Y(j202_soc_core_j22_cpu_rf_N2922) );
  sky130_fd_sc_hd__o22ai_1 U32319 ( .A1(n27389), .A2(n26894), .B1(n27839), 
        .B2(n12246), .Y(j202_soc_core_j22_cpu_rf_N2932) );
  sky130_fd_sc_hd__nand2_1 U32320 ( .A(n27764), .B(n27809), .Y(n27387) );
  sky130_fd_sc_hd__o211ai_1 U32321 ( .A1(n27389), .A2(n27388), .B1(n27387), 
        .C1(n24292), .Y(j202_soc_core_j22_cpu_ml_N332) );
  sky130_fd_sc_hd__nand2_1 U32322 ( .A(n27994), .B(j202_soc_core_uart_div0[4]), 
        .Y(n27390) );
  sky130_fd_sc_hd__o21ai_1 U32323 ( .A1(n27994), .A2(n27391), .B1(n27390), .Y(
        n68) );
  sky130_fd_sc_hd__o22ai_1 U32324 ( .A1(n27395), .A2(n28316), .B1(n27392), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U32325 ( .A1(n27395), .A2(n28064), .B1(n27393), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U32326 ( .A1(n27395), .A2(n28553), .B1(n27394), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U32327 ( .A1(n27658), .A2(n27396), .B1(n29062), 
        .B2(n27656), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U32328 ( .A1(n28235), .A2(n27397), .B1(n29062), 
        .B2(n28233), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__a21oi_1 U32329 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[31]), .B1(n28326), .Y(n27406) );
  sky130_fd_sc_hd__nand2_1 U32330 ( .A(n28236), .B(
        j202_soc_core_intc_core_00_rg_ie[28]), .Y(n27401) );
  sky130_fd_sc_hd__a22oi_1 U32331 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[23]), .B1(n27398), .B2(
        j202_soc_core_intc_core_00_rg_itgt[7]), .Y(n27400) );
  sky130_fd_sc_hd__nand2_1 U32332 ( .A(n28331), .B(
        j202_soc_core_intc_core_00_rg_itgt[15]), .Y(n27399) );
  sky130_fd_sc_hd__nand3_1 U32333 ( .A(n27401), .B(n27400), .C(n27399), .Y(
        n27402) );
  sky130_fd_sc_hd__a21oi_1 U32334 ( .A1(n28330), .A2(
        j202_soc_core_intc_core_00_rg_ipr[60]), .B1(n27402), .Y(n27405) );
  sky130_fd_sc_hd__a22oi_1 U32335 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[28]), .B1(n28329), .B2(
        j202_soc_core_intc_core_00_rg_ipr[124]), .Y(n27404) );
  sky130_fd_sc_hd__nand2_1 U32336 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[92]), .Y(n27403) );
  sky130_fd_sc_hd__nand4_1 U32337 ( .A(n27406), .B(n27405), .C(n27404), .D(
        n27403), .Y(j202_soc_core_ahb2apb_01_N156) );
  sky130_fd_sc_hd__a22o_1 U32338 ( .A1(n28026), .A2(
        j202_soc_core_wbqspiflash_00_spi_out[28]), .B1(n28025), .B2(n27407), 
        .X(j202_soc_core_wbqspiflash_00_N695) );
  sky130_fd_sc_hd__nand2_1 U32339 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[5]), .Y(n27408) );
  sky130_fd_sc_hd__o21ai_1 U32340 ( .A1(n27409), .A2(n28545), .B1(n27408), .Y(
        n52) );
  sky130_fd_sc_hd__o22ai_1 U32341 ( .A1(n29159), .A2(n28310), .B1(n27410), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U32342 ( .A1(n29159), .A2(n28313), .B1(n27411), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U32343 ( .A1(n29159), .A2(n28316), .B1(n27412), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U32344 ( .A1(n29159), .A2(n29082), .B1(n27413), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__nor2_1 U32345 ( .A(j202_soc_core_intc_core_00_bs_addr[8]), 
        .B(j202_soc_core_intc_core_00_bs_addr[7]), .Y(n27415) );
  sky130_fd_sc_hd__nand3_1 U32346 ( .A(n27416), .B(n27415), .C(n27414), .Y(
        n29413) );
  sky130_fd_sc_hd__nor2_1 U32347 ( .A(n29414), .B(n29413), .Y(n29409) );
  sky130_fd_sc_hd__nand4_1 U32348 ( .A(n29409), .B(n29406), .C(n29408), .D(
        n27417), .Y(n27425) );
  sky130_fd_sc_hd__nand2_1 U32349 ( .A(n27418), .B(j202_soc_core_pwrite[1]), 
        .Y(n29079) );
  sky130_fd_sc_hd__nand2_1 U32350 ( .A(n29079), .B(n29828), .Y(n29077) );
  sky130_fd_sc_hd__o22ai_1 U32351 ( .A1(n29159), .A2(n29079), .B1(n27419), 
        .B2(n29077), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U32352 ( .A1(n29159), .A2(n29076), .B1(n27420), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__a22o_1 U32353 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[57]), .B1(n28331), .B2(
        j202_soc_core_intc_core_00_rg_itgt[41]), .X(n27424) );
  sky130_fd_sc_hd__a22oi_1 U32354 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[5]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[5]), .Y(n27422) );
  sky130_fd_sc_hd__a22oi_1 U32355 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[49]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[33]), .Y(n27421) );
  sky130_fd_sc_hd__nand3_1 U32356 ( .A(n27422), .B(n28238), .C(n27421), .Y(
        n27423) );
  sky130_fd_sc_hd__a211oi_1 U32357 ( .A1(j202_soc_core_intc_core_00_rg_ipr[69]), .A2(n28321), .B1(n27424), .C1(n27423), .Y(n27428) );
  sky130_fd_sc_hd__a22oi_1 U32358 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[5]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[37]), .B2(n28330), .Y(n27427) );
  sky130_fd_sc_hd__nor2_1 U32359 ( .A(n29088), .B(n27425), .Y(n28319) );
  sky130_fd_sc_hd__a22oi_1 U32360 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[101]), .B1(n28319), .B2(
        j202_soc_core_intc_core_00_rg_eimk[5]), .Y(n27426) );
  sky130_fd_sc_hd__nand3_1 U32361 ( .A(n27428), .B(n27427), .C(n27426), .Y(
        j202_soc_core_ahb2apb_01_N133) );
  sky130_fd_sc_hd__a211oi_1 U32362 ( .A1(n27431), .A2(n27430), .B1(n27429), 
        .C1(n28026), .Y(n28336) );
  sky130_fd_sc_hd__nor2_1 U32363 ( .A(n27432), .B(n28336), .Y(
        j202_soc_core_wbqspiflash_00_N672) );
  sky130_fd_sc_hd__mux2i_1 U32364 ( .A0(n27433), .A1(n11189), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N308) );
  sky130_fd_sc_hd__a21oi_1 U32365 ( .A1(n27479), .A2(
        j202_soc_core_cmt_core_00_cnt0[4]), .B1(
        j202_soc_core_cmt_core_00_cnt0[5]), .Y(n27436) );
  sky130_fd_sc_hd__a22oi_1 U32366 ( .A1(n27486), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[5]), .B1(n29169), .B2(
        j202_soc_core_cmt_core_00_cnt0[5]), .Y(n27435) );
  sky130_fd_sc_hd__o31ai_1 U32367 ( .A1(n27484), .A2(n27437), .A3(n27436), 
        .B1(n27435), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[5])
         );
  sky130_fd_sc_hd__a21oi_1 U32368 ( .A1(n27437), .A2(n27477), .B1(
        j202_soc_core_cmt_core_00_cnt0[6]), .Y(n27439) );
  sky130_fd_sc_hd__o22ai_1 U32369 ( .A1(n27482), .A2(n27465), .B1(n27439), 
        .B2(n27438), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[6])
         );
  sky130_fd_sc_hd__a22oi_1 U32370 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[6]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[6]), .Y(
        n27443) );
  sky130_fd_sc_hd__a22oi_1 U32371 ( .A1(n28297), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[6]), 
        .B1(n28299), .B2(j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[6]), .Y(
        n27442) );
  sky130_fd_sc_hd__nand2_1 U32372 ( .A(n28301), .B(
        j202_soc_core_cmt_core_00_const0[6]), .Y(n27441) );
  sky130_fd_sc_hd__nand2_1 U32373 ( .A(n28300), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[6]), .Y(n27440) );
  sky130_fd_sc_hd__nand4_1 U32374 ( .A(n27443), .B(n27442), .C(n27441), .D(
        n27440), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[6]) );
  sky130_fd_sc_hd__nand2_1 U32375 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[6]), .Y(n27444) );
  sky130_fd_sc_hd__o21ai_1 U32376 ( .A1(n27445), .A2(n28545), .B1(n27444), .Y(
        n53) );
  sky130_fd_sc_hd__o22ai_1 U32377 ( .A1(n29158), .A2(n28310), .B1(n27446), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U32378 ( .A1(n29158), .A2(n28313), .B1(n27447), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U32379 ( .A1(n29158), .A2(n28316), .B1(n27448), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U32380 ( .A1(n29158), .A2(n29082), .B1(n27449), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U32381 ( .A1(n29158), .A2(n29079), .B1(n27450), 
        .B2(n29077), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U32382 ( .A1(n29158), .A2(n29076), .B1(n27451), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__a22o_1 U32383 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[89]), .B1(n28331), .B2(
        j202_soc_core_intc_core_00_rg_itgt[73]), .X(n27455) );
  sky130_fd_sc_hd__a22oi_1 U32384 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[6]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[6]), .Y(n27453) );
  sky130_fd_sc_hd__a22oi_1 U32385 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[81]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[65]), .Y(n27452) );
  sky130_fd_sc_hd__nand3_1 U32386 ( .A(n27453), .B(n28238), .C(n27452), .Y(
        n27454) );
  sky130_fd_sc_hd__a211oi_1 U32387 ( .A1(j202_soc_core_intc_core_00_rg_ipr[70]), .A2(n28321), .B1(n27455), .C1(n27454), .Y(n27458) );
  sky130_fd_sc_hd__a22oi_1 U32388 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[6]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[38]), .B2(n28330), .Y(n27457) );
  sky130_fd_sc_hd__a22oi_1 U32389 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[102]), .B1(n28319), .B2(
        j202_soc_core_intc_core_00_rg_eimk[6]), .Y(n27456) );
  sky130_fd_sc_hd__nand3_1 U32390 ( .A(n27458), .B(n27457), .C(n27456), .Y(
        j202_soc_core_ahb2apb_01_N134) );
  sky130_fd_sc_hd__nor2_1 U32391 ( .A(n27459), .B(n28336), .Y(
        j202_soc_core_wbqspiflash_00_N673) );
  sky130_fd_sc_hd__o22ai_1 U32392 ( .A1(n27461), .A2(n25983), .B1(n27838), 
        .B2(n12471), .Y(j202_soc_core_j22_cpu_rf_N3054) );
  sky130_fd_sc_hd__mux2i_1 U32393 ( .A0(n27461), .A1(n11191), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N309) );
  sky130_fd_sc_hd__nand2_1 U32394 ( .A(n28055), .B(n27462), .Y(n27463) );
  sky130_fd_sc_hd__nand2_1 U32395 ( .A(n27463), .B(n12203), .Y(
        j202_soc_core_j22_cpu_ml_machj[6]) );
  sky130_fd_sc_hd__nand2_1 U32396 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[6]), .Y(n27464) );
  sky130_fd_sc_hd__o21ai_1 U32397 ( .A1(n27465), .A2(n28291), .B1(n27464), .Y(
        n111) );
  sky130_fd_sc_hd__nand2_1 U32398 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[13]), .Y(n27466) );
  sky130_fd_sc_hd__o21ai_1 U32399 ( .A1(n27723), .A2(n28291), .B1(n27466), .Y(
        n132) );
  sky130_fd_sc_hd__nand2_1 U32400 ( .A(n29168), .B(
        j202_soc_core_cmt_core_00_cnt0[0]), .Y(n27468) );
  sky130_fd_sc_hd__a222oi_1 U32401 ( .A1(n27468), .A2(n27467), .B1(n27486), 
        .B2(j202_soc_core_cmt_core_00_wdata_cnt0[0]), .C1(
        j202_soc_core_cmt_core_00_cnt0[0]), .C2(n29169), .Y(n27469) );
  sky130_fd_sc_hd__xor2_1 U32402 ( .A(j202_soc_core_cmt_core_00_cnt0[1]), .B(
        j202_soc_core_cmt_core_00_cnt0[0]), .X(n27470) );
  sky130_fd_sc_hd__a222oi_1 U32403 ( .A1(n27477), .A2(n27470), .B1(n27486), 
        .B2(j202_soc_core_cmt_core_00_wdata_cnt0[1]), .C1(n29169), .C2(
        j202_soc_core_cmt_core_00_cnt0[1]), .Y(n27471) );
  sky130_fd_sc_hd__nand2_1 U32404 ( .A(n29169), .B(
        j202_soc_core_cmt_core_00_cnt0[2]), .Y(n27475) );
  sky130_fd_sc_hd__nand2_1 U32405 ( .A(n27486), .B(
        j202_soc_core_cmt_core_00_wdata_cnt0[2]), .Y(n27474) );
  sky130_fd_sc_hd__o211ai_1 U32406 ( .A1(n27472), .A2(
        j202_soc_core_cmt_core_00_cnt0[2]), .B1(n27477), .C1(n27476), .Y(
        n27473) );
  sky130_fd_sc_hd__nand3_1 U32407 ( .A(n27475), .B(n27474), .C(n27473), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[2]) );
  sky130_fd_sc_hd__a21oi_1 U32408 ( .A1(n27478), .A2(n27477), .B1(
        j202_soc_core_cmt_core_00_cnt0[3]), .Y(n27481) );
  sky130_fd_sc_hd__o22ai_1 U32410 ( .A1(n27482), .A2(n27674), .B1(n27481), 
        .B2(n27488), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[3])
         );
  sky130_fd_sc_hd__nor3_1 U32411 ( .A(n27484), .B(
        j202_soc_core_cmt_core_00_cnt0[4]), .C(n27483), .Y(n27485) );
  sky130_fd_sc_hd__a21oi_1 U32412 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[4]), .A2(n27486), .B1(n27485), 
        .Y(n27487) );
  sky130_fd_sc_hd__o21ai_1 U32413 ( .A1(n27489), .A2(n27488), .B1(n27487), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[4]) );
  sky130_fd_sc_hd__a22oi_1 U32414 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[4]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[4]), .Y(
        n27493) );
  sky130_fd_sc_hd__a22oi_1 U32415 ( .A1(n28297), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[4]), 
        .B1(n28299), .B2(j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[4]), .Y(
        n27492) );
  sky130_fd_sc_hd__nand2_1 U32416 ( .A(n28301), .B(
        j202_soc_core_cmt_core_00_const0[4]), .Y(n27491) );
  sky130_fd_sc_hd__nand2_1 U32417 ( .A(n28300), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[4]), .Y(n27490) );
  sky130_fd_sc_hd__nand4_1 U32418 ( .A(n27493), .B(n27492), .C(n27491), .D(
        n27490), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[4]) );
  sky130_fd_sc_hd__nand2_1 U32419 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[4]), .Y(n27494) );
  sky130_fd_sc_hd__o21ai_1 U32420 ( .A1(n27495), .A2(n28545), .B1(n27494), .Y(
        n51) );
  sky130_fd_sc_hd__o22ai_1 U32421 ( .A1(n29160), .A2(n28316), .B1(n27496), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U32422 ( .A1(n29160), .A2(n28553), .B1(n27497), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U32423 ( .A1(n29160), .A2(n29079), .B1(n27498), 
        .B2(n29077), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U32424 ( .A1(n28235), .A2(n27499), .B1(n28931), 
        .B2(n28233), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__a22o_1 U32425 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[25]), .B1(
        j202_soc_core_intc_core_00_rg_itgt[9]), .B2(n28331), .X(n27503) );
  sky130_fd_sc_hd__a22oi_1 U32426 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[4]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[4]), .Y(n27501) );
  sky130_fd_sc_hd__a22oi_1 U32427 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[17]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[1]), .Y(n27500) );
  sky130_fd_sc_hd__nand3_1 U32428 ( .A(n27501), .B(n28238), .C(n27500), .Y(
        n27502) );
  sky130_fd_sc_hd__a211oi_1 U32429 ( .A1(n28321), .A2(
        j202_soc_core_intc_core_00_rg_ipr[68]), .B1(n27503), .C1(n27502), .Y(
        n27506) );
  sky130_fd_sc_hd__a22oi_1 U32430 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[4]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[36]), .B2(n28330), .Y(n27505) );
  sky130_fd_sc_hd__a22oi_1 U32431 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[100]), .B1(n28319), .B2(
        j202_soc_core_intc_core_00_rg_eimk[4]), .Y(n27504) );
  sky130_fd_sc_hd__nand3_1 U32432 ( .A(n27506), .B(n27505), .C(n27504), .Y(
        j202_soc_core_ahb2apb_01_N132) );
  sky130_fd_sc_hd__nor2_1 U32433 ( .A(n28806), .B(n28336), .Y(
        j202_soc_core_wbqspiflash_00_N671) );
  sky130_fd_sc_hd__o22ai_1 U32434 ( .A1(n28059), .A2(n27859), .B1(n27858), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N3314) );
  sky130_fd_sc_hd__mux2i_1 U32435 ( .A0(n12344), .A1(n28059), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3274) );
  sky130_fd_sc_hd__a22oi_1 U32436 ( .A1(n27507), .A2(n27862), .B1(n28508), 
        .B2(n27861), .Y(n27508) );
  sky130_fd_sc_hd__o21ai_0 U32437 ( .A1(n27648), .A2(n12344), .B1(n27508), .Y(
        j202_soc_core_j22_cpu_rf_N3349) );
  sky130_fd_sc_hd__a21oi_1 U32438 ( .A1(j202_soc_core_intr_level__0_), .A2(
        n27578), .B1(n27577), .Y(n27511) );
  sky130_fd_sc_hd__inv_1 U32439 ( .A(n27363), .Y(n27509) );
  sky130_fd_sc_hd__nand2_1 U32440 ( .A(n27509), .B(n27576), .Y(n27510) );
  sky130_fd_sc_hd__o211ai_1 U32441 ( .A1(n28059), .A2(n27580), .B1(n27511), 
        .C1(n27510), .Y(j202_soc_core_j22_cpu_rf_N3386) );
  sky130_fd_sc_hd__nand2_1 U32442 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[9]), .Y(n27512) );
  sky130_fd_sc_hd__o21ai_1 U32443 ( .A1(n27928), .A2(n28289), .B1(n27512), .Y(
        n30) );
  sky130_fd_sc_hd__nand2_1 U32444 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[8]), .Y(n27513) );
  sky130_fd_sc_hd__o21ai_1 U32445 ( .A1(n27964), .A2(n28289), .B1(n27513), .Y(
        n123) );
  sky130_fd_sc_hd__o21ai_1 U32446 ( .A1(n27516), .A2(n27515), .B1(n27514), .Y(
        n27518) );
  sky130_fd_sc_hd__a22oi_1 U32447 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[0]), .A2(n27544), .B1(n29171), 
        .B2(j202_soc_core_cmt_core_00_cnt1[0]), .Y(n27517) );
  sky130_fd_sc_hd__nand2_1 U32448 ( .A(n27518), .B(n27517), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[0]) );
  sky130_fd_sc_hd__nand2_1 U32450 ( .A(n27521), .B(
        j202_soc_core_cmt_core_00_cnt1[1]), .Y(n27520) );
  sky130_fd_sc_hd__nor2_1 U32451 ( .A(n27540), .B(
        j202_soc_core_cmt_core_00_cnt1[1]), .Y(n27522) );
  sky130_fd_sc_hd__a22oi_1 U32452 ( .A1(j202_soc_core_cmt_core_00_cnt1[0]), 
        .A2(n27522), .B1(n27544), .B2(j202_soc_core_cmt_core_00_wdata_cnt0[1]), 
        .Y(n27519) );
  sky130_fd_sc_hd__nand2_1 U32453 ( .A(n27520), .B(n27519), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[1]) );
  sky130_fd_sc_hd__o21ai_1 U32454 ( .A1(n27522), .A2(n27521), .B1(
        j202_soc_core_cmt_core_00_cnt1[2]), .Y(n27526) );
  sky130_fd_sc_hd__nor2_1 U32455 ( .A(n27540), .B(n27523), .Y(n27527) );
  sky130_fd_sc_hd__a22oi_1 U32456 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[2]), .A2(n27544), .B1(n27527), 
        .B2(n27524), .Y(n27525) );
  sky130_fd_sc_hd__nand2_1 U32457 ( .A(n27526), .B(n27525), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[2]) );
  sky130_fd_sc_hd__nand3_1 U32458 ( .A(n27532), .B(
        j202_soc_core_cmt_core_00_cnt1[2]), .C(n27527), .Y(n27529) );
  sky130_fd_sc_hd__nand2_1 U32460 ( .A(n27531), .B(
        j202_soc_core_cmt_core_00_cnt1[3]), .Y(n27528) );
  sky130_fd_sc_hd__o211ai_1 U32461 ( .A1(n27530), .A2(n27674), .B1(n27529), 
        .C1(n27528), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[3])
         );
  sky130_fd_sc_hd__nand2_1 U32462 ( .A(n27531), .B(
        j202_soc_core_cmt_core_00_cnt1[4]), .Y(n27535) );
  sky130_fd_sc_hd__nor3_1 U32463 ( .A(n27540), .B(
        j202_soc_core_cmt_core_00_cnt1[4]), .C(n27532), .Y(n27533) );
  sky130_fd_sc_hd__a21oi_1 U32464 ( .A1(n27544), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[4]), .B1(n27533), .Y(n27534) );
  sky130_fd_sc_hd__nand2_1 U32465 ( .A(n27535), .B(n27534), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[4]) );
  sky130_fd_sc_hd__a21oi_1 U32466 ( .A1(n27537), .A2(
        j202_soc_core_cmt_core_00_cnt1[4]), .B1(
        j202_soc_core_cmt_core_00_cnt1[5]), .Y(n27538) );
  sky130_fd_sc_hd__nor3_1 U32467 ( .A(n27540), .B(n27539), .C(n27538), .Y(
        n27541) );
  sky130_fd_sc_hd__a21oi_1 U32468 ( .A1(n27544), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[5]), .B1(n27541), .Y(n27542) );
  sky130_fd_sc_hd__nand2_1 U32470 ( .A(n27544), .B(
        j202_soc_core_cmt_core_00_wdata_cnt0[7]), .Y(n27547) );
  sky130_fd_sc_hd__nand2_1 U32471 ( .A(n27545), .B(
        j202_soc_core_cmt_core_00_cnt1[7]), .Y(n27546) );
  sky130_fd_sc_hd__o211ai_1 U32472 ( .A1(j202_soc_core_cmt_core_00_cnt1[7]), 
        .A2(n27548), .B1(n27547), .C1(n27546), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[7]) );
  sky130_fd_sc_hd__nand2_1 U32473 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[7]), .Y(n27549) );
  sky130_fd_sc_hd__nand2_1 U32476 ( .A(n27552), .B(n27551), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_nxt_latch_status_0_) );
  sky130_fd_sc_hd__a22oi_1 U32477 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[7]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[7]), .Y(
        n27556) );
  sky130_fd_sc_hd__a22oi_1 U32478 ( .A1(n28297), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[7]), 
        .B1(n28299), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_0_), .Y(
        n27555) );
  sky130_fd_sc_hd__nand2_1 U32479 ( .A(n28301), .B(
        j202_soc_core_cmt_core_00_const0[7]), .Y(n27554) );
  sky130_fd_sc_hd__nand2_1 U32480 ( .A(n28300), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_0_), .Y(
        n27553) );
  sky130_fd_sc_hd__nand4_1 U32481 ( .A(n27556), .B(n27555), .C(n27554), .D(
        n27553), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[7]) );
  sky130_fd_sc_hd__nand2_1 U32482 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[7]), .Y(n27557) );
  sky130_fd_sc_hd__o21ai_1 U32483 ( .A1(n27558), .A2(n28545), .B1(n27557), .Y(
        n54) );
  sky130_fd_sc_hd__o22ai_1 U32484 ( .A1(n29157), .A2(n28310), .B1(n27559), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U32485 ( .A1(n29157), .A2(n28313), .B1(n27560), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U32486 ( .A1(n29157), .A2(n28316), .B1(n27561), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U32487 ( .A1(n29157), .A2(n29082), .B1(n27562), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U32488 ( .A1(n29157), .A2(n29079), .B1(n27563), 
        .B2(n29077), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U32489 ( .A1(n29157), .A2(n29076), .B1(n27564), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__a22o_1 U32490 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[121]), .B1(n28331), .B2(
        j202_soc_core_intc_core_00_rg_itgt[105]), .X(n27568) );
  sky130_fd_sc_hd__a22oi_1 U32491 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[7]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[7]), .Y(n27566) );
  sky130_fd_sc_hd__a22oi_1 U32492 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[113]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[97]), .Y(n27565) );
  sky130_fd_sc_hd__nand3_1 U32493 ( .A(n27566), .B(n28238), .C(n27565), .Y(
        n27567) );
  sky130_fd_sc_hd__a211oi_1 U32494 ( .A1(j202_soc_core_intc_core_00_rg_ipr[71]), .A2(n28321), .B1(n27568), .C1(n27567), .Y(n27571) );
  sky130_fd_sc_hd__a22oi_1 U32495 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[7]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[39]), .B2(n28330), .Y(n27570) );
  sky130_fd_sc_hd__a22oi_1 U32496 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[103]), .B1(n28319), .B2(
        j202_soc_core_intc_core_00_rg_eimk[7]), .Y(n27569) );
  sky130_fd_sc_hd__nand3_1 U32497 ( .A(n27571), .B(n27570), .C(n27569), .Y(
        j202_soc_core_ahb2apb_01_N135) );
  sky130_fd_sc_hd__nor2_1 U32498 ( .A(n28829), .B(n28336), .Y(
        j202_soc_core_wbqspiflash_00_N674) );
  sky130_fd_sc_hd__o22ai_1 U32499 ( .A1(n26894), .A2(n12264), .B1(n27839), 
        .B2(n11115), .Y(j202_soc_core_j22_cpu_rf_N2917) );
  sky130_fd_sc_hd__mux2i_1 U32500 ( .A0(n11115), .A1(n27572), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3287) );
  sky130_fd_sc_hd__o22ai_1 U32501 ( .A1(n29161), .A2(n27575), .B1(n27574), 
        .B2(n27573), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__a21oi_1 U32502 ( .A1(j202_soc_core_intr_level__3_), .A2(
        n27578), .B1(n27577), .Y(n27579) );
  sky130_fd_sc_hd__o21a_1 U32503 ( .A1(n27580), .A2(n11180), .B1(n27579), .X(
        n27581) );
  sky130_fd_sc_hd__o21ai_1 U32504 ( .A1(n27582), .A2(n27988), .B1(n27581), .Y(
        j202_soc_core_j22_cpu_rf_N3392) );
  sky130_fd_sc_hd__nand2_1 U32505 ( .A(n27584), .B(n24832), .Y(n27585) );
  sky130_fd_sc_hd__o21ai_1 U32506 ( .A1(n24832), .A2(n27586), .B1(n27585), .Y(
        j202_soc_core_j22_cpu_rf_N3305) );
  sky130_fd_sc_hd__a22oi_1 U32507 ( .A1(n27587), .A2(n27862), .B1(n12260), 
        .B2(n27861), .Y(n27590) );
  sky130_fd_sc_hd__nand2_1 U32508 ( .A(n27588), .B(n27860), .Y(n27589) );
  sky130_fd_sc_hd__o211ai_1 U32509 ( .A1(n27648), .A2(n27591), .B1(n27590), 
        .C1(n27589), .Y(j202_soc_core_j22_cpu_rf_N3379) );
  sky130_fd_sc_hd__nand2_1 U32510 ( .A(n27994), .B(j202_soc_core_uart_div0[7]), 
        .Y(n27592) );
  sky130_fd_sc_hd__o22ai_1 U32512 ( .A1(n27601), .A2(n28310), .B1(n27594), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U32513 ( .A1(n27601), .A2(n28313), .B1(n27595), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U32514 ( .A1(n27601), .A2(n28316), .B1(n27596), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U32515 ( .A1(n27601), .A2(n28064), .B1(n27597), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U32516 ( .A1(n27601), .A2(n28553), .B1(n27598), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U32517 ( .A1(n27601), .A2(n29082), .B1(n27599), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U32518 ( .A1(n27601), .A2(n29076), .B1(n27600), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__a21oi_1 U32519 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[127]), .B1(n28326), .Y(n27609) );
  sky130_fd_sc_hd__nand2_1 U32520 ( .A(n28236), .B(
        j202_soc_core_intc_core_00_rg_ie[31]), .Y(n27604) );
  sky130_fd_sc_hd__a22oi_1 U32521 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[119]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[103]), .Y(n27603) );
  sky130_fd_sc_hd__nand2_1 U32522 ( .A(n28331), .B(
        j202_soc_core_intc_core_00_rg_itgt[111]), .Y(n27602) );
  sky130_fd_sc_hd__nand3_1 U32523 ( .A(n27604), .B(n27603), .C(n27602), .Y(
        n27605) );
  sky130_fd_sc_hd__a21oi_1 U32524 ( .A1(j202_soc_core_intc_core_00_rg_ipr[63]), 
        .A2(n28330), .B1(n27605), .Y(n27608) );
  sky130_fd_sc_hd__a22oi_1 U32525 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[31]), .B1(n28329), .B2(
        j202_soc_core_intc_core_00_rg_ipr[127]), .Y(n27607) );
  sky130_fd_sc_hd__nand2_1 U32526 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[95]), .Y(n27606) );
  sky130_fd_sc_hd__nand4_1 U32527 ( .A(n27609), .B(n27608), .C(n27607), .D(
        n27606), .Y(j202_soc_core_ahb2apb_01_N159) );
  sky130_fd_sc_hd__a22oi_1 U32528 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[0]), .A2(n27611), .B1(
        j202_soc_core_wbqspiflash_00_spi_out[31]), .B2(n28026), .Y(n27612) );
  sky130_fd_sc_hd__o22ai_1 U32530 ( .A1(n11180), .A2(n26894), .B1(n27839), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N2908) );
  sky130_fd_sc_hd__o22ai_1 U32531 ( .A1(n11180), .A2(n25983), .B1(n27838), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N3056) );
  sky130_fd_sc_hd__o22ai_1 U32532 ( .A1(n11180), .A2(n25979), .B1(n28112), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N3204) );
  sky130_fd_sc_hd__o22ai_1 U32533 ( .A1(n11180), .A2(n25981), .B1(n27836), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N3167) );
  sky130_fd_sc_hd__o22ai_1 U32534 ( .A1(n11180), .A2(n25989), .B1(n27846), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N2760) );
  sky130_fd_sc_hd__o22ai_1 U32535 ( .A1(n11180), .A2(n25984), .B1(n27840), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N2723) );
  sky130_fd_sc_hd__o22ai_1 U32536 ( .A1(n11180), .A2(n25988), .B1(n27845), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N2834) );
  sky130_fd_sc_hd__o22ai_1 U32537 ( .A1(n11180), .A2(n25980), .B1(n27835), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N2797) );
  sky130_fd_sc_hd__o22ai_1 U32538 ( .A1(n11180), .A2(n25986), .B1(n27843), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N2982) );
  sky130_fd_sc_hd__o22ai_1 U32539 ( .A1(n11180), .A2(n25982), .B1(n27837), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N3019) );
  sky130_fd_sc_hd__o22ai_1 U32540 ( .A1(n11180), .A2(n25985), .B1(n27842), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N3093) );
  sky130_fd_sc_hd__o22ai_1 U32541 ( .A1(n11180), .A2(n25987), .B1(n27844), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N3130) );
  sky130_fd_sc_hd__o22ai_1 U32542 ( .A1(n11180), .A2(n25978), .B1(n27834), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N2945) );
  sky130_fd_sc_hd__mux2i_1 U32543 ( .A0(n11180), .A1(n27616), .S(n27615), .Y(
        j202_soc_core_j22_cpu_ml_N310) );
  sky130_fd_sc_hd__nand2_1 U32544 ( .A(n28055), .B(n27617), .Y(n27620) );
  sky130_fd_sc_hd__nand2_1 U32545 ( .A(n28056), .B(n27618), .Y(n27619) );
  sky130_fd_sc_hd__nand3_1 U32546 ( .A(n27620), .B(n12203), .C(n27619), .Y(
        j202_soc_core_j22_cpu_ml_machj[7]) );
  sky130_fd_sc_hd__nand2_1 U32547 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[23]), .Y(n27621) );
  sky130_fd_sc_hd__o21ai_1 U32548 ( .A1(n27622), .A2(n28545), .B1(n27621), .Y(
        n46) );
  sky130_fd_sc_hd__nand2_1 U32549 ( .A(n27624), .B(j202_soc_core_uart_div1[7]), 
        .Y(n27623) );
  sky130_fd_sc_hd__o21ai_1 U32550 ( .A1(n27625), .A2(n27624), .B1(n27623), .Y(
        n97) );
  sky130_fd_sc_hd__o22ai_1 U32551 ( .A1(n27633), .A2(n28310), .B1(n27626), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U32552 ( .A1(n27633), .A2(n28313), .B1(n27627), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U32553 ( .A1(n27633), .A2(n28316), .B1(n27628), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U32554 ( .A1(n27633), .A2(n28064), .B1(n27629), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U32555 ( .A1(n27633), .A2(n28553), .B1(n27630), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U32556 ( .A1(n27633), .A2(n29082), .B1(n27631), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U32557 ( .A1(n27633), .A2(n29076), .B1(n27632), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__a21oi_1 U32558 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[125]), .B1(n28326), .Y(n27641) );
  sky130_fd_sc_hd__nand2_1 U32559 ( .A(n28236), .B(
        j202_soc_core_intc_core_00_rg_ie[23]), .Y(n27636) );
  sky130_fd_sc_hd__a22oi_1 U32560 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[117]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[101]), .Y(n27635) );
  sky130_fd_sc_hd__nand2_1 U32561 ( .A(n28331), .B(
        j202_soc_core_intc_core_00_rg_itgt[109]), .Y(n27634) );
  sky130_fd_sc_hd__nand3_1 U32562 ( .A(n27636), .B(n27635), .C(n27634), .Y(
        n27637) );
  sky130_fd_sc_hd__a21oi_1 U32563 ( .A1(j202_soc_core_intc_core_00_rg_ipr[55]), 
        .A2(n28330), .B1(n27637), .Y(n27640) );
  sky130_fd_sc_hd__a22oi_1 U32564 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[23]), .B1(n28329), .B2(
        j202_soc_core_intc_core_00_rg_ipr[119]), .Y(n27639) );
  sky130_fd_sc_hd__nand2_1 U32565 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[87]), .Y(n27638) );
  sky130_fd_sc_hd__nand4_1 U32566 ( .A(n27641), .B(n27640), .C(n27639), .D(
        n27638), .Y(j202_soc_core_ahb2apb_01_N151) );
  sky130_fd_sc_hd__o22ai_1 U32567 ( .A1(n26894), .A2(n27642), .B1(n27839), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N2933) );
  sky130_fd_sc_hd__o22ai_1 U32568 ( .A1(n25980), .A2(n27642), .B1(n27835), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N2822) );
  sky130_fd_sc_hd__o22ai_1 U32569 ( .A1(n25983), .A2(n27642), .B1(n27838), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N3081) );
  sky130_fd_sc_hd__o22ai_1 U32570 ( .A1(n25979), .A2(n27642), .B1(n28112), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N3229) );
  sky130_fd_sc_hd__o22ai_1 U32571 ( .A1(n25981), .A2(n27642), .B1(n27836), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N3192) );
  sky130_fd_sc_hd__o22ai_1 U32572 ( .A1(n25986), .A2(n27642), .B1(n27843), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N3007) );
  sky130_fd_sc_hd__o22ai_1 U32573 ( .A1(n25982), .A2(n27642), .B1(n27837), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N3044) );
  sky130_fd_sc_hd__o22ai_1 U32574 ( .A1(n25985), .A2(n27642), .B1(n27842), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N3118) );
  sky130_fd_sc_hd__o22ai_1 U32575 ( .A1(n25987), .A2(n27642), .B1(n27844), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N3155) );
  sky130_fd_sc_hd__o22ai_1 U32576 ( .A1(n25989), .A2(n27642), .B1(n27846), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N2785) );
  sky130_fd_sc_hd__o22ai_1 U32577 ( .A1(n25984), .A2(n27642), .B1(n27840), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N2748) );
  sky130_fd_sc_hd__o22ai_1 U32578 ( .A1(n25988), .A2(n27642), .B1(n27845), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N2859) );
  sky130_fd_sc_hd__o22ai_1 U32579 ( .A1(n25978), .A2(n27642), .B1(n27834), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N2970) );
  sky130_fd_sc_hd__o22ai_1 U32580 ( .A1(n25977), .A2(n27642), .B1(n28061), 
        .B2(n27643), .Y(j202_soc_core_j22_cpu_rf_N2896) );
  sky130_fd_sc_hd__o22ai_1 U32581 ( .A1(n27668), .A2(n27859), .B1(n27858), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N3307) );
  sky130_fd_sc_hd__nor2_1 U32582 ( .A(n27644), .B(n27669), .Y(
        j202_soc_core_j22_cpu_rf_N2642) );
  sky130_fd_sc_hd__o22ai_1 U32583 ( .A1(n27668), .A2(n27841), .B1(n24712), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N3233) );
  sky130_fd_sc_hd__o22ai_1 U32584 ( .A1(n27668), .A2(n25977), .B1(n28061), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N2863) );
  sky130_fd_sc_hd__o22ai_1 U32585 ( .A1(n27668), .A2(n25978), .B1(n27834), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N2937) );
  sky130_fd_sc_hd__o22ai_1 U32586 ( .A1(n27668), .A2(n25979), .B1(n28112), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N3196) );
  sky130_fd_sc_hd__o22ai_1 U32587 ( .A1(n27668), .A2(n25980), .B1(n27835), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N2789) );
  sky130_fd_sc_hd__o22ai_1 U32588 ( .A1(n27668), .A2(n25981), .B1(n27836), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N3159) );
  sky130_fd_sc_hd__o22ai_1 U32589 ( .A1(n27668), .A2(n25982), .B1(n27837), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N3011) );
  sky130_fd_sc_hd__o22ai_1 U32590 ( .A1(n27668), .A2(n25983), .B1(n27838), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N3048) );
  sky130_fd_sc_hd__o22ai_1 U32591 ( .A1(n27668), .A2(n25984), .B1(n27840), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N2715) );
  sky130_fd_sc_hd__o22ai_1 U32592 ( .A1(n27668), .A2(n25985), .B1(n27842), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N3085) );
  sky130_fd_sc_hd__o22ai_1 U32593 ( .A1(n27668), .A2(n25986), .B1(n27843), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N2974) );
  sky130_fd_sc_hd__o22ai_1 U32594 ( .A1(n27668), .A2(n25987), .B1(n27844), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N3122) );
  sky130_fd_sc_hd__o22ai_1 U32595 ( .A1(n27668), .A2(n25988), .B1(n27845), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N2826) );
  sky130_fd_sc_hd__o22ai_1 U32596 ( .A1(n27668), .A2(n25989), .B1(n27846), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N2752) );
  sky130_fd_sc_hd__o22ai_1 U32597 ( .A1(n27668), .A2(n25964), .B1(n27847), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N2678) );
  sky130_fd_sc_hd__a22oi_1 U32598 ( .A1(j202_soc_core_j22_cpu_pc[0]), .A2(
        n27862), .B1(n11442), .B2(n27861), .Y(n27647) );
  sky130_fd_sc_hd__nand2_1 U32599 ( .A(n27645), .B(n27772), .Y(n27646) );
  sky130_fd_sc_hd__o211ai_1 U32600 ( .A1(n27649), .A2(n27648), .B1(n27647), 
        .C1(n27646), .Y(j202_soc_core_j22_cpu_rf_N3345) );
  sky130_fd_sc_hd__nand2_1 U32601 ( .A(n27994), .B(j202_soc_core_uart_div0[0]), 
        .Y(n27650) );
  sky130_fd_sc_hd__o22ai_1 U32603 ( .A1(n27655), .A2(n28316), .B1(n27652), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U32604 ( .A1(n27655), .A2(n28064), .B1(n27653), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U32605 ( .A1(n27655), .A2(n28553), .B1(n27654), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U32606 ( .A1(n27658), .A2(n27657), .B1(n29054), 
        .B2(n27656), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U32607 ( .A1(n28235), .A2(n27659), .B1(n29054), 
        .B2(n28233), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__a21oi_1 U32608 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[30]), .B1(n28326), .Y(n27667) );
  sky130_fd_sc_hd__nand2_1 U32609 ( .A(n28318), .B(
        j202_soc_core_intc_core_00_rg_ie[24]), .Y(n27662) );
  sky130_fd_sc_hd__a22oi_1 U32610 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[22]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[6]), .Y(n27661) );
  sky130_fd_sc_hd__nand2_1 U32611 ( .A(n28331), .B(
        j202_soc_core_intc_core_00_rg_itgt[14]), .Y(n27660) );
  sky130_fd_sc_hd__nand3_1 U32612 ( .A(n27662), .B(n27661), .C(n27660), .Y(
        n27663) );
  sky130_fd_sc_hd__a21oi_1 U32613 ( .A1(j202_soc_core_intc_core_00_rg_ipr[56]), 
        .A2(n28330), .B1(n27663), .Y(n27666) );
  sky130_fd_sc_hd__a22oi_1 U32614 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[24]), .B1(n28329), .B2(
        j202_soc_core_intc_core_00_rg_ipr[120]), .Y(n27665) );
  sky130_fd_sc_hd__nand2_1 U32615 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[88]), .Y(n27664) );
  sky130_fd_sc_hd__nand4_1 U32616 ( .A(n27667), .B(n27666), .C(n27665), .D(
        n27664), .Y(j202_soc_core_ahb2apb_01_N152) );
  sky130_fd_sc_hd__o22ai_1 U32617 ( .A1(n27668), .A2(n26894), .B1(n27839), 
        .B2(n27669), .Y(j202_soc_core_j22_cpu_rf_N2900) );
  sky130_fd_sc_hd__mux2i_1 U32618 ( .A0(n27669), .A1(n27668), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3270) );
  sky130_fd_sc_hd__mux2i_1 U32619 ( .A0(n24791), .A1(n24788), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3271) );
  sky130_fd_sc_hd__nand2_1 U32620 ( .A(n28287), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[3]), .Y(n27670) );
  sky130_fd_sc_hd__o21ai_1 U32621 ( .A1(n27674), .A2(n28287), .B1(n27670), .Y(
        n78) );
  sky130_fd_sc_hd__nand2_1 U32622 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[3]), .Y(n27671) );
  sky130_fd_sc_hd__o21ai_1 U32623 ( .A1(n27674), .A2(n28289), .B1(n27671), .Y(
        n80) );
  sky130_fd_sc_hd__nand2_1 U32624 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[3]), .Y(n27672) );
  sky130_fd_sc_hd__o21ai_1 U32625 ( .A1(n27674), .A2(n28291), .B1(n27672), .Y(
        n79) );
  sky130_fd_sc_hd__nand2_1 U32626 ( .A(n28293), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[3]), .Y(n27673) );
  sky130_fd_sc_hd__a22oi_1 U32628 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[3]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[3]), .Y(
        n27678) );
  sky130_fd_sc_hd__a22oi_1 U32629 ( .A1(n28297), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[3]), 
        .B1(n28299), .B2(j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[3]), .Y(
        n27677) );
  sky130_fd_sc_hd__nand2_1 U32630 ( .A(n28301), .B(
        j202_soc_core_cmt_core_00_const0[3]), .Y(n27676) );
  sky130_fd_sc_hd__nand2_1 U32631 ( .A(n28300), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[3]), .Y(n27675) );
  sky130_fd_sc_hd__nand4_1 U32632 ( .A(n27678), .B(n27677), .C(n27676), .D(
        n27675), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[3]) );
  sky130_fd_sc_hd__nand2_1 U32633 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[3]), .Y(n27679) );
  sky130_fd_sc_hd__o21ai_1 U32634 ( .A1(n27680), .A2(n28545), .B1(n27679), .Y(
        n50) );
  sky130_fd_sc_hd__o22ai_1 U32635 ( .A1(n29161), .A2(n28310), .B1(n27681), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U32636 ( .A1(n29161), .A2(n28313), .B1(n27682), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U32637 ( .A1(n29161), .A2(n28316), .B1(n27683), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U32638 ( .A1(n29161), .A2(n28553), .B1(n27684), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U32639 ( .A1(n29161), .A2(n29082), .B1(n27685), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U32640 ( .A1(n29161), .A2(n29079), .B1(n27686), 
        .B2(n29077), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U32641 ( .A1(n29161), .A2(n29076), .B1(n27687), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__a22o_1 U32642 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[120]), .B1(n28331), .B2(
        j202_soc_core_intc_core_00_rg_itgt[104]), .X(n27691) );
  sky130_fd_sc_hd__a22oi_1 U32643 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[3]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[3]), .Y(n27689) );
  sky130_fd_sc_hd__a22oi_1 U32644 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[112]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[96]), .Y(n27688) );
  sky130_fd_sc_hd__nand3_1 U32645 ( .A(n27689), .B(n28238), .C(n27688), .Y(
        n27690) );
  sky130_fd_sc_hd__a211oi_1 U32646 ( .A1(n28321), .A2(
        j202_soc_core_intc_core_00_rg_ipr[67]), .B1(n27691), .C1(n27690), .Y(
        n27694) );
  sky130_fd_sc_hd__a22oi_1 U32647 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[3]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[35]), .B2(n28330), .Y(n27693) );
  sky130_fd_sc_hd__a22oi_1 U32648 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[99]), .B1(n28319), .B2(
        j202_soc_core_intc_core_00_rg_eimk[3]), .Y(n27692) );
  sky130_fd_sc_hd__nand3_1 U32649 ( .A(n27694), .B(n27693), .C(n27692), .Y(
        j202_soc_core_ahb2apb_01_N131) );
  sky130_fd_sc_hd__nor2_1 U32650 ( .A(n28898), .B(n27695), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N361) );
  sky130_fd_sc_hd__nor2_1 U32651 ( .A(n28798), .B(n28336), .Y(
        j202_soc_core_wbqspiflash_00_N670) );
  sky130_fd_sc_hd__o22ai_1 U32652 ( .A1(n29150), .A2(n28064), .B1(n27710), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__nand2_1 U32653 ( .A(n27696), .B(n28201), .Y(n27697) );
  sky130_fd_sc_hd__mux2_2 U32654 ( .A0(j202_soc_core_bldc_core_00_wdata[0]), 
        .A1(j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_), .S(
        n27697), .X(n40) );
  sky130_fd_sc_hd__a21oi_1 U32656 ( .A1(n29585), .A2(n28209), .B1(n27698), .Y(
        n39) );
  sky130_fd_sc_hd__nor2_1 U32657 ( .A(
        j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_2), .B(n27699), 
        .Y(n27700) );
  sky130_fd_sc_hd__a22oi_1 U32658 ( .A1(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_0_), .A2(n27701), .B1(n27700), .B2(
        j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1), .Y(n27702)
         );
  sky130_fd_sc_hd__o21ai_1 U32659 ( .A1(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_0_), .A2(
        n27703), .B1(n27702), .Y(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_nxt_latch_status_0_) );
  sky130_fd_sc_hd__nor2_1 U32660 ( .A(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_wen), .B(
        n27703), .Y(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_nxt_bldc_int) );
  sky130_fd_sc_hd__nand2_1 U32661 ( .A(n27704), .B(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[1]), .Y(n27708) );
  sky130_fd_sc_hd__nor2_1 U32662 ( .A(j202_soc_core_intc_core_00_rg_irqc[19]), 
        .B(n29088), .Y(n27707) );
  sky130_fd_sc_hd__nor2_1 U32663 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[19]), 
        .B(n27705), .Y(n27706) );
  sky130_fd_sc_hd__a31oi_1 U32664 ( .A1(n27708), .A2(
        j202_soc_core_intc_core_00_in_intreq[19]), .A3(n27707), .B1(n27706), 
        .Y(n27709) );
  sky130_fd_sc_hd__nor2_1 U32665 ( .A(n27710), .B(n27709), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N22) );
  sky130_fd_sc_hd__o21ai_1 U32666 ( .A1(n27713), .A2(n27712), .B1(n27711), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N6) );
  sky130_fd_sc_hd__nand3_1 U32667 ( .A(n27716), .B(n27715), .C(n27714), .Y(
        n27718) );
  sky130_fd_sc_hd__nand2_1 U32668 ( .A(n27718), .B(n27717), .Y(n27719) );
  sky130_fd_sc_hd__nand3_1 U32669 ( .A(n27721), .B(n27720), .C(n27719), .Y(
        n10655) );
  sky130_fd_sc_hd__nand2_1 U32670 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[13]), .Y(n27722) );
  sky130_fd_sc_hd__o21ai_1 U32671 ( .A1(n27723), .A2(n28289), .B1(n27722), .Y(
        n126) );
  sky130_fd_sc_hd__a22oi_1 U32672 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[13]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[13]), 
        .Y(n27725) );
  sky130_fd_sc_hd__a22oi_1 U32673 ( .A1(n28297), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[13]), 
        .B1(n28301), .B2(j202_soc_core_cmt_core_00_const0[13]), .Y(n27724) );
  sky130_fd_sc_hd__nand2_1 U32674 ( .A(n27725), .B(n27724), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[13]) );
  sky130_fd_sc_hd__nand2_1 U32675 ( .A(n27901), .B(n27740), .Y(n27733) );
  sky130_fd_sc_hd__nand2_1 U32676 ( .A(n27980), .B(n28267), .Y(n27732) );
  sky130_fd_sc_hd__inv_1 U32678 ( .A(n27736), .Y(n27738) );
  sky130_fd_sc_hd__nor2_1 U32679 ( .A(n27738), .B(n27737), .Y(n28138) );
  sky130_fd_sc_hd__o211ai_1 U32680 ( .A1(n12332), .A2(n11395), .B1(n27742), 
        .C1(n27741), .Y(n27744) );
  sky130_fd_sc_hd__nor2_1 U32681 ( .A(n27747), .B(n27746), .Y(n27748) );
  sky130_fd_sc_hd__nand4_1 U32682 ( .A(n27749), .B(n30202), .C(n28138), .D(
        n27748), .Y(n27750) );
  sky130_fd_sc_hd__nand2_1 U32683 ( .A(n27750), .B(n28417), .Y(n27752) );
  sky130_fd_sc_hd__nand2_1 U32684 ( .A(n27752), .B(n27912), .Y(n10632) );
  sky130_fd_sc_hd__mux2i_1 U32685 ( .A0(n24791), .A1(n24788), .S(n27753), .Y(
        j202_soc_core_j22_cpu_rf_N2628) );
  sky130_fd_sc_hd__nand2_1 U32686 ( .A(n29746), .B(n27755), .Y(n27758) );
  sky130_fd_sc_hd__nand4_1 U32688 ( .A(n27757), .B(
        j202_soc_core_j22_cpu_macop_MAC_[1]), .C(n29746), .D(n27756), .Y(
        n27759) );
  sky130_fd_sc_hd__nand3_1 U32689 ( .A(n27759), .B(n28422), .C(n27758), .Y(
        j202_soc_core_j22_cpu_ml_N192) );
  sky130_fd_sc_hd__a21oi_1 U32690 ( .A1(n27761), .A2(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[4]), .B1(n13325), .Y(n27762) );
  sky130_fd_sc_hd__o21ai_1 U32691 ( .A1(n27763), .A2(n28052), .B1(n27762), .Y(
        j202_soc_core_j22_cpu_ml_N156) );
  sky130_fd_sc_hd__a22oi_1 U32692 ( .A1(n27788), .A2(n27764), .B1(n28470), 
        .B2(n28425), .Y(n27765) );
  sky130_fd_sc_hd__nand2_1 U32693 ( .A(n24292), .B(n27765), .Y(
        j202_soc_core_j22_cpu_ml_N330) );
  sky130_fd_sc_hd__a21oi_1 U32694 ( .A1(n27768), .A2(n27767), .B1(n27766), .Y(
        n27769) );
  sky130_fd_sc_hd__o21ai_1 U32695 ( .A1(n27783), .A2(n27770), .B1(n27769), .Y(
        j202_soc_core_j22_cpu_ml_maclj[26]) );
  sky130_fd_sc_hd__o22ai_1 U32696 ( .A1(n26965), .A2(n27859), .B1(n27858), 
        .B2(n27771), .Y(j202_soc_core_j22_cpu_rf_N3321) );
  sky130_fd_sc_hd__mux2i_1 U32697 ( .A0(n27771), .A1(n26965), .S(n23749), .Y(
        j202_soc_core_j22_cpu_rf_N3281) );
  sky130_fd_sc_hd__nand2_1 U32698 ( .A(n27773), .B(n27772), .Y(n27780) );
  sky130_fd_sc_hd__o22ai_1 U32699 ( .A1(n27776), .A2(n27775), .B1(n27774), 
        .B2(n26965), .Y(n27777) );
  sky130_fd_sc_hd__a21oi_1 U32700 ( .A1(n27860), .A2(n27778), .B1(n27777), .Y(
        n27779) );
  sky130_fd_sc_hd__nand2_1 U32701 ( .A(n27780), .B(n27779), .Y(
        j202_soc_core_j22_cpu_rf_N3356) );
  sky130_fd_sc_hd__a21oi_1 U32702 ( .A1(n27783), .A2(n27782), .B1(n26926), .Y(
        n27830) );
  sky130_fd_sc_hd__nand2_1 U32703 ( .A(n27784), .B(n27830), .Y(n27833) );
  sky130_fd_sc_hd__nand2_1 U32705 ( .A(n27853), .B(n27789), .Y(n27821) );
  sky130_fd_sc_hd__a21oi_1 U32706 ( .A1(n28471), .A2(n27791), .B1(n27790), .Y(
        n27792) );
  sky130_fd_sc_hd__o22a_1 U32707 ( .A1(n28471), .A2(n27793), .B1(n27825), .B2(
        n27792), .X(n27794) );
  sky130_fd_sc_hd__o22ai_1 U32709 ( .A1(n27800), .A2(n27799), .B1(n27798), 
        .B2(n27797), .Y(n27801) );
  sky130_fd_sc_hd__nor2_1 U32710 ( .A(n27802), .B(n27801), .Y(n27813) );
  sky130_fd_sc_hd__a2bb2oi_1 U32711 ( .B1(n27806), .B2(n27805), .A1_N(n27804), 
        .A2_N(n27803), .Y(n27812) );
  sky130_fd_sc_hd__a22oi_1 U32712 ( .A1(n27810), .A2(n27809), .B1(n27808), 
        .B2(n27807), .Y(n27811) );
  sky130_fd_sc_hd__nand4_1 U32713 ( .A(n27814), .B(n27813), .C(n27812), .D(
        n27811), .Y(n27819) );
  sky130_fd_sc_hd__o22ai_1 U32714 ( .A1(n27851), .A2(n27817), .B1(n27816), 
        .B2(n27815), .Y(n27818) );
  sky130_fd_sc_hd__nor2_1 U32715 ( .A(n27819), .B(n27818), .Y(n27820) );
  sky130_fd_sc_hd__nand2_1 U32716 ( .A(n27821), .B(n27820), .Y(n27822) );
  sky130_fd_sc_hd__a21oi_1 U32717 ( .A1(n28470), .A2(n27823), .B1(n27822), .Y(
        n27824) );
  sky130_fd_sc_hd__nand4_1 U32718 ( .A(n27829), .B(n27828), .C(n27827), .D(
        n27826), .Y(n27831) );
  sky130_fd_sc_hd__nand2_1 U32719 ( .A(n27831), .B(n27830), .Y(n27832) );
  sky130_fd_sc_hd__o22ai_1 U32720 ( .A1(n25977), .A2(n27897), .B1(n28061), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N2892) );
  sky130_fd_sc_hd__o22ai_1 U32721 ( .A1(n25978), .A2(n27897), .B1(n27834), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N2966) );
  sky130_fd_sc_hd__o22ai_1 U32722 ( .A1(n25979), .A2(n27897), .B1(n28112), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N3225) );
  sky130_fd_sc_hd__o22ai_1 U32723 ( .A1(n25980), .A2(n27897), .B1(n27835), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N2818) );
  sky130_fd_sc_hd__o22ai_1 U32724 ( .A1(n25981), .A2(n27897), .B1(n27836), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N3188) );
  sky130_fd_sc_hd__o22ai_1 U32725 ( .A1(n25983), .A2(n27897), .B1(n27838), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N3077) );
  sky130_fd_sc_hd__o22ai_1 U32726 ( .A1(n26894), .A2(n27897), .B1(n27839), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N2929) );
  sky130_fd_sc_hd__o22ai_1 U32727 ( .A1(n25984), .A2(n27897), .B1(n27840), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N2744) );
  sky130_fd_sc_hd__o22ai_1 U32728 ( .A1(n27841), .A2(n27897), .B1(n24712), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N3262) );
  sky130_fd_sc_hd__o22ai_1 U32729 ( .A1(n25985), .A2(n27897), .B1(n27842), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N3114) );
  sky130_fd_sc_hd__o22ai_1 U32730 ( .A1(n25986), .A2(n27897), .B1(n27843), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N3003) );
  sky130_fd_sc_hd__o22ai_1 U32731 ( .A1(n25987), .A2(n27897), .B1(n27844), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N3151) );
  sky130_fd_sc_hd__o22ai_1 U32732 ( .A1(n25988), .A2(n27897), .B1(n27845), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N2855) );
  sky130_fd_sc_hd__o22ai_1 U32733 ( .A1(n25989), .A2(n27897), .B1(n27846), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N2781) );
  sky130_fd_sc_hd__o22ai_1 U32734 ( .A1(n25964), .A2(n27897), .B1(n27847), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N2707) );
  sky130_fd_sc_hd__o22ai_1 U32735 ( .A1(n27851), .A2(n27850), .B1(n27849), 
        .B2(n27848), .Y(n27852) );
  sky130_fd_sc_hd__a21oi_1 U32736 ( .A1(n27853), .A2(n26068), .B1(n27852), .Y(
        n27854) );
  sky130_fd_sc_hd__o21ai_0 U32737 ( .A1(n27855), .A2(n27897), .B1(n27854), .Y(
        j202_soc_core_j22_cpu_rf_N324) );
  sky130_fd_sc_hd__o22ai_1 U32738 ( .A1(n27859), .A2(n27897), .B1(n27858), 
        .B2(n27857), .Y(j202_soc_core_j22_cpu_rf_N3338) );
  sky130_fd_sc_hd__nand2_1 U32739 ( .A(n27896), .B(n27860), .Y(n27865) );
  sky130_fd_sc_hd__a22oi_1 U32740 ( .A1(n27863), .A2(n27862), .B1(n28470), 
        .B2(n27861), .Y(n27864) );
  sky130_fd_sc_hd__nand2_1 U32741 ( .A(n27865), .B(n27864), .Y(
        j202_soc_core_j22_cpu_rf_N3374) );
  sky130_fd_sc_hd__nand2_1 U32742 ( .A(n27994), .B(j202_soc_core_uart_div0[2]), 
        .Y(n27866) );
  sky130_fd_sc_hd__o22ai_1 U32744 ( .A1(n27875), .A2(n28310), .B1(n27868), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U32745 ( .A1(n27875), .A2(n28313), .B1(n27869), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U32746 ( .A1(n27875), .A2(n28316), .B1(n27870), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U32747 ( .A1(n27875), .A2(n28064), .B1(n27871), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U32748 ( .A1(n27875), .A2(n28553), .B1(n27872), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U32749 ( .A1(n27875), .A2(n29082), .B1(n27873), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U32750 ( .A1(n27875), .A2(n29076), .B1(n27874), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__a21oi_1 U32751 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[94]), .B1(n28326), .Y(n27883) );
  sky130_fd_sc_hd__nand2_1 U32752 ( .A(n28236), .B(
        j202_soc_core_intc_core_00_rg_ie[26]), .Y(n27878) );
  sky130_fd_sc_hd__a22oi_1 U32753 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[86]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[70]), .Y(n27877) );
  sky130_fd_sc_hd__nand2_1 U32754 ( .A(n28331), .B(
        j202_soc_core_intc_core_00_rg_itgt[78]), .Y(n27876) );
  sky130_fd_sc_hd__nand3_1 U32755 ( .A(n27878), .B(n27877), .C(n27876), .Y(
        n27879) );
  sky130_fd_sc_hd__a21oi_1 U32756 ( .A1(j202_soc_core_intc_core_00_rg_ipr[58]), 
        .A2(n28330), .B1(n27879), .Y(n27882) );
  sky130_fd_sc_hd__a22oi_1 U32757 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[26]), .B1(n28329), .B2(
        j202_soc_core_intc_core_00_rg_ipr[122]), .Y(n27881) );
  sky130_fd_sc_hd__nand2_1 U32758 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[90]), .Y(n27880) );
  sky130_fd_sc_hd__nand4_1 U32759 ( .A(n27883), .B(n27882), .C(n27881), .D(
        n27880), .Y(j202_soc_core_ahb2apb_01_N154) );
  sky130_fd_sc_hd__nand3_1 U32760 ( .A(n11173), .B(n27886), .C(n12219), .Y(
        n27887) );
  sky130_fd_sc_hd__nor2_1 U32761 ( .A(n27887), .B(n28033), .Y(n27889) );
  sky130_fd_sc_hd__nand4_1 U32762 ( .A(n24594), .B(n27890), .C(n27889), .D(
        n24592), .Y(n27891) );
  sky130_fd_sc_hd__nand2_1 U32763 ( .A(n27891), .B(n28417), .Y(n27895) );
  sky130_fd_sc_hd__nand2_1 U32764 ( .A(n28198), .B(
        j202_soc_core_j22_cpu_opst[0]), .Y(n28144) );
  sky130_fd_sc_hd__and4_1 U32765 ( .A(n28144), .B(n28155), .C(n28352), .D(
        n27892), .X(n27893) );
  sky130_fd_sc_hd__nand3_1 U32766 ( .A(n27895), .B(n27894), .C(n27893), .Y(
        n10621) );
  sky130_fd_sc_hd__a21boi_1 U32767 ( .A1(n28027), .A2(n11646), .B1_N(n27898), 
        .Y(n27903) );
  sky130_fd_sc_hd__nand2_1 U32768 ( .A(n11729), .B(n27900), .Y(n27902) );
  sky130_fd_sc_hd__nand4_1 U32769 ( .A(n27903), .B(n28387), .C(n12235), .D(
        n27902), .Y(n27907) );
  sky130_fd_sc_hd__nor2_1 U32770 ( .A(n29587), .B(n11007), .Y(n28120) );
  sky130_fd_sc_hd__nor3_1 U32771 ( .A(n27907), .B(n28120), .C(n27906), .Y(
        n27908) );
  sky130_fd_sc_hd__nand4_1 U32773 ( .A(n27913), .B(n27912), .C(n28394), .D(
        n28144), .Y(n10629) );
  sky130_fd_sc_hd__nand2_1 U32774 ( .A(n27915), .B(n27914), .Y(n27917) );
  sky130_fd_sc_hd__nor2_1 U32775 ( .A(n29301), .B(n29278), .Y(n27923) );
  sky130_fd_sc_hd__a21oi_1 U32776 ( .A1(n29301), .A2(n29278), .B1(n27923), .Y(
        n23) );
  sky130_fd_sc_hd__nand2_1 U32777 ( .A(n28910), .B(j202_soc_core_uart_WRTXD1), 
        .Y(n27924) );
  sky130_fd_sc_hd__a21oi_1 U32778 ( .A1(n27921), .A2(n27924), .B1(n27920), .Y(
        n99) );
  sky130_fd_sc_hd__a21o_1 U32779 ( .A1(j202_soc_core_uart_TOP_tx_fifo_wp[1]), 
        .A2(n27922), .B1(n29880), .X(n98) );
  sky130_fd_sc_hd__xor2_1 U32780 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[1]), 
        .B(n27923), .X(n22) );
  sky130_fd_sc_hd__a211o_1 U32781 ( .A1(n27925), .A2(n28584), .B1(n27924), 
        .C1(n28586), .X(n27926) );
  sky130_fd_sc_hd__nor2_1 U32782 ( .A(n29088), .B(n27926), .Y(
        j202_soc_core_uart_TOP_tx_fifo_N42) );
  sky130_fd_sc_hd__nand3_1 U32783 ( .A(n27926), .B(n29301), .C(n29745), .Y(
        j202_soc_core_uart_TOP_tx_fifo_N41) );
  sky130_fd_sc_hd__nand2_1 U32784 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[9]), .Y(n27927) );
  sky130_fd_sc_hd__a22oi_1 U32786 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[9]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[9]), .Y(
        n27930) );
  sky130_fd_sc_hd__a22oi_1 U32787 ( .A1(n28297), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[9]), 
        .B1(n28301), .B2(j202_soc_core_cmt_core_00_const0[9]), .Y(n27929) );
  sky130_fd_sc_hd__nand2_1 U32788 ( .A(n27930), .B(n27929), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[9]) );
  sky130_fd_sc_hd__nand2_1 U32789 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[9]), .Y(n27931) );
  sky130_fd_sc_hd__o22ai_1 U32791 ( .A1(n29148), .A2(n28310), .B1(n27933), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U32792 ( .A1(n29148), .A2(n28313), .B1(n27934), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U32793 ( .A1(n29148), .A2(n28316), .B1(n27935), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U32794 ( .A1(n29148), .A2(n28553), .B1(n27936), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U32795 ( .A1(n29148), .A2(n29082), .B1(n27937), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U32796 ( .A1(n29148), .A2(n29076), .B1(n27938), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__a22oi_1 U32797 ( .A1(n28318), .A2(
        j202_soc_core_intc_core_00_rg_ie[9]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[9]), .Y(n27940) );
  sky130_fd_sc_hd__a22oi_1 U32798 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[50]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[34]), .Y(n27939) );
  sky130_fd_sc_hd__nand3_1 U32799 ( .A(n27940), .B(n28238), .C(n27939), .Y(
        n27941) );
  sky130_fd_sc_hd__a21oi_1 U32800 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[105]), .B1(n27941), .Y(n27945) );
  sky130_fd_sc_hd__a22oi_1 U32801 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[58]), .B1(n28331), .B2(
        j202_soc_core_intc_core_00_rg_itgt[42]), .Y(n27944) );
  sky130_fd_sc_hd__a22oi_1 U32802 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[9]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[41]), .B2(n28330), .Y(n27943) );
  sky130_fd_sc_hd__nand2_1 U32803 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[73]), .Y(n27942) );
  sky130_fd_sc_hd__nand4_1 U32804 ( .A(n27945), .B(n27944), .C(n27943), .D(
        n27942), .Y(j202_soc_core_ahb2apb_01_N137) );
  sky130_fd_sc_hd__o22ai_1 U32805 ( .A1(n28911), .A2(n28257), .B1(n28964), 
        .B2(n29311), .Y(n27946) );
  sky130_fd_sc_hd__a21oi_1 U32806 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[9]), .A2(n29391), .B1(
        n27946), .Y(n27948) );
  sky130_fd_sc_hd__a22oi_1 U32807 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[9]), .A2(n29390), .B1(
        n29389), .B2(la_data_out[9]), .Y(n27947) );
  sky130_fd_sc_hd__o211ai_1 U32808 ( .A1(n29310), .A2(io_oeb[29]), .B1(n27948), 
        .C1(n27947), .Y(j202_soc_core_ahb2apb_02_N137) );
  sky130_fd_sc_hd__nand2_1 U32809 ( .A(n28079), .B(n12669), .Y(n27949) );
  sky130_fd_sc_hd__nand2_1 U32810 ( .A(n28081), .B(n27949), .Y(n10531) );
  sky130_fd_sc_hd__nor2_1 U32811 ( .A(n27951), .B(n27950), .Y(
        j202_soc_core_ahb2aqu_00_N98) );
  sky130_fd_sc_hd__a21oi_1 U32812 ( .A1(n27957), .A2(n27961), .B1(n27952), .Y(
        n105) );
  sky130_fd_sc_hd__a21o_1 U32814 ( .A1(j202_soc_core_uart_TOP_rx_fifo_wp[1]), 
        .A2(n27954), .B1(n29870), .X(n25) );
  sky130_fd_sc_hd__nor2_1 U32815 ( .A(n27955), .B(n27957), .Y(n27956) );
  sky130_fd_sc_hd__a21oi_1 U32816 ( .A1(n27960), .A2(n27957), .B1(n27956), .Y(
        n27959) );
  sky130_fd_sc_hd__o211ai_1 U32817 ( .A1(j202_soc_core_uart_TOP_rx_fifo_wp[0]), 
        .A2(n27960), .B1(n27959), .C1(n27958), .Y(n27962) );
  sky130_fd_sc_hd__nor2_1 U32818 ( .A(n29088), .B(n27962), .Y(
        j202_soc_core_uart_TOP_rx_fifo_N42) );
  sky130_fd_sc_hd__nand3_1 U32819 ( .A(n27962), .B(n29827), .C(n27961), .Y(
        j202_soc_core_uart_TOP_rx_fifo_N41) );
  sky130_fd_sc_hd__nand2_1 U32820 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[8]), .Y(n27963) );
  sky130_fd_sc_hd__o21ai_1 U32821 ( .A1(n27964), .A2(n28291), .B1(n27963), .Y(
        n129) );
  sky130_fd_sc_hd__a22oi_1 U32822 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[8]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[8]), .Y(
        n27966) );
  sky130_fd_sc_hd__a22oi_1 U32823 ( .A1(n28297), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[8]), 
        .B1(n28301), .B2(j202_soc_core_cmt_core_00_const0[8]), .Y(n27965) );
  sky130_fd_sc_hd__nand2_1 U32824 ( .A(n27966), .B(n27965), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[8]) );
  sky130_fd_sc_hd__nand2_1 U32825 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[8]), .Y(n27967) );
  sky130_fd_sc_hd__o21ai_1 U32826 ( .A1(n27968), .A2(n28545), .B1(n27967), .Y(
        n55) );
  sky130_fd_sc_hd__o22ai_1 U32827 ( .A1(n29146), .A2(n28316), .B1(n27969), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U32828 ( .A1(n29146), .A2(n28553), .B1(n27970), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U32829 ( .A1(n28235), .A2(n27971), .B1(n28959), 
        .B2(n28233), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__a22oi_1 U32830 ( .A1(n28318), .A2(
        j202_soc_core_intc_core_00_rg_ie[8]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[8]), .Y(n27973) );
  sky130_fd_sc_hd__a22oi_1 U32831 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[18]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[2]), .Y(n27972) );
  sky130_fd_sc_hd__nand3_1 U32832 ( .A(n27973), .B(n28238), .C(n27972), .Y(
        n27974) );
  sky130_fd_sc_hd__a21oi_1 U32833 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[104]), .B1(n27974), .Y(n27978) );
  sky130_fd_sc_hd__a22oi_1 U32834 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[26]), .B1(
        j202_soc_core_intc_core_00_rg_itgt[10]), .B2(n28331), .Y(n27977) );
  sky130_fd_sc_hd__a22oi_1 U32835 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[8]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[40]), .B2(n28330), .Y(n27976) );
  sky130_fd_sc_hd__nand2_1 U32836 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[72]), .Y(n27975) );
  sky130_fd_sc_hd__nand4_1 U32837 ( .A(n27978), .B(n27977), .C(n27976), .D(
        n27975), .Y(j202_soc_core_ahb2apb_01_N136) );
  sky130_fd_sc_hd__nand2_1 U32838 ( .A(n27980), .B(n27979), .Y(n28135) );
  sky130_fd_sc_hd__nand4_1 U32839 ( .A(n30202), .B(n27983), .C(n28135), .D(
        n27982), .Y(n27985) );
  sky130_fd_sc_hd__nand2_1 U32840 ( .A(n27985), .B(n28417), .Y(n27987) );
  sky130_fd_sc_hd__nand2_1 U32841 ( .A(n27987), .B(n27986), .Y(n10637) );
  sky130_fd_sc_hd__o22ai_1 U32842 ( .A1(n11180), .A2(n25977), .B1(n28061), 
        .B2(n27988), .Y(j202_soc_core_j22_cpu_rf_N2871) );
  sky130_fd_sc_hd__nand2_1 U32843 ( .A(n28079), .B(n29593), .Y(n27989) );
  sky130_fd_sc_hd__nand2_1 U32844 ( .A(n27994), .B(j202_soc_core_uart_div0[6]), 
        .Y(n27992) );
  sky130_fd_sc_hd__o21ai_1 U32845 ( .A1(n27994), .A2(n27993), .B1(n27992), .Y(
        n69) );
  sky130_fd_sc_hd__o22ai_1 U32846 ( .A1(n28002), .A2(n28310), .B1(n27995), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U32847 ( .A1(n28002), .A2(n28313), .B1(n27996), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U32848 ( .A1(n28002), .A2(n28316), .B1(n27997), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U32849 ( .A1(n28002), .A2(n28064), .B1(n27998), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U32850 ( .A1(n28002), .A2(n28553), .B1(n27999), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U32851 ( .A1(n28002), .A2(n29082), .B1(n28000), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U32852 ( .A1(n28002), .A2(n29076), .B1(n28001), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__a21oi_1 U32853 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[95]), .B1(n28326), .Y(n28010) );
  sky130_fd_sc_hd__nand2_1 U32854 ( .A(n28236), .B(
        j202_soc_core_intc_core_00_rg_ie[30]), .Y(n28005) );
  sky130_fd_sc_hd__a22oi_1 U32855 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[87]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[71]), .Y(n28004) );
  sky130_fd_sc_hd__nand2_1 U32856 ( .A(n28331), .B(
        j202_soc_core_intc_core_00_rg_itgt[79]), .Y(n28003) );
  sky130_fd_sc_hd__nand3_1 U32857 ( .A(n28005), .B(n28004), .C(n28003), .Y(
        n28006) );
  sky130_fd_sc_hd__a21oi_1 U32858 ( .A1(j202_soc_core_intc_core_00_rg_ipr[62]), 
        .A2(n28330), .B1(n28006), .Y(n28009) );
  sky130_fd_sc_hd__a22oi_1 U32859 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[30]), .B1(n28329), .B2(
        j202_soc_core_intc_core_00_rg_ipr[126]), .Y(n28008) );
  sky130_fd_sc_hd__nand2_1 U32860 ( .A(n28321), .B(
        j202_soc_core_intc_core_00_rg_ipr[94]), .Y(n28007) );
  sky130_fd_sc_hd__nand4_1 U32861 ( .A(n28010), .B(n28009), .C(n28008), .D(
        n28007), .Y(j202_soc_core_ahb2apb_01_N158) );
  sky130_fd_sc_hd__nand2_1 U32862 ( .A(n28731), .B(n29830), .Y(
        j202_soc_core_wbqspiflash_00_N720) );
  sky130_fd_sc_hd__xor2_1 U32863 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[4]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]), .X(n28014) );
  sky130_fd_sc_hd__xor2_1 U32864 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[5]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]), .X(n28013) );
  sky130_fd_sc_hd__xor2_1 U32865 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[1]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]), .X(n28012) );
  sky130_fd_sc_hd__xor2_1 U32866 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[2]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .X(n28011) );
  sky130_fd_sc_hd__nor4_1 U32867 ( .A(n28014), .B(n28013), .C(n28012), .D(
        n28011), .Y(n28020) );
  sky130_fd_sc_hd__xor2_1 U32868 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[3]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .X(n28016) );
  sky130_fd_sc_hd__xor2_1 U32869 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[0]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]), .X(n28015) );
  sky130_fd_sc_hd__nor3_1 U32870 ( .A(n28016), .B(n28015), .C(n28731), .Y(
        n28019) );
  sky130_fd_sc_hd__xnor2_1 U32871 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[6]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .Y(n28018) );
  sky130_fd_sc_hd__xnor2_1 U32872 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[7]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]), .Y(n28017) );
  sky130_fd_sc_hd__nand4_1 U32873 ( .A(n28020), .B(n28019), .C(n28018), .D(
        n28017), .Y(n28021) );
  sky130_fd_sc_hd__nand2_1 U32874 ( .A(n28022), .B(n28021), .Y(
        j202_soc_core_wbqspiflash_00_N719) );
  sky130_fd_sc_hd__nor2_1 U32875 ( .A(n28895), .B(n28024), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N352) );
  sky130_fd_sc_hd__a22o_1 U32876 ( .A1(n28026), .A2(
        j202_soc_core_wbqspiflash_00_spi_out[30]), .B1(n28025), .B2(
        j202_soc_core_wbqspiflash_00_dirty_sector), .X(
        j202_soc_core_wbqspiflash_00_N697) );
  sky130_fd_sc_hd__nand2_1 U32877 ( .A(n11175), .B(n28027), .Y(n28028) );
  sky130_fd_sc_hd__nand3_1 U32878 ( .A(n28030), .B(n28417), .C(n11384), .Y(
        n28034) );
  sky130_fd_sc_hd__nand2b_1 U32879 ( .A_N(n28155), .B(n28085), .Y(n28390) );
  sky130_fd_sc_hd__nand2b_1 U32880 ( .A_N(n28031), .B(n28390), .Y(n28032) );
  sky130_fd_sc_hd__nand2_1 U32881 ( .A(n28037), .B(n28036), .Y(n28134) );
  sky130_fd_sc_hd__nand2_1 U32882 ( .A(n28134), .B(n11389), .Y(n28039) );
  sky130_fd_sc_hd__nand2_1 U32883 ( .A(n28416), .B(n28039), .Y(n28040) );
  sky130_fd_sc_hd__nand2_1 U32884 ( .A(n28040), .B(n28417), .Y(n28041) );
  sky130_fd_sc_hd__o21a_1 U32885 ( .A1(n28379), .A2(n28344), .B1(n28390), .X(
        n28420) );
  sky130_fd_sc_hd__nand2_1 U32886 ( .A(n28041), .B(n28420), .Y(n10626) );
  sky130_fd_sc_hd__o22ai_1 U32888 ( .A1(n28044), .A2(n28043), .B1(n28042), 
        .B2(n28052), .Y(j202_soc_core_j22_cpu_ml_N155) );
  sky130_fd_sc_hd__a22oi_1 U32889 ( .A1(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]), .A2(n28045), .B1(n28050), 
        .B2(j202_soc_core_j22_cpu_ml_M_macop_MAC_[2]), .Y(n28046) );
  sky130_fd_sc_hd__o21ai_1 U32890 ( .A1(n28424), .A2(n28052), .B1(n28046), .Y(
        j202_soc_core_j22_cpu_ml_N154) );
  sky130_fd_sc_hd__a21oi_1 U32892 ( .A1(n28050), .A2(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .B1(n28049), .Y(n28051) );
  sky130_fd_sc_hd__o21ai_1 U32893 ( .A1(n28053), .A2(n28052), .B1(n28051), .Y(
        j202_soc_core_j22_cpu_ml_N153) );
  sky130_fd_sc_hd__nand2_1 U32894 ( .A(n28055), .B(n28054), .Y(n28058) );
  sky130_fd_sc_hd__nand2_1 U32895 ( .A(n28056), .B(
        j202_soc_core_j22_cpu_ml_bufa[4]), .Y(n28057) );
  sky130_fd_sc_hd__nand3_1 U32896 ( .A(n28058), .B(n12203), .C(n28057), .Y(
        j202_soc_core_j22_cpu_ml_machj[4]) );
  sky130_fd_sc_hd__o22ai_1 U32897 ( .A1(n28059), .A2(n25977), .B1(n28061), 
        .B2(n12344), .Y(j202_soc_core_j22_cpu_rf_N2867) );
  sky130_fd_sc_hd__o22ai_1 U32898 ( .A1(n25977), .A2(n28537), .B1(n28061), 
        .B2(n12256), .Y(j202_soc_core_j22_cpu_rf_N2881) );
  sky130_fd_sc_hd__o22ai_1 U32899 ( .A1(n29155), .A2(n28064), .B1(n28068), 
        .B2(n28063), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__nand2_1 U32900 ( .A(n28066), .B(n28065), .Y(n28067) );
  sky130_fd_sc_hd__nand4b_1 U32901 ( .A_N(
        j202_soc_core_intc_core_00_rg_irqc[11]), .B(n28067), .C(
        j202_soc_core_intc_core_00_in_intreq[11]), .D(n12069), .Y(n28070) );
  sky130_fd_sc_hd__nand2b_1 U32902 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[11]), 
        .B(n29590), .Y(n28069) );
  sky130_fd_sc_hd__a21oi_1 U32903 ( .A1(n28070), .A2(n28069), .B1(n28068), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N14) );
  sky130_fd_sc_hd__o21ai_1 U32904 ( .A1(j202_soc_core_j22_cpu_opst[2]), .A2(
        n28072), .B1(n28071), .Y(n28354) );
  sky130_fd_sc_hd__nand2_1 U32905 ( .A(n28360), .B(n28354), .Y(n28073) );
  sky130_fd_sc_hd__nand2_1 U32906 ( .A(n28074), .B(n28073), .Y(n28075) );
  sky130_fd_sc_hd__a21oi_1 U32907 ( .A1(n28076), .A2(n28417), .B1(n28075), .Y(
        n28077) );
  sky130_fd_sc_hd__nand2_1 U32908 ( .A(n28078), .B(n28077), .Y(n10541) );
  sky130_fd_sc_hd__nand2_1 U32909 ( .A(n28079), .B(n23549), .Y(n28080) );
  sky130_fd_sc_hd__nand2_1 U32910 ( .A(n28081), .B(n28080), .Y(n10529) );
  sky130_fd_sc_hd__inv_1 U32911 ( .A(n29591), .Y(n10591) );
  sky130_fd_sc_hd__nand2_1 U32912 ( .A(n28083), .B(n28082), .Y(n28088) );
  sky130_fd_sc_hd__nand3_1 U32913 ( .A(n28087), .B(n28086), .C(n28085), .Y(
        n28370) );
  sky130_fd_sc_hd__o21a_1 U32914 ( .A1(n28417), .A2(n28088), .B1(n28370), .X(
        n28101) );
  sky130_fd_sc_hd__nand2_1 U32915 ( .A(n28093), .B(n30061), .Y(n28094) );
  sky130_fd_sc_hd__nand2_1 U32916 ( .A(n28099), .B(n13048), .Y(n28100) );
  sky130_fd_sc_hd__nand2_1 U32917 ( .A(n28101), .B(n28100), .Y(n28110) );
  sky130_fd_sc_hd__a21oi_1 U32918 ( .A1(n28105), .A2(n28104), .B1(n28103), .Y(
        n28108) );
  sky130_fd_sc_hd__nand3_1 U32919 ( .A(n28109), .B(n28108), .C(n28107), .Y(
        n28364) );
  sky130_fd_sc_hd__nand2_1 U32920 ( .A(n28110), .B(n28364), .Y(n10608) );
  sky130_fd_sc_hd__o22ai_1 U32921 ( .A1(n28113), .A2(n25979), .B1(n28112), 
        .B2(n28111), .Y(j202_soc_core_j22_cpu_rf_N3208) );
  sky130_fd_sc_hd__inv_1 U32922 ( .A(n29592), .Y(n10583) );
  sky130_fd_sc_hd__nand3_1 U32924 ( .A(n28118), .B(n28367), .C(n28117), .Y(
        n28119) );
  sky130_fd_sc_hd__nor2_1 U32925 ( .A(n28120), .B(n28119), .Y(n28122) );
  sky130_fd_sc_hd__nand2_1 U32926 ( .A(n28126), .B(n28125), .Y(n28128) );
  sky130_fd_sc_hd__nand2_1 U32927 ( .A(n28128), .B(n28127), .Y(n10620) );
  sky130_fd_sc_hd__nand2_1 U32928 ( .A(n12669), .B(n29593), .Y(n28408) );
  sky130_fd_sc_hd__nor2_1 U32929 ( .A(n29595), .B(n28129), .Y(n28131) );
  sky130_fd_sc_hd__o2bb2ai_1 U32930 ( .B1(n12395), .B2(n28408), .A1_N(n28131), 
        .A2_N(n11423), .Y(n28132) );
  sky130_fd_sc_hd__a21oi_1 U32931 ( .A1(n11175), .A2(n28133), .B1(n28132), .Y(
        n28137) );
  sky130_fd_sc_hd__nand4_1 U32932 ( .A(n28138), .B(n28137), .C(n28136), .D(
        n28135), .Y(n28139) );
  sky130_fd_sc_hd__nor2_1 U32933 ( .A(n28139), .B(n28140), .Y(n28141) );
  sky130_fd_sc_hd__nand2_1 U32934 ( .A(n28141), .B(n28142), .Y(n28143) );
  sky130_fd_sc_hd__nand2_1 U32935 ( .A(n28143), .B(n28417), .Y(n28146) );
  sky130_fd_sc_hd__nand3_1 U32936 ( .A(n28146), .B(n28145), .C(n28144), .Y(
        n10633) );
  sky130_fd_sc_hd__inv_1 U32937 ( .A(n29596), .Y(n10586) );
  sky130_fd_sc_hd__nand2_1 U32939 ( .A(n28153), .B(n28417), .Y(n28156) );
  sky130_fd_sc_hd__nand3_1 U32940 ( .A(n28156), .B(n28155), .C(n28154), .Y(
        n10630) );
  sky130_fd_sc_hd__a21oi_1 U32941 ( .A1(n28160), .A2(n28159), .B1(n28158), .Y(
        n138) );
  sky130_fd_sc_hd__nand3_1 U32942 ( .A(n28165), .B(n28164), .C(n28163), .Y(
        n28281) );
  sky130_fd_sc_hd__nand2_1 U32943 ( .A(n28281), .B(
        j202_soc_core_bldc_core_00_comm[2]), .Y(n28166) );
  sky130_fd_sc_hd__o21ai_1 U32944 ( .A1(n28178), .A2(n28281), .B1(n28166), .Y(
        n41) );
  sky130_fd_sc_hd__nand2_1 U32945 ( .A(n28287), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[2]), .Y(n28167) );
  sky130_fd_sc_hd__nand2_1 U32947 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[2]), .Y(n28168) );
  sky130_fd_sc_hd__o21ai_1 U32948 ( .A1(n28171), .A2(n28289), .B1(n28168), .Y(
        n85) );
  sky130_fd_sc_hd__nand2_1 U32949 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[2]), .Y(n28169) );
  sky130_fd_sc_hd__o21ai_1 U32950 ( .A1(n28171), .A2(n28291), .B1(n28169), .Y(
        n84) );
  sky130_fd_sc_hd__nand2_1 U32951 ( .A(n28293), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[2]), .Y(n28170) );
  sky130_fd_sc_hd__o21ai_1 U32952 ( .A1(n28171), .A2(n28293), .B1(n28170), .Y(
        n82) );
  sky130_fd_sc_hd__a22oi_1 U32953 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[2]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[2]), .Y(
        n28175) );
  sky130_fd_sc_hd__a22oi_1 U32954 ( .A1(n28297), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[2]), 
        .B1(n28299), .B2(j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[2]), .Y(
        n28174) );
  sky130_fd_sc_hd__nand2_1 U32955 ( .A(n28301), .B(
        j202_soc_core_cmt_core_00_const0[2]), .Y(n28173) );
  sky130_fd_sc_hd__nand2_1 U32956 ( .A(n28300), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[2]), .Y(n28172) );
  sky130_fd_sc_hd__nand4_1 U32957 ( .A(n28175), .B(n28174), .C(n28173), .D(
        n28172), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[2]) );
  sky130_fd_sc_hd__nand2_1 U32958 ( .A(n28177), .B(
        j202_soc_core_bldc_core_00_pwm_period[2]), .Y(n28176) );
  sky130_fd_sc_hd__o21ai_1 U32959 ( .A1(n28178), .A2(n28177), .B1(n28176), .Y(
        n49) );
  sky130_fd_sc_hd__o22ai_1 U32960 ( .A1(n29162), .A2(n28310), .B1(n28179), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U32961 ( .A1(n29162), .A2(n28313), .B1(n28180), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U32962 ( .A1(n29162), .A2(n28316), .B1(n28181), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U32963 ( .A1(n29162), .A2(n28553), .B1(n28182), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U32964 ( .A1(n29162), .A2(n29082), .B1(n28183), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U32965 ( .A1(n29162), .A2(n29079), .B1(n28184), 
        .B2(n29077), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U32966 ( .A1(n29162), .A2(n29076), .B1(n28185), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__a22o_1 U32967 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[88]), .B1(n28331), .B2(
        j202_soc_core_intc_core_00_rg_itgt[72]), .X(n28189) );
  sky130_fd_sc_hd__a22oi_1 U32968 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[2]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[2]), .Y(n28187) );
  sky130_fd_sc_hd__a22oi_1 U32969 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[80]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[64]), .Y(n28186) );
  sky130_fd_sc_hd__nand3_1 U32970 ( .A(n28187), .B(n28238), .C(n28186), .Y(
        n28188) );
  sky130_fd_sc_hd__a211oi_1 U32971 ( .A1(n28321), .A2(
        j202_soc_core_intc_core_00_rg_ipr[66]), .B1(n28189), .C1(n28188), .Y(
        n28192) );
  sky130_fd_sc_hd__a22oi_1 U32972 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[2]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[34]), .B2(n28330), .Y(n28191) );
  sky130_fd_sc_hd__a22oi_1 U32973 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[98]), .B1(n28319), .B2(
        j202_soc_core_intc_core_00_rg_eimk[2]), .Y(n28190) );
  sky130_fd_sc_hd__nand3_1 U32974 ( .A(n28192), .B(n28191), .C(n28190), .Y(
        j202_soc_core_ahb2apb_01_N130) );
  sky130_fd_sc_hd__nor2_1 U32975 ( .A(n28898), .B(n28193), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N360) );
  sky130_fd_sc_hd__nor2_1 U32976 ( .A(n29086), .B(n28336), .Y(
        j202_soc_core_wbqspiflash_00_N669) );
  sky130_fd_sc_hd__a22oi_1 U32977 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[2]), .A2(n29394), 
        .B1(n29389), .B2(la_data_out[2]), .Y(n28196) );
  sky130_fd_sc_hd__a22o_1 U32978 ( .A1(gpio_en_o[2]), .A2(n29393), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[2]), .B2(n29390), .X(
        n28194) );
  sky130_fd_sc_hd__a21oi_1 U32979 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[2]), .A2(n29391), .B1(
        n28194), .Y(n28195) );
  sky130_fd_sc_hd__o211ai_1 U32980 ( .A1(n29311), .A2(n28916), .B1(n28196), 
        .C1(n28195), .Y(j202_soc_core_ahb2apb_02_N130) );
  sky130_fd_sc_hd__a22oi_1 U32981 ( .A1(n28198), .A2(n28355), .B1(n28197), 
        .B2(n28417), .Y(n28199) );
  sky130_fd_sc_hd__nand2_1 U32982 ( .A(n28200), .B(n28199), .Y(n10631) );
  sky130_fd_sc_hd__nand4_1 U32983 ( .A(n28204), .B(n28203), .C(n28202), .D(
        n28201), .Y(n28277) );
  sky130_fd_sc_hd__nand2_1 U32984 ( .A(n28277), .B(
        j202_soc_core_bldc_core_00_pwm_en), .Y(n28205) );
  sky130_fd_sc_hd__nand2_1 U32986 ( .A(n29599), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[0]), .Y(n28206) );
  sky130_fd_sc_hd__nand2_1 U32988 ( .A(n28281), .B(
        j202_soc_core_bldc_core_00_comm[0]), .Y(n28208) );
  sky130_fd_sc_hd__o21ai_1 U32989 ( .A1(n28209), .A2(n28281), .B1(n28208), .Y(
        n42) );
  sky130_fd_sc_hd__nor2_1 U32990 ( .A(n28211), .B(n28210), .Y(n28284) );
  sky130_fd_sc_hd__nand2_1 U32991 ( .A(n28284), .B(
        j202_soc_core_cmt_core_00_wdata_cnt0[0]), .Y(n28212) );
  sky130_fd_sc_hd__nand2_1 U32993 ( .A(n28287), .B(
        j202_soc_core_cmt_core_00_cks1[0]), .Y(n28214) );
  sky130_fd_sc_hd__nand2_1 U32995 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[0]), .Y(n28215) );
  sky130_fd_sc_hd__o21ai_1 U32996 ( .A1(n28218), .A2(n28289), .B1(n28215), .Y(
        n91) );
  sky130_fd_sc_hd__nand2_1 U32997 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[0]), .Y(n28216) );
  sky130_fd_sc_hd__o21ai_1 U32998 ( .A1(n28218), .A2(n28291), .B1(n28216), .Y(
        n90) );
  sky130_fd_sc_hd__nand2_1 U32999 ( .A(n28293), .B(
        j202_soc_core_cmt_core_00_cks0[0]), .Y(n28217) );
  sky130_fd_sc_hd__o21ai_1 U33000 ( .A1(n28218), .A2(n28293), .B1(n28217), .Y(
        n88) );
  sky130_fd_sc_hd__a22oi_1 U33001 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[0]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[0]), .Y(
        n28226) );
  sky130_fd_sc_hd__and3_1 U33002 ( .A(n28222), .B(n28221), .C(n28220), .X(
        n28298) );
  sky130_fd_sc_hd__a22oi_1 U33003 ( .A1(n28298), .A2(
        j202_soc_core_cmt_core_00_str0), .B1(n28297), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[0]), .Y(
        n28225) );
  sky130_fd_sc_hd__a22oi_1 U33004 ( .A1(n28300), .A2(
        j202_soc_core_cmt_core_00_cks1[0]), .B1(n28299), .B2(
        j202_soc_core_cmt_core_00_cks0[0]), .Y(n28224) );
  sky130_fd_sc_hd__nand2_1 U33005 ( .A(n28301), .B(
        j202_soc_core_cmt_core_00_const0[0]), .Y(n28223) );
  sky130_fd_sc_hd__nand4_1 U33006 ( .A(n28226), .B(n28225), .C(n28224), .D(
        n28223), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[0]) );
  sky130_fd_sc_hd__nand2_1 U33007 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[0]), .Y(n28227) );
  sky130_fd_sc_hd__o21ai_1 U33008 ( .A1(n28228), .A2(n28545), .B1(n28227), .Y(
        n47) );
  sky130_fd_sc_hd__o22ai_1 U33009 ( .A1(n29165), .A2(n28316), .B1(n28229), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U33010 ( .A1(n28231), .A2(n29399), .B1(n28230), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U33011 ( .A1(n29165), .A2(n29079), .B1(n28232), 
        .B2(n29077), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U33012 ( .A1(n28235), .A2(n28234), .B1(n28246), 
        .B2(n28233), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__a22o_1 U33013 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[24]), .B1(
        j202_soc_core_intc_core_00_rg_itgt[8]), .B2(n28331), .X(n28241) );
  sky130_fd_sc_hd__a22oi_1 U33014 ( .A1(n28236), .A2(
        j202_soc_core_intc_core_00_rg_ie[0]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[0]), .Y(n28239) );
  sky130_fd_sc_hd__a22oi_1 U33015 ( .A1(n28322), .A2(
        j202_soc_core_intc_core_00_rg_itgt[16]), .B1(n28328), .B2(
        j202_soc_core_intc_core_00_rg_itgt[0]), .Y(n28237) );
  sky130_fd_sc_hd__nand3_1 U33016 ( .A(n28239), .B(n28238), .C(n28237), .Y(
        n28240) );
  sky130_fd_sc_hd__a211oi_1 U33017 ( .A1(n28321), .A2(
        j202_soc_core_intc_core_00_rg_ipr[64]), .B1(n28241), .C1(n28240), .Y(
        n28244) );
  sky130_fd_sc_hd__a22oi_1 U33018 ( .A1(n28323), .A2(
        j202_soc_core_intc_core_00_rg_ipr[0]), .B1(
        j202_soc_core_intc_core_00_rg_ipr[32]), .B2(n28330), .Y(n28243) );
  sky130_fd_sc_hd__a22oi_1 U33019 ( .A1(n28329), .A2(
        j202_soc_core_intc_core_00_rg_ipr[96]), .B1(n28319), .B2(
        j202_soc_core_intc_core_00_rg_eimk[0]), .Y(n28242) );
  sky130_fd_sc_hd__nand3_1 U33020 ( .A(n28244), .B(n28243), .C(n28242), .Y(
        j202_soc_core_ahb2apb_01_N128) );
  sky130_fd_sc_hd__nor2_1 U33021 ( .A(n28780), .B(n28336), .Y(
        j202_soc_core_wbqspiflash_00_N667) );
  sky130_fd_sc_hd__a21oi_1 U33022 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[0]), .A2(n29830), .B1(
        n29598), .Y(n28249) );
  sky130_fd_sc_hd__o21ai_1 U33023 ( .A1(n28250), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[0]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[0]), .Y(n28245) );
  sky130_fd_sc_hd__a21o_1 U33024 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[0]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[0]), .B1(n28245), 
        .X(n28248) );
  sky130_fd_sc_hd__o31ai_1 U33026 ( .A1(gpio_en_o[0]), .A2(n28249), .A3(n28248), .B1(n28247), .Y(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N40) );
  sky130_fd_sc_hd__o22ai_1 U33027 ( .A1(n28250), .A2(n29311), .B1(io_oeb[0]), 
        .B2(n29310), .Y(n28251) );
  sky130_fd_sc_hd__a21oi_1 U33028 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[0]), .A2(n29390), .B1(
        n28251), .Y(n28252) );
  sky130_fd_sc_hd__o21ai_1 U33029 ( .A1(n28254), .A2(n28253), .B1(n28252), .Y(
        n28255) );
  sky130_fd_sc_hd__a21oi_1 U33030 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[0]), .A2(n29391), .B1(
        n28255), .Y(n28256) );
  sky130_fd_sc_hd__nand2_1 U33032 ( .A(n28260), .B(n28259), .Y(n28265) );
  sky130_fd_sc_hd__nand2_1 U33033 ( .A(n28262), .B(n28261), .Y(n28263) );
  sky130_fd_sc_hd__nor3_1 U33034 ( .A(n28265), .B(n28264), .C(n28263), .Y(
        n28269) );
  sky130_fd_sc_hd__nand2_1 U33035 ( .A(n28271), .B(n28417), .Y(n28273) );
  sky130_fd_sc_hd__nand2_1 U33036 ( .A(n28273), .B(n28272), .Y(n10635) );
  sky130_fd_sc_hd__o21ai_1 U33037 ( .A1(n28275), .A2(n28274), .B1(n12069), .Y(
        n10578) );
  sky130_fd_sc_hd__nand2_1 U33038 ( .A(n28277), .B(
        j202_soc_core_bldc_core_00_adc_en), .Y(n28276) );
  sky130_fd_sc_hd__o21ai_1 U33039 ( .A1(n28282), .A2(n28277), .B1(n28276), .Y(
        n44) );
  sky130_fd_sc_hd__nand2_1 U33040 ( .A(n29599), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[1]), .Y(n28278) );
  sky130_fd_sc_hd__o21ai_1 U33041 ( .A1(n29599), .A2(n28279), .B1(n28278), .Y(
        n136) );
  sky130_fd_sc_hd__nand2_1 U33042 ( .A(n28281), .B(
        j202_soc_core_bldc_core_00_comm[1]), .Y(n28280) );
  sky130_fd_sc_hd__o21ai_1 U33043 ( .A1(n28282), .A2(n28281), .B1(n28280), .Y(
        n43) );
  sky130_fd_sc_hd__nand2_1 U33044 ( .A(n28284), .B(
        j202_soc_core_cmt_core_00_wdata_cnt0[1]), .Y(n28283) );
  sky130_fd_sc_hd__nand2_1 U33046 ( .A(n28287), .B(
        j202_soc_core_cmt_core_00_cks1[1]), .Y(n28286) );
  sky130_fd_sc_hd__o21ai_1 U33047 ( .A1(n28294), .A2(n28287), .B1(n28286), .Y(
        n117) );
  sky130_fd_sc_hd__nand2_1 U33048 ( .A(n28289), .B(
        j202_soc_core_cmt_core_00_const1[1]), .Y(n28288) );
  sky130_fd_sc_hd__o21ai_1 U33049 ( .A1(n28294), .A2(n28289), .B1(n28288), .Y(
        n119) );
  sky130_fd_sc_hd__nand2_1 U33050 ( .A(n28291), .B(
        j202_soc_core_cmt_core_00_const0[1]), .Y(n28290) );
  sky130_fd_sc_hd__o21ai_1 U33051 ( .A1(n28294), .A2(n28291), .B1(n28290), .Y(
        n118) );
  sky130_fd_sc_hd__nand2_1 U33052 ( .A(n28293), .B(
        j202_soc_core_cmt_core_00_cks0[1]), .Y(n28292) );
  sky130_fd_sc_hd__o21ai_1 U33053 ( .A1(n28294), .A2(n28293), .B1(n28292), .Y(
        n116) );
  sky130_fd_sc_hd__a22oi_1 U33054 ( .A1(n28296), .A2(
        j202_soc_core_cmt_core_00_const1[1]), .B1(n28295), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[1]), .Y(
        n28305) );
  sky130_fd_sc_hd__a22oi_1 U33055 ( .A1(n28298), .A2(
        j202_soc_core_cmt_core_00_str1), .B1(n28297), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[1]), .Y(
        n28304) );
  sky130_fd_sc_hd__a22oi_1 U33056 ( .A1(n28300), .A2(
        j202_soc_core_cmt_core_00_cks1[1]), .B1(n28299), .B2(
        j202_soc_core_cmt_core_00_cks0[1]), .Y(n28303) );
  sky130_fd_sc_hd__nand2_1 U33057 ( .A(n28301), .B(
        j202_soc_core_cmt_core_00_const0[1]), .Y(n28302) );
  sky130_fd_sc_hd__nand4_1 U33058 ( .A(n28305), .B(n28304), .C(n28303), .D(
        n28302), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[1]) );
  sky130_fd_sc_hd__nand2_1 U33059 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[1]), .Y(n28306) );
  sky130_fd_sc_hd__o21ai_1 U33060 ( .A1(n28307), .A2(n28545), .B1(n28306), .Y(
        n48) );
  sky130_fd_sc_hd__o22ai_1 U33061 ( .A1(n29163), .A2(n28310), .B1(n28309), 
        .B2(n28308), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U33062 ( .A1(n29163), .A2(n28313), .B1(n28312), 
        .B2(n28311), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U33063 ( .A1(n29163), .A2(n28316), .B1(n28315), 
        .B2(n28314), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__a22oi_1 U33064 ( .A1(n28318), .A2(
        j202_soc_core_intc_core_00_rg_ie[1]), .B1(n28317), .B2(
        j202_soc_core_intc_core_00_in_intreq[1]), .Y(n28335) );
  sky130_fd_sc_hd__a22oi_1 U33065 ( .A1(n28320), .A2(
        j202_soc_core_intc_core_00_rg_itgt[56]), .B1(n28319), .B2(
        j202_soc_core_intc_core_00_rg_eimk[1]), .Y(n28325) );
  sky130_fd_sc_hd__a222oi_1 U33066 ( .A1(j202_soc_core_intc_core_00_rg_ipr[1]), 
        .A2(n28323), .B1(n28322), .B2(j202_soc_core_intc_core_00_rg_itgt[48]), 
        .C1(n28321), .C2(j202_soc_core_intc_core_00_rg_ipr[65]), .Y(n28324) );
  sky130_fd_sc_hd__nand2_1 U33067 ( .A(n28325), .B(n28324), .Y(n28327) );
  sky130_fd_sc_hd__a211oi_1 U33068 ( .A1(n28328), .A2(
        j202_soc_core_intc_core_00_rg_itgt[32]), .B1(n28327), .C1(n28326), .Y(
        n28334) );
  sky130_fd_sc_hd__a22oi_1 U33069 ( .A1(n28330), .A2(
        j202_soc_core_intc_core_00_rg_ipr[33]), .B1(n28329), .B2(
        j202_soc_core_intc_core_00_rg_ipr[97]), .Y(n28333) );
  sky130_fd_sc_hd__nand2_1 U33070 ( .A(n28331), .B(
        j202_soc_core_intc_core_00_rg_itgt[40]), .Y(n28332) );
  sky130_fd_sc_hd__nand4_1 U33071 ( .A(n28335), .B(n28334), .C(n28333), .D(
        n28332), .Y(j202_soc_core_ahb2apb_01_N129) );
  sky130_fd_sc_hd__nor2_1 U33072 ( .A(n29084), .B(n28336), .Y(
        j202_soc_core_wbqspiflash_00_N668) );
  sky130_fd_sc_hd__a22oi_1 U33073 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[1]), .A2(n29391), .B1(
        n29389), .B2(la_data_out[1]), .Y(n28339) );
  sky130_fd_sc_hd__a22o_1 U33074 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[1]), .A2(n29392), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[1]), .B2(n29390), .X(
        n28337) );
  sky130_fd_sc_hd__a21oi_1 U33075 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]), .A2(n29394), 
        .B1(n28337), .Y(n28338) );
  sky130_fd_sc_hd__o211ai_1 U33076 ( .A1(n29310), .A2(io_oeb[1]), .B1(n28339), 
        .C1(n28338), .Y(j202_soc_core_ahb2apb_02_N129) );
  sky130_fd_sc_hd__nor2_1 U33077 ( .A(n28341), .B(n28405), .Y(n28343) );
  sky130_fd_sc_hd__nor2_1 U33078 ( .A(n28343), .B(n28342), .Y(n28382) );
  sky130_fd_sc_hd__nand2_1 U33079 ( .A(n28345), .B(n28344), .Y(n28400) );
  sky130_fd_sc_hd__nand2_1 U33080 ( .A(n28400), .B(n28417), .Y(n28351) );
  sky130_fd_sc_hd__nand3_1 U33081 ( .A(n28394), .B(n28346), .C(n28370), .Y(
        n28347) );
  sky130_fd_sc_hd__a21oi_1 U33082 ( .A1(n28348), .A2(n28417), .B1(n28347), .Y(
        n28350) );
  sky130_fd_sc_hd__nand4_1 U33083 ( .A(n28382), .B(n28351), .C(n28350), .D(
        n28349), .Y(n10607) );
  sky130_fd_sc_hd__a31oi_1 U33084 ( .A1(n28360), .A2(n28355), .A3(n28354), 
        .B1(n28353), .Y(n28356) );
  sky130_fd_sc_hd__nand2_1 U33085 ( .A(n28358), .B(n28417), .Y(n28362) );
  sky130_fd_sc_hd__nand2_1 U33086 ( .A(n28360), .B(n28359), .Y(n28374) );
  sky130_fd_sc_hd__nand3_1 U33087 ( .A(n28362), .B(n28361), .C(n28374), .Y(
        n28363) );
  sky130_fd_sc_hd__nand2_1 U33088 ( .A(n28370), .B(n28364), .Y(n28406) );
  sky130_fd_sc_hd__nand2_1 U33089 ( .A(n28363), .B(n28396), .Y(n28371) );
  sky130_fd_sc_hd__nand2_1 U33090 ( .A(n28364), .B(n29088), .Y(n28369) );
  sky130_fd_sc_hd__or3_1 U33091 ( .A(j202_soc_core_intr_vec__0_), .B(
        j202_soc_core_intr_vec__3_), .C(j202_soc_core_intr_vec__4_), .X(n28365) );
  sky130_fd_sc_hd__or3_1 U33092 ( .A(j202_soc_core_intr_vec__2_), .B(
        j202_soc_core_intr_vec__6_), .C(n28365), .X(n28372) );
  sky130_fd_sc_hd__nor2_1 U33093 ( .A(n28366), .B(n28372), .Y(n28368) );
  sky130_fd_sc_hd__o21ai_1 U33094 ( .A1(n28368), .A2(n28370), .B1(n28367), .Y(
        n28395) );
  sky130_fd_sc_hd__a21o_1 U33095 ( .A1(n28370), .A2(n28369), .B1(n28395), .X(
        n28404) );
  sky130_fd_sc_hd__nand2_1 U33096 ( .A(n28371), .B(n28404), .Y(n10604) );
  sky130_fd_sc_hd__nor3_1 U33097 ( .A(j202_soc_core_intr_vec__1_), .B(n28373), 
        .C(n28372), .Y(n28375) );
  sky130_fd_sc_hd__nor2_1 U33098 ( .A(n28375), .B(n28374), .Y(
        j202_soc_core_j22_cpu_id_idec_N822) );
  sky130_fd_sc_hd__a211oi_1 U33099 ( .A1(n28377), .A2(n28376), .B1(
        j202_soc_core_intc_core_00_cp_intack_all_0_), .C1(n29073), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_req_N3) );
  sky130_fd_sc_hd__inv_1 U33100 ( .A(n29600), .Y(n10590) );
  sky130_fd_sc_hd__nor2_1 U33101 ( .A(n28379), .B(n28406), .Y(n28410) );
  sky130_fd_sc_hd__nand3_1 U33102 ( .A(n28411), .B(n28410), .C(n28380), .Y(
        n28381) );
  sky130_fd_sc_hd__o211ai_1 U33103 ( .A1(n28406), .A2(n28382), .B1(n28404), 
        .C1(n28381), .Y(j202_soc_core_j22_cpu_id_idec_N894) );
  sky130_fd_sc_hd__a31oi_1 U33104 ( .A1(n28385), .A2(n29830), .A3(n28384), 
        .B1(n28383), .Y(n10579) );
  sky130_fd_sc_hd__nand4b_1 U33105 ( .A_N(n28388), .B(n28387), .C(n28415), .D(
        n28386), .Y(n28389) );
  sky130_fd_sc_hd__nand2_1 U33106 ( .A(n28389), .B(n28417), .Y(n28391) );
  sky130_fd_sc_hd__nand2_1 U33107 ( .A(n28391), .B(n28390), .Y(n10625) );
  sky130_fd_sc_hd__nand2_1 U33108 ( .A(n24594), .B(n11172), .Y(n28392) );
  sky130_fd_sc_hd__o21ai_1 U33109 ( .A1(n28393), .A2(n28392), .B1(n28410), .Y(
        n28399) );
  sky130_fd_sc_hd__a21oi_1 U33110 ( .A1(n28397), .A2(n28396), .B1(n28395), .Y(
        n28398) );
  sky130_fd_sc_hd__nand2_1 U33111 ( .A(n28399), .B(n28398), .Y(n10606) );
  sky130_fd_sc_hd__nand2_1 U33112 ( .A(n28400), .B(n28410), .Y(n28414) );
  sky130_fd_sc_hd__a21oi_1 U33113 ( .A1(n28403), .A2(n28402), .B1(n28401), .Y(
        n28407) );
  sky130_fd_sc_hd__o31a_1 U33114 ( .A1(n28407), .A2(n28406), .A3(n28405), .B1(
        n28404), .X(n28413) );
  sky130_fd_sc_hd__nand4_1 U33115 ( .A(n28411), .B(n28410), .C(n28409), .D(
        n28408), .Y(n28412) );
  sky130_fd_sc_hd__nand3_1 U33116 ( .A(n28414), .B(n28413), .C(n28412), .Y(
        n10605) );
  sky130_fd_sc_hd__o21ai_1 U33117 ( .A1(n28419), .A2(n28418), .B1(n28417), .Y(
        n28421) );
  sky130_fd_sc_hd__nand2_1 U33118 ( .A(n28421), .B(n28420), .Y(n10627) );
  sky130_fd_sc_hd__o21ai_1 U33119 ( .A1(n28424), .A2(n28423), .B1(n28422), .Y(
        j202_soc_core_j22_cpu_ml_N193) );
  sky130_fd_sc_hd__nand3_1 U33120 ( .A(n12260), .B(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[3]), .C(n28425), .Y(n28427) );
  sky130_fd_sc_hd__o211ai_1 U33121 ( .A1(n28429), .A2(n28428), .B1(n28427), 
        .C1(n24292), .Y(j202_soc_core_j22_cpu_ml_N336) );
  sky130_fd_sc_hd__a22oi_1 U33122 ( .A1(n28533), .A2(n28431), .B1(n12260), 
        .B2(n28524), .Y(n28433) );
  sky130_fd_sc_hd__nand2_1 U33123 ( .A(n28433), .B(n28535), .Y(
        j202_soc_core_j22_cpu_ml_N370) );
  sky130_fd_sc_hd__nor2_1 U33124 ( .A(n28435), .B(n28434), .Y(n28436) );
  sky130_fd_sc_hd__mux2i_1 U33125 ( .A0(n28437), .A1(n28436), .S(n13325), .Y(
        n28440) );
  sky130_fd_sc_hd__nand3_1 U33126 ( .A(n28443), .B(n28438), .C(n28540), .Y(
        n28439) );
  sky130_fd_sc_hd__nand2_1 U33127 ( .A(n28440), .B(n28439), .Y(
        j202_soc_core_j22_cpu_ml_N429) );
  sky130_fd_sc_hd__nand2_1 U33128 ( .A(n28441), .B(n28512), .Y(n28491) );
  sky130_fd_sc_hd__nand2_1 U33129 ( .A(n28442), .B(n28539), .Y(n28445) );
  sky130_fd_sc_hd__a22oi_1 U33130 ( .A1(j202_soc_core_j22_cpu_ml_bufb[31]), 
        .A2(n13325), .B1(n28443), .B2(n28540), .Y(n28444) );
  sky130_fd_sc_hd__nand2_1 U33131 ( .A(n28445), .B(n28444), .Y(
        j202_soc_core_j22_cpu_ml_N427) );
  sky130_fd_sc_hd__nand2_1 U33132 ( .A(n28446), .B(n28533), .Y(n28447) );
  sky130_fd_sc_hd__o211ai_1 U33133 ( .A1(n28538), .A2(n28448), .B1(n28447), 
        .C1(n28535), .Y(j202_soc_core_j22_cpu_ml_N369) );
  sky130_fd_sc_hd__a22oi_1 U33134 ( .A1(j202_soc_core_j22_cpu_ml_bufb[30]), 
        .A2(n13325), .B1(n28449), .B2(n28540), .Y(n28450) );
  sky130_fd_sc_hd__o21ai_1 U33135 ( .A1(n28491), .A2(n26896), .B1(n28450), .Y(
        j202_soc_core_j22_cpu_ml_N426) );
  sky130_fd_sc_hd__o22a_1 U33136 ( .A1(n28451), .A2(n28512), .B1(n28538), .B2(
        n27642), .X(n28452) );
  sky130_fd_sc_hd__nand2_1 U33137 ( .A(n28535), .B(n28452), .Y(
        j202_soc_core_j22_cpu_ml_N368) );
  sky130_fd_sc_hd__nand2_1 U33138 ( .A(n28453), .B(n28539), .Y(n28456) );
  sky130_fd_sc_hd__a22oi_1 U33139 ( .A1(j202_soc_core_j22_cpu_ml_bufb[29]), 
        .A2(n13325), .B1(n28454), .B2(n28540), .Y(n28455) );
  sky130_fd_sc_hd__nand2_1 U33140 ( .A(n28456), .B(n28455), .Y(
        j202_soc_core_j22_cpu_ml_N425) );
  sky130_fd_sc_hd__o22a_1 U33141 ( .A1(n28457), .A2(n28512), .B1(n28538), .B2(
        n27389), .X(n28458) );
  sky130_fd_sc_hd__nand2_1 U33142 ( .A(n28535), .B(n28458), .Y(
        j202_soc_core_j22_cpu_ml_N367) );
  sky130_fd_sc_hd__nand2_1 U33143 ( .A(n28459), .B(n28539), .Y(n28462) );
  sky130_fd_sc_hd__a22oi_1 U33144 ( .A1(j202_soc_core_j22_cpu_ml_bufb[28]), 
        .A2(n13325), .B1(n28460), .B2(n28540), .Y(n28461) );
  sky130_fd_sc_hd__nand2_1 U33145 ( .A(n28462), .B(n28461), .Y(
        j202_soc_core_j22_cpu_ml_N424) );
  sky130_fd_sc_hd__nand2_1 U33146 ( .A(n28463), .B(n28533), .Y(n28464) );
  sky130_fd_sc_hd__o211ai_1 U33147 ( .A1(n28538), .A2(n27019), .B1(n28535), 
        .C1(n28464), .Y(j202_soc_core_j22_cpu_ml_N366) );
  sky130_fd_sc_hd__nand2_1 U33148 ( .A(n28466), .B(n28539), .Y(n28469) );
  sky130_fd_sc_hd__a22oi_1 U33149 ( .A1(j202_soc_core_j22_cpu_ml_bufb[27]), 
        .A2(n13325), .B1(n28467), .B2(n28540), .Y(n28468) );
  sky130_fd_sc_hd__nand2_1 U33150 ( .A(n28469), .B(n28468), .Y(
        j202_soc_core_j22_cpu_ml_N423) );
  sky130_fd_sc_hd__a22oi_1 U33151 ( .A1(n28533), .A2(n28471), .B1(n28470), 
        .B2(n28524), .Y(n28472) );
  sky130_fd_sc_hd__nand2_1 U33152 ( .A(n28535), .B(n28472), .Y(
        j202_soc_core_j22_cpu_ml_N365) );
  sky130_fd_sc_hd__a22oi_1 U33153 ( .A1(j202_soc_core_j22_cpu_ml_bufb[26]), 
        .A2(n13325), .B1(n28473), .B2(n28540), .Y(n28474) );
  sky130_fd_sc_hd__o21ai_1 U33154 ( .A1(n28491), .A2(n26965), .B1(n28474), .Y(
        j202_soc_core_j22_cpu_ml_N422) );
  sky130_fd_sc_hd__nand2_1 U33155 ( .A(n28475), .B(n28533), .Y(n28476) );
  sky130_fd_sc_hd__o211ai_1 U33156 ( .A1(n28538), .A2(n28477), .B1(n28476), 
        .C1(n28535), .Y(j202_soc_core_j22_cpu_ml_N364) );
  sky130_fd_sc_hd__a22oi_1 U33157 ( .A1(j202_soc_core_j22_cpu_ml_bufb[25]), 
        .A2(n13325), .B1(n28478), .B2(n28540), .Y(n28479) );
  sky130_fd_sc_hd__o21ai_0 U33158 ( .A1(n28491), .A2(n28480), .B1(n28479), .Y(
        j202_soc_core_j22_cpu_ml_N421) );
  sky130_fd_sc_hd__o22a_1 U33159 ( .A1(n28481), .A2(n28512), .B1(n28538), .B2(
        n26456), .X(n28482) );
  sky130_fd_sc_hd__nand2_1 U33160 ( .A(n28535), .B(n28482), .Y(
        j202_soc_core_j22_cpu_ml_N363) );
  sky130_fd_sc_hd__nand2_1 U33161 ( .A(n28483), .B(n28539), .Y(n28486) );
  sky130_fd_sc_hd__a22oi_1 U33162 ( .A1(j202_soc_core_j22_cpu_ml_bufb[24]), 
        .A2(n13325), .B1(n28484), .B2(n28540), .Y(n28485) );
  sky130_fd_sc_hd__nand2_1 U33163 ( .A(n28486), .B(n28485), .Y(
        j202_soc_core_j22_cpu_ml_N420) );
  sky130_fd_sc_hd__o22a_1 U33164 ( .A1(n28487), .A2(n28512), .B1(n28538), .B2(
        n25245), .X(n28488) );
  sky130_fd_sc_hd__nand2_1 U33165 ( .A(n28535), .B(n28488), .Y(
        j202_soc_core_j22_cpu_ml_N362) );
  sky130_fd_sc_hd__a22oi_1 U33166 ( .A1(j202_soc_core_j22_cpu_ml_bufb[23]), 
        .A2(n13325), .B1(n28489), .B2(n28540), .Y(n28490) );
  sky130_fd_sc_hd__o21ai_1 U33167 ( .A1(n28491), .A2(n11180), .B1(n28490), .Y(
        j202_soc_core_j22_cpu_ml_N419) );
  sky130_fd_sc_hd__a22oi_1 U33168 ( .A1(n28533), .A2(n28493), .B1(n12396), 
        .B2(n28524), .Y(n28494) );
  sky130_fd_sc_hd__nand2_1 U33169 ( .A(n28535), .B(n28494), .Y(
        j202_soc_core_j22_cpu_ml_N361) );
  sky130_fd_sc_hd__nand2_1 U33170 ( .A(n12402), .B(n28539), .Y(n28497) );
  sky130_fd_sc_hd__a22oi_1 U33171 ( .A1(j202_soc_core_j22_cpu_ml_bufb[22]), 
        .A2(n13325), .B1(n28495), .B2(n28540), .Y(n28496) );
  sky130_fd_sc_hd__nand2_1 U33172 ( .A(n28497), .B(n28496), .Y(
        j202_soc_core_j22_cpu_ml_N418) );
  sky130_fd_sc_hd__a22oi_1 U33173 ( .A1(n28533), .A2(n28499), .B1(n12222), 
        .B2(n28524), .Y(n28500) );
  sky130_fd_sc_hd__nand2_1 U33174 ( .A(n28535), .B(n28500), .Y(
        j202_soc_core_j22_cpu_ml_N360) );
  sky130_fd_sc_hd__nand2_1 U33175 ( .A(n28501), .B(n28539), .Y(n28504) );
  sky130_fd_sc_hd__a22oi_1 U33176 ( .A1(j202_soc_core_j22_cpu_ml_bufb[21]), 
        .A2(n13325), .B1(n28502), .B2(n28540), .Y(n28503) );
  sky130_fd_sc_hd__nand2_1 U33177 ( .A(n28504), .B(n28503), .Y(
        j202_soc_core_j22_cpu_ml_N417) );
  sky130_fd_sc_hd__o22a_1 U33178 ( .A1(n28506), .A2(n28512), .B1(n28538), .B2(
        n28505), .X(n28507) );
  sky130_fd_sc_hd__nand2_1 U33179 ( .A(n28535), .B(n28507), .Y(
        j202_soc_core_j22_cpu_ml_N359) );
  sky130_fd_sc_hd__nand2_1 U33180 ( .A(n28508), .B(n28539), .Y(n28511) );
  sky130_fd_sc_hd__a22oi_1 U33181 ( .A1(j202_soc_core_j22_cpu_ml_bufb[20]), 
        .A2(n13325), .B1(n28509), .B2(n28540), .Y(n28510) );
  sky130_fd_sc_hd__nand2_1 U33182 ( .A(n28511), .B(n28510), .Y(
        j202_soc_core_j22_cpu_ml_N416) );
  sky130_fd_sc_hd__o22a_1 U33183 ( .A1(n28513), .A2(n28512), .B1(n28538), .B2(
        n25720), .X(n28514) );
  sky130_fd_sc_hd__nand2_1 U33184 ( .A(n28535), .B(n28514), .Y(
        j202_soc_core_j22_cpu_ml_N357) );
  sky130_fd_sc_hd__a22oi_1 U33185 ( .A1(j202_soc_core_j22_cpu_ml_bufb[19]), 
        .A2(n13325), .B1(n28515), .B2(n28540), .Y(n28516) );
  sky130_fd_sc_hd__nand2_1 U33186 ( .A(n28517), .B(n28516), .Y(
        j202_soc_core_j22_cpu_ml_N415) );
  sky130_fd_sc_hd__a22oi_1 U33187 ( .A1(n28533), .A2(n28519), .B1(n28518), 
        .B2(n28524), .Y(n28520) );
  sky130_fd_sc_hd__nand2_1 U33188 ( .A(n28535), .B(n28520), .Y(
        j202_soc_core_j22_cpu_ml_N356) );
  sky130_fd_sc_hd__a22oi_1 U33189 ( .A1(j202_soc_core_j22_cpu_ml_bufb[18]), 
        .A2(n13325), .B1(n28521), .B2(n28540), .Y(n28522) );
  sky130_fd_sc_hd__nand2_1 U33190 ( .A(n28523), .B(n28522), .Y(
        j202_soc_core_j22_cpu_ml_N414) );
  sky130_fd_sc_hd__a22oi_1 U33191 ( .A1(n28533), .A2(n28526), .B1(n28525), 
        .B2(n28524), .Y(n28527) );
  sky130_fd_sc_hd__nand2_1 U33192 ( .A(n28535), .B(n28527), .Y(
        j202_soc_core_j22_cpu_ml_N355) );
  sky130_fd_sc_hd__nand2_1 U33193 ( .A(n12431), .B(n28539), .Y(n28531) );
  sky130_fd_sc_hd__a22oi_1 U33194 ( .A1(j202_soc_core_j22_cpu_ml_bufb[17]), 
        .A2(n13325), .B1(n12354), .B2(n28540), .Y(n28530) );
  sky130_fd_sc_hd__nand2_1 U33195 ( .A(n28531), .B(n28530), .Y(
        j202_soc_core_j22_cpu_ml_N413) );
  sky130_fd_sc_hd__nand2_1 U33196 ( .A(n28534), .B(n28533), .Y(n28536) );
  sky130_fd_sc_hd__o211ai_1 U33197 ( .A1(n28538), .A2(n28537), .B1(n28536), 
        .C1(n28535), .Y(j202_soc_core_j22_cpu_ml_N354) );
  sky130_fd_sc_hd__nand2_1 U33198 ( .A(n11442), .B(n28539), .Y(n28543) );
  sky130_fd_sc_hd__a22oi_1 U33199 ( .A1(j202_soc_core_j22_cpu_ml_bufb[16]), 
        .A2(n13325), .B1(n28541), .B2(n28540), .Y(n28542) );
  sky130_fd_sc_hd__nand2_1 U33200 ( .A(n28543), .B(n28542), .Y(
        j202_soc_core_j22_cpu_ml_N412) );
  sky130_fd_sc_hd__nand2_1 U33201 ( .A(n28545), .B(
        j202_soc_core_bldc_core_00_wdata[10]), .Y(n28544) );
  sky130_fd_sc_hd__o21ai_1 U33202 ( .A1(n28546), .A2(n28545), .B1(n28544), .Y(
        n56) );
  sky130_fd_sc_hd__nand2_1 U33203 ( .A(n28547), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[11]), .Y(n28550) );
  sky130_fd_sc_hd__nand2_1 U33204 ( .A(n28548), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .Y(n28549) );
  sky130_fd_sc_hd__xor2_1 U33205 ( .A(n28550), .B(n28549), .X(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[11]) );
  sky130_fd_sc_hd__o22ai_1 U33206 ( .A1(n29163), .A2(n28553), .B1(n28552), 
        .B2(n28551), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__nand2_1 U33208 ( .A(n29169), .B(n28555), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[0]) );
  sky130_fd_sc_hd__a211oi_1 U33209 ( .A1(n28558), .A2(n28557), .B1(n28556), 
        .C1(n28564), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[5])
         );
  sky130_fd_sc_hd__a211oi_1 U33210 ( .A1(n28561), .A2(n28560), .B1(n28564), 
        .C1(n28559), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[7])
         );
  sky130_fd_sc_hd__xor2_1 U33211 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[9]), .B(n28562), .X(
        n28563) );
  sky130_fd_sc_hd__nor2_1 U33212 ( .A(n28564), .B(n28563), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[9]) );
  sky130_fd_sc_hd__nand2_1 U33214 ( .A(n29171), .B(n28565), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[0]) );
  sky130_fd_sc_hd__a211oi_1 U33215 ( .A1(n28567), .A2(n28566), .B1(n28568), 
        .C1(n28583), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[1])
         );
  sky130_fd_sc_hd__o21ai_1 U33216 ( .A1(n28568), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[2]), .B1(n28570), .Y(
        n28569) );
  sky130_fd_sc_hd__nor2_1 U33217 ( .A(n28569), .B(n28583), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[2]) );
  sky130_fd_sc_hd__a211oi_1 U33218 ( .A1(n28571), .A2(n28570), .B1(n28572), 
        .C1(n28583), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[3])
         );
  sky130_fd_sc_hd__o21ai_1 U33219 ( .A1(n28572), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[4]), .B1(n28574), .Y(
        n28573) );
  sky130_fd_sc_hd__nor2_1 U33220 ( .A(n28573), .B(n28583), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[4]) );
  sky130_fd_sc_hd__a211oi_1 U33221 ( .A1(n28575), .A2(n28574), .B1(n28576), 
        .C1(n28583), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[5])
         );
  sky130_fd_sc_hd__nor2_1 U33223 ( .A(n28583), .B(n28577), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[6]) );
  sky130_fd_sc_hd__a211oi_1 U33224 ( .A1(n28580), .A2(n28579), .B1(n28583), 
        .C1(n28578), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[7])
         );
  sky130_fd_sc_hd__xor2_1 U33225 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[9]), .B(n28581), .X(
        n28582) );
  sky130_fd_sc_hd__nor2_1 U33226 ( .A(n28583), .B(n28582), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[9]) );
  sky130_fd_sc_hd__nand4_1 U33227 ( .A(n28586), .B(j202_soc_core_uart_sio_ce), 
        .C(n28585), .D(n28584), .Y(n28587) );
  sky130_fd_sc_hd__nand2_1 U33228 ( .A(n28587), .B(n29828), .Y(
        j202_soc_core_uart_TOP_N16) );
  sky130_fd_sc_hd__nand2_1 U33229 ( .A(n12069), .B(n29099), .Y(n10717) );
  sky130_fd_sc_hd__nand2b_1 U33230 ( .A_N(j202_soc_core_uart_TOP_rxd_s), .B(
        j202_soc_core_uart_TOP_rxd_r), .Y(n28588) );
  sky130_fd_sc_hd__o211ai_1 U33231 ( .A1(j202_soc_core_uart_TOP_rx_go), .A2(
        n28588), .B1(n28593), .C1(n29830), .Y(j202_soc_core_uart_TOP_N85) );
  sky130_fd_sc_hd__a21oi_1 U33232 ( .A1(n29172), .A2(
        j202_soc_core_uart_TOP_rx_bit_cnt[1]), .B1(n28589), .Y(n28590) );
  sky130_fd_sc_hd__o21ai_1 U33233 ( .A1(n28593), .A2(n28590), .B1(n29830), .Y(
        j202_soc_core_uart_TOP_N87) );
  sky130_fd_sc_hd__xor2_1 U33234 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[3]), 
        .B(n28591), .X(n28592) );
  sky130_fd_sc_hd__o21ai_1 U33235 ( .A1(n28593), .A2(n28592), .B1(n29828), .Y(
        j202_soc_core_uart_TOP_N89) );
  sky130_fd_sc_hd__nand2_1 U33237 ( .A(n29306), .B(n29828), .Y(
        j202_soc_core_uart_TOP_N57) );
  sky130_fd_sc_hd__xor2_1 U33238 ( .A(n28594), .B(
        j202_soc_core_uart_TOP_tx_bit_cnt[3]), .X(n28596) );
  sky130_fd_sc_hd__o21ai_1 U33239 ( .A1(n28596), .A2(n28595), .B1(n29827), .Y(
        j202_soc_core_uart_TOP_N61) );
  sky130_fd_sc_hd__nand2_1 U33240 ( .A(n28597), .B(n12069), .Y(
        j202_soc_core_uart_BRG_N55) );
  sky130_fd_sc_hd__nor2_1 U33241 ( .A(j202_soc_core_uart_BRG_cnt[1]), .B(
        n28598), .Y(n28599) );
  sky130_fd_sc_hd__nor2_1 U33242 ( .A(n28599), .B(n29602), .Y(n28600) );
  sky130_fd_sc_hd__nor2_1 U33243 ( .A(n29609), .B(n28600), .Y(
        j202_soc_core_uart_BRG_N57) );
  sky130_fd_sc_hd__nand2_1 U33244 ( .A(j202_soc_core_uart_BRG_ps[1]), .B(
        j202_soc_core_uart_BRG_ps[0]), .Y(n28603) );
  sky130_fd_sc_hd__o21ai_1 U33245 ( .A1(j202_soc_core_uart_BRG_ps[1]), .A2(
        j202_soc_core_uart_BRG_ps[0]), .B1(n28603), .Y(n28602) );
  sky130_fd_sc_hd__nand2_1 U33246 ( .A(n28601), .B(n29745), .Y(n28623) );
  sky130_fd_sc_hd__nor2_1 U33247 ( .A(n28602), .B(n28623), .Y(
        j202_soc_core_uart_BRG_N13) );
  sky130_fd_sc_hd__nor2_1 U33248 ( .A(j202_soc_core_uart_BRG_ps[0]), .B(n28623), .Y(j202_soc_core_uart_BRG_N12) );
  sky130_fd_sc_hd__nor2_1 U33249 ( .A(n28604), .B(n28603), .Y(n28608) );
  sky130_fd_sc_hd__o21ai_1 U33250 ( .A1(n28606), .A2(
        j202_soc_core_uart_BRG_ps[2]), .B1(n28605), .Y(n28607) );
  sky130_fd_sc_hd__nor2_1 U33251 ( .A(n28607), .B(n28623), .Y(
        j202_soc_core_uart_BRG_N14) );
  sky130_fd_sc_hd__nand2_1 U33252 ( .A(j202_soc_core_uart_BRG_ps[3]), .B(
        n28608), .Y(n28610) );
  sky130_fd_sc_hd__o21ai_1 U33253 ( .A1(j202_soc_core_uart_BRG_ps[3]), .A2(
        n28608), .B1(n28610), .Y(n28609) );
  sky130_fd_sc_hd__nor2_1 U33254 ( .A(n28609), .B(n28623), .Y(
        j202_soc_core_uart_BRG_N15) );
  sky130_fd_sc_hd__nor2_1 U33255 ( .A(n28611), .B(n28610), .Y(n28615) );
  sky130_fd_sc_hd__o21ai_1 U33256 ( .A1(n28613), .A2(
        j202_soc_core_uart_BRG_ps[4]), .B1(n28612), .Y(n28614) );
  sky130_fd_sc_hd__nor2_1 U33257 ( .A(n28614), .B(n28623), .Y(
        j202_soc_core_uart_BRG_N16) );
  sky130_fd_sc_hd__nand2_1 U33258 ( .A(j202_soc_core_uart_BRG_ps[5]), .B(
        n28615), .Y(n28617) );
  sky130_fd_sc_hd__o21ai_1 U33259 ( .A1(j202_soc_core_uart_BRG_ps[5]), .A2(
        n28615), .B1(n28617), .Y(n28616) );
  sky130_fd_sc_hd__nor2_1 U33260 ( .A(n28616), .B(n28623), .Y(
        j202_soc_core_uart_BRG_N17) );
  sky130_fd_sc_hd__nor2_1 U33261 ( .A(n28618), .B(n28617), .Y(n29176) );
  sky130_fd_sc_hd__nor2_1 U33263 ( .A(n28621), .B(n28623), .Y(
        j202_soc_core_uart_BRG_N18) );
  sky130_fd_sc_hd__nand2_1 U33264 ( .A(j202_soc_core_uart_BRG_br_cnt[1]), .B(
        j202_soc_core_uart_BRG_br_cnt[0]), .Y(n28643) );
  sky130_fd_sc_hd__nor2_1 U33265 ( .A(n28632), .B(n28643), .Y(n28631) );
  sky130_fd_sc_hd__nand2_1 U33266 ( .A(j202_soc_core_uart_BRG_br_cnt[3]), .B(
        n28631), .Y(n28625) );
  sky130_fd_sc_hd__nand3_1 U33268 ( .A(n28624), .B(
        j202_soc_core_uart_BRG_ps_clr), .C(n29745), .Y(n29177) );
  sky130_fd_sc_hd__nor2_1 U33269 ( .A(n28622), .B(n29177), .Y(
        j202_soc_core_uart_BRG_N38) );
  sky130_fd_sc_hd__nand2_1 U33270 ( .A(n29174), .B(n28624), .Y(n10716) );
  sky130_fd_sc_hd__nor2_1 U33271 ( .A(n28626), .B(n28625), .Y(n28627) );
  sky130_fd_sc_hd__a211oi_1 U33272 ( .A1(n28626), .A2(n28625), .B1(n28627), 
        .C1(n29177), .Y(j202_soc_core_uart_BRG_N39) );
  sky130_fd_sc_hd__nand2_1 U33273 ( .A(j202_soc_core_uart_BRG_br_cnt[5]), .B(
        n28627), .Y(n28629) );
  sky130_fd_sc_hd__o21ai_1 U33274 ( .A1(j202_soc_core_uart_BRG_br_cnt[5]), 
        .A2(n28627), .B1(n28629), .Y(n28628) );
  sky130_fd_sc_hd__nor2_1 U33275 ( .A(n28628), .B(n29177), .Y(
        j202_soc_core_uart_BRG_N40) );
  sky130_fd_sc_hd__nor2_1 U33276 ( .A(n28630), .B(n28629), .Y(n29180) );
  sky130_fd_sc_hd__a211oi_1 U33277 ( .A1(n28630), .A2(n28629), .B1(n29180), 
        .C1(n29177), .Y(j202_soc_core_uart_BRG_N41) );
  sky130_fd_sc_hd__nor2_1 U33278 ( .A(j202_soc_core_uart_BRG_br_cnt[0]), .B(
        n29177), .Y(j202_soc_core_uart_BRG_N35) );
  sky130_fd_sc_hd__a211oi_1 U33279 ( .A1(n28632), .A2(n28643), .B1(n28631), 
        .C1(n29177), .Y(j202_soc_core_uart_BRG_N37) );
  sky130_fd_sc_hd__xnor2_1 U33280 ( .A(j202_soc_core_uart_div1[2]), .B(
        j202_soc_core_uart_BRG_br_cnt[2]), .Y(n28636) );
  sky130_fd_sc_hd__xnor2_1 U33281 ( .A(j202_soc_core_uart_div1[6]), .B(
        j202_soc_core_uart_BRG_br_cnt[6]), .Y(n28635) );
  sky130_fd_sc_hd__xnor2_1 U33282 ( .A(j202_soc_core_uart_div1[4]), .B(
        j202_soc_core_uart_BRG_br_cnt[4]), .Y(n28634) );
  sky130_fd_sc_hd__xnor2_1 U33283 ( .A(j202_soc_core_uart_div1[7]), .B(
        j202_soc_core_uart_BRG_br_cnt[7]), .Y(n28633) );
  sky130_fd_sc_hd__nand4_1 U33284 ( .A(n28636), .B(n28635), .C(n28634), .D(
        n28633), .Y(n28642) );
  sky130_fd_sc_hd__xnor2_1 U33285 ( .A(j202_soc_core_uart_div1[5]), .B(
        j202_soc_core_uart_BRG_br_cnt[5]), .Y(n28640) );
  sky130_fd_sc_hd__xnor2_1 U33286 ( .A(j202_soc_core_uart_div1[1]), .B(
        j202_soc_core_uart_BRG_br_cnt[1]), .Y(n28639) );
  sky130_fd_sc_hd__xnor2_1 U33287 ( .A(j202_soc_core_uart_div1[3]), .B(
        j202_soc_core_uart_BRG_br_cnt[3]), .Y(n28638) );
  sky130_fd_sc_hd__xnor2_1 U33288 ( .A(j202_soc_core_uart_div1[0]), .B(
        j202_soc_core_uart_BRG_br_cnt[0]), .Y(n28637) );
  sky130_fd_sc_hd__nand4_1 U33289 ( .A(n28640), .B(n28639), .C(n28638), .D(
        n28637), .Y(n28641) );
  sky130_fd_sc_hd__nor2_1 U33290 ( .A(n28642), .B(n28641), .Y(
        j202_soc_core_uart_BRG_N47) );
  sky130_fd_sc_hd__o21ai_1 U33291 ( .A1(j202_soc_core_uart_BRG_br_cnt[1]), 
        .A2(j202_soc_core_uart_BRG_br_cnt[0]), .B1(n28643), .Y(n28644) );
  sky130_fd_sc_hd__nor2_1 U33292 ( .A(n28644), .B(n29177), .Y(
        j202_soc_core_uart_BRG_N36) );
  sky130_fd_sc_hd__nand2_1 U33293 ( .A(n28645), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[4]), .Y(n28646) );
  sky130_fd_sc_hd__a31oi_1 U33294 ( .A1(n28646), .A2(
        j202_soc_core_wbqspiflash_00_state[0]), .A3(n28648), .B1(n28651), .Y(
        j202_soc_core_wbqspiflash_00_N618) );
  sky130_fd_sc_hd__a21oi_1 U33295 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[5]), .A2(n28648), .B1(
        n28647), .Y(n28649) );
  sky130_fd_sc_hd__a21oi_1 U33296 ( .A1(n28649), .A2(n28650), .B1(n28651), .Y(
        j202_soc_core_wbqspiflash_00_N619) );
  sky130_fd_sc_hd__nand2_1 U33297 ( .A(n28650), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[6]), .Y(n28652) );
  sky130_fd_sc_hd__a31oi_1 U33298 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), 
        .A2(n28653), .A3(n28652), .B1(n28651), .Y(
        j202_soc_core_wbqspiflash_00_N620) );
  sky130_fd_sc_hd__a22oi_1 U33299 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[28]), .B1(n28887), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]), .Y(n28660) );
  sky130_fd_sc_hd__nand2_1 U33300 ( .A(n28836), .B(n28655), .Y(n28672) );
  sky130_fd_sc_hd__nand3_1 U33301 ( .A(n28672), .B(n28656), .C(n28671), .Y(
        n28657) );
  sky130_fd_sc_hd__a21oi_1 U33302 ( .A1(j202_soc_core_qspi_wb_addr[2]), .A2(
        n28677), .B1(n28657), .Y(n28659) );
  sky130_fd_sc_hd__nand2_1 U33303 ( .A(n28888), .B(
        j202_soc_core_qspi_wb_addr[20]), .Y(n28658) );
  sky130_fd_sc_hd__nand4_1 U33304 ( .A(n28661), .B(n28660), .C(n28659), .D(
        n28658), .Y(n10547) );
  sky130_fd_sc_hd__a21oi_1 U33305 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[30]), .B1(n28662), .Y(n28665)
         );
  sky130_fd_sc_hd__nand2_1 U33306 ( .A(n28887), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .Y(n28664) );
  sky130_fd_sc_hd__nand2_1 U33307 ( .A(n28888), .B(
        j202_soc_core_qspi_wb_addr[22]), .Y(n28663) );
  sky130_fd_sc_hd__nand4_1 U33308 ( .A(n28666), .B(n28665), .C(n28664), .D(
        n28663), .Y(n10545) );
  sky130_fd_sc_hd__a21oi_1 U33309 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[29]), .B1(n28668), .Y(n28681)
         );
  sky130_fd_sc_hd__nand3_1 U33310 ( .A(n28669), .B(
        j202_soc_core_wbqspiflash_00_state[2]), .C(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]), .Y(n28670) );
  sky130_fd_sc_hd__nand2_1 U33311 ( .A(n28671), .B(n28670), .Y(n28674) );
  sky130_fd_sc_hd__nor2_1 U33312 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .B(n28672), .Y(n28673)
         );
  sky130_fd_sc_hd__a211oi_1 U33313 ( .A1(j202_soc_core_qspi_wb_addr[21]), .A2(
        n28675), .B1(n28674), .C1(n28673), .Y(n28680) );
  sky130_fd_sc_hd__nand2_1 U33314 ( .A(n28677), .B(n28676), .Y(n28678) );
  sky130_fd_sc_hd__nand4_1 U33315 ( .A(n28681), .B(n28680), .C(n28679), .D(
        n28678), .Y(n10546) );
  sky130_fd_sc_hd__nand2_1 U33316 ( .A(n28683), .B(n28682), .Y(
        j202_soc_core_wbqspiflash_00_N86) );
  sky130_fd_sc_hd__nand3_1 U33317 ( .A(n28686), .B(n28685), .C(n28684), .Y(
        j202_soc_core_wbqspiflash_00_N594) );
  sky130_fd_sc_hd__a21oi_1 U33318 ( .A1(n28688), .A2(
        j202_soc_core_wbqspiflash_00_state[4]), .B1(n28687), .Y(n28689) );
  sky130_fd_sc_hd__a21oi_1 U33319 ( .A1(n28690), .A2(n28689), .B1(
        j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N747) );
  sky130_fd_sc_hd__a211o_1 U33320 ( .A1(U7_RSOP_1495_C3_DATA3_2), .A2(n29270), 
        .B1(n28714), .C1(n29603), .X(
        j202_soc_core_wbqspiflash_00_lldriver_N427) );
  sky130_fd_sc_hd__nand3_1 U33321 ( .A(n28693), .B(n28692), .C(n28691), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N424) );
  sky130_fd_sc_hd__nor3_1 U33322 ( .A(n29184), .B(n28695), .C(n28694), .Y(
        DP_OP_1508J1_126_2326_n6) );
  sky130_fd_sc_hd__nand2_1 U33323 ( .A(n28714), .B(n28727), .Y(n28699) );
  sky130_fd_sc_hd__nand2_1 U33324 ( .A(n28699), .B(n13045), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N426) );
  sky130_fd_sc_hd__o211ai_1 U33325 ( .A1(n28701), .A2(n28700), .B1(n28699), 
        .C1(n28698), .Y(j202_soc_core_wbqspiflash_00_lldriver_N425) );
  sky130_fd_sc_hd__o22ai_1 U33326 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_len[0]), .A2(n28898), .B1(n28703), 
        .B2(n28702), .Y(n28704) );
  sky130_fd_sc_hd__nor2_1 U33327 ( .A(n28704), .B(DP_OP_1508J1_126_2326_n3), 
        .Y(n28709) );
  sky130_fd_sc_hd__a21oi_1 U33328 ( .A1(DP_OP_1508J1_126_2326_n3), .A2(n28704), 
        .B1(n28709), .Y(n28707) );
  sky130_fd_sc_hd__nor2_1 U33329 ( .A(j202_soc_core_wbqspiflash_00_spi_len[0]), 
        .B(j202_soc_core_wbqspiflash_00_lldriver_N311), .Y(n28705) );
  sky130_fd_sc_hd__a21oi_1 U33330 ( .A1(n28714), .A2(
        j202_soc_core_wbqspiflash_00_spi_len[0]), .B1(n28705), .Y(n28706) );
  sky130_fd_sc_hd__o21ai_1 U33331 ( .A1(n28721), .A2(n28707), .B1(n28706), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N428) );
  sky130_fd_sc_hd__nor2_1 U33332 ( .A(n28717), .B(n28708), .Y(n28713) );
  sky130_fd_sc_hd__a22oi_1 U33333 ( .A1(n28713), .A2(n29603), .B1(n29270), 
        .B2(j202_soc_core_wbqspiflash_00_lldriver_spi_len[4]), .Y(n28710) );
  sky130_fd_sc_hd__nand2_1 U33334 ( .A(n28709), .B(n28710), .Y(n28719) );
  sky130_fd_sc_hd__a21oi_1 U33335 ( .A1(n28719), .A2(n28709), .B1(n28721), .Y(
        n28712) );
  sky130_fd_sc_hd__nand2_1 U33336 ( .A(n28719), .B(n28710), .Y(n28711) );
  sky130_fd_sc_hd__nand2_1 U33337 ( .A(n28712), .B(n28711), .Y(n28716) );
  sky130_fd_sc_hd__a22oi_1 U33338 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_len[1]), .A2(n28714), .B1(n29257), 
        .B2(n28713), .Y(n28715) );
  sky130_fd_sc_hd__nand2_1 U33339 ( .A(n28716), .B(n28715), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N429) );
  sky130_fd_sc_hd__a22oi_1 U33340 ( .A1(n28717), .A2(n29603), .B1(n29270), 
        .B2(j202_soc_core_wbqspiflash_00_lldriver_spi_len[5]), .Y(n28718) );
  sky130_fd_sc_hd__xnor2_1 U33341 ( .A(n28719), .B(n28718), .Y(n28720) );
  sky130_fd_sc_hd__o22ai_1 U33342 ( .A1(n28722), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B1(n28721), .B2(n28720), 
        .Y(j202_soc_core_wbqspiflash_00_lldriver_N430) );
  sky130_fd_sc_hd__nor2_1 U33343 ( .A(n28723), .B(n28724), .Y(
        j202_soc_core_wbqspiflash_00_N628) );
  sky130_fd_sc_hd__nor2_1 U33344 ( .A(n29139), .B(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N391) );
  sky130_fd_sc_hd__nor2_1 U33345 ( .A(n28725), .B(n28724), .Y(
        j202_soc_core_wbqspiflash_00_N629) );
  sky130_fd_sc_hd__nand2_1 U33346 ( .A(n29267), .B(n28727), .Y(n29261) );
  sky130_fd_sc_hd__a222oi_1 U33347 ( .A1(n29265), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[0]), .B1(n29264), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[0]), .C1(n29257), .C2(
        j202_soc_core_wbqspiflash_00_spi_in[1]), .Y(n28728) );
  sky130_fd_sc_hd__nand2_1 U33348 ( .A(n28730), .B(n28729), .Y(n28732) );
  sky130_fd_sc_hd__nand2_1 U33349 ( .A(n28732), .B(n28731), .Y(n28831) );
  sky130_fd_sc_hd__a222oi_1 U33350 ( .A1(n28831), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[4]), .B1(n28847), .B2(
        j202_soc_core_qspi_wb_addr[4]), .C1(n28886), .C2(
        j202_soc_core_wbqspiflash_00_spif_data[4]), .Y(n28733) );
  sky130_fd_sc_hd__nand2_1 U33351 ( .A(n28831), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[5]), .Y(n28736) );
  sky130_fd_sc_hd__nand2_1 U33352 ( .A(n28817), .B(n28734), .Y(n28743) );
  sky130_fd_sc_hd__a21oi_1 U33353 ( .A1(n28744), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[5]), .B1(n28743), .Y(n28735) );
  sky130_fd_sc_hd__o211ai_1 U33354 ( .A1(n28737), .A2(n28747), .B1(n28736), 
        .C1(n28735), .Y(n10570) );
  sky130_fd_sc_hd__a22oi_1 U33355 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[2]), .B1(n28831), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .Y(n28738) );
  sky130_fd_sc_hd__o21ai_1 U33356 ( .A1(n28739), .A2(n28751), .B1(n28738), .Y(
        n10573) );
  sky130_fd_sc_hd__a222oi_1 U33357 ( .A1(n29265), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[1]), .B1(n29264), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[1]), .C1(n29257), .C2(
        j202_soc_core_wbqspiflash_00_spi_in[2]), .Y(n28740) );
  sky130_fd_sc_hd__a222oi_1 U33358 ( .A1(n28831), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[6]), .B1(n28847), .B2(
        j202_soc_core_qspi_wb_addr[6]), .C1(n28886), .C2(
        j202_soc_core_wbqspiflash_00_spif_data[6]), .Y(n28741) );
  sky130_fd_sc_hd__a222oi_1 U33359 ( .A1(n28831), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .B1(n28886), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[3]), .C1(
        j202_soc_core_qspi_wb_addr[3]), .C2(n28847), .Y(n28742) );
  sky130_fd_sc_hd__nand2_1 U33360 ( .A(n28831), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[7]), .Y(n28746) );
  sky130_fd_sc_hd__a21oi_1 U33361 ( .A1(n28744), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[7]), .B1(n28743), .Y(n28745) );
  sky130_fd_sc_hd__o211ai_1 U33362 ( .A1(n28748), .A2(n28747), .B1(n28746), 
        .C1(n28745), .Y(n10568) );
  sky130_fd_sc_hd__a22o_1 U33363 ( .A1(n28848), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[0]), .B1(n28886), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[8]), .X(n28749) );
  sky130_fd_sc_hd__a21oi_1 U33364 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[8]), .A2(n28831), .B1(n28749), 
        .Y(n28750) );
  sky130_fd_sc_hd__o21ai_1 U33365 ( .A1(n28782), .A2(n28751), .B1(n28750), .Y(
        n10567) );
  sky130_fd_sc_hd__nand2_1 U33366 ( .A(n28847), .B(
        j202_soc_core_qspi_wb_addr[9]), .Y(n28755) );
  sky130_fd_sc_hd__nand2_1 U33367 ( .A(n28831), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[9]), .Y(n28754) );
  sky130_fd_sc_hd__nand2_1 U33368 ( .A(n28886), .B(
        j202_soc_core_wbqspiflash_00_spif_data[9]), .Y(n28752) );
  sky130_fd_sc_hd__nand4_1 U33369 ( .A(n28755), .B(n28754), .C(n28753), .D(
        n28752), .Y(n10566) );
  sky130_fd_sc_hd__nand2_1 U33370 ( .A(n28847), .B(
        j202_soc_core_qspi_wb_addr[10]), .Y(n28759) );
  sky130_fd_sc_hd__a22oi_1 U33371 ( .A1(n28848), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[2]), .B1(n28888), .B2(
        j202_soc_core_qspi_wb_addr[2]), .Y(n28758) );
  sky130_fd_sc_hd__a22oi_1 U33372 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[10]), .B1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .B2(n28887), .Y(n28757)
         );
  sky130_fd_sc_hd__nand2_1 U33373 ( .A(n28831), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[10]), .Y(n28756) );
  sky130_fd_sc_hd__nand4_1 U33374 ( .A(n28759), .B(n28758), .C(n28757), .D(
        n28756), .Y(n10565) );
  sky130_fd_sc_hd__nand2_1 U33375 ( .A(n28847), .B(
        j202_soc_core_qspi_wb_addr[11]), .Y(n28763) );
  sky130_fd_sc_hd__a22oi_1 U33376 ( .A1(n28848), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[3]), .B1(n28888), .B2(
        j202_soc_core_qspi_wb_addr[3]), .Y(n28762) );
  sky130_fd_sc_hd__a22oi_1 U33377 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[11]), .B1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .B2(n28887), .Y(n28761)
         );
  sky130_fd_sc_hd__nand2_1 U33378 ( .A(n28831), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[11]), .Y(n28760) );
  sky130_fd_sc_hd__nand4_1 U33379 ( .A(n28763), .B(n28762), .C(n28761), .D(
        n28760), .Y(n10564) );
  sky130_fd_sc_hd__nand2_1 U33380 ( .A(n28847), .B(
        j202_soc_core_qspi_wb_addr[12]), .Y(n28767) );
  sky130_fd_sc_hd__a22oi_1 U33381 ( .A1(n28848), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[4]), .B1(n28888), .B2(
        j202_soc_core_qspi_wb_addr[4]), .Y(n28766) );
  sky130_fd_sc_hd__a22oi_1 U33382 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[12]), .B1(n28887), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[4]), .Y(n28765) );
  sky130_fd_sc_hd__nand2_1 U33383 ( .A(n28831), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[12]), .Y(n28764) );
  sky130_fd_sc_hd__nand4_1 U33384 ( .A(n28767), .B(n28766), .C(n28765), .D(
        n28764), .Y(n10563) );
  sky130_fd_sc_hd__nand2_1 U33385 ( .A(n28847), .B(
        j202_soc_core_qspi_wb_addr[13]), .Y(n28771) );
  sky130_fd_sc_hd__a22oi_1 U33386 ( .A1(n28848), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[5]), .B1(n28888), .B2(
        j202_soc_core_qspi_wb_addr[5]), .Y(n28770) );
  sky130_fd_sc_hd__a22oi_1 U33387 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[13]), .B1(n28887), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[5]), .Y(n28769) );
  sky130_fd_sc_hd__nand2_1 U33388 ( .A(n28831), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[13]), .Y(n28768) );
  sky130_fd_sc_hd__nand4_1 U33389 ( .A(n28771), .B(n28770), .C(n28769), .D(
        n28768), .Y(n10562) );
  sky130_fd_sc_hd__nand2_1 U33390 ( .A(n28847), .B(
        j202_soc_core_qspi_wb_addr[14]), .Y(n28775) );
  sky130_fd_sc_hd__a22oi_1 U33391 ( .A1(n28848), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[6]), .B1(n28888), .B2(
        j202_soc_core_qspi_wb_addr[6]), .Y(n28774) );
  sky130_fd_sc_hd__a22oi_1 U33392 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[14]), .B1(n28887), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[6]), .Y(n28773) );
  sky130_fd_sc_hd__nand2_1 U33393 ( .A(n28831), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]), .Y(n28772) );
  sky130_fd_sc_hd__nand4_1 U33394 ( .A(n28775), .B(n28774), .C(n28773), .D(
        n28772), .Y(n10561) );
  sky130_fd_sc_hd__nand2_1 U33395 ( .A(n28847), .B(
        j202_soc_core_qspi_wb_addr[15]), .Y(n28779) );
  sky130_fd_sc_hd__a22oi_1 U33396 ( .A1(n28848), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[7]), .B1(n28888), .B2(
        j202_soc_core_qspi_wb_addr[7]), .Y(n28778) );
  sky130_fd_sc_hd__a22oi_1 U33397 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[15]), .B1(n28887), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[7]), .Y(n28777) );
  sky130_fd_sc_hd__nand2_1 U33398 ( .A(n28831), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[15]), .Y(n28776) );
  sky130_fd_sc_hd__nand4_1 U33399 ( .A(n28779), .B(n28778), .C(n28777), .D(
        n28776), .Y(n10560) );
  sky130_fd_sc_hd__nand2_1 U33400 ( .A(n28828), .B(
        j202_soc_core_wbqspiflash_00_spif_data[0]), .Y(n28785) );
  sky130_fd_sc_hd__o21ai_1 U33401 ( .A1(n29087), .A2(n28780), .B1(n28785), .Y(
        j202_soc_core_wbqspiflash_00_N605) );
  sky130_fd_sc_hd__a22oi_1 U33402 ( .A1(n28814), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[14]), .B1(n28886), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[16]), .Y(n28781) );
  sky130_fd_sc_hd__o21ai_1 U33403 ( .A1(n28817), .A2(n28782), .B1(n28781), .Y(
        n28783) );
  sky130_fd_sc_hd__a21oi_1 U33404 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]), .A2(n28831), .B1(n28783), .Y(n28787) );
  sky130_fd_sc_hd__a22oi_1 U33405 ( .A1(n28848), .A2(
        j202_soc_core_wbqspiflash_00_last_status[0]), .B1(n28887), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[8]), .Y(n28786) );
  sky130_fd_sc_hd__nand2_1 U33406 ( .A(n28847), .B(
        j202_soc_core_qspi_wb_addr[16]), .Y(n28784) );
  sky130_fd_sc_hd__nand4_1 U33407 ( .A(n28787), .B(n28786), .C(n28785), .D(
        n28784), .Y(n10559) );
  sky130_fd_sc_hd__a22o_1 U33408 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]), .A2(n28831), .B1(n28887), .B2(j202_soc_core_wbqspiflash_00_w_spif_addr[9]), .X(n28788) );
  sky130_fd_sc_hd__a21oi_1 U33409 ( .A1(n28848), .A2(
        j202_soc_core_wbqspiflash_00_last_status[1]), .B1(n28788), .Y(n28792)
         );
  sky130_fd_sc_hd__a22o_1 U33410 ( .A1(n28814), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[15]), .B1(n28886), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[17]), .X(n28789) );
  sky130_fd_sc_hd__a21oi_1 U33411 ( .A1(n28888), .A2(
        j202_soc_core_qspi_wb_addr[9]), .B1(n28789), .Y(n28791) );
  sky130_fd_sc_hd__nand2_1 U33412 ( .A(n28828), .B(
        j202_soc_core_wbqspiflash_00_spif_data[1]), .Y(n29083) );
  sky130_fd_sc_hd__nand2_1 U33413 ( .A(n28847), .B(
        j202_soc_core_qspi_wb_addr[17]), .Y(n28790) );
  sky130_fd_sc_hd__nand4_1 U33414 ( .A(n28792), .B(n28791), .C(n29083), .D(
        n28790), .Y(n10558) );
  sky130_fd_sc_hd__a22o_1 U33415 ( .A1(n28887), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[10]), .B1(n28847), .B2(
        j202_soc_core_qspi_wb_addr[18]), .X(n28793) );
  sky130_fd_sc_hd__a21oi_1 U33416 ( .A1(n28848), .A2(
        j202_soc_core_wbqspiflash_00_last_status[2]), .B1(n28793), .Y(n28797)
         );
  sky130_fd_sc_hd__a22o_1 U33417 ( .A1(n28814), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[16]), .B1(n28886), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[18]), .X(n28794) );
  sky130_fd_sc_hd__a21oi_1 U33418 ( .A1(n28888), .A2(
        j202_soc_core_qspi_wb_addr[10]), .B1(n28794), .Y(n28796) );
  sky130_fd_sc_hd__nand2_1 U33419 ( .A(n28828), .B(
        j202_soc_core_wbqspiflash_00_spif_data[2]), .Y(n29085) );
  sky130_fd_sc_hd__nand2_1 U33420 ( .A(n28831), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .Y(n28795) );
  sky130_fd_sc_hd__nand4_1 U33421 ( .A(n28797), .B(n28796), .C(n29085), .D(
        n28795), .Y(n10557) );
  sky130_fd_sc_hd__nand2_1 U33422 ( .A(n28828), .B(
        j202_soc_core_wbqspiflash_00_spif_data[3]), .Y(n28803) );
  sky130_fd_sc_hd__o21ai_1 U33423 ( .A1(n29087), .A2(n28798), .B1(n28803), .Y(
        j202_soc_core_wbqspiflash_00_N608) );
  sky130_fd_sc_hd__a22oi_1 U33424 ( .A1(n28814), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[17]), .B1(n28886), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[19]), .Y(n28799) );
  sky130_fd_sc_hd__o21ai_1 U33425 ( .A1(n28817), .A2(n28800), .B1(n28799), .Y(
        n28801) );
  sky130_fd_sc_hd__a21oi_1 U33426 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .A2(n28831), .B1(n28801), .Y(n28805) );
  sky130_fd_sc_hd__a22oi_1 U33427 ( .A1(n28848), .A2(
        j202_soc_core_wbqspiflash_00_last_status[3]), .B1(n28887), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[11]), .Y(n28804) );
  sky130_fd_sc_hd__nand2_1 U33428 ( .A(n28847), .B(
        j202_soc_core_qspi_wb_addr[19]), .Y(n28802) );
  sky130_fd_sc_hd__nand4_1 U33429 ( .A(n28805), .B(n28804), .C(n28803), .D(
        n28802), .Y(n10556) );
  sky130_fd_sc_hd__nand2_1 U33430 ( .A(n28828), .B(
        j202_soc_core_wbqspiflash_00_spif_data[4]), .Y(n28811) );
  sky130_fd_sc_hd__o21ai_1 U33431 ( .A1(n29087), .A2(n28806), .B1(n28811), .Y(
        j202_soc_core_wbqspiflash_00_N609) );
  sky130_fd_sc_hd__a22oi_1 U33432 ( .A1(n28814), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[18]), .B1(n28886), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[20]), .Y(n28807) );
  sky130_fd_sc_hd__o21ai_1 U33433 ( .A1(n28817), .A2(n28808), .B1(n28807), .Y(
        n28809) );
  sky130_fd_sc_hd__a21oi_1 U33434 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]), .A2(n28831), .B1(n28809), .Y(n28813) );
  sky130_fd_sc_hd__a22oi_1 U33435 ( .A1(n28848), .A2(
        j202_soc_core_wbqspiflash_00_last_status[4]), .B1(n28887), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[12]), .Y(n28812) );
  sky130_fd_sc_hd__nand2_1 U33436 ( .A(n28847), .B(
        j202_soc_core_qspi_wb_addr[20]), .Y(n28810) );
  sky130_fd_sc_hd__nand4_1 U33437 ( .A(n28813), .B(n28812), .C(n28811), .D(
        n28810), .Y(n10555) );
  sky130_fd_sc_hd__a22oi_1 U33438 ( .A1(n28814), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[19]), .B1(n28886), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[21]), .Y(n28815) );
  sky130_fd_sc_hd__o21ai_1 U33439 ( .A1(n28817), .A2(n28816), .B1(n28815), .Y(
        n28818) );
  sky130_fd_sc_hd__a21oi_1 U33440 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]), .A2(n28831), .B1(n28818), .Y(n28822) );
  sky130_fd_sc_hd__a22oi_1 U33441 ( .A1(n28848), .A2(
        j202_soc_core_wbqspiflash_00_last_status[5]), .B1(n28887), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[13]), .Y(n28821) );
  sky130_fd_sc_hd__nand2_1 U33442 ( .A(n28847), .B(
        j202_soc_core_qspi_wb_addr[21]), .Y(n28819) );
  sky130_fd_sc_hd__nand4_1 U33443 ( .A(n28822), .B(n28821), .C(n28820), .D(
        n28819), .Y(n10554) );
  sky130_fd_sc_hd__a22o_1 U33444 ( .A1(
        j202_soc_core_wbqspiflash_00_last_status[6]), .A2(n28848), .B1(n28888), 
        .B2(j202_soc_core_qspi_wb_addr[14]), .X(n28823) );
  sky130_fd_sc_hd__a21oi_1 U33445 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .A2(n28831), .B1(n28823), .Y(n28827) );
  sky130_fd_sc_hd__a22oi_1 U33446 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[22]), .B1(n28887), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]), .Y(n28826) );
  sky130_fd_sc_hd__nand2_1 U33447 ( .A(n28847), .B(
        j202_soc_core_qspi_wb_addr[22]), .Y(n28824) );
  sky130_fd_sc_hd__nand4_1 U33448 ( .A(n28827), .B(n28826), .C(n28825), .D(
        n28824), .Y(n10553) );
  sky130_fd_sc_hd__nand2_1 U33449 ( .A(n28828), .B(
        j202_soc_core_wbqspiflash_00_spif_data[7]), .Y(n28833) );
  sky130_fd_sc_hd__a22o_1 U33451 ( .A1(n28848), .A2(
        j202_soc_core_wbqspiflash_00_last_status[7]), .B1(n28888), .B2(
        j202_soc_core_qspi_wb_addr[15]), .X(n28830) );
  sky130_fd_sc_hd__a21oi_1 U33452 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]), .A2(n28831), .B1(n28830), .Y(n28835) );
  sky130_fd_sc_hd__a22oi_1 U33453 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[23]), .B1(n28887), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[15]), .Y(n28834) );
  sky130_fd_sc_hd__nand2_1 U33454 ( .A(n28847), .B(
        j202_soc_core_qspi_wb_addr[23]), .Y(n28832) );
  sky130_fd_sc_hd__nand4_1 U33455 ( .A(n28835), .B(n28834), .C(n28833), .D(
        n28832), .Y(n10552) );
  sky130_fd_sc_hd__a22oi_1 U33456 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[24]), .B1(n28887), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]), .Y(n28856) );
  sky130_fd_sc_hd__nand2_1 U33457 ( .A(n28837), .B(n28836), .Y(n28855) );
  sky130_fd_sc_hd__and3_1 U33458 ( .A(n28841), .B(n28840), .C(n28839), .X(
        n28880) );
  sky130_fd_sc_hd__nand2_1 U33459 ( .A(n28843), .B(n28842), .Y(n28845) );
  sky130_fd_sc_hd__nand3_1 U33460 ( .A(n28845), .B(n28844), .C(n29276), .Y(
        n28877) );
  sky130_fd_sc_hd__a21o_1 U33461 ( .A1(j202_soc_core_qspi_wb_addr[16]), .A2(
        n28880), .B1(n28877), .X(n28846) );
  sky130_fd_sc_hd__nor4_1 U33462 ( .A(n28849), .B(n28848), .C(n28847), .D(
        n28846), .Y(n28854) );
  sky130_fd_sc_hd__nand3_1 U33463 ( .A(n28852), .B(n28851), .C(n28850), .Y(
        n28853) );
  sky130_fd_sc_hd__nand4_1 U33464 ( .A(n28856), .B(n28855), .C(n28854), .D(
        n28853), .Y(n10551) );
  sky130_fd_sc_hd__nor3_1 U33465 ( .A(n28859), .B(n28858), .C(n28857), .Y(
        n28860) );
  sky130_fd_sc_hd__a211oi_1 U33466 ( .A1(n28888), .A2(
        j202_soc_core_qspi_wb_addr[17]), .B1(n28879), .C1(n28860), .Y(n28875)
         );
  sky130_fd_sc_hd__nor2_1 U33467 ( .A(n28861), .B(n28878), .Y(n28862) );
  sky130_fd_sc_hd__o21a_1 U33468 ( .A1(n28864), .A2(n28863), .B1(n28862), .X(
        n28874) );
  sky130_fd_sc_hd__a211oi_1 U33469 ( .A1(j202_soc_core_qspi_wb_addr[24]), .A2(
        n28867), .B1(n28866), .C1(n28865), .Y(n28868) );
  sky130_fd_sc_hd__a21oi_1 U33470 ( .A1(
        j202_soc_core_wbqspiflash_00_spif_data[25]), .A2(n28869), .B1(n28868), 
        .Y(n28873) );
  sky130_fd_sc_hd__nand3_1 U33471 ( .A(n28871), .B(n28870), .C(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]), .Y(n28872) );
  sky130_fd_sc_hd__nand4_1 U33472 ( .A(n28875), .B(n28874), .C(n28873), .D(
        n28872), .Y(n10550) );
  sky130_fd_sc_hd__a22o_1 U33473 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[26]), .B1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .B2(n28887), .X(n28876)
         );
  sky130_fd_sc_hd__nor3_1 U33474 ( .A(n28878), .B(n28877), .C(n28876), .Y(
        n28883) );
  sky130_fd_sc_hd__a21oi_1 U33475 ( .A1(j202_soc_core_qspi_wb_addr[18]), .A2(
        n28880), .B1(n28879), .Y(n28881) );
  sky130_fd_sc_hd__nand3_1 U33476 ( .A(n28883), .B(n28882), .C(n28881), .Y(
        n10549) );
  sky130_fd_sc_hd__a21oi_1 U33477 ( .A1(n28886), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[27]), .B1(n28885), .Y(n28891)
         );
  sky130_fd_sc_hd__nand2_1 U33478 ( .A(n28887), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .Y(n28890) );
  sky130_fd_sc_hd__nand2_1 U33479 ( .A(n28888), .B(
        j202_soc_core_qspi_wb_addr[19]), .Y(n28889) );
  sky130_fd_sc_hd__nand4_1 U33480 ( .A(n28892), .B(n28891), .C(n28890), .D(
        n28889), .Y(n10548) );
  sky130_fd_sc_hd__nor2_1 U33481 ( .A(n28895), .B(n28894), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N353) );
  sky130_fd_sc_hd__o22ai_1 U33482 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[30]), .B1(n28896), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[27]), .Y(n28897) );
  sky130_fd_sc_hd__nor2_1 U33483 ( .A(n28898), .B(n28897), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N389) );
  sky130_fd_sc_hd__nand2_1 U33484 ( .A(n28910), .B(j202_soc_core_uart_din_i[0]), .Y(n28899) );
  sky130_fd_sc_hd__o21ai_1 U33485 ( .A1(n28900), .A2(n28910), .B1(n28899), .Y(
        n92) );
  sky130_fd_sc_hd__nand2_1 U33486 ( .A(n28910), .B(j202_soc_core_uart_din_i[1]), .Y(n28901) );
  sky130_fd_sc_hd__nand2_1 U33488 ( .A(n28910), .B(j202_soc_core_uart_din_i[2]), .Y(n28903) );
  sky130_fd_sc_hd__o21ai_1 U33489 ( .A1(n28915), .A2(n28910), .B1(n28903), .Y(
        n86) );
  sky130_fd_sc_hd__nand2_1 U33490 ( .A(n28910), .B(j202_soc_core_uart_din_i[3]), .Y(n28904) );
  sky130_fd_sc_hd__o21ai_1 U33491 ( .A1(n28922), .A2(n28910), .B1(n28904), .Y(
        n81) );
  sky130_fd_sc_hd__nand2_1 U33492 ( .A(n28910), .B(j202_soc_core_uart_din_i[4]), .Y(n28905) );
  sky130_fd_sc_hd__o21ai_1 U33493 ( .A1(n28906), .A2(n28910), .B1(n28905), .Y(
        n76) );
  sky130_fd_sc_hd__nand2_1 U33494 ( .A(n28910), .B(j202_soc_core_uart_din_i[5]), .Y(n28907) );
  sky130_fd_sc_hd__o21ai_1 U33495 ( .A1(n28935), .A2(n28910), .B1(n28907), .Y(
        n102) );
  sky130_fd_sc_hd__nand2_1 U33496 ( .A(n28910), .B(j202_soc_core_uart_din_i[6]), .Y(n28908) );
  sky130_fd_sc_hd__o21ai_1 U33497 ( .A1(n28942), .A2(n28910), .B1(n28908), .Y(
        n101) );
  sky130_fd_sc_hd__nand2_1 U33498 ( .A(n28910), .B(j202_soc_core_uart_din_i[7]), .Y(n28909) );
  sky130_fd_sc_hd__o21ai_1 U33499 ( .A1(n28949), .A2(n28910), .B1(n28909), .Y(
        n100) );
  sky130_fd_sc_hd__nor2_1 U33500 ( .A(n29088), .B(n28911), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N12) );
  sky130_fd_sc_hd__nor2_1 U33501 ( .A(n29088), .B(n28912), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N13) );
  sky130_fd_sc_hd__nor2_1 U33502 ( .A(n29088), .B(n28913), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N14) );
  sky130_fd_sc_hd__nand2_1 U33503 ( .A(n29827), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[12]), .Y(n28986) );
  sky130_fd_sc_hd__nand2_1 U33504 ( .A(n29830), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[17]), .Y(n29023) );
  sky130_fd_sc_hd__nand2_1 U33505 ( .A(n28914), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[19]), .Y(n29037) );
  sky130_fd_sc_hd__a21oi_1 U33506 ( .A1(n29827), .A2(n28915), .B1(n29061), .Y(
        n28920) );
  sky130_fd_sc_hd__o22ai_1 U33507 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[2]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[2]), .B1(n28916), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[2]), .Y(n28917)
         );
  sky130_fd_sc_hd__a21oi_1 U33508 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[2]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[2]), .B1(n28917), 
        .Y(n28918) );
  sky130_fd_sc_hd__nand4_1 U33509 ( .A(n28918), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[2]), .C(n29745), .D(
        io_oeb[2]), .Y(n28919) );
  sky130_fd_sc_hd__o21ai_1 U33510 ( .A1(n28921), .A2(n28920), .B1(n28919), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N42) );
  sky130_fd_sc_hd__a21oi_1 U33511 ( .A1(n29827), .A2(n28922), .B1(n29061), .Y(
        n28926) );
  sky130_fd_sc_hd__clkinv_1 U33512 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[3]), .Y(n29312) );
  sky130_fd_sc_hd__o22ai_1 U33513 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[3]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]), .B1(n29312), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[3]), .Y(n28923)
         );
  sky130_fd_sc_hd__a21oi_1 U33514 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[3]), .B1(n28923), 
        .Y(n28924) );
  sky130_fd_sc_hd__nand4_1 U33515 ( .A(n28924), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[3]), .C(n29745), .D(
        io_oeb[3]), .Y(n28925) );
  sky130_fd_sc_hd__nor2_1 U33517 ( .A(n29088), .B(n28928), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N7) );
  sky130_fd_sc_hd__a21oi_1 U33518 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[4]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[4]), .B1(n29088), 
        .Y(n28929) );
  sky130_fd_sc_hd__o21ai_1 U33519 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[4]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[4]), .B1(n28929), .Y(
        n28934) );
  sky130_fd_sc_hd__o211ai_1 U33520 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[4]), .A2(n28930), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_ier[4]), .C1(io_oeb[4]), 
        .Y(n28933) );
  sky130_fd_sc_hd__o21ai_1 U33522 ( .A1(n28934), .A2(n28933), .B1(n28932), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N44) );
  sky130_fd_sc_hd__a21oi_1 U33523 ( .A1(n29827), .A2(n28935), .B1(n29061), .Y(
        n28940) );
  sky130_fd_sc_hd__clkinv_1 U33524 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[5]), .Y(n28936) );
  sky130_fd_sc_hd__o22ai_1 U33525 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[5]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]), .B1(n28936), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[5]), .Y(n28937)
         );
  sky130_fd_sc_hd__a21oi_1 U33526 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[5]), .B1(n28937), 
        .Y(n28938) );
  sky130_fd_sc_hd__nand4_1 U33527 ( .A(n28938), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[5]), .C(n29745), .D(
        io_oeb[7]), .Y(n28939) );
  sky130_fd_sc_hd__o21ai_1 U33528 ( .A1(n28941), .A2(n28940), .B1(n28939), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N45) );
  sky130_fd_sc_hd__a21oi_1 U33529 ( .A1(n29745), .A2(n28942), .B1(n29061), .Y(
        n28947) );
  sky130_fd_sc_hd__clkinv_1 U33530 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[6]), .Y(n28943) );
  sky130_fd_sc_hd__o22ai_1 U33531 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[6]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]), .B1(n28943), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[6]), .Y(n28944)
         );
  sky130_fd_sc_hd__a21oi_1 U33532 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[6]), .B1(n28944), 
        .Y(n28945) );
  sky130_fd_sc_hd__nand4_1 U33533 ( .A(n28945), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[6]), .C(n29745), .D(
        io_oeb[26]), .Y(n28946) );
  sky130_fd_sc_hd__o21ai_1 U33534 ( .A1(n28948), .A2(n28947), .B1(n28946), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N46) );
  sky130_fd_sc_hd__a21oi_1 U33535 ( .A1(n29830), .A2(n28949), .B1(n29061), .Y(
        n28954) );
  sky130_fd_sc_hd__clkinv_1 U33536 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[7]), .Y(n28950) );
  sky130_fd_sc_hd__o22ai_1 U33537 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[7]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]), .B1(n28950), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[7]), .Y(n28951)
         );
  sky130_fd_sc_hd__a21oi_1 U33538 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[7]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]), .B1(n28951), 
        .Y(n28952) );
  sky130_fd_sc_hd__nand4_1 U33539 ( .A(n28952), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[7]), .C(n29830), .D(
        io_oeb[27]), .Y(n28953) );
  sky130_fd_sc_hd__o21ai_1 U33540 ( .A1(n28955), .A2(n28954), .B1(n28953), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N47) );
  sky130_fd_sc_hd__nor2_1 U33541 ( .A(n29088), .B(n28956), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N11) );
  sky130_fd_sc_hd__a21oi_1 U33542 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[8]), .B1(
        j202_soc_core_rst), .Y(n28957) );
  sky130_fd_sc_hd__o21ai_1 U33543 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[8]), .B1(n28957), .Y(
        n28962) );
  sky130_fd_sc_hd__o211ai_1 U33544 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[8]), .A2(n28958), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_ier[8]), .C1(io_oeb[28]), 
        .Y(n28961) );
  sky130_fd_sc_hd__o21ai_1 U33546 ( .A1(n28962), .A2(n28961), .B1(n28960), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N48) );
  sky130_fd_sc_hd__a21oi_1 U33547 ( .A1(n29827), .A2(n28963), .B1(n29061), .Y(
        n28968) );
  sky130_fd_sc_hd__o22ai_1 U33548 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[9]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[9]), .B1(n28964), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[9]), .Y(n28965)
         );
  sky130_fd_sc_hd__a21oi_1 U33549 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[9]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[9]), .B1(n28965), 
        .Y(n28966) );
  sky130_fd_sc_hd__nand4_1 U33550 ( .A(n28966), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[9]), .C(n29745), .D(
        io_oeb[29]), .Y(n28967) );
  sky130_fd_sc_hd__o21ai_1 U33551 ( .A1(n28969), .A2(n28968), .B1(n28967), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N49) );
  sky130_fd_sc_hd__a21oi_1 U33552 ( .A1(n29827), .A2(n28970), .B1(n29061), .Y(
        n28975) );
  sky130_fd_sc_hd__o22ai_1 U33553 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[10]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[10]), .B1(n28971), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[10]), .Y(n28972)
         );
  sky130_fd_sc_hd__a21oi_1 U33554 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[10]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[10]), .B1(n28972), 
        .Y(n28973) );
  sky130_fd_sc_hd__nand4_1 U33555 ( .A(n28973), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[10]), .C(n29827), .D(
        io_oeb[30]), .Y(n28974) );
  sky130_fd_sc_hd__o21ai_1 U33556 ( .A1(n28976), .A2(n28975), .B1(n28974), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N50) );
  sky130_fd_sc_hd__a21oi_1 U33557 ( .A1(n29830), .A2(n28977), .B1(n29061), .Y(
        n28982) );
  sky130_fd_sc_hd__o22ai_1 U33558 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[11]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[11]), .B1(n28978), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[11]), .Y(n28979)
         );
  sky130_fd_sc_hd__a21oi_1 U33559 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[11]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[11]), .B1(n28979), 
        .Y(n28980) );
  sky130_fd_sc_hd__nand4_1 U33560 ( .A(n28980), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[11]), .C(n29830), .D(
        io_oeb[31]), .Y(n28981) );
  sky130_fd_sc_hd__a21oi_1 U33564 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[12]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[12]), .B1(n28985), 
        .Y(n28989) );
  sky130_fd_sc_hd__nand3_1 U33566 ( .A(n28989), .B(n28988), .C(io_oeb[32]), 
        .Y(n28990) );
  sky130_fd_sc_hd__nand2_1 U33567 ( .A(n28991), .B(n28990), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N52) );
  sky130_fd_sc_hd__a21oi_1 U33568 ( .A1(n29745), .A2(n28992), .B1(n29061), .Y(
        n28997) );
  sky130_fd_sc_hd__clkinv_1 U33569 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[13]), .Y(n28993) );
  sky130_fd_sc_hd__o22ai_1 U33570 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[13]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13]), .B1(n28993), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[13]), .Y(n28994)
         );
  sky130_fd_sc_hd__a21oi_1 U33571 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[13]), .B1(n28994), 
        .Y(n28995) );
  sky130_fd_sc_hd__nand4_1 U33572 ( .A(n28995), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[13]), .C(n29827), .D(
        io_oeb[33]), .Y(n28996) );
  sky130_fd_sc_hd__o21ai_1 U33573 ( .A1(n28998), .A2(n28997), .B1(n28996), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N53) );
  sky130_fd_sc_hd__a21oi_1 U33574 ( .A1(n29827), .A2(n28999), .B1(n29061), .Y(
        n29004) );
  sky130_fd_sc_hd__clkinv_1 U33575 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[14]), .Y(n29000) );
  sky130_fd_sc_hd__o22ai_1 U33576 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[14]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14]), .B1(n29000), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[14]), .Y(n29001)
         );
  sky130_fd_sc_hd__a21oi_1 U33577 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[14]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14]), .B1(n29001), 
        .Y(n29002) );
  sky130_fd_sc_hd__nand4_1 U33578 ( .A(n29002), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[14]), .C(n29828), .D(
        io_oeb[34]), .Y(n29003) );
  sky130_fd_sc_hd__o21ai_1 U33579 ( .A1(n29005), .A2(n29004), .B1(n29003), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N54) );
  sky130_fd_sc_hd__a21oi_1 U33580 ( .A1(n29745), .A2(n29006), .B1(n29061), .Y(
        n29011) );
  sky130_fd_sc_hd__clkinv_1 U33581 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[15]), .Y(n29007) );
  sky130_fd_sc_hd__o22ai_1 U33582 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[15]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15]), .B1(n29007), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[15]), .Y(n29008)
         );
  sky130_fd_sc_hd__a21oi_1 U33583 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[15]), .B1(n29008), 
        .Y(n29009) );
  sky130_fd_sc_hd__nand4_1 U33584 ( .A(n29009), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[15]), .C(n29745), .D(
        io_oeb[35]), .Y(n29010) );
  sky130_fd_sc_hd__nor2_1 U33586 ( .A(n29088), .B(n29013), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N19) );
  sky130_fd_sc_hd__a21oi_1 U33587 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[16]), .B1(n29088), 
        .Y(n29014) );
  sky130_fd_sc_hd__o21ai_1 U33588 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[16]), .B1(n29014), .Y(
        n29019) );
  sky130_fd_sc_hd__o211ai_1 U33589 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[16]), .A2(n29015), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_ier[16]), .C1(io_oeb[36]), 
        .Y(n29018) );
  sky130_fd_sc_hd__clkinv_1 U33592 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[17]), .Y(n29020) );
  sky130_fd_sc_hd__a21oi_1 U33593 ( .A1(n29020), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[17]), .B1(
        gpio_en_o[17]), .Y(n29021) );
  sky130_fd_sc_hd__nand2_1 U33594 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[17]), .B(n29021), .Y(
        n29022) );
  sky130_fd_sc_hd__a21oi_1 U33595 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[17]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[17]), .B1(n29022), .Y(
        n29027) );
  sky130_fd_sc_hd__o21ai_1 U33596 ( .A1(n29088), .A2(n29024), .B1(n29023), .Y(
        n29026) );
  sky130_fd_sc_hd__o21ai_1 U33597 ( .A1(n29088), .A2(
        j202_soc_core_qspi_wb_wdat[17]), .B1(n29039), .Y(n29025) );
  sky130_fd_sc_hd__a22o_1 U33598 ( .A1(n29027), .A2(n29026), .B1(n29025), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[17]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N57) );
  sky130_fd_sc_hd__a21oi_1 U33599 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[18]), .A2(n12069), 
        .B1(n29604), .Y(n29028) );
  sky130_fd_sc_hd__nor2_1 U33600 ( .A(gpio_en_o[18]), .B(n29028), .Y(n29033)
         );
  sky130_fd_sc_hd__clkinv_1 U33601 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[18]), .Y(n29029) );
  sky130_fd_sc_hd__a21oi_1 U33603 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[18]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[18]), .B1(n29030), 
        .Y(n29032) );
  sky130_fd_sc_hd__a22o_1 U33605 ( .A1(n29033), .A2(n29032), .B1(n29031), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[18]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N58) );
  sky130_fd_sc_hd__a21oi_1 U33606 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[19]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[19]), .B1(gpio_en_o[19]), 
        .Y(n29034) );
  sky130_fd_sc_hd__nand2_1 U33607 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[19]), .B(n29034), .Y(
        n29035) );
  sky130_fd_sc_hd__a21oi_1 U33608 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[19]), .A2(n29036), 
        .B1(n29035), .Y(n29042) );
  sky130_fd_sc_hd__o21ai_1 U33609 ( .A1(n29088), .A2(n29038), .B1(n29037), .Y(
        n29041) );
  sky130_fd_sc_hd__o21ai_1 U33610 ( .A1(j202_soc_core_rst), .A2(
        j202_soc_core_qspi_wb_wdat[19]), .B1(n29039), .Y(n29040) );
  sky130_fd_sc_hd__a22o_1 U33611 ( .A1(n29042), .A2(n29041), .B1(n29040), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[19]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N59) );
  sky130_fd_sc_hd__nor2_1 U33612 ( .A(j202_soc_core_rst), .B(n29043), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N23) );
  sky130_fd_sc_hd__nand2_1 U33613 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[20]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[20]), .Y(n29044) );
  sky130_fd_sc_hd__o211ai_1 U33614 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[20]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[20]), .B1(n29745), 
        .C1(n29044), .Y(n29050) );
  sky130_fd_sc_hd__clkinv_1 U33615 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[20]), .Y(n29046) );
  sky130_fd_sc_hd__clkinv_1 U33616 ( .A(gpio_en_o[20]), .Y(n29045) );
  sky130_fd_sc_hd__o211ai_1 U33617 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[20]), .A2(n29046), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[20]), .C1(n29045), .Y(
        n29049) );
  sky130_fd_sc_hd__o21ai_1 U33618 ( .A1(n29047), .A2(n29061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[20]), .Y(n29048) );
  sky130_fd_sc_hd__o21ai_1 U33619 ( .A1(n29050), .A2(n29049), .B1(n29048), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N60) );
  sky130_fd_sc_hd__a21oi_1 U33620 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[24]), .A2(n12069), 
        .B1(n29605), .Y(n29057) );
  sky130_fd_sc_hd__o2bb2ai_1 U33621 ( .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[24]), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[24]), .A1_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[24]), .A2_N(n29051), .Y(
        n29053) );
  sky130_fd_sc_hd__nand3_1 U33622 ( .A(n29053), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[24]), .C(n29052), .Y(
        n29056) );
  sky130_fd_sc_hd__a21oi_1 U33625 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[28]), .A2(n29745), 
        .B1(n29606), .Y(n29065) );
  sky130_fd_sc_hd__o2bb2ai_1 U33626 ( .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[28]), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[28]), .A1_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[28]), .A2_N(n29058), .Y(
        n29060) );
  sky130_fd_sc_hd__nand3_1 U33627 ( .A(n29060), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[28]), .C(n29059), .Y(
        n29064) );
  sky130_fd_sc_hd__o21ai_1 U33629 ( .A1(n29065), .A2(n29064), .B1(n29063), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N68) );
  sky130_fd_sc_hd__o22ai_1 U33630 ( .A1(n29073), .A2(n29067), .B1(n29066), 
        .B2(n29070), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N9) );
  sky130_fd_sc_hd__o22ai_1 U33631 ( .A1(n29073), .A2(n29069), .B1(n29068), 
        .B2(n29070), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N7) );
  sky130_fd_sc_hd__o22ai_1 U33632 ( .A1(n29073), .A2(n29072), .B1(n29071), 
        .B2(n29070), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N6) );
  sky130_fd_sc_hd__o22ai_1 U33633 ( .A1(n29163), .A2(n29076), .B1(n29075), 
        .B2(n29074), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U33634 ( .A1(n29163), .A2(n29079), .B1(n29078), 
        .B2(n29077), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U33635 ( .A1(n29163), .A2(n29082), .B1(n29081), 
        .B2(n29080), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o21ai_1 U33637 ( .A1(n29087), .A2(n29086), .B1(n29085), .Y(
        j202_soc_core_wbqspiflash_00_N607) );
  sky130_fd_sc_hd__xnor2_1 U33638 ( .A(j202_soc_core_uart_TOP_rxd_s), .B(
        j202_soc_core_uart_TOP_rxd_r), .Y(n29089) );
  sky130_fd_sc_hd__nor2_1 U33639 ( .A(n29088), .B(n29089), .Y(
        j202_soc_core_uart_TOP_N102) );
  sky130_fd_sc_hd__nand3_1 U33640 ( .A(n29089), .B(n29827), .C(n29095), .Y(
        j202_soc_core_uart_TOP_N101) );
  sky130_fd_sc_hd__nand2_1 U33641 ( .A(n29607), .B(
        j202_soc_core_uart_TOP_change), .Y(n29091) );
  sky130_fd_sc_hd__nor2_1 U33642 ( .A(j202_soc_core_uart_TOP_change), .B(
        j202_soc_core_uart_TOP_dpll_state[0]), .Y(n29093) );
  sky130_fd_sc_hd__nand2_1 U33643 ( .A(n29093), .B(
        j202_soc_core_uart_sio_ce_x4), .Y(n29090) );
  sky130_fd_sc_hd__o211ai_1 U33644 ( .A1(j202_soc_core_uart_sio_ce_x4), .A2(
        n29092), .B1(n29091), .C1(n29090), .Y(n27) );
  sky130_fd_sc_hd__nor2_1 U33647 ( .A(j202_soc_core_uart_TOP_shift_en), .B(
        j202_soc_core_uart_TOP_shift_en_r), .Y(n29097) );
  sky130_fd_sc_hd__nor2_1 U33648 ( .A(j202_soc_core_uart_TOP_hold_reg[0]), .B(
        n29097), .Y(n29098) );
  sky130_fd_sc_hd__xnor2_1 U33650 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[8]), .Y(n29103) );
  sky130_fd_sc_hd__xnor2_1 U33651 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[1]), .Y(n29102) );
  sky130_fd_sc_hd__xnor2_1 U33652 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[0]), .Y(n29101) );
  sky130_fd_sc_hd__xnor2_1 U33653 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[2]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[2]), .Y(n29100) );
  sky130_fd_sc_hd__nand4_1 U33654 ( .A(n29103), .B(n29102), .C(n29101), .D(
        n29100), .Y(n29114) );
  sky130_fd_sc_hd__xnor2_1 U33655 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[7]), .Y(n29107) );
  sky130_fd_sc_hd__xnor2_1 U33656 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[11]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[11]), .Y(n29106) );
  sky130_fd_sc_hd__xnor2_1 U33657 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[9]), .Y(n29105) );
  sky130_fd_sc_hd__xnor2_1 U33658 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[6]), .Y(n29104) );
  sky130_fd_sc_hd__nand4_1 U33659 ( .A(n29107), .B(n29106), .C(n29105), .D(
        n29104), .Y(n29113) );
  sky130_fd_sc_hd__xnor2_1 U33660 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[4]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[4]), .Y(n29111) );
  sky130_fd_sc_hd__xnor2_1 U33661 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[3]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[3]), .Y(n29110) );
  sky130_fd_sc_hd__xnor2_1 U33662 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[10]), .Y(n29109) );
  sky130_fd_sc_hd__xnor2_1 U33663 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[5]), .Y(n29108) );
  sky130_fd_sc_hd__nand4_1 U33664 ( .A(n29111), .B(n29110), .C(n29109), .D(
        n29108), .Y(n29112) );
  sky130_fd_sc_hd__nor3_1 U33665 ( .A(n29114), .B(n29113), .C(n29112), .Y(
        n29118) );
  sky130_fd_sc_hd__nand2_1 U33666 ( .A(n29115), .B(
        j202_soc_core_bldc_core_00_pwm_en), .Y(n29116) );
  sky130_fd_sc_hd__o22ai_1 U33667 ( .A1(n29118), .A2(n29117), .B1(n29116), 
        .B2(io_in[25]), .Y(n31) );
  sky130_fd_sc_hd__nand4_1 U33668 ( .A(n29119), .B(n29121), .C(
        j202_soc_core_bldc_core_00_comm[0]), .D(
        j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld), .Y(n29123) );
  sky130_fd_sc_hd__o21ai_1 U33669 ( .A1(j202_soc_core_bldc_core_00_comm[0]), 
        .A2(n29120), .B1(n29123), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posa) );
  sky130_fd_sc_hd__nand3_1 U33670 ( .A(n29121), .B(
        j202_soc_core_bldc_core_00_comm[2]), .C(
        j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld), .Y(n29125) );
  sky130_fd_sc_hd__nand2_1 U33671 ( .A(n29608), .B(
        j202_soc_core_bldc_core_00_comm[0]), .Y(n29122) );
  sky130_fd_sc_hd__o21ai_1 U33672 ( .A1(j202_soc_core_bldc_core_00_comm[0]), 
        .A2(n29125), .B1(n29122), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posb) );
  sky130_fd_sc_hd__nand4_1 U33673 ( .A(n29126), .B(
        j202_soc_core_bldc_core_00_comm[1]), .C(
        j202_soc_core_bldc_core_00_comm[2]), .D(
        j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld), .Y(n29124) );
  sky130_fd_sc_hd__nand2_1 U33674 ( .A(n29123), .B(n29124), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_negb) );
  sky130_fd_sc_hd__o21ai_1 U33675 ( .A1(n29126), .A2(n29125), .B1(n29124), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posc) );
  sky130_fd_sc_hd__a21o_1 U33676 ( .A1(n29262), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[28]), .B1(n29266), .X(
        n29128) );
  sky130_fd_sc_hd__nand2_1 U33677 ( .A(j202_soc_core_wbqspiflash_00_spi_in[31]), .B(n29267), .Y(n29272) );
  sky130_fd_sc_hd__o22ai_1 U33678 ( .A1(j202_soc_core_wbqspiflash_00_spi_spd), 
        .A2(n29272), .B1(n29196), .B2(n29256), .Y(n29127) );
  sky130_fd_sc_hd__a211o_1 U33679 ( .A1(n29265), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[31]), .B1(n29128), .C1(
        n29127), .X(j202_soc_core_wbqspiflash_00_lldriver_N316) );
  sky130_fd_sc_hd__a22oi_1 U33680 ( .A1(n29265), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[30]), .B1(n29262), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[27]), .Y(n29129) );
  sky130_fd_sc_hd__a21oi_1 U33682 ( .A1(n29264), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[30]), .B1(n29131), .Y(n29132) );
  sky130_fd_sc_hd__a22oi_1 U33684 ( .A1(n29265), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[27]), .B1(n29262), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[24]), .Y(n29134) );
  sky130_fd_sc_hd__o21ai_1 U33685 ( .A1(n29196), .A2(n29135), .B1(n29134), .Y(
        n29136) );
  sky130_fd_sc_hd__a21oi_1 U33686 ( .A1(n29264), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[27]), .B1(n29136), .Y(n29137) );
  sky130_fd_sc_hd__a22oi_1 U33688 ( .A1(n29265), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[3]), .B1(n29262), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[0]), .Y(n29138) );
  sky130_fd_sc_hd__a21oi_1 U33690 ( .A1(n29264), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[3]), .B1(n29140), .Y(n29141) );
  sky130_fd_sc_hd__a222oi_1 U33692 ( .A1(n29265), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[2]), .B1(n29264), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[2]), .C1(n29257), .C2(
        j202_soc_core_wbqspiflash_00_spi_in[3]), .Y(n29142) );
  sky130_fd_sc_hd__nand2_1 U33693 ( .A(n29143), .B(
        j202_soc_core_intc_core_00_bs_addr[7]), .Y(n29164) );
  sky130_fd_sc_hd__nor2_1 U33694 ( .A(n29144), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N17) );
  sky130_fd_sc_hd__nor2_1 U33695 ( .A(n29145), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N16) );
  sky130_fd_sc_hd__nor2_1 U33696 ( .A(n29146), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N11) );
  sky130_fd_sc_hd__nor2_1 U33697 ( .A(n29147), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N15) );
  sky130_fd_sc_hd__nor2_1 U33698 ( .A(n29148), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N12) );
  sky130_fd_sc_hd__nor2_1 U33699 ( .A(n29149), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N20) );
  sky130_fd_sc_hd__nor2_1 U33700 ( .A(n29150), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N22) );
  sky130_fd_sc_hd__nor2_1 U33701 ( .A(n29151), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N19) );
  sky130_fd_sc_hd__nor2_1 U33702 ( .A(n29152), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N23) );
  sky130_fd_sc_hd__nor2_1 U33703 ( .A(n29153), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N21) );
  sky130_fd_sc_hd__nor2_1 U33704 ( .A(n29154), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N18) );
  sky130_fd_sc_hd__nor2_1 U33705 ( .A(n29155), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N14) );
  sky130_fd_sc_hd__nor2_1 U33706 ( .A(n29156), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N13) );
  sky130_fd_sc_hd__nor2_1 U33707 ( .A(n29157), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N10) );
  sky130_fd_sc_hd__nor2_1 U33708 ( .A(n29158), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N9) );
  sky130_fd_sc_hd__nor2_1 U33709 ( .A(n29159), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N8) );
  sky130_fd_sc_hd__nor2_1 U33710 ( .A(n29160), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N7) );
  sky130_fd_sc_hd__nor2_1 U33711 ( .A(n29161), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N6) );
  sky130_fd_sc_hd__nor2_1 U33712 ( .A(n29162), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N5) );
  sky130_fd_sc_hd__nor2_1 U33713 ( .A(n29163), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N4) );
  sky130_fd_sc_hd__nor2_1 U33714 ( .A(n29165), .B(n29164), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand3_1 U33715 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B(n29167), .C(n29166), 
        .Y(j202_soc_core_wbqspiflash_00_lldriver_N354) );
  sky130_fd_sc_hd__or3_1 U33716 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[0]), .C(n28896), .X(io_oeb[11]) );
  sky130_fd_sc_hd__nor2_1 U33717 ( .A(n29169), .B(n29168), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt0_to1) );
  sky130_fd_sc_hd__nor2_1 U33718 ( .A(n29171), .B(n29170), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt1_to1) );
  sky130_fd_sc_hd__nor2b_1 U33719 ( .B_N(j202_soc_core_uart_TOP_rx_sio_ce_r1), 
        .A(j202_soc_core_uart_TOP_rx_sio_ce_r2), .Y(
        j202_soc_core_uart_TOP_N118) );
  sky130_fd_sc_hd__nor2_1 U33720 ( .A(j202_soc_core_uart_TOP_shift_en), .B(
        j202_soc_core_uart_TOP_txf_empty_r), .Y(j202_soc_core_uart_TOP_N137)
         );
  sky130_fd_sc_hd__nand3_1 U33721 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[1]), 
        .B(n29173), .C(n29172), .Y(j202_soc_core_uart_TOP_N128) );
  sky130_fd_sc_hd__nor2b_1 U33722 ( .B_N(n29609), .A(
        j202_soc_core_uart_BRG_sio_ce_r), .Y(j202_soc_core_uart_BRG_N59) );
  sky130_fd_sc_hd__o21ai_1 U33723 ( .A1(j202_soc_core_uart_BRG_ps[7]), .A2(
        n29176), .B1(n29174), .Y(n29175) );
  sky130_fd_sc_hd__a21oi_1 U33724 ( .A1(j202_soc_core_uart_BRG_ps[7]), .A2(
        n29176), .B1(n29175), .Y(j202_soc_core_uart_BRG_N19) );
  sky130_fd_sc_hd__a21oi_1 U33726 ( .A1(j202_soc_core_uart_BRG_br_cnt[7]), 
        .A2(n29180), .B1(n29179), .Y(j202_soc_core_uart_BRG_N42) );
  sky130_fd_sc_hd__a31oi_1 U33727 ( .A1(n29610), .A2(wbs_we_i), .A3(
        wbs_sel_i[0]), .B1(wb_rst_i), .Y(n29181) );
  sky130_fd_sc_hd__nand2_1 U33728 ( .A(start_n_reg[1]), .B(n29181), .Y(n10) );
  sky130_fd_sc_hd__nand2_1 U33729 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .B(
        j202_soc_core_wbqspiflash_00_alt_ctrl), .Y(n29182) );
  sky130_fd_sc_hd__o21ai_0 U33730 ( .A1(n29183), .A2(
        j202_soc_core_wbqspiflash_00_spif_override), .B1(n29182), .Y(io_out[9]) );
  sky130_fd_sc_hd__a22o_1 U33731 ( .A1(n29184), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_dir), .B1(n29263), .B2(
        j202_soc_core_wbqspiflash_00_spi_dir), .X(
        j202_soc_core_wbqspiflash_00_lldriver_N355) );
  sky130_fd_sc_hd__a22oi_1 U33732 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[4]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[1]), .B2(n29262), .Y(
        n29186) );
  sky130_fd_sc_hd__a22oi_1 U33733 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[1]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[5]), .Y(n29185) );
  sky130_fd_sc_hd__o211ai_1 U33734 ( .A1(n29261), .A2(n29195), .B1(n29186), 
        .C1(n29185), .Y(j202_soc_core_wbqspiflash_00_lldriver_N396) );
  sky130_fd_sc_hd__a22oi_1 U33735 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[5]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[2]), .B2(n29262), .Y(
        n29189) );
  sky130_fd_sc_hd__a22oi_1 U33736 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[2]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[6]), .Y(n29188) );
  sky130_fd_sc_hd__nand2_1 U33737 ( .A(j202_soc_core_wbqspiflash_00_spi_in[5]), 
        .B(n29264), .Y(n29187) );
  sky130_fd_sc_hd__nand3_1 U33738 ( .A(n29189), .B(n29188), .C(n29187), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N397) );
  sky130_fd_sc_hd__a22oi_1 U33739 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[6]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[3]), .B2(n29262), .Y(
        n29192) );
  sky130_fd_sc_hd__a22oi_1 U33740 ( .A1(n29264), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[6]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[7]), .Y(n29191) );
  sky130_fd_sc_hd__nand2_1 U33741 ( .A(n29263), .B(
        j202_soc_core_wbqspiflash_00_spi_in[3]), .Y(n29190) );
  sky130_fd_sc_hd__nand3_1 U33742 ( .A(n29192), .B(n29191), .C(n29190), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N398) );
  sky130_fd_sc_hd__a22oi_1 U33743 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[7]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[4]), .B2(n29262), .Y(
        n29194) );
  sky130_fd_sc_hd__a22oi_1 U33744 ( .A1(n29264), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[7]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[8]), .Y(n29193) );
  sky130_fd_sc_hd__o211ai_1 U33745 ( .A1(n29196), .A2(n29195), .B1(n29194), 
        .C1(n29193), .Y(j202_soc_core_wbqspiflash_00_lldriver_N399) );
  sky130_fd_sc_hd__a22oi_1 U33746 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[8]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[5]), .B2(n29262), .Y(
        n29199) );
  sky130_fd_sc_hd__a22oi_1 U33747 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[5]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[9]), .Y(n29198) );
  sky130_fd_sc_hd__nand2_1 U33748 ( .A(j202_soc_core_wbqspiflash_00_spi_in[8]), 
        .B(n29264), .Y(n29197) );
  sky130_fd_sc_hd__nand3_1 U33749 ( .A(n29199), .B(n29198), .C(n29197), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N400) );
  sky130_fd_sc_hd__a22oi_1 U33750 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[9]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[6]), .B2(n29262), .Y(
        n29202) );
  sky130_fd_sc_hd__a22oi_1 U33751 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[6]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[10]), .Y(n29201) );
  sky130_fd_sc_hd__nand2_1 U33752 ( .A(j202_soc_core_wbqspiflash_00_spi_in[9]), 
        .B(n29264), .Y(n29200) );
  sky130_fd_sc_hd__nand3_1 U33753 ( .A(n29202), .B(n29201), .C(n29200), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N401) );
  sky130_fd_sc_hd__a22oi_1 U33754 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[10]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[7]), .B2(n29262), .Y(
        n29205) );
  sky130_fd_sc_hd__a22oi_1 U33755 ( .A1(n29264), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[10]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[11]), .Y(n29204) );
  sky130_fd_sc_hd__nand2_1 U33756 ( .A(n29263), .B(
        j202_soc_core_wbqspiflash_00_spi_in[7]), .Y(n29203) );
  sky130_fd_sc_hd__nand3_1 U33757 ( .A(n29205), .B(n29204), .C(n29203), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N402) );
  sky130_fd_sc_hd__a22oi_1 U33758 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[11]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[8]), .B2(n29262), .Y(
        n29208) );
  sky130_fd_sc_hd__a22oi_1 U33759 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[8]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[11]), .B2(n29264), .Y(n29207) );
  sky130_fd_sc_hd__nand2_1 U33760 ( .A(n29257), .B(
        j202_soc_core_wbqspiflash_00_spi_in[12]), .Y(n29206) );
  sky130_fd_sc_hd__nand3_1 U33761 ( .A(n29208), .B(n29207), .C(n29206), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N403) );
  sky130_fd_sc_hd__a22oi_1 U33762 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[12]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[9]), .B2(n29262), .Y(
        n29211) );
  sky130_fd_sc_hd__a22oi_1 U33763 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[9]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[12]), .B2(n29264), .Y(n29210) );
  sky130_fd_sc_hd__nand2_1 U33764 ( .A(n29257), .B(
        j202_soc_core_wbqspiflash_00_spi_in[13]), .Y(n29209) );
  sky130_fd_sc_hd__nand3_1 U33765 ( .A(n29211), .B(n29210), .C(n29209), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N404) );
  sky130_fd_sc_hd__a22oi_1 U33766 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[13]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[10]), .B2(n29262), .Y(
        n29214) );
  sky130_fd_sc_hd__a22oi_1 U33767 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[10]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[14]), .Y(n29213) );
  sky130_fd_sc_hd__nand2_1 U33768 ( .A(j202_soc_core_wbqspiflash_00_spi_in[13]), .B(n29264), .Y(n29212) );
  sky130_fd_sc_hd__nand3_1 U33769 ( .A(n29214), .B(n29213), .C(n29212), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N405) );
  sky130_fd_sc_hd__a22oi_1 U33770 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[14]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[11]), .B2(n29262), .Y(
        n29217) );
  sky130_fd_sc_hd__a22oi_1 U33771 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[11]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[14]), .B2(n29264), .Y(n29216) );
  sky130_fd_sc_hd__nand2_1 U33772 ( .A(n29257), .B(
        j202_soc_core_wbqspiflash_00_spi_in[15]), .Y(n29215) );
  sky130_fd_sc_hd__nand3_1 U33773 ( .A(n29217), .B(n29216), .C(n29215), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N406) );
  sky130_fd_sc_hd__a22oi_1 U33774 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[15]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[12]), .B2(n29262), .Y(
        n29220) );
  sky130_fd_sc_hd__a22oi_1 U33775 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[12]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[15]), .B2(n29264), .Y(n29219) );
  sky130_fd_sc_hd__nand2_1 U33776 ( .A(n29257), .B(
        j202_soc_core_wbqspiflash_00_spi_in[16]), .Y(n29218) );
  sky130_fd_sc_hd__nand3_1 U33777 ( .A(n29220), .B(n29219), .C(n29218), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N407) );
  sky130_fd_sc_hd__a22oi_1 U33778 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[16]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[13]), .B2(n29262), .Y(
        n29223) );
  sky130_fd_sc_hd__a22oi_1 U33779 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[13]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[17]), .Y(n29222) );
  sky130_fd_sc_hd__nand2_1 U33780 ( .A(j202_soc_core_wbqspiflash_00_spi_in[16]), .B(n29264), .Y(n29221) );
  sky130_fd_sc_hd__nand3_1 U33781 ( .A(n29223), .B(n29222), .C(n29221), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N408) );
  sky130_fd_sc_hd__a22oi_1 U33782 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[17]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[14]), .B2(n29262), .Y(
        n29226) );
  sky130_fd_sc_hd__a22oi_1 U33783 ( .A1(n29264), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[17]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[18]), .Y(n29225) );
  sky130_fd_sc_hd__nand2_1 U33784 ( .A(n29263), .B(
        j202_soc_core_wbqspiflash_00_spi_in[14]), .Y(n29224) );
  sky130_fd_sc_hd__nand3_1 U33785 ( .A(n29226), .B(n29225), .C(n29224), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N409) );
  sky130_fd_sc_hd__a22oi_1 U33786 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[18]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[15]), .B2(n29262), .Y(
        n29229) );
  sky130_fd_sc_hd__a22oi_1 U33787 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[15]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[19]), .Y(n29228) );
  sky130_fd_sc_hd__nand2_1 U33788 ( .A(j202_soc_core_wbqspiflash_00_spi_in[18]), .B(n29264), .Y(n29227) );
  sky130_fd_sc_hd__nand3_1 U33789 ( .A(n29229), .B(n29228), .C(n29227), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N410) );
  sky130_fd_sc_hd__a22oi_1 U33790 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[19]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[16]), .B2(n29262), .Y(
        n29232) );
  sky130_fd_sc_hd__a22oi_1 U33791 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[16]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[19]), .B2(n29264), .Y(n29231) );
  sky130_fd_sc_hd__nand2_1 U33792 ( .A(n29257), .B(
        j202_soc_core_wbqspiflash_00_spi_in[20]), .Y(n29230) );
  sky130_fd_sc_hd__nand3_1 U33793 ( .A(n29232), .B(n29231), .C(n29230), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N411) );
  sky130_fd_sc_hd__a22oi_1 U33794 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[20]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[17]), .B2(n29262), .Y(
        n29235) );
  sky130_fd_sc_hd__a22oi_1 U33795 ( .A1(n29264), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[20]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[21]), .Y(n29234) );
  sky130_fd_sc_hd__nand2_1 U33796 ( .A(n29263), .B(
        j202_soc_core_wbqspiflash_00_spi_in[17]), .Y(n29233) );
  sky130_fd_sc_hd__nand3_1 U33797 ( .A(n29235), .B(n29234), .C(n29233), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N412) );
  sky130_fd_sc_hd__a22oi_1 U33798 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[21]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[18]), .B2(n29262), .Y(
        n29238) );
  sky130_fd_sc_hd__a22oi_1 U33799 ( .A1(n29264), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[21]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[22]), .Y(n29237) );
  sky130_fd_sc_hd__nand2_1 U33800 ( .A(n29263), .B(
        j202_soc_core_wbqspiflash_00_spi_in[18]), .Y(n29236) );
  sky130_fd_sc_hd__nand3_1 U33801 ( .A(n29238), .B(n29237), .C(n29236), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N413) );
  sky130_fd_sc_hd__a22oi_1 U33802 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[22]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[19]), .B2(n29262), .Y(
        n29241) );
  sky130_fd_sc_hd__a22oi_1 U33803 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[19]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[22]), .B2(n29264), .Y(n29240) );
  sky130_fd_sc_hd__nand2_1 U33804 ( .A(n29257), .B(
        j202_soc_core_wbqspiflash_00_spi_in[23]), .Y(n29239) );
  sky130_fd_sc_hd__nand3_1 U33805 ( .A(n29241), .B(n29240), .C(n29239), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N414) );
  sky130_fd_sc_hd__a22oi_1 U33806 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[23]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[20]), .B2(n29262), .Y(
        n29244) );
  sky130_fd_sc_hd__a22oi_1 U33807 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[20]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[23]), .B2(n29264), .Y(n29243) );
  sky130_fd_sc_hd__nand2_1 U33808 ( .A(n29257), .B(
        j202_soc_core_wbqspiflash_00_spi_in[24]), .Y(n29242) );
  sky130_fd_sc_hd__nand3_1 U33809 ( .A(n29244), .B(n29243), .C(n29242), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N415) );
  sky130_fd_sc_hd__a22oi_1 U33810 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[24]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[21]), .B2(n29262), .Y(
        n29247) );
  sky130_fd_sc_hd__a22oi_1 U33811 ( .A1(n29264), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[24]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[25]), .Y(n29246) );
  sky130_fd_sc_hd__nand2_1 U33812 ( .A(n29263), .B(
        j202_soc_core_wbqspiflash_00_spi_in[21]), .Y(n29245) );
  sky130_fd_sc_hd__nand3_1 U33813 ( .A(n29247), .B(n29246), .C(n29245), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N416) );
  sky130_fd_sc_hd__a22oi_1 U33814 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[25]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[22]), .B2(n29262), .Y(
        n29250) );
  sky130_fd_sc_hd__a22oi_1 U33815 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[22]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[26]), .Y(n29249) );
  sky130_fd_sc_hd__nand2_1 U33816 ( .A(j202_soc_core_wbqspiflash_00_spi_in[25]), .B(n29264), .Y(n29248) );
  sky130_fd_sc_hd__nand3_1 U33817 ( .A(n29250), .B(n29249), .C(n29248), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N417) );
  sky130_fd_sc_hd__a22oi_1 U33818 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[26]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[23]), .B2(n29262), .Y(
        n29253) );
  sky130_fd_sc_hd__a22oi_1 U33819 ( .A1(n29264), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[26]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[27]), .Y(n29252) );
  sky130_fd_sc_hd__nand2_1 U33820 ( .A(n29263), .B(
        j202_soc_core_wbqspiflash_00_spi_in[23]), .Y(n29251) );
  sky130_fd_sc_hd__nand3_1 U33821 ( .A(n29253), .B(n29252), .C(n29251), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N418) );
  sky130_fd_sc_hd__a22oi_1 U33822 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[28]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[25]), .B2(n29262), .Y(
        n29255) );
  sky130_fd_sc_hd__a22oi_1 U33823 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[25]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[29]), .Y(n29254) );
  sky130_fd_sc_hd__o211ai_1 U33824 ( .A1(n29261), .A2(n29256), .B1(n29255), 
        .C1(n29254), .Y(j202_soc_core_wbqspiflash_00_lldriver_N420) );
  sky130_fd_sc_hd__a22oi_1 U33825 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[29]), .A2(n29265), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[26]), .B2(n29262), .Y(
        n29259) );
  sky130_fd_sc_hd__a22oi_1 U33826 ( .A1(n29263), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[26]), .B1(n29257), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[30]), .Y(n29258) );
  sky130_fd_sc_hd__o211ai_1 U33827 ( .A1(n29261), .A2(n29260), .B1(n29259), 
        .C1(n29258), .Y(j202_soc_core_wbqspiflash_00_lldriver_N421) );
  sky130_fd_sc_hd__a22o_1 U33828 ( .A1(j202_soc_core_wbqspiflash_00_spi_in[29]), .A2(n29263), .B1(n29262), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[29]), .X(
        j202_soc_core_wbqspiflash_00_lldriver_N317) );
  sky130_fd_sc_hd__or3_1 U33829 ( .A(n29266), .B(n29265), .C(n29264), .X(
        n29273) );
  sky130_fd_sc_hd__a21oi_1 U33830 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[30]), .A2(n29270), .B1(
        n29273), .Y(n29269) );
  sky130_fd_sc_hd__nand2_1 U33831 ( .A(j202_soc_core_wbqspiflash_00_spi_in[30]), .B(n29267), .Y(n29268) );
  sky130_fd_sc_hd__nand2_1 U33832 ( .A(n29269), .B(n29268), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N318) );
  sky130_fd_sc_hd__nand2_1 U33833 ( .A(n29270), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[31]), .Y(n29271) );
  sky130_fd_sc_hd__nand3b_1 U33834 ( .A_N(n29273), .B(n29272), .C(n29271), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N319) );
  sky130_fd_sc_hd__a21oi_1 U33835 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[0]), .A2(
        j202_soc_core_wbqspiflash_00_reset_counter[1]), .B1(n29274), .Y(n29275) );
  sky130_fd_sc_hd__nor2_1 U33836 ( .A(n29276), .B(n29275), .Y(
        j202_soc_core_wbqspiflash_00_N615) );
  sky130_fd_sc_hd__nor2_1 U33837 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[0]), 
        .B(j202_soc_core_uart_TOP_tx_fifo_rp[1]), .Y(n29305) );
  sky130_fd_sc_hd__a22oi_1 U33838 ( .A1(n29305), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[24]), .B1(n29302), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[0]), .Y(n29280) );
  sky130_fd_sc_hd__nor2_1 U33839 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[0]), 
        .B(n29277), .Y(n29304) );
  sky130_fd_sc_hd__nor2_1 U33840 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[1]), 
        .B(n29278), .Y(n29303) );
  sky130_fd_sc_hd__a22oi_1 U33841 ( .A1(n29304), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[8]), .B1(n29303), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[16]), .Y(n29279) );
  sky130_fd_sc_hd__a21oi_1 U33842 ( .A1(n29280), .A2(n29279), .B1(n29301), .Y(
        n29281) );
  sky130_fd_sc_hd__a21o_1 U33843 ( .A1(j202_soc_core_uart_TOP_hold_reg[2]), 
        .A2(n29300), .B1(n29281), .X(j202_soc_core_uart_TOP_N26) );
  sky130_fd_sc_hd__a22oi_1 U33844 ( .A1(n29303), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[17]), .B1(n29302), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[1]), .Y(n29283) );
  sky130_fd_sc_hd__a22oi_1 U33845 ( .A1(n29304), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[9]), .B1(n29305), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[25]), .Y(n29282) );
  sky130_fd_sc_hd__a21oi_1 U33846 ( .A1(n29283), .A2(n29282), .B1(n29301), .Y(
        n29284) );
  sky130_fd_sc_hd__a21o_1 U33847 ( .A1(j202_soc_core_uart_TOP_hold_reg[3]), 
        .A2(n29300), .B1(n29284), .X(j202_soc_core_uart_TOP_N27) );
  sky130_fd_sc_hd__a22oi_1 U33848 ( .A1(n29304), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[10]), .B1(n29305), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[26]), .Y(n29286) );
  sky130_fd_sc_hd__a22oi_1 U33849 ( .A1(n29303), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[18]), .B1(n29302), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[2]), .Y(n29285) );
  sky130_fd_sc_hd__a21oi_1 U33850 ( .A1(n29286), .A2(n29285), .B1(n29301), .Y(
        n29287) );
  sky130_fd_sc_hd__a21o_1 U33851 ( .A1(j202_soc_core_uart_TOP_hold_reg[4]), 
        .A2(n29300), .B1(n29287), .X(j202_soc_core_uart_TOP_N28) );
  sky130_fd_sc_hd__a22oi_1 U33852 ( .A1(n29303), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[19]), .B1(n29305), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[27]), .Y(n29289) );
  sky130_fd_sc_hd__a22oi_1 U33853 ( .A1(n29304), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[11]), .B1(n29302), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[3]), .Y(n29288) );
  sky130_fd_sc_hd__a21oi_1 U33854 ( .A1(n29289), .A2(n29288), .B1(n29301), .Y(
        n29290) );
  sky130_fd_sc_hd__a21o_1 U33855 ( .A1(j202_soc_core_uart_TOP_hold_reg[5]), 
        .A2(n29300), .B1(n29290), .X(j202_soc_core_uart_TOP_N29) );
  sky130_fd_sc_hd__a22oi_1 U33856 ( .A1(n29303), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[20]), .B1(n29305), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[28]), .Y(n29292) );
  sky130_fd_sc_hd__a22oi_1 U33857 ( .A1(n29304), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[12]), .B1(n29302), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[4]), .Y(n29291) );
  sky130_fd_sc_hd__a21oi_1 U33858 ( .A1(n29292), .A2(n29291), .B1(n29301), .Y(
        n29293) );
  sky130_fd_sc_hd__a21o_1 U33859 ( .A1(j202_soc_core_uart_TOP_hold_reg[6]), 
        .A2(n29300), .B1(n29293), .X(j202_soc_core_uart_TOP_N30) );
  sky130_fd_sc_hd__a22oi_1 U33860 ( .A1(n29304), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[13]), .B1(n29302), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[5]), .Y(n29295) );
  sky130_fd_sc_hd__a22oi_1 U33861 ( .A1(n29303), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[21]), .B1(n29305), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[29]), .Y(n29294) );
  sky130_fd_sc_hd__a21oi_1 U33862 ( .A1(n29295), .A2(n29294), .B1(n29301), .Y(
        n29296) );
  sky130_fd_sc_hd__a21o_1 U33863 ( .A1(j202_soc_core_uart_TOP_hold_reg[7]), 
        .A2(n29300), .B1(n29296), .X(j202_soc_core_uart_TOP_N31) );
  sky130_fd_sc_hd__a22oi_1 U33864 ( .A1(n29304), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[14]), .B1(n29302), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[6]), .Y(n29298) );
  sky130_fd_sc_hd__a22oi_1 U33865 ( .A1(n29303), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[22]), .B1(n29305), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[30]), .Y(n29297) );
  sky130_fd_sc_hd__a21oi_1 U33866 ( .A1(n29298), .A2(n29297), .B1(n29301), .Y(
        n29299) );
  sky130_fd_sc_hd__a21o_1 U33867 ( .A1(j202_soc_core_uart_TOP_hold_reg[8]), 
        .A2(n29300), .B1(n29299), .X(j202_soc_core_uart_TOP_N32) );
  sky130_fd_sc_hd__a21oi_1 U33868 ( .A1(n29302), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[7]), .B1(n29301), .Y(n29309) );
  sky130_fd_sc_hd__a22oi_1 U33869 ( .A1(n29304), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[15]), .B1(n29303), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[23]), .Y(n29308) );
  sky130_fd_sc_hd__nand2_1 U33870 ( .A(n29305), .B(
        j202_soc_core_uart_TOP_tx_fifo_mem[31]), .Y(n29307) );
  sky130_fd_sc_hd__a31oi_1 U33871 ( .A1(n29309), .A2(n29308), .A3(n29307), 
        .B1(n29306), .Y(j202_soc_core_uart_TOP_N33) );
  sky130_fd_sc_hd__a22oi_1 U33872 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]), .A2(n29394), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_ier[3]), .B2(n29391), .Y(
        n29316) );
  sky130_fd_sc_hd__o22ai_1 U33873 ( .A1(n29312), .A2(n29311), .B1(io_oeb[3]), 
        .B2(n29310), .Y(n29313) );
  sky130_fd_sc_hd__a21oi_1 U33874 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[3]), .A2(n29390), .B1(
        n29313), .Y(n29315) );
  sky130_fd_sc_hd__nand2_1 U33875 ( .A(n29389), .B(la_data_out[3]), .Y(n29314)
         );
  sky130_fd_sc_hd__nand3_1 U33876 ( .A(n29316), .B(n29315), .C(n29314), .Y(
        j202_soc_core_ahb2apb_02_N131) );
  sky130_fd_sc_hd__a22oi_1 U33877 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[4]), .A2(n29394), 
        .B1(n29389), .B2(la_data_out[4]), .Y(n29319) );
  sky130_fd_sc_hd__a22oi_1 U33878 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[4]), .A2(n29392), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[4]), .B2(n29391), .Y(
        n29318) );
  sky130_fd_sc_hd__a22oi_1 U33879 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[4]), .A2(n29390), .B1(
        gpio_en_o[4]), .B2(n29393), .Y(n29317) );
  sky130_fd_sc_hd__nand3_1 U33880 ( .A(n29319), .B(n29318), .C(n29317), .Y(
        j202_soc_core_ahb2apb_02_N132) );
  sky130_fd_sc_hd__a22oi_1 U33881 ( .A1(gpio_en_o[5]), .A2(n29393), .B1(n29389), .B2(la_data_out[5]), .Y(n29322) );
  sky130_fd_sc_hd__a22oi_1 U33882 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[5]), .A2(n29392), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[5]), .B2(n29391), .Y(
        n29321) );
  sky130_fd_sc_hd__a22oi_1 U33883 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[5]), .A2(n29390), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]), .B2(n29394), 
        .Y(n29320) );
  sky130_fd_sc_hd__nand3_1 U33884 ( .A(n29322), .B(n29321), .C(n29320), .Y(
        j202_soc_core_ahb2apb_02_N133) );
  sky130_fd_sc_hd__a22oi_1 U33885 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[6]), .A2(n29390), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[6]), .B2(n29392), .Y(
        n29325) );
  sky130_fd_sc_hd__a22oi_1 U33886 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]), .A2(n29394), 
        .B1(gpio_en_o[6]), .B2(n29393), .Y(n29324) );
  sky130_fd_sc_hd__a22oi_1 U33887 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[6]), .A2(n29391), .B1(
        n29389), .B2(la_data_out[6]), .Y(n29323) );
  sky130_fd_sc_hd__nand3_1 U33888 ( .A(n29325), .B(n29324), .C(n29323), .Y(
        j202_soc_core_ahb2apb_02_N134) );
  sky130_fd_sc_hd__a22oi_1 U33889 ( .A1(gpio_en_o[7]), .A2(n29393), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[7]), .B2(n29391), .Y(
        n29328) );
  sky130_fd_sc_hd__a22oi_1 U33890 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[7]), .A2(n29390), .B1(
        n29389), .B2(la_data_out[7]), .Y(n29327) );
  sky130_fd_sc_hd__a22oi_1 U33891 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[7]), .A2(n29392), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]), .B2(n29394), 
        .Y(n29326) );
  sky130_fd_sc_hd__nand3_1 U33892 ( .A(n29328), .B(n29327), .C(n29326), .Y(
        j202_soc_core_ahb2apb_02_N135) );
  sky130_fd_sc_hd__a22oi_1 U33893 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[8]), .A2(n29392), .B1(
        gpio_en_o[8]), .B2(n29393), .Y(n29331) );
  sky130_fd_sc_hd__a22oi_1 U33894 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]), .A2(n29394), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_ier[8]), .B2(n29391), .Y(
        n29330) );
  sky130_fd_sc_hd__a22oi_1 U33895 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[8]), .A2(n29390), .B1(
        n29389), .B2(la_data_out[8]), .Y(n29329) );
  sky130_fd_sc_hd__nand3_1 U33896 ( .A(n29331), .B(n29330), .C(n29329), .Y(
        j202_soc_core_ahb2apb_02_N136) );
  sky130_fd_sc_hd__a22oi_1 U33897 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[12]), .A2(n29394), 
        .B1(n29389), .B2(la_data_out[12]), .Y(n29334) );
  sky130_fd_sc_hd__a22oi_1 U33898 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[12]), .A2(n29390), .B1(
        gpio_en_o[12]), .B2(n29393), .Y(n29333) );
  sky130_fd_sc_hd__a22oi_1 U33899 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[12]), .A2(n29392), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[12]), .B2(n29391), .Y(
        n29332) );
  sky130_fd_sc_hd__nand3_1 U33900 ( .A(n29334), .B(n29333), .C(n29332), .Y(
        j202_soc_core_ahb2apb_02_N140) );
  sky130_fd_sc_hd__a22oi_1 U33901 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[13]), .A2(n29392), .B1(
        n29389), .B2(la_data_out[13]), .Y(n29337) );
  sky130_fd_sc_hd__a22oi_1 U33902 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[13]), .A2(n29390), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[13]), .B2(n29391), .Y(
        n29336) );
  sky130_fd_sc_hd__a22oi_1 U33903 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13]), .A2(n29394), 
        .B1(gpio_en_o[13]), .B2(n29393), .Y(n29335) );
  sky130_fd_sc_hd__nand3_1 U33904 ( .A(n29337), .B(n29336), .C(n29335), .Y(
        j202_soc_core_ahb2apb_02_N141) );
  sky130_fd_sc_hd__a22oi_1 U33905 ( .A1(gpio_en_o[14]), .A2(n29393), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[14]), .B2(n29391), .Y(
        n29340) );
  sky130_fd_sc_hd__a22oi_1 U33906 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[14]), .A2(n29390), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[14]), .B2(n29392), .Y(
        n29339) );
  sky130_fd_sc_hd__a22oi_1 U33907 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14]), .A2(n29394), 
        .B1(n29389), .B2(la_data_out[14]), .Y(n29338) );
  sky130_fd_sc_hd__nand3_1 U33908 ( .A(n29340), .B(n29339), .C(n29338), .Y(
        j202_soc_core_ahb2apb_02_N142) );
  sky130_fd_sc_hd__a22oi_1 U33909 ( .A1(gpio_en_o[15]), .A2(n29393), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[15]), .B2(n29391), .Y(
        n29343) );
  sky130_fd_sc_hd__a22oi_1 U33910 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[15]), .A2(n29390), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15]), .B2(n29394), 
        .Y(n29342) );
  sky130_fd_sc_hd__a22oi_1 U33911 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[15]), .A2(n29392), .B1(
        n29389), .B2(la_data_out[15]), .Y(n29341) );
  sky130_fd_sc_hd__nand3_1 U33912 ( .A(n29343), .B(n29342), .C(n29341), .Y(
        j202_soc_core_ahb2apb_02_N143) );
  sky130_fd_sc_hd__a22oi_1 U33913 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[16]), .A2(n29390), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[16]), .B2(n29392), .Y(
        n29346) );
  sky130_fd_sc_hd__a22oi_1 U33914 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[16]), .A2(n29391), .B1(
        n29389), .B2(la_data_out[16]), .Y(n29345) );
  sky130_fd_sc_hd__a22oi_1 U33915 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16]), .A2(n29394), 
        .B1(gpio_en_o[16]), .B2(n29393), .Y(n29344) );
  sky130_fd_sc_hd__nand3_1 U33916 ( .A(n29346), .B(n29345), .C(n29344), .Y(
        j202_soc_core_ahb2apb_02_N144) );
  sky130_fd_sc_hd__a22oi_1 U33917 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[17]), .A2(n29394), 
        .B1(gpio_en_o[17]), .B2(n29393), .Y(n29349) );
  sky130_fd_sc_hd__a22oi_1 U33918 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[17]), .A2(n29390), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[17]), .B2(n29392), .Y(
        n29348) );
  sky130_fd_sc_hd__a22oi_1 U33919 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[17]), .A2(n29391), .B1(
        n29389), .B2(la_data_out[17]), .Y(n29347) );
  sky130_fd_sc_hd__nand3_1 U33920 ( .A(n29349), .B(n29348), .C(n29347), .Y(
        j202_soc_core_ahb2apb_02_N145) );
  sky130_fd_sc_hd__a22oi_1 U33921 ( .A1(n29389), .A2(la_data_out[18]), .B1(
        n29390), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_isr[18]), .Y(
        n29352) );
  sky130_fd_sc_hd__a22oi_1 U33922 ( .A1(n29393), .A2(gpio_en_o[18]), .B1(
        n29392), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_dtr[18]), .Y(
        n29351) );
  sky130_fd_sc_hd__a22oi_1 U33923 ( .A1(n29394), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[18]), .B1(n29391), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_ier[18]), .Y(n29350) );
  sky130_fd_sc_hd__nand3_1 U33924 ( .A(n29352), .B(n29351), .C(n29350), .Y(
        j202_soc_core_ahb2apb_02_N146) );
  sky130_fd_sc_hd__a22oi_1 U33925 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[19]), .A2(n29394), 
        .B1(n29389), .B2(la_data_out[19]), .Y(n29355) );
  sky130_fd_sc_hd__a22oi_1 U33926 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[19]), .A2(n29391), .B1(
        gpio_en_o[19]), .B2(n29393), .Y(n29354) );
  sky130_fd_sc_hd__a22oi_1 U33927 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[19]), .A2(n29390), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[19]), .B2(n29392), .Y(
        n29353) );
  sky130_fd_sc_hd__nand3_1 U33928 ( .A(n29355), .B(n29354), .C(n29353), .Y(
        j202_soc_core_ahb2apb_02_N147) );
  sky130_fd_sc_hd__a22oi_1 U33929 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[20]), .A2(n29392), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[20]), .B2(n29394), 
        .Y(n29358) );
  sky130_fd_sc_hd__a22oi_1 U33930 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[20]), .A2(n29391), .B1(
        n29389), .B2(la_data_out[20]), .Y(n29357) );
  sky130_fd_sc_hd__a22oi_1 U33931 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[20]), .A2(n29390), .B1(
        gpio_en_o[20]), .B2(n29393), .Y(n29356) );
  sky130_fd_sc_hd__nand3_1 U33932 ( .A(n29358), .B(n29357), .C(n29356), .Y(
        j202_soc_core_ahb2apb_02_N148) );
  sky130_fd_sc_hd__a22oi_1 U33933 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[21]), .A2(n29394), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_ier[21]), .B2(n29391), .Y(
        n29361) );
  sky130_fd_sc_hd__a22oi_1 U33934 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[21]), .A2(n29390), .B1(
        gpio_en_o[21]), .B2(n29393), .Y(n29360) );
  sky130_fd_sc_hd__a22oi_1 U33935 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[21]), .A2(n29392), .B1(
        n29389), .B2(la_data_out[21]), .Y(n29359) );
  sky130_fd_sc_hd__nand3_1 U33936 ( .A(n29361), .B(n29360), .C(n29359), .Y(
        j202_soc_core_ahb2apb_02_N149) );
  sky130_fd_sc_hd__a22oi_1 U33937 ( .A1(n29389), .A2(la_data_out[22]), .B1(
        n29390), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_isr[22]), .Y(
        n29364) );
  sky130_fd_sc_hd__a22oi_1 U33938 ( .A1(n29394), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[22]), .B1(n29393), 
        .B2(gpio_en_o[22]), .Y(n29363) );
  sky130_fd_sc_hd__a22oi_1 U33939 ( .A1(n29392), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[22]), .B1(n29391), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[22]), .Y(n29362) );
  sky130_fd_sc_hd__nand3_1 U33940 ( .A(n29364), .B(n29363), .C(n29362), .Y(
        j202_soc_core_ahb2apb_02_N150) );
  sky130_fd_sc_hd__a22oi_1 U33941 ( .A1(n29393), .A2(gpio_en_o[23]), .B1(
        n29392), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_dtr[23]), .Y(
        n29367) );
  sky130_fd_sc_hd__a22oi_1 U33942 ( .A1(n29389), .A2(la_data_out[23]), .B1(
        n29391), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_ier[23]), .Y(
        n29366) );
  sky130_fd_sc_hd__a22oi_1 U33943 ( .A1(n29394), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[23]), .B1(n29390), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_isr[23]), .Y(n29365) );
  sky130_fd_sc_hd__nand3_1 U33944 ( .A(n29367), .B(n29366), .C(n29365), .Y(
        j202_soc_core_ahb2apb_02_N151) );
  sky130_fd_sc_hd__a22oi_1 U33945 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[24]), .A2(n29390), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[24]), .B2(n29392), .Y(
        n29370) );
  sky130_fd_sc_hd__a22oi_1 U33946 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[24]), .A2(n29394), 
        .B1(gpio_en_o[24]), .B2(n29393), .Y(n29369) );
  sky130_fd_sc_hd__a22oi_1 U33947 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[24]), .A2(n29391), .B1(
        n29389), .B2(la_data_out[24]), .Y(n29368) );
  sky130_fd_sc_hd__nand3_1 U33948 ( .A(n29370), .B(n29369), .C(n29368), .Y(
        j202_soc_core_ahb2apb_02_N152) );
  sky130_fd_sc_hd__a22oi_1 U33949 ( .A1(gpio_en_o[25]), .A2(n29393), .B1(
        n29389), .B2(la_data_out[25]), .Y(n29373) );
  sky130_fd_sc_hd__a22oi_1 U33950 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[25]), .A2(n29390), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[25]), .B2(n29394), 
        .Y(n29372) );
  sky130_fd_sc_hd__a22oi_1 U33951 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[25]), .A2(n29392), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[25]), .B2(n29391), .Y(
        n29371) );
  sky130_fd_sc_hd__nand3_1 U33952 ( .A(n29373), .B(n29372), .C(n29371), .Y(
        j202_soc_core_ahb2apb_02_N153) );
  sky130_fd_sc_hd__a22oi_1 U33953 ( .A1(n29394), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[26]), .B1(n29392), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_dtr[26]), .Y(n29376) );
  sky130_fd_sc_hd__a22oi_1 U33954 ( .A1(n29393), .A2(gpio_en_o[26]), .B1(
        n29390), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_isr[26]), .Y(
        n29375) );
  sky130_fd_sc_hd__a22oi_1 U33955 ( .A1(n29389), .A2(la_data_out[26]), .B1(
        n29391), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_ier[26]), .Y(
        n29374) );
  sky130_fd_sc_hd__nand3_1 U33956 ( .A(n29376), .B(n29375), .C(n29374), .Y(
        j202_soc_core_ahb2apb_02_N154) );
  sky130_fd_sc_hd__a22oi_1 U33957 ( .A1(n29393), .A2(gpio_en_o[27]), .B1(
        n29390), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_isr[27]), .Y(
        n29379) );
  sky130_fd_sc_hd__a22oi_1 U33958 ( .A1(n29394), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[27]), .B1(n29391), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_ier[27]), .Y(n29378) );
  sky130_fd_sc_hd__a22oi_1 U33959 ( .A1(n29389), .A2(la_data_out[27]), .B1(
        n29392), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_dtr[27]), .Y(
        n29377) );
  sky130_fd_sc_hd__nand3_1 U33960 ( .A(n29379), .B(n29378), .C(n29377), .Y(
        j202_soc_core_ahb2apb_02_N155) );
  sky130_fd_sc_hd__a22oi_1 U33961 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[28]), .A2(n29390), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[28]), .B2(n29392), .Y(
        n29382) );
  sky130_fd_sc_hd__a22oi_1 U33962 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[28]), .A2(n29394), 
        .B1(gpio_en_o[28]), .B2(n29393), .Y(n29381) );
  sky130_fd_sc_hd__a22oi_1 U33963 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[28]), .A2(n29391), .B1(
        n29389), .B2(la_data_out[28]), .Y(n29380) );
  sky130_fd_sc_hd__nand3_1 U33964 ( .A(n29382), .B(n29381), .C(n29380), .Y(
        j202_soc_core_ahb2apb_02_N156) );
  sky130_fd_sc_hd__a22oi_1 U33965 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[29]), .A2(n29394), 
        .B1(n29389), .B2(la_data_out[29]), .Y(n29385) );
  sky130_fd_sc_hd__a22oi_1 U33966 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[29]), .A2(n29390), .B1(
        gpio_en_o[29]), .B2(n29393), .Y(n29384) );
  sky130_fd_sc_hd__a22oi_1 U33967 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[29]), .A2(n29392), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[29]), .B2(n29391), .Y(
        n29383) );
  sky130_fd_sc_hd__nand3_1 U33968 ( .A(n29385), .B(n29384), .C(n29383), .Y(
        j202_soc_core_ahb2apb_02_N157) );
  sky130_fd_sc_hd__a22oi_1 U33969 ( .A1(gpio_en_o[30]), .A2(n29393), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[30]), .B2(n29391), .Y(
        n29388) );
  sky130_fd_sc_hd__a22oi_1 U33970 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[30]), .A2(n29394), 
        .B1(n29389), .B2(la_data_out[30]), .Y(n29387) );
  sky130_fd_sc_hd__a22oi_1 U33971 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[30]), .A2(n29390), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[30]), .B2(n29392), .Y(
        n29386) );
  sky130_fd_sc_hd__nand3_1 U33972 ( .A(n29388), .B(n29387), .C(n29386), .Y(
        j202_soc_core_ahb2apb_02_N158) );
  sky130_fd_sc_hd__a22oi_1 U33973 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[31]), .A2(n29390), .B1(
        n29389), .B2(la_data_out[31]), .Y(n29397) );
  sky130_fd_sc_hd__a22oi_1 U33974 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[31]), .A2(n29392), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[31]), .B2(n29391), .Y(
        n29396) );
  sky130_fd_sc_hd__a22oi_1 U33975 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[31]), .A2(n29394), 
        .B1(gpio_en_o[31]), .B2(n29393), .Y(n29395) );
  sky130_fd_sc_hd__nand3_1 U33976 ( .A(n29397), .B(n29396), .C(n29395), .Y(
        j202_soc_core_ahb2apb_02_N159) );
  sky130_fd_sc_hd__nor2_1 U33977 ( .A(n29400), .B(n29399), .Y(n29404) );
  sky130_fd_sc_hd__nand2_1 U33978 ( .A(n29404), .B(
        j202_soc_core_intc_core_00_bs_addr[3]), .Y(n29417) );
  sky130_fd_sc_hd__nand2_1 U33979 ( .A(j202_soc_core_intc_core_00_bs_addr[6]), 
        .B(j202_soc_core_intc_core_00_bs_addr[4]), .Y(n29411) );
  sky130_fd_sc_hd__nand2_1 U33980 ( .A(n29409), .B(n29401), .Y(n29407) );
  sky130_fd_sc_hd__nor2_1 U33981 ( .A(n29417), .B(n29407), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_15__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand2_1 U33982 ( .A(n29405), .B(n29402), .Y(n29418) );
  sky130_fd_sc_hd__nor2_1 U33983 ( .A(n29418), .B(n29407), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_14__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand2_1 U33984 ( .A(n29404), .B(n29403), .Y(n29419) );
  sky130_fd_sc_hd__nor2_1 U33985 ( .A(n29407), .B(n29419), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_13__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand2_1 U33986 ( .A(n29406), .B(n29405), .Y(n29421) );
  sky130_fd_sc_hd__nor2_1 U33987 ( .A(n29407), .B(n29421), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_12__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33988 ( .A(j202_soc_core_intc_core_00_bs_addr[4]), 
        .B(n29408), .Y(n29415) );
  sky130_fd_sc_hd__nand2_1 U33989 ( .A(n29409), .B(n29415), .Y(n29410) );
  sky130_fd_sc_hd__nor2_1 U33990 ( .A(n29417), .B(n29410), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_11__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33991 ( .A(n29418), .B(n29410), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_10__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33992 ( .A(n29419), .B(n29410), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_9__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33993 ( .A(n29421), .B(n29410), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_8__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__or3_1 U33994 ( .A(j202_soc_core_intc_core_00_bs_addr[5]), 
        .B(n29411), .C(n29413), .X(n29412) );
  sky130_fd_sc_hd__nor2_1 U33995 ( .A(n29417), .B(n29412), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_7__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33996 ( .A(n29418), .B(n29412), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_6__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33997 ( .A(n29419), .B(n29412), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_5__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33998 ( .A(n29421), .B(n29412), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_4__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand3_1 U33999 ( .A(n29416), .B(n29415), .C(n29414), .Y(
        n29420) );
  sky130_fd_sc_hd__nor2_1 U34000 ( .A(n29417), .B(n29420), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_3__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U34001 ( .A(n29418), .B(n29420), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_2__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U34002 ( .A(n29419), .B(n29420), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_1__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U34003 ( .A(n29421), .B(n29420), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_0__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__or3_1 U34004 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[2]), .C(n28896), .X(io_out[12]) );
  sky130_fd_sc_hd__or3_1 U34005 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[3]), .C(n28896), .X(io_out[13]) );
  sky130_fd_sc_hd__nand2_1 U34006 ( .A(n29610), .B(wbs_dat_i[0]), .Y(n29422)
         );
  sky130_fd_sc_hd__nand2_1 U34007 ( .A(n470), .B(n29422), .Y(n11) );
  sky130_fd_sc_hd__xor2_1 U34008 ( .A(j202_soc_core_uart_BRG_ps[4]), .B(
        j202_soc_core_uart_div0[4]), .X(n29424) );
  sky130_fd_sc_hd__xor2_1 U34009 ( .A(j202_soc_core_uart_BRG_ps[5]), .B(
        j202_soc_core_uart_div0[5]), .X(n29423) );
  sky130_fd_sc_hd__nor2_1 U34010 ( .A(n29424), .B(n29423), .Y(n29434) );
  sky130_fd_sc_hd__xor2_1 U34011 ( .A(j202_soc_core_uart_BRG_ps[6]), .B(
        j202_soc_core_uart_div0[6]), .X(n29426) );
  sky130_fd_sc_hd__xor2_1 U34012 ( .A(j202_soc_core_uart_BRG_ps[3]), .B(
        j202_soc_core_uart_div0[3]), .X(n29425) );
  sky130_fd_sc_hd__nor2_1 U34013 ( .A(n29426), .B(n29425), .Y(n29433) );
  sky130_fd_sc_hd__xor2_1 U34014 ( .A(j202_soc_core_uart_BRG_ps[7]), .B(
        j202_soc_core_uart_div0[7]), .X(n29428) );
  sky130_fd_sc_hd__xor2_1 U34015 ( .A(j202_soc_core_uart_BRG_ps[1]), .B(
        j202_soc_core_uart_div0[1]), .X(n29427) );
  sky130_fd_sc_hd__nor2_1 U34016 ( .A(n29428), .B(n29427), .Y(n29432) );
  sky130_fd_sc_hd__xor2_1 U34017 ( .A(j202_soc_core_uart_BRG_ps[2]), .B(
        j202_soc_core_uart_div0[2]), .X(n29430) );
  sky130_fd_sc_hd__xor2_1 U34018 ( .A(j202_soc_core_uart_BRG_ps[0]), .B(
        j202_soc_core_uart_div0[0]), .X(n29429) );
  sky130_fd_sc_hd__nor2_1 U34019 ( .A(n29430), .B(n29429), .Y(n29431) );
  sky130_fd_sc_hd__and4_1 U34020 ( .A(n29434), .B(n29433), .C(n29432), .D(
        n29431), .X(j202_soc_core_uart_BRG_N21) );
  sky130_fd_sc_hd__nand3_2 U17503 ( .A(n12232), .B(n23408), .C(n27728), .Y(
        n28092) );
  sky130_fd_sc_hd__nand3_2 U16930 ( .A(n13035), .B(n30047), .C(n13034), .Y(
        n29588) );
  sky130_fd_sc_hd__nand2_4 U17446 ( .A(n11621), .B(n23421), .Y(n27899) );
  sky130_fd_sc_hd__nor2_2 U20468 ( .A(n13403), .B(n13408), .Y(n14525) );
  sky130_fd_sc_hd__nand3_2 U13415 ( .A(n13584), .B(n13583), .C(n13110), .Y(
        n28495) );
  sky130_fd_sc_hd__a22oi_2 U18025 ( .A1(n21924), .A2(n28446), .B1(n25141), 
        .B2(n17225), .Y(n17065) );
  sky130_fd_sc_hd__and4_1 U20671 ( .A(n13570), .B(n13569), .C(n13568), .D(
        n13567), .X(n13571) );
  sky130_fd_sc_hd__nand2_1 U20670 ( .A(n11200), .B(
        j202_soc_core_j22_cpu_rf_gpr[102]), .Y(n13567) );
  sky130_fd_sc_hd__nand2_2 U20467 ( .A(j202_soc_core_j22_cpu_regop_Rm__1_), 
        .B(j202_soc_core_j22_cpu_regop_Rm__0_), .Y(n13403) );
  sky130_fd_sc_hd__o21ai_1 U20989 ( .A1(n16088), .A2(n26937), .B1(n13921), .Y(
        n13924) );
  sky130_fd_sc_hd__nand2_2 U13384 ( .A(n12729), .B(n12728), .Y(n29479) );
  sky130_fd_sc_hd__inv_2 U18333 ( .A(n13819), .Y(n13726) );
  sky130_fd_sc_hd__nand2_2 U20478 ( .A(n13412), .B(
        j202_soc_core_j22_cpu_regop_Rm__1_), .Y(n13409) );
  sky130_fd_sc_hd__o21ai_1 U21442 ( .A1(n22748), .A2(n22751), .B1(n22749), .Y(
        n21342) );
  sky130_fd_sc_hd__nand2_1 U21324 ( .A(n23787), .B(
        j202_soc_core_j22_cpu_rf_gpr[454]), .Y(n14267) );
  sky130_fd_sc_hd__nor2_2 U26700 ( .A(n20896), .B(n12328), .Y(n20898) );
  sky130_fd_sc_hd__nand2_2 U19145 ( .A(n27092), .B(n27093), .Y(n27918) );
  sky130_fd_sc_hd__nand3_2 U17094 ( .A(n23438), .B(n11489), .C(n23437), .Y(
        n11488) );
  sky130_fd_sc_hd__nor2_2 U19237 ( .A(n24563), .B(n12524), .Y(n24607) );
  sky130_fd_sc_hd__inv_4 U17936 ( .A(n23378), .Y(n23421) );
  sky130_fd_sc_hd__nand2_2 U17316 ( .A(n12575), .B(n19855), .Y(n12816) );
  sky130_fd_sc_hd__nor2_1 U20990 ( .A(n13923), .B(n13924), .Y(n17219) );
  sky130_fd_sc_hd__nand2_1 U20134 ( .A(n17250), .B(n15684), .Y(n19120) );
  sky130_fd_sc_hd__o211ai_1 U25887 ( .A1(n19530), .A2(n19726), .B1(n19529), 
        .C1(n19528), .Y(n19531) );
  sky130_fd_sc_hd__nand2_2 U17028 ( .A(n11174), .B(n11176), .Y(n11724) );
  sky130_fd_sc_hd__nand2_1 U28386 ( .A(n23194), .B(n23193), .Y(n23203) );
  sky130_fd_sc_hd__nand2_2 U13657 ( .A(n20090), .B(n11928), .Y(n20888) );
  sky130_fd_sc_hd__nand3_2 U14078 ( .A(n12510), .B(n12509), .C(n22266), .Y(
        n22560) );
  sky130_fd_sc_hd__nand2_1 U13693 ( .A(n12430), .B(n11726), .Y(n22008) );
  sky130_fd_sc_hd__nand3_1 U16997 ( .A(n11382), .B(n11015), .C(n21174), .Y(
        n23386) );
  sky130_fd_sc_hd__inv_1 U17005 ( .A(n11383), .Y(n12518) );
  sky130_fd_sc_hd__nor2_4 U20095 ( .A(n21816), .B(n15198), .Y(n21020) );
  sky130_fd_sc_hd__nor2_2 U19076 ( .A(n22007), .B(n23447), .Y(n23405) );
  sky130_fd_sc_hd__inv_4 U14580 ( .A(n12351), .Y(n11183) );
  sky130_fd_sc_hd__inv_2 U13621 ( .A(n11133), .Y(n10990) );
  sky130_fd_sc_hd__inv_2 U18771 ( .A(n14209), .Y(n14993) );
  sky130_fd_sc_hd__nor2_2 U20408 ( .A(n12032), .B(n12034), .Y(n13483) );
  sky130_fd_sc_hd__nand2_1 U13483 ( .A(n21938), .B(n11401), .Y(n19243) );
  sky130_fd_sc_hd__nand2_2 U15957 ( .A(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[0]), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .Y(n23492) );
  sky130_fd_sc_hd__nand3_1 U17190 ( .A(n12017), .B(n12018), .C(n20453), .Y(
        n11666) );
  sky130_fd_sc_hd__o22ai_1 U21554 ( .A1(n16501), .A2(n26322), .B1(n26430), 
        .B2(n16500), .Y(n14575) );
  sky130_fd_sc_hd__o22ai_1 U24836 ( .A1(n22365), .A2(n22764), .B1(n21708), 
        .B2(n11561), .Y(n21703) );
  sky130_fd_sc_hd__nand2_2 U13642 ( .A(n25890), .B(n24452), .Y(n27122) );
  sky130_fd_sc_hd__o22ai_1 U23074 ( .A1(n16501), .A2(n27026), .B1(n27804), 
        .B2(n16500), .Y(n16023) );
  sky130_fd_sc_hd__nor2_2 U20520 ( .A(n12034), .B(n12033), .Y(n13481) );
  sky130_fd_sc_hd__nand2b_4 U29065 ( .A_N(n12466), .B(n30189), .Y(n23989) );
  sky130_fd_sc_hd__nor2_1 U13399 ( .A(n17041), .B(n16194), .Y(n16718) );
  sky130_fd_sc_hd__nand3_2 U14242 ( .A(n21482), .B(n21481), .C(n21480), .Y(
        n21836) );
  sky130_fd_sc_hd__nand3_2 U16939 ( .A(n12822), .B(n12453), .C(n12248), .Y(
        n24543) );
  sky130_fd_sc_hd__nand2_1 U17505 ( .A(n11684), .B(n11673), .Y(n19853) );
  sky130_fd_sc_hd__nor2_2 U28618 ( .A(n23543), .B(n23542), .Y(n25557) );
  sky130_fd_sc_hd__a21oi_2 U27642 ( .A1(n22214), .A2(n22213), .B1(n22212), .Y(
        n22219) );
  sky130_fd_sc_hd__buf_6 U24307 ( .A(n17460), .X(n18079) );
  sky130_fd_sc_hd__clkinv_1 U19058 ( .A(n12644), .Y(n12643) );
  sky130_fd_sc_hd__a21boi_1 U26048 ( .A1(n21691), .A2(n21917), .B1_N(n19846), 
        .Y(n19847) );
  sky130_fd_sc_hd__inv_2 U13879 ( .A(n12253), .Y(n12254) );
  sky130_fd_sc_hd__buf_2 U19031 ( .A(n30088), .X(n12417) );
  sky130_fd_sc_hd__nand2_2 U14509 ( .A(n12597), .B(n11550), .Y(n24578) );
  sky130_fd_sc_hd__nand2_2 U16950 ( .A(n12623), .B(n12630), .Y(n12324) );
  sky130_fd_sc_hd__nand3_2 U13522 ( .A(n27898), .B(n24695), .C(n10962), .Y(
        n22010) );
  sky130_fd_sc_hd__nand2_1 U13491 ( .A(n23395), .B(n12434), .Y(n23400) );
  sky130_fd_sc_hd__nand3_2 U14151 ( .A(n12559), .B(n12571), .C(n12558), .Y(
        n12565) );
  sky130_fd_sc_hd__nand2_1 U17547 ( .A(n11712), .B(n11207), .Y(n11710) );
  sky130_fd_sc_hd__xnor2_2 U13442 ( .A(j202_soc_core_j22_cpu_ml_bufa[18]), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .Y(n17729) );
  sky130_fd_sc_hd__buf_4 U28530 ( .A(n23405), .X(n24560) );
  sky130_fd_sc_hd__nor2_2 U18359 ( .A(n13157), .B(n13156), .Y(n21490) );
  sky130_fd_sc_hd__nand2_1 U14014 ( .A(n11927), .B(n12332), .Y(n24401) );
  sky130_fd_sc_hd__nor2_1 U17270 ( .A(n24399), .B(n28411), .Y(n12452) );
  sky130_fd_sc_hd__nor2_1 U13967 ( .A(n18665), .B(n18666), .Y(n22190) );
  sky130_fd_sc_hd__nand3_1 U17650 ( .A(n21922), .B(n21921), .C(n21923), .Y(
        n11794) );
  sky130_fd_sc_hd__nand2_2 U14021 ( .A(n11768), .B(n26377), .Y(n11765) );
  sky130_fd_sc_hd__nor2_1 U18947 ( .A(n12446), .B(n12443), .Y(n24404) );
  sky130_fd_sc_hd__nor2_8 U15294 ( .A(n13161), .B(n15198), .Y(n21633) );
  sky130_fd_sc_hd__nor2_4 U17186 ( .A(j202_soc_core_memory0_ram_dout0_sel[14]), 
        .B(n13148), .Y(n12156) );
  sky130_fd_sc_hd__nor2_8 U16977 ( .A(j202_soc_core_j22_cpu_pc[1]), .B(n19430), 
        .Y(n21917) );
  sky130_fd_sc_hd__nand2_1 U17575 ( .A(n24405), .B(n12152), .Y(n28148) );
  sky130_fd_sc_hd__a22oi_1 U26050 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__15_), .B1(n21916), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__15_), .Y(n19854) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_rf_vbr_reg_27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3339), .DE(n13071), .CLK(wb_clk_i), .Q(
        n30074), .Q_N(n30075) );
  sky130_fd_sc_hd__inv_2 U13878 ( .A(n25941), .Y(n11139) );
  sky130_fd_sc_hd__clkinv_1 U28661 ( .A(n24690), .Y(n23598) );
  sky130_fd_sc_hd__and3_1 U13962 ( .A(n23994), .B(n24591), .C(n23947), .X(
        n23399) );
  sky130_fd_sc_hd__and4_1 U15043 ( .A(n21646), .B(n21645), .C(n21644), .D(
        n21643), .X(n21647) );
  sky130_fd_sc_hd__nor2_2 U14698 ( .A(n18656), .B(n18655), .Y(n21957) );
  sky130_fd_sc_hd__a21oi_1 U19755 ( .A1(n23036), .A2(n22017), .B1(n23021), .Y(
        n23022) );
  sky130_fd_sc_hd__a22oi_2 U14413 ( .A1(n24467), .A2(n27720), .B1(n27716), 
        .B2(n24446), .Y(n24448) );
  sky130_fd_sc_hd__inv_1 U15553 ( .A(n17402), .Y(n17425) );
  sky130_fd_sc_hd__nor2_1 U27911 ( .A(n22593), .B(n22602), .Y(n22595) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__11_ ( 
        .D(n10530), .DE(n12363), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__11_), .Q_N(n30012) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__9_ ( 
        .D(n10532), .DE(n12363), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__9_), .Q_N(n30027) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__3_ ( 
        .D(n10538), .DE(n12363), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__3_), .Q_N(n30017) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__12_ ( 
        .D(n10529), .DE(n12363), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__12_), .Q_N(n30011) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__2_ ( 
        .D(n10539), .DE(n12363), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__2_), .Q_N(n30018) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_7_ ( .D(
        n29530), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[23]) );
  sky130_fd_sc_hd__buf_4 U24163 ( .A(n17341), .X(n18993) );
  sky130_fd_sc_hd__buf_4 U13480 ( .A(n17337), .X(n18533) );
  sky130_fd_sc_hd__buf_4 U13474 ( .A(n17368), .X(n19002) );
  sky130_fd_sc_hd__fa_1 U24336 ( .A(n17477), .B(n17476), .CIN(n17475), .COUT(
        n17532), .SUM(n17820) );
  sky130_fd_sc_hd__fa_1 U24378 ( .A(n17511), .B(n17510), .CIN(n17509), .COUT(
        n17531), .SUM(n17527) );
  sky130_fd_sc_hd__fa_1 U19751 ( .A(n18114), .B(n18113), .CIN(n18112), .COUT(
        n18173), .SUM(n18160) );
  sky130_fd_sc_hd__nand3_1 U19744 ( .A(n14510), .B(n12106), .C(n14509), .Y(
        n26064) );
  sky130_fd_sc_hd__a21oi_2 U14980 ( .A1(n21797), .A2(n16523), .B1(n13756), .Y(
        n26240) );
  sky130_fd_sc_hd__fa_1 U24406 ( .A(n17547), .B(n17548), .CIN(n17549), .COUT(
        n17578), .SUM(n17559) );
  sky130_fd_sc_hd__fa_1 U19806 ( .A(n17932), .B(n17931), .CIN(n17930), .COUT(
        n17921), .SUM(n17950) );
  sky130_fd_sc_hd__fa_1 U13476 ( .A(n18554), .B(n18553), .CIN(n18552), .COUT(
        n18563), .SUM(n18581) );
  sky130_fd_sc_hd__nor2_2 U18113 ( .A(n13168), .B(n13172), .Y(n20457) );
  sky130_fd_sc_hd__nor2_2 U18360 ( .A(n13150), .B(n13149), .Y(n21496) );
  sky130_fd_sc_hd__nand2_1 U14332 ( .A(n21689), .B(n21917), .Y(n11713) );
  sky130_fd_sc_hd__nand2_1 U14196 ( .A(n13086), .B(n19061), .Y(n22918) );
  sky130_fd_sc_hd__nand3_1 U27430 ( .A(n21920), .B(n21919), .C(n21918), .Y(
        n21921) );
  sky130_fd_sc_hd__nand3_1 U17889 ( .A(n12462), .B(n15389), .C(n15390), .Y(
        n29437) );
  sky130_fd_sc_hd__clkbuf_1 U13471 ( .A(n22872), .X(n11403) );
  sky130_fd_sc_hd__o21a_1 U27648 ( .A1(n22225), .A2(n22224), .B1(n22223), .X(
        n22231) );
  sky130_fd_sc_hd__nand3_2 U14135 ( .A(n11851), .B(n11850), .C(n11849), .Y(
        n12184) );
  sky130_fd_sc_hd__nand3b_1 U13468 ( .A_N(n23508), .B(
        j202_soc_core_j22_cpu_ma_M_address[1]), .C(n23510), .Y(n23513) );
  sky130_fd_sc_hd__a2bb2oi_1 U13372 ( .B1(n26034), .B2(n28451), .A1_N(n26926), 
        .A2_N(n25444), .Y(n25445) );
  sky130_fd_sc_hd__clkbuf_1 U17306 ( .A(n29490), .X(n11520) );
  sky130_fd_sc_hd__nor2_1 U19325 ( .A(n29595), .B(n24128), .Y(n12597) );
  sky130_fd_sc_hd__nor2_1 U17097 ( .A(n23947), .B(n27743), .Y(n12844) );
  sky130_fd_sc_hd__clkbuf_1 U13597 ( .A(n29437), .X(n12353) );
  sky130_fd_sc_hd__clkbuf_1 U26842 ( .A(n21693), .X(n29486) );
  sky130_fd_sc_hd__and2_1 U13493 ( .A(n12368), .B(n26189), .X(n26196) );
  sky130_fd_sc_hd__clkbuf_1 U28557 ( .A(n23551), .X(n24574) );
  sky130_fd_sc_hd__nand2_2 U13712 ( .A(n28095), .B(n24691), .Y(n24421) );
  sky130_fd_sc_hd__inv_4 U13685 ( .A(n28492), .Y(n25632) );
  sky130_fd_sc_hd__clkbuf_1 U13458 ( .A(n12798), .X(n12284) );
  sky130_fd_sc_hd__buf_2 U13578 ( .A(n26159), .X(n27047) );
  sky130_fd_sc_hd__nor2_1 U17824 ( .A(n25816), .B(n12279), .Y(n25845) );
  sky130_fd_sc_hd__clkbuf_1 U13361 ( .A(n28528), .X(n12431) );
  sky130_fd_sc_hd__clkbuf_1 U27318 ( .A(n23484), .X(n24153) );
  sky130_fd_sc_hd__inv_2 U13358 ( .A(n11442), .Y(n27668) );
  sky130_fd_sc_hd__and2_2 U13954 ( .A(n25103), .B(n30077), .X(n11114) );
  sky130_fd_sc_hd__a21oi_1 U14025 ( .A1(n28498), .A2(n23539), .B1(n23538), .Y(
        n25563) );
  sky130_fd_sc_hd__o21a_1 U28527 ( .A1(n23421), .A2(n23946), .B1(n27736), .X(
        n24583) );
  sky130_fd_sc_hd__nand2_1 U14658 ( .A(n27775), .B(n27648), .Y(n27774) );
  sky130_fd_sc_hd__a21oi_1 U13466 ( .A1(n12046), .A2(n26446), .B1(n26445), .Y(
        n26447) );
  sky130_fd_sc_hd__clkbuf_1 U26429 ( .A(n12220), .X(n29491) );
  sky130_fd_sc_hd__clkbuf_1 U26937 ( .A(n10994), .X(n29559) );
  sky130_fd_sc_hd__nand3_1 U13488 ( .A(n24956), .B(n24955), .C(n24954), .Y(
        n26978) );
  sky130_fd_sc_hd__nand2b_1 U28832 ( .A_N(n23841), .B(n23776), .Y(n23780) );
  sky130_fd_sc_hd__nand2b_1 U28834 ( .A_N(n23841), .B(n23781), .Y(n23785) );
  sky130_fd_sc_hd__inv_1 U30155 ( .A(n25478), .Y(n25023) );
  sky130_fd_sc_hd__and4_1 U14123 ( .A(n30046), .B(n20892), .C(n20891), .D(
        n20890), .X(n12127) );
  sky130_fd_sc_hd__clkinv_1 U13622 ( .A(n11133), .Y(n10993) );
  sky130_fd_sc_hd__nand2_2 U19787 ( .A(n26450), .B(n27591), .Y(n27584) );
  sky130_fd_sc_hd__nand2_1 U28820 ( .A(n23759), .B(n23758), .Y(n25978) );
  sky130_fd_sc_hd__nand2_1 U28824 ( .A(n23764), .B(n23763), .Y(n25980) );
  sky130_fd_sc_hd__nand2_1 U28845 ( .A(n23800), .B(n23799), .Y(n25983) );
  sky130_fd_sc_hd__nand2_1 U28848 ( .A(n23806), .B(n23805), .Y(n25977) );
  sky130_fd_sc_hd__nand2_1 U28853 ( .A(n23817), .B(n23816), .Y(n25986) );
  sky130_fd_sc_hd__nand2_1 U19122 ( .A(n12428), .B(n12427), .Y(n25893) );
  sky130_fd_sc_hd__nand2_1 U13450 ( .A(n29502), .B(n11853), .Y(n24471) );
  sky130_fd_sc_hd__inv_1 U13588 ( .A(n11133), .Y(n10992) );
  sky130_fd_sc_hd__and2_0 U18759 ( .A(n27124), .B(n27123), .X(n12087) );
  sky130_fd_sc_hd__nand2_2 U30652 ( .A(n25427), .B(n25425), .Y(n25555) );
  sky130_fd_sc_hd__nand2_1 U29984 ( .A(n27044), .B(n27047), .Y(n27019) );
  sky130_fd_sc_hd__buf_4 U13673 ( .A(n23979), .X(n11137) );
  sky130_fd_sc_hd__buf_4 U18991 ( .A(n24297), .X(n24307) );
  sky130_fd_sc_hd__inv_2 U13333 ( .A(n29821), .Y(n12371) );
  sky130_fd_sc_hd__clkinv_2 U19827 ( .A(n25893), .Y(n27113) );
  sky130_fd_sc_hd__clkinv_2 U30901 ( .A(n25709), .Y(n25719) );
  sky130_fd_sc_hd__clkinv_2 U18181 ( .A(n12281), .Y(n27669) );
  sky130_fd_sc_hd__clkinv_2 U14075 ( .A(n11475), .Y(n27988) );
  sky130_fd_sc_hd__nor2_1 U18350 ( .A(n13170), .B(n13169), .Y(n20456) );
  sky130_fd_sc_hd__nor2_4 U16976 ( .A(n15199), .B(n15198), .Y(n21488) );
  sky130_fd_sc_hd__inv_2 U14251 ( .A(n16294), .Y(n20462) );
  sky130_fd_sc_hd__nand2_1 U13593 ( .A(n24179), .B(n22739), .Y(n17068) );
  sky130_fd_sc_hd__nand2_1 U14213 ( .A(n12567), .B(n22230), .Y(n12566) );
  sky130_fd_sc_hd__a21oi_1 U19024 ( .A1(n23036), .A2(n21762), .B1(n21761), .Y(
        n21763) );
  sky130_fd_sc_hd__xnor2_1 U16917 ( .A(n12108), .B(n11348), .Y(n12673) );
  sky130_fd_sc_hd__o21a_1 U18970 ( .A1(n26158), .A2(n12279), .B1(n30077), .X(
        n28470) );
  sky130_fd_sc_hd__o211ai_1 U27943 ( .A1(n27052), .A2(n23579), .B1(n22638), 
        .C1(n22637), .Y(n25817) );
  sky130_fd_sc_hd__and2b_1 U13957 ( .B(n29545), .A_N(n25024), .X(n23986) );
  sky130_fd_sc_hd__nand3_1 U31185 ( .A(n25993), .B(n25992), .C(n25991), .Y(
        n26025) );
  sky130_fd_sc_hd__a21oi_1 U17819 ( .A1(n11950), .A2(n25853), .B1(n11947), .Y(
        n25857) );
  sky130_fd_sc_hd__inv_2 U13591 ( .A(n12369), .Y(n11133) );
  sky130_fd_sc_hd__o21a_1 U31490 ( .A1(n26449), .A2(n26448), .B1(n26447), .X(
        n27591) );
  sky130_fd_sc_hd__nor2_1 U13653 ( .A(n23978), .B(n12466), .Y(n23979) );
  sky130_fd_sc_hd__nand2_1 U13322 ( .A(n11978), .B(n12459), .Y(n30150) );
  sky130_fd_sc_hd__clkinv_1 U13323 ( .A(n30149), .Y(n12461) );
  sky130_fd_sc_hd__nand3_1 U13324 ( .A(n12892), .B(n11100), .C(n12893), .Y(
        n11348) );
  sky130_fd_sc_hd__nand3_1 U13327 ( .A(n17057), .B(n17058), .C(n17095), .Y(
        n30149) );
  sky130_fd_sc_hd__inv_6 U13350 ( .A(n22107), .Y(n23030) );
  sky130_fd_sc_hd__nand2_1 U13354 ( .A(n30159), .B(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n21689) );
  sky130_fd_sc_hd__nand2_1 U13357 ( .A(n24297), .B(n29830), .Y(n30052) );
  sky130_fd_sc_hd__nand2_1 U13363 ( .A(n24297), .B(n29830), .Y(
        j202_soc_core_ahb2apb_02_N22) );
  sky130_fd_sc_hd__inv_4 U13365 ( .A(n26454), .Y(n26453) );
  sky130_fd_sc_hd__inv_2 U13375 ( .A(n29821), .Y(n12370) );
  sky130_fd_sc_hd__clkinv_2 U13377 ( .A(n27087), .Y(n27089) );
  sky130_fd_sc_hd__inv_2 U13383 ( .A(n30180), .Y(n30193) );
  sky130_fd_sc_hd__inv_2 U13385 ( .A(n30182), .Y(n30195) );
  sky130_fd_sc_hd__inv_2 U13386 ( .A(n30183), .Y(n30196) );
  sky130_fd_sc_hd__buf_2 U13387 ( .A(n24957), .X(n26972) );
  sky130_fd_sc_hd__clkinv_1 U13389 ( .A(n30181), .Y(n30192) );
  sky130_fd_sc_hd__clkinv_1 U13390 ( .A(n30186), .Y(n30191) );
  sky130_fd_sc_hd__clkbuf_1 U13392 ( .A(n16100), .X(n30058) );
  sky130_fd_sc_hd__inv_8 U13404 ( .A(n12386), .Y(n11135) );
  sky130_fd_sc_hd__inv_2 U13408 ( .A(n10992), .Y(n30099) );
  sky130_fd_sc_hd__nor2_1 U13426 ( .A(n21317), .B(n12359), .Y(n29551) );
  sky130_fd_sc_hd__nand3_1 U13446 ( .A(n22688), .B(n19313), .C(n19312), .Y(
        n29499) );
  sky130_fd_sc_hd__a21oi_1 U13452 ( .A1(n12361), .A2(n24952), .B1(n24951), .Y(
        n24955) );
  sky130_fd_sc_hd__nand2_1 U13454 ( .A(n25417), .B(n25416), .Y(n25418) );
  sky130_fd_sc_hd__nand3_1 U13459 ( .A(n12459), .B(n12461), .C(n30046), .Y(
        n12328) );
  sky130_fd_sc_hd__nand2_1 U13461 ( .A(n22121), .B(n22120), .Y(n22147) );
  sky130_fd_sc_hd__o21ai_1 U13462 ( .A1(n21764), .A2(n12349), .B1(n21763), .Y(
        n12887) );
  sky130_fd_sc_hd__nor2_1 U13470 ( .A(n30164), .B(n30163), .Y(n30162) );
  sky130_fd_sc_hd__nand3_1 U13479 ( .A(n17068), .B(n17063), .C(n16566), .Y(
        n16567) );
  sky130_fd_sc_hd__nand2_1 U13481 ( .A(n11852), .B(n22739), .Y(n17066) );
  sky130_fd_sc_hd__a21o_1 U13486 ( .A1(n17040), .A2(n16028), .B1(n16027), .X(
        n30158) );
  sky130_fd_sc_hd__nand2_1 U13495 ( .A(n18668), .B(n22193), .Y(n18670) );
  sky130_fd_sc_hd__nor2_1 U13511 ( .A(n13018), .B(n13013), .Y(n13012) );
  sky130_fd_sc_hd__o21ai_1 U13514 ( .A1(n21232), .A2(n21235), .B1(n21236), .Y(
        n21866) );
  sky130_fd_sc_hd__inv_6 U13515 ( .A(n24912), .Y(n28109) );
  sky130_fd_sc_hd__xor2_1 U13520 ( .A(n12508), .B(n30041), .X(n18538) );
  sky130_fd_sc_hd__and2_1 U13521 ( .A(n18868), .B(n13431), .X(n11093) );
  sky130_fd_sc_hd__nor2_1 U13524 ( .A(j202_soc_core_j22_cpu_regop_Rm__3_), .B(
        j202_soc_core_j22_cpu_regop_Rm__2_), .Y(n13385) );
  sky130_fd_sc_hd__clkinv_1 U13529 ( .A(j202_soc_core_j22_cpu_ml_bufa[12]), 
        .Y(n17452) );
  sky130_fd_sc_hd__o21ai_0 U13530 ( .A1(n16820), .A2(n16819), .B1(n16818), .Y(
        n16821) );
  sky130_fd_sc_hd__o21ai_0 U13531 ( .A1(n15159), .A2(n15270), .B1(n15532), .Y(
        n15160) );
  sky130_fd_sc_hd__o21ai_0 U13533 ( .A1(n15330), .A2(n15329), .B1(n21103), .Y(
        n15331) );
  sky130_fd_sc_hd__clkinv_1 U13539 ( .A(n19203), .Y(n16634) );
  sky130_fd_sc_hd__o21ai_0 U13541 ( .A1(n16844), .A2(n16843), .B1(n19394), .Y(
        n16855) );
  sky130_fd_sc_hd__o21ai_0 U13546 ( .A1(n16850), .A2(n16763), .B1(n16747), .Y(
        n16748) );
  sky130_fd_sc_hd__clkinv_1 U13550 ( .A(n16942), .Y(n15719) );
  sky130_fd_sc_hd__inv_2 U13552 ( .A(n20126), .Y(n15111) );
  sky130_fd_sc_hd__o21ai_0 U13556 ( .A1(n18396), .A2(n18397), .B1(n18395), .Y(
        n30036) );
  sky130_fd_sc_hd__clkinv_1 U13558 ( .A(n30119), .Y(n30114) );
  sky130_fd_sc_hd__o21ai_0 U13559 ( .A1(n22047), .A2(n22784), .B1(n22046), .Y(
        n22048) );
  sky130_fd_sc_hd__clkinv_1 U13560 ( .A(n15339), .Y(n15569) );
  sky130_fd_sc_hd__o21ai_0 U13561 ( .A1(n15294), .A2(n15293), .B1(n21103), .Y(
        n15298) );
  sky130_fd_sc_hd__clkinv_1 U13580 ( .A(n15148), .Y(n15570) );
  sky130_fd_sc_hd__clkinv_1 U13583 ( .A(n14619), .Y(n14698) );
  sky130_fd_sc_hd__o21ai_0 U13584 ( .A1(n14677), .A2(n14676), .B1(n17242), .Y(
        n14679) );
  sky130_fd_sc_hd__o21ai_0 U13592 ( .A1(n15299), .A2(n15291), .B1(n17237), .Y(
        n15144) );
  sky130_fd_sc_hd__clkinv_1 U13594 ( .A(n20809), .Y(n19184) );
  sky130_fd_sc_hd__clkinv_1 U13596 ( .A(n17100), .Y(n15668) );
  sky130_fd_sc_hd__clkinv_1 U13601 ( .A(n16959), .Y(n16641) );
  sky130_fd_sc_hd__o21ai_0 U13602 ( .A1(n16772), .A2(n16152), .B1(n20368), .Y(
        n16172) );
  sky130_fd_sc_hd__o21ai_0 U13607 ( .A1(n16134), .A2(n16133), .B1(n20393), .Y(
        n16146) );
  sky130_fd_sc_hd__o21ai_0 U13608 ( .A1(n16814), .A2(n16795), .B1(n20374), .Y(
        n16796) );
  sky130_fd_sc_hd__o21ai_0 U13609 ( .A1(n19184), .A2(n21101), .B1(n16858), .Y(
        n16272) );
  sky130_fd_sc_hd__o21ai_0 U13610 ( .A1(n15294), .A2(n15211), .B1(n17237), .Y(
        n15104) );
  sky130_fd_sc_hd__o21ai_0 U13611 ( .A1(n17762), .A2(n11145), .B1(n17375), .Y(
        n17403) );
  sky130_fd_sc_hd__clkinv_1 U13613 ( .A(n18277), .Y(n12178) );
  sky130_fd_sc_hd__o21ai_0 U13615 ( .A1(n24934), .A2(n24933), .B1(n26414), .Y(
        n24937) );
  sky130_fd_sc_hd__o21ai_0 U13616 ( .A1(n21687), .A2(n18340), .B1(n18339), .Y(
        n18481) );
  sky130_fd_sc_hd__o21ai_0 U13618 ( .A1(n23026), .A2(n23031), .B1(n23027), .Y(
        n22506) );
  sky130_fd_sc_hd__or2_0 U13624 ( .A(n17561), .B(n18471), .X(n30082) );
  sky130_fd_sc_hd__nor2b_1 U13626 ( .B_N(n18470), .A(n18474), .Y(n17487) );
  sky130_fd_sc_hd__clkinv_1 U13630 ( .A(n22543), .Y(n22674) );
  sky130_fd_sc_hd__o22ai_1 U13632 ( .A1(n18474), .A2(n17416), .B1(n17429), 
        .B2(n18471), .Y(n18413) );
  sky130_fd_sc_hd__buf_2 U13639 ( .A(j202_soc_core_j22_cpu_ml_bufb[13]), .X(
        n18994) );
  sky130_fd_sc_hd__o21ai_0 U13645 ( .A1(n16676), .A2(n16675), .B1(n17099), .Y(
        n16709) );
  sky130_fd_sc_hd__o21ai_0 U13648 ( .A1(n17161), .A2(n20515), .B1(n19571), .Y(
        n17163) );
  sky130_fd_sc_hd__o21ai_0 U13651 ( .A1(n15355), .A2(n15354), .B1(n17237), .Y(
        n15356) );
  sky130_fd_sc_hd__o21ai_0 U13654 ( .A1(n15285), .A2(n15284), .B1(n17237), .Y(
        n15286) );
  sky130_fd_sc_hd__clkinv_1 U13655 ( .A(n19763), .Y(n13235) );
  sky130_fd_sc_hd__o21ai_0 U13656 ( .A1(n16373), .A2(n16942), .B1(n16980), .Y(
        n16379) );
  sky130_fd_sc_hd__o21ai_0 U13661 ( .A1(n16118), .A2(n16782), .B1(n20393), .Y(
        n16119) );
  sky130_fd_sc_hd__o21ai_0 U13662 ( .A1(n20626), .A2(n19165), .B1(n20833), .Y(
        n19166) );
  sky130_fd_sc_hd__o21ai_0 U13663 ( .A1(n16278), .A2(n16277), .B1(n20368), .Y(
        n16279) );
  sky130_fd_sc_hd__clkinv_1 U13664 ( .A(n15684), .Y(n20810) );
  sky130_fd_sc_hd__o21ai_0 U13670 ( .A1(n18982), .A2(n11145), .B1(n18981), .Y(
        n19039) );
  sky130_fd_sc_hd__o21ai_0 U13671 ( .A1(n21745), .A2(n11145), .B1(n18974), .Y(
        n19003) );
  sky130_fd_sc_hd__o21ai_0 U13672 ( .A1(n15597), .A2(n15232), .B1(n17237), .Y(
        n15233) );
  sky130_fd_sc_hd__o21ai_0 U13675 ( .A1(n15227), .A2(n15226), .B1(n19804), .Y(
        n15235) );
  sky130_fd_sc_hd__o21ai_0 U13678 ( .A1(n15501), .A2(n15205), .B1(n19804), .Y(
        n15206) );
  sky130_fd_sc_hd__o21ai_0 U13681 ( .A1(n18619), .A2(n18623), .B1(n18620), .Y(
        n18507) );
  sky130_fd_sc_hd__clkinv_1 U13683 ( .A(n18416), .Y(n18354) );
  sky130_fd_sc_hd__o21ai_0 U13684 ( .A1(n12668), .A2(n17612), .B1(n17611), .Y(
        n12666) );
  sky130_fd_sc_hd__clkinv_1 U13692 ( .A(n22335), .Y(n22336) );
  sky130_fd_sc_hd__o21ai_0 U13696 ( .A1(n18433), .A2(n18432), .B1(n12504), .Y(
        n12503) );
  sky130_fd_sc_hd__o21ai_0 U13697 ( .A1(n15605), .A2(n15604), .B1(n19816), .Y(
        n15606) );
  sky130_fd_sc_hd__o21ai_0 U13699 ( .A1(n15512), .A2(n15511), .B1(n19816), .Y(
        n15513) );
  sky130_fd_sc_hd__o21ai_0 U13703 ( .A1(n16223), .A2(n14671), .B1(n20368), .Y(
        n14691) );
  sky130_fd_sc_hd__o21ai_0 U13705 ( .A1(n14615), .A2(n16743), .B1(n20393), .Y(
        n14616) );
  sky130_fd_sc_hd__clkinv_1 U13711 ( .A(n17108), .Y(n20673) );
  sky130_fd_sc_hd__o21ai_0 U13715 ( .A1(n26347), .A2(n26346), .B1(n26345), .Y(
        n26349) );
  sky130_fd_sc_hd__o21ai_0 U13726 ( .A1(n27023), .A2(n23531), .B1(n21202), .Y(
        n21208) );
  sky130_fd_sc_hd__o21ai_0 U13727 ( .A1(n20044), .A2(n20043), .B1(n20113), .Y(
        n20045) );
  sky130_fd_sc_hd__clkinv_1 U13731 ( .A(n19579), .Y(n19610) );
  sky130_fd_sc_hd__o21ai_0 U13732 ( .A1(n18735), .A2(n18734), .B1(n20225), .Y(
        n18736) );
  sky130_fd_sc_hd__clkinv_1 U13734 ( .A(n20804), .Y(n20846) );
  sky130_fd_sc_hd__clkinv_1 U13762 ( .A(n20623), .Y(n19178) );
  sky130_fd_sc_hd__clkinv_1 U13763 ( .A(n20625), .Y(n20496) );
  sky130_fd_sc_hd__o21ai_0 U13764 ( .A1(n20304), .A2(n20303), .B1(n20302), .Y(
        n20305) );
  sky130_fd_sc_hd__inv_2 U13765 ( .A(n13179), .Y(n21359) );
  sky130_fd_sc_hd__clkinv_1 U13771 ( .A(n19571), .Y(n19607) );
  sky130_fd_sc_hd__clkinv_1 U13772 ( .A(n19779), .Y(n19513) );
  sky130_fd_sc_hd__o21ai_0 U13774 ( .A1(n19444), .A2(n19470), .B1(n19816), .Y(
        n13216) );
  sky130_fd_sc_hd__o21ai_0 U13776 ( .A1(n16320), .A2(n16976), .B1(n16980), .Y(
        n16329) );
  sky130_fd_sc_hd__or2_0 U13785 ( .A(n19148), .B(n19130), .X(n16986) );
  sky130_fd_sc_hd__o21ai_0 U13793 ( .A1(n16130), .A2(n16129), .B1(n16770), .Y(
        n16176) );
  sky130_fd_sc_hd__o21ai_0 U13801 ( .A1(j202_soc_core_j22_cpu_id_op2_inst__12_), .A2(j202_soc_core_j22_cpu_id_op2_inst__13_), .B1(
        j202_soc_core_j22_cpu_id_op2_v_), .Y(n19859) );
  sky130_fd_sc_hd__o21ai_0 U13810 ( .A1(n15757), .A2(n16995), .B1(n17099), .Y(
        n15767) );
  sky130_fd_sc_hd__clkinv_1 U13814 ( .A(n15409), .Y(n19728) );
  sky130_fd_sc_hd__o21ai_0 U13821 ( .A1(n11860), .A2(n18235), .B1(n18234), .Y(
        n11858) );
  sky130_fd_sc_hd__o21ai_0 U13822 ( .A1(n25872), .A2(n26226), .B1(n24834), .Y(
        n24840) );
  sky130_fd_sc_hd__o21ai_0 U13837 ( .A1(n18556), .A2(n18557), .B1(n18555), .Y(
        n11881) );
  sky130_fd_sc_hd__o21ai_0 U13846 ( .A1(n22599), .A2(n22603), .B1(n22600), .Y(
        n22511) );
  sky130_fd_sc_hd__or2_0 U13849 ( .A(n17761), .B(n17760), .X(n17764) );
  sky130_fd_sc_hd__o21ai_0 U13854 ( .A1(n18307), .A2(n18306), .B1(n18305), .Y(
        n30136) );
  sky130_fd_sc_hd__o21ai_0 U13859 ( .A1(n21961), .A2(n21957), .B1(n21958), .Y(
        n18657) );
  sky130_fd_sc_hd__o21ai_0 U13864 ( .A1(n18630), .A2(n18632), .B1(n18629), .Y(
        n18559) );
  sky130_fd_sc_hd__o21ai_0 U13869 ( .A1(n26435), .A2(n27803), .B1(n25445), .Y(
        n25447) );
  sky130_fd_sc_hd__o21ai_0 U13871 ( .A1(n26285), .A2(n26932), .B1(n21941), .Y(
        n21952) );
  sky130_fd_sc_hd__o21ai_0 U13872 ( .A1(n27796), .A2(n27795), .B1(n27794), .Y(
        n27802) );
  sky130_fd_sc_hd__o21ai_0 U13874 ( .A1(n19818), .A2(n19817), .B1(n19816), .Y(
        n19834) );
  sky130_fd_sc_hd__o21ai_0 U13876 ( .A1(n18757), .A2(n20206), .B1(n20210), .Y(
        n18758) );
  sky130_fd_sc_hd__o21ai_0 U13877 ( .A1(n19970), .A2(n18746), .B1(n20225), .Y(
        n18761) );
  sky130_fd_sc_hd__o21ai_0 U13883 ( .A1(n20764), .A2(n20763), .B1(n20833), .Y(
        n20783) );
  sky130_fd_sc_hd__o21ai_0 U13884 ( .A1(n21580), .A2(n21419), .B1(n17290), .Y(
        n17297) );
  sky130_fd_sc_hd__clkinv_1 U13889 ( .A(n20381), .Y(n20277) );
  sky130_fd_sc_hd__o21ai_0 U13893 ( .A1(n23327), .A2(n23328), .B1(n23323), .Y(
        n23303) );
  sky130_fd_sc_hd__clkinv_1 U13896 ( .A(n16994), .Y(n17001) );
  sky130_fd_sc_hd__o21ai_0 U13914 ( .A1(n16968), .A2(n16967), .B1(n16980), .Y(
        n16971) );
  sky130_fd_sc_hd__o21ai_0 U13917 ( .A1(n16257), .A2(n16256), .B1(n16840), .Y(
        n16285) );
  sky130_fd_sc_hd__o21ai_0 U13920 ( .A1(n15448), .A2(n15447), .B1(n17237), .Y(
        n15460) );
  sky130_fd_sc_hd__and2_0 U13924 ( .A(n19855), .B(n21917), .X(n13082) );
  sky130_fd_sc_hd__nand2_1 U13927 ( .A(j202_soc_core_memory0_ram_dout0[445]), 
        .B(n12156), .Y(n12447) );
  sky130_fd_sc_hd__a2bb2oi_1 U13928 ( .B1(n15577), .B2(n15217), .A1_N(n19728), 
        .A2_N(n15216), .Y(n15239) );
  sky130_fd_sc_hd__clkinv_1 U13931 ( .A(n22196), .Y(n22198) );
  sky130_fd_sc_hd__o21ai_0 U13933 ( .A1(n21007), .A2(n21011), .B1(n21012), .Y(
        n14406) );
  sky130_fd_sc_hd__o21ai_0 U13947 ( .A1(n25682), .A2(n26331), .B1(n25636), .Y(
        n25637) );
  sky130_fd_sc_hd__a2bb2oi_1 U13953 ( .B1(n27810), .B2(n25697), .A1_N(n25872), 
        .A2_N(n26230), .Y(n25298) );
  sky130_fd_sc_hd__and2_0 U13956 ( .A(n22017), .B(n22512), .X(n22514) );
  sky130_fd_sc_hd__o21ai_0 U13963 ( .A1(n17624), .A2(n17623), .B1(n17622), .Y(
        n17626) );
  sky130_fd_sc_hd__o21ai_0 U13964 ( .A1(n17874), .A2(n17875), .B1(n17877), .Y(
        n17805) );
  sky130_fd_sc_hd__o21ai_0 U13965 ( .A1(n22920), .A2(n22921), .B1(n22919), .Y(
        n22922) );
  sky130_fd_sc_hd__clkinv_1 U13970 ( .A(n27803), .Y(n26942) );
  sky130_fd_sc_hd__o21ai_0 U13974 ( .A1(n26926), .A2(n22456), .B1(n21861), .Y(
        n21862) );
  sky130_fd_sc_hd__o21ai_0 U13977 ( .A1(n26049), .A2(n26048), .B1(n26047), .Y(
        n26053) );
  sky130_fd_sc_hd__o21ai_0 U13979 ( .A1(n21619), .A2(n21618), .B1(n21617), .Y(
        n21620) );
  sky130_fd_sc_hd__o21ai_0 U13983 ( .A1(n21557), .A2(n21618), .B1(n21603), .Y(
        n21558) );
  sky130_fd_sc_hd__inv_2 U13991 ( .A(n19058), .Y(n21903) );
  sky130_fd_sc_hd__o21ai_0 U13997 ( .A1(n14618), .A2(n16129), .B1(n16770), .Y(
        n14720) );
  sky130_fd_sc_hd__inv_2 U14000 ( .A(n11142), .Y(n11184) );
  sky130_fd_sc_hd__o21ai_0 U14009 ( .A1(n20650), .A2(n20686), .B1(n20833), .Y(
        n20671) );
  sky130_fd_sc_hd__clkinv_1 U14043 ( .A(n21580), .Y(n21610) );
  sky130_fd_sc_hd__o21ai_0 U14045 ( .A1(n19482), .A2(n19704), .B1(n19804), .Y(
        n19501) );
  sky130_fd_sc_hd__o21ai_0 U14059 ( .A1(n19438), .A2(n19805), .B1(n19816), .Y(
        n19455) );
  sky130_fd_sc_hd__o21ai_0 U14063 ( .A1(n20212), .A2(n20211), .B1(n20210), .Y(
        n20233) );
  sky130_fd_sc_hd__o21ai_0 U14070 ( .A1(n20136), .A2(n20135), .B1(n20227), .Y(
        n20161) );
  sky130_fd_sc_hd__clkinv_1 U14080 ( .A(n12316), .Y(n11579) );
  sky130_fd_sc_hd__o21ai_0 U14106 ( .A1(n19671), .A2(n19670), .B1(n20368), .Y(
        n19672) );
  sky130_fd_sc_hd__o21ai_0 U14107 ( .A1(n20282), .A2(n19553), .B1(n20393), .Y(
        n19569) );
  sky130_fd_sc_hd__clkinv_1 U14109 ( .A(n20140), .Y(n20003) );
  sky130_fd_sc_hd__o21ai_0 U14117 ( .A1(n19867), .A2(n20198), .B1(n20227), .Y(
        n19868) );
  sky130_fd_sc_hd__o21ai_0 U14122 ( .A1(n20835), .A2(n20834), .B1(n20833), .Y(
        n20861) );
  sky130_fd_sc_hd__o21ai_0 U14124 ( .A1(n17260), .A2(n21107), .B1(n21598), .Y(
        n17261) );
  sky130_fd_sc_hd__o21ai_0 U14136 ( .A1(n20395), .A2(n20394), .B1(n20393), .Y(
        n20396) );
  sky130_fd_sc_hd__o21ai_0 U14148 ( .A1(n20283), .A2(n20282), .B1(n20393), .Y(
        n20284) );
  sky130_fd_sc_hd__o21ai_0 U14149 ( .A1(n17116), .A2(n19317), .B1(n20374), .Y(
        n17117) );
  sky130_fd_sc_hd__o21ai_0 U14163 ( .A1(n13210), .A2(n19797), .B1(n19816), .Y(
        n13212) );
  sky130_fd_sc_hd__o21ai_0 U14171 ( .A1(n16982), .A2(n16981), .B1(n16980), .Y(
        n17000) );
  sky130_fd_sc_hd__o21ai_0 U14173 ( .A1(n19209), .A2(n20646), .B1(n20856), .Y(
        n19210) );
  sky130_fd_sc_hd__o21ai_0 U14188 ( .A1(n22199), .A2(n22198), .B1(n22197), .Y(
        n22200) );
  sky130_fd_sc_hd__fa_1 U14195 ( .A(n18301), .B(n18300), .CIN(n18299), .COUT(
        n17999), .SUM(n18310) );
  sky130_fd_sc_hd__o21ai_0 U14217 ( .A1(n21273), .A2(n21268), .B1(n21269), .Y(
        n22959) );
  sky130_fd_sc_hd__o21ai_0 U14222 ( .A1(n17573), .A2(n17574), .B1(n17572), .Y(
        n12413) );
  sky130_fd_sc_hd__clkinv_1 U14231 ( .A(n13446), .Y(n14200) );
  sky130_fd_sc_hd__o21ai_0 U14244 ( .A1(n16552), .A2(n16551), .B1(n16550), .Y(
        n16553) );
  sky130_fd_sc_hd__o21ai_0 U14291 ( .A1(n26411), .A2(n26929), .B1(n27787), .Y(
        n19257) );
  sky130_fd_sc_hd__o21ai_0 U14326 ( .A1(j202_soc_core_j22_cpu_regop_other__2_), 
        .A2(n13428), .B1(j202_soc_core_j22_cpu_regop_Rs__0_), .Y(n13301) );
  sky130_fd_sc_hd__clkinv_1 U14339 ( .A(n12032), .Y(n12033) );
  sky130_fd_sc_hd__clkinv_1 U14355 ( .A(n22915), .Y(n22917) );
  sky130_fd_sc_hd__clkinv_1 U14372 ( .A(j202_soc_core_j22_cpu_regop_Ra__1_), 
        .Y(n13477) );
  sky130_fd_sc_hd__o21ai_0 U14381 ( .A1(n17031), .A2(n17041), .B1(n17042), .Y(
        n16720) );
  sky130_fd_sc_hd__o21ai_0 U14382 ( .A1(n21832), .A2(n21831), .B1(n22232), .Y(
        n21834) );
  sky130_fd_sc_hd__o21ai_0 U14384 ( .A1(n15640), .A2(n15184), .B1(n15185), .Y(
        n15080) );
  sky130_fd_sc_hd__o21ai_0 U14391 ( .A1(n16893), .A2(n16901), .B1(n16902), .Y(
        n16019) );
  sky130_fd_sc_hd__clkinv_1 U14393 ( .A(n30042), .Y(n11540) );
  sky130_fd_sc_hd__clkinv_1 U14404 ( .A(n28409), .Y(n12217) );
  sky130_fd_sc_hd__o21ai_0 U14405 ( .A1(n26926), .A2(n22387), .B1(n18851), .Y(
        n18852) );
  sky130_fd_sc_hd__o21ai_0 U14408 ( .A1(n21133), .A2(n21523), .B1(n21603), .Y(
        n21134) );
  sky130_fd_sc_hd__o21ai_0 U14409 ( .A1(n21090), .A2(n21530), .B1(n21610), .Y(
        n21091) );
  sky130_fd_sc_hd__clkinv_1 U14412 ( .A(n29437), .Y(n17057) );
  sky130_fd_sc_hd__o21ai_0 U14414 ( .A1(n15490), .A2(n15384), .B1(n15385), .Y(
        n15180) );
  sky130_fd_sc_hd__clkinv_1 U14421 ( .A(n19853), .Y(n11748) );
  sky130_fd_sc_hd__and2_0 U14428 ( .A(n23421), .B(n12861), .X(n12153) );
  sky130_fd_sc_hd__o21ai_0 U14431 ( .A1(n20596), .A2(n20536), .B1(n20833), .Y(
        n20537) );
  sky130_fd_sc_hd__o21ai_0 U14432 ( .A1(n20500), .A2(n20499), .B1(n20833), .Y(
        n20501) );
  sky130_fd_sc_hd__o21ai_0 U14443 ( .A1(n21412), .A2(n17300), .B1(n17299), .Y(
        n17301) );
  sky130_fd_sc_hd__o21ai_0 U14454 ( .A1(n19375), .A2(n19374), .B1(n20368), .Y(
        n19385) );
  sky130_fd_sc_hd__o21ai_0 U14463 ( .A1(n19331), .A2(n19620), .B1(n20374), .Y(
        n19332) );
  sky130_fd_sc_hd__inv_2 U14467 ( .A(n11855), .Y(n11886) );
  sky130_fd_sc_hd__clkinv_1 U14471 ( .A(n12858), .Y(n12634) );
  sky130_fd_sc_hd__o21ai_0 U14476 ( .A1(n13781), .A2(n16490), .B1(n13780), .Y(
        n13783) );
  sky130_fd_sc_hd__nor2_1 U14479 ( .A(j202_soc_core_j22_cpu_regop_other__0_), 
        .B(n18859), .Y(n13429) );
  sky130_fd_sc_hd__and2_0 U14485 ( .A(n24631), .B(n24630), .X(n11113) );
  sky130_fd_sc_hd__clkinv_1 U14490 ( .A(n22190), .Y(n22192) );
  sky130_fd_sc_hd__o21ai_0 U14493 ( .A1(n16543), .A2(n25692), .B1(n14928), .Y(
        n15073) );
  sky130_fd_sc_hd__nor2_1 U14496 ( .A(n18316), .B(n18317), .Y(n21969) );
  sky130_fd_sc_hd__o21ai_0 U14503 ( .A1(n16088), .A2(n27816), .B1(n14353), .Y(
        n14395) );
  sky130_fd_sc_hd__o21ai_0 U14507 ( .A1(n16543), .A2(n28460), .B1(n14071), .Y(
        n14401) );
  sky130_fd_sc_hd__o21ai_0 U14511 ( .A1(n11123), .A2(n26009), .B1(n26922), .Y(
        n25958) );
  sky130_fd_sc_hd__o21ai_0 U14512 ( .A1(n22837), .A2(n12349), .B1(n22836), .Y(
        n22838) );
  sky130_fd_sc_hd__buf_1 U14519 ( .A(n21964), .X(n11349) );
  sky130_fd_sc_hd__o21ai_0 U14538 ( .A1(n11471), .A2(n22961), .B1(n22960), .Y(
        n22963) );
  sky130_fd_sc_hd__o21ai_0 U14550 ( .A1(n22552), .A2(n12349), .B1(n22551), .Y(
        n22553) );
  sky130_fd_sc_hd__o21ai_0 U14563 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[5]), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[9]), .B1(n24009), .Y(
        n24010) );
  sky130_fd_sc_hd__o21ai_0 U14564 ( .A1(n16543), .A2(n28493), .B1(n15037), .Y(
        n15079) );
  sky130_fd_sc_hd__o21ai_0 U14566 ( .A1(n16088), .A2(n26276), .B1(n15895), .Y(
        n16016) );
  sky130_fd_sc_hd__o21ai_0 U14570 ( .A1(n16543), .A2(n25825), .B1(n15977), .Y(
        n16024) );
  sky130_fd_sc_hd__o21ai_0 U14581 ( .A1(n11866), .A2(n22075), .B1(n22074), .Y(
        n22076) );
  sky130_fd_sc_hd__o21ai_0 U14596 ( .A1(n26926), .A2(n22421), .B1(n21725), .Y(
        n21726) );
  sky130_fd_sc_hd__o21a_1 U14605 ( .A1(n12279), .A2(n24179), .B1(n30077), .X(
        n28430) );
  sky130_fd_sc_hd__clkinv_1 U14635 ( .A(n16524), .Y(n16493) );
  sky130_fd_sc_hd__o21ai_0 U14644 ( .A1(n11123), .A2(n26050), .B1(n26922), .Y(
        n25401) );
  sky130_fd_sc_hd__clkinv_1 U14645 ( .A(n22199), .Y(n21810) );
  sky130_fd_sc_hd__clkinv_1 U14649 ( .A(n11941), .Y(n23949) );
  sky130_fd_sc_hd__clkinv_1 U14655 ( .A(n27886), .Y(n11730) );
  sky130_fd_sc_hd__clkinv_1 U14656 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .Y(n18809) );
  sky130_fd_sc_hd__o21ai_0 U14661 ( .A1(n16088), .A2(n28451), .B1(n16087), .Y(
        n16090) );
  sky130_fd_sc_hd__o21ai_0 U14678 ( .A1(n25682), .A2(n27807), .B1(n25636), .Y(
        n24166) );
  sky130_fd_sc_hd__clkinv_1 U14710 ( .A(n27781), .Y(n27784) );
  sky130_fd_sc_hd__o21ai_0 U14737 ( .A1(n16543), .A2(n25230), .B1(n14873), .Y(
        n15085) );
  sky130_fd_sc_hd__o21ai_0 U14795 ( .A1(n26926), .A2(n22407), .B1(n22255), .Y(
        n22256) );
  sky130_fd_sc_hd__clkinv_1 U14815 ( .A(n23221), .Y(n23223) );
  sky130_fd_sc_hd__o21ai_0 U15065 ( .A1(n26761), .A2(n27342), .B1(n23289), .Y(
        n23317) );
  sky130_fd_sc_hd__o21ai_0 U15093 ( .A1(n16543), .A2(n28495), .B1(n13588), .Y(
        n13934) );
  sky130_fd_sc_hd__o21ai_0 U15117 ( .A1(n16088), .A2(n26285), .B1(n14488), .Y(
        n14578) );
  sky130_fd_sc_hd__clkinv_1 U15124 ( .A(n26379), .Y(n26384) );
  sky130_fd_sc_hd__o21ai_0 U15157 ( .A1(n16543), .A2(n28499), .B1(n15067), .Y(
        n15077) );
  sky130_fd_sc_hd__clkinv_1 U15166 ( .A(n15629), .Y(n15630) );
  sky130_fd_sc_hd__clkinv_1 U15192 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .Y(n17264) );
  sky130_fd_sc_hd__o21ai_0 U15202 ( .A1(n20164), .A2(n19969), .B1(n20225), .Y(
        n19990) );
  sky130_fd_sc_hd__nor2_1 U15217 ( .A(n13176), .B(n13175), .Y(n20459) );
  sky130_fd_sc_hd__o21ai_0 U15331 ( .A1(n19337), .A2(n19600), .B1(n19336), .Y(
        n19338) );
  sky130_fd_sc_hd__o21ai_0 U15335 ( .A1(j202_soc_core_intc_core_00_rg_ipr[83]), 
        .A2(n23369), .B1(n23338), .Y(n23340) );
  sky130_fd_sc_hd__o21ai_0 U15470 ( .A1(
        j202_soc_core_wbqspiflash_00_write_protect), .A2(
        j202_soc_core_wbqspiflash_00_spif_ctrl), .B1(n26535), .Y(n26537) );
  sky130_fd_sc_hd__o21ai_0 U15561 ( .A1(n16543), .A2(n28519), .B1(n14582), .Y(
        n14584) );
  sky130_fd_sc_hd__o21ai_0 U15563 ( .A1(n16543), .A2(n28446), .B1(n16542), .Y(
        n16547) );
  sky130_fd_sc_hd__nand2_1 U15633 ( .A(j202_soc_core_memory0_ram_dout0[44]), 
        .B(n21633), .Y(n20904) );
  sky130_fd_sc_hd__and2_0 U15644 ( .A(n21025), .B(n11637), .X(n11097) );
  sky130_fd_sc_hd__clkinv_1 U15679 ( .A(n21042), .Y(n17074) );
  sky130_fd_sc_hd__clkinv_1 U15718 ( .A(n23492), .Y(n13323) );
  sky130_fd_sc_hd__inv_2 U15768 ( .A(n11201), .Y(n16525) );
  sky130_fd_sc_hd__inv_2 U15812 ( .A(n30157), .Y(n12459) );
  sky130_fd_sc_hd__and2_0 U15820 ( .A(n11395), .B(n28417), .X(n11922) );
  sky130_fd_sc_hd__nand2_1 U15868 ( .A(n25349), .B(n22739), .Y(n15191) );
  sky130_fd_sc_hd__o21ai_0 U15896 ( .A1(n12435), .A2(n22210), .B1(n22209), .Y(
        n22212) );
  sky130_fd_sc_hd__clkinv_1 U15986 ( .A(n15489), .Y(n15491) );
  sky130_fd_sc_hd__buf_1 U16034 ( .A(n21684), .X(n12221) );
  sky130_fd_sc_hd__clkinv_1 U16045 ( .A(n22693), .Y(n22695) );
  sky130_fd_sc_hd__clkinv_1 U16060 ( .A(n22976), .Y(n21881) );
  sky130_fd_sc_hd__o21ai_0 U16247 ( .A1(n26926), .A2(n25928), .B1(n25927), .Y(
        n25929) );
  sky130_fd_sc_hd__clkinv_1 U16250 ( .A(n21189), .Y(n21191) );
  sky130_fd_sc_hd__clkinv_1 U16350 ( .A(n22953), .Y(n22955) );
  sky130_fd_sc_hd__clkinv_1 U16441 ( .A(n18683), .Y(n18685) );
  sky130_fd_sc_hd__nor2_1 U16467 ( .A(n19109), .B(n21235), .Y(n22207) );
  sky130_fd_sc_hd__clkinv_1 U16486 ( .A(n23482), .Y(n23490) );
  sky130_fd_sc_hd__or2_0 U16514 ( .A(n19239), .B(n19238), .X(n19241) );
  sky130_fd_sc_hd__o21ai_0 U16568 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[7]), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[3]), .B1(
        j202_soc_core_cmt_core_00_cks0[0]), .Y(n24014) );
  sky130_fd_sc_hd__o21ai_0 U16617 ( .A1(n15639), .A2(n15636), .B1(n15640), .Y(
        n15182) );
  sky130_fd_sc_hd__o21ai_0 U16715 ( .A1(n23972), .A2(n29581), .B1(n23971), .Y(
        n23975) );
  sky130_fd_sc_hd__clkinv_1 U16759 ( .A(n13837), .Y(n14053) );
  sky130_fd_sc_hd__o21ai_0 U16760 ( .A1(n24763), .A2(n24765), .B1(n22633), .Y(
        n22636) );
  sky130_fd_sc_hd__o21ai_0 U16773 ( .A1(n16526), .A2(n16525), .B1(n16524), .Y(
        n16530) );
  sky130_fd_sc_hd__clkinv_1 U16774 ( .A(n18138), .Y(n21939) );
  sky130_fd_sc_hd__inv_2 U16775 ( .A(n18832), .Y(n17357) );
  sky130_fd_sc_hd__clkinv_1 U16776 ( .A(n23384), .Y(n10981) );
  sky130_fd_sc_hd__a21boi_0 U16777 ( .A1(n25280), .A2(n25281), .B1_N(n12392), 
        .Y(n11414) );
  sky130_fd_sc_hd__o21ai_0 U16778 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[5]), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[9]), .B1(n23908), .Y(
        n23909) );
  sky130_fd_sc_hd__o21ai_0 U16779 ( .A1(n26411), .A2(n27788), .B1(n27787), .Y(
        n27823) );
  sky130_fd_sc_hd__o21ai_0 U16780 ( .A1(n16898), .A2(n17036), .B1(n16897), .Y(
        n16899) );
  sky130_fd_sc_hd__o21ai_0 U16781 ( .A1(n21749), .A2(n22735), .B1(n21748), .Y(
        n21750) );
  sky130_fd_sc_hd__nand2_1 U16782 ( .A(n20720), .B(n20719), .Y(n26165) );
  sky130_fd_sc_hd__o21ai_0 U16783 ( .A1(j202_soc_core_intc_core_00_rg_ipr[73]), 
        .A2(n27339), .B1(n23300), .Y(n23327) );
  sky130_fd_sc_hd__clkinv_1 U16784 ( .A(n21833), .Y(n21483) );
  sky130_fd_sc_hd__nand2_1 U16785 ( .A(n30184), .B(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n21025) );
  sky130_fd_sc_hd__clkinv_1 U16786 ( .A(j202_soc_core_memory0_ram_dout0[496]), 
        .Y(n30159) );
  sky130_fd_sc_hd__clkinv_1 U16787 ( .A(n11531), .Y(n11378) );
  sky130_fd_sc_hd__and4_1 U16788 ( .A(n20724), .B(n20723), .C(n20722), .D(
        n20721), .X(n30194) );
  sky130_fd_sc_hd__o21ai_0 U16789 ( .A1(n27339), .A2(n27341), .B1(n29830), .Y(
        n27340) );
  sky130_fd_sc_hd__o21ai_0 U16790 ( .A1(n27196), .A2(n27195), .B1(n27194), .Y(
        n27200) );
  sky130_fd_sc_hd__o21ai_0 U16791 ( .A1(j202_soc_core_qspi_wb_addr[2]), .A2(
        n27294), .B1(n27229), .Y(n23873) );
  sky130_fd_sc_hd__clkinv_1 U16792 ( .A(io_in[15]), .Y(n17093) );
  sky130_fd_sc_hd__o21ai_0 U16793 ( .A1(n11424), .A2(n27745), .B1(n11609), .Y(
        n27746) );
  sky130_fd_sc_hd__clkinv_1 U16794 ( .A(n11494), .Y(n11659) );
  sky130_fd_sc_hd__clkinv_1 U16795 ( .A(n11013), .Y(n11014) );
  sky130_fd_sc_hd__clkinv_1 U16796 ( .A(j202_soc_core_j22_cpu_regop_Rb__1_), 
        .Y(n13426) );
  sky130_fd_sc_hd__clkinv_1 U16797 ( .A(n12399), .Y(n28098) );
  sky130_fd_sc_hd__o21ai_0 U16798 ( .A1(n28987), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[12]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[12]), .Y(n28985) );
  sky130_fd_sc_hd__o21ai_0 U16799 ( .A1(n11123), .A2(n28518), .B1(n25867), .Y(
        n25888) );
  sky130_fd_sc_hd__o21ai_0 U16800 ( .A1(n22753), .A2(n22752), .B1(n22751), .Y(
        n22754) );
  sky130_fd_sc_hd__nand2_1 U16801 ( .A(n23476), .B(n24452), .Y(n25908) );
  sky130_fd_sc_hd__clkinv_1 U16802 ( .A(n24953), .Y(n26175) );
  sky130_fd_sc_hd__o21ai_0 U16803 ( .A1(n28842), .A2(n26585), .B1(n28843), .Y(
        n26586) );
  sky130_fd_sc_hd__o21ai_0 U16804 ( .A1(n22968), .A2(n22967), .B1(n22966), .Y(
        n22969) );
  sky130_fd_sc_hd__o21ai_0 U16805 ( .A1(n21271), .A2(n22967), .B1(n21272), .Y(
        n19305) );
  sky130_fd_sc_hd__and2_0 U16806 ( .A(n24147), .B(n24155), .X(n11101) );
  sky130_fd_sc_hd__nand2_1 U16807 ( .A(n18679), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .Y(n17359) );
  sky130_fd_sc_hd__xnor2_1 U16808 ( .A(n26206), .B(n25806), .Y(n26417) );
  sky130_fd_sc_hd__o21ai_0 U16809 ( .A1(n26411), .A2(n26416), .B1(n27787), .Y(
        n26446) );
  sky130_fd_sc_hd__o21ai_0 U16810 ( .A1(n25443), .A2(n25442), .B1(n25441), .Y(
        n25459) );
  sky130_fd_sc_hd__clkinv_1 U16811 ( .A(n21705), .Y(n11143) );
  sky130_fd_sc_hd__clkinv_1 U16812 ( .A(n12565), .Y(n12560) );
  sky130_fd_sc_hd__clkinv_1 U16813 ( .A(n24628), .Y(n11172) );
  sky130_fd_sc_hd__o21ai_0 U16814 ( .A1(n26926), .A2(n26061), .B1(n26060), .Y(
        n26062) );
  sky130_fd_sc_hd__o21ai_0 U16815 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[7]), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[3]), .B1(
        j202_soc_core_cmt_core_00_cks1[0]), .Y(n23913) );
  sky130_fd_sc_hd__o211a_2 U16816 ( .A1(n26323), .A2(n11186), .B1(n14787), 
        .C1(n14786), .X(n15091) );
  sky130_fd_sc_hd__o21ai_0 U16817 ( .A1(n21344), .A2(n22752), .B1(n21343), .Y(
        n22692) );
  sky130_fd_sc_hd__nand3_1 U16818 ( .A(n18793), .B(n18792), .C(n18791), .Y(
        n19852) );
  sky130_fd_sc_hd__clkinv_1 U16819 ( .A(n11625), .Y(n12884) );
  sky130_fd_sc_hd__and2_0 U16820 ( .A(n20416), .B(n20415), .X(n30200) );
  sky130_fd_sc_hd__o21ai_0 U16821 ( .A1(n26617), .A2(n28730), .B1(io_out[8]), 
        .Y(n26618) );
  sky130_fd_sc_hd__o21ai_0 U16822 ( .A1(
        j202_soc_core_wbqspiflash_00_last_status[5]), .A2(
        j202_soc_core_wbqspiflash_00_last_status[6]), .B1(n27239), .Y(n27283)
         );
  sky130_fd_sc_hd__o21ai_0 U16823 ( .A1(n28506), .A2(n22745), .B1(n15378), .Y(
        n15379) );
  sky130_fd_sc_hd__o21ai_0 U16824 ( .A1(n19928), .A2(n21819), .B1(n21919), .Y(
        n19933) );
  sky130_fd_sc_hd__clkinv_1 U16825 ( .A(n11623), .Y(n12883) );
  sky130_fd_sc_hd__nand3_1 U16826 ( .A(n30199), .B(n11645), .C(n11641), .Y(
        n30148) );
  sky130_fd_sc_hd__clkinv_1 U16827 ( .A(n27979), .Y(n24099) );
  sky130_fd_sc_hd__clkinv_1 U16828 ( .A(n28114), .Y(n28124) );
  sky130_fd_sc_hd__clkinv_1 U16829 ( .A(n10577), .Y(n13145) );
  sky130_fd_sc_hd__o21ai_0 U16830 ( .A1(n11478), .A2(n28048), .B1(n28047), .Y(
        n28049) );
  sky130_fd_sc_hd__o21ai_0 U16831 ( .A1(n29196), .A2(n29130), .B1(n29129), .Y(
        n29131) );
  sky130_fd_sc_hd__o21ai_0 U16832 ( .A1(n29196), .A2(n29139), .B1(n29138), .Y(
        n29140) );
  sky130_fd_sc_hd__o21ai_0 U16833 ( .A1(n29088), .A2(n28987), .B1(n28986), .Y(
        n28988) );
  sky130_fd_sc_hd__clkinv_1 U16834 ( .A(n12419), .Y(n30146) );
  sky130_fd_sc_hd__o21ai_0 U16835 ( .A1(n29029), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[18]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[18]), .Y(n29030) );
  sky130_fd_sc_hd__o21ai_0 U16836 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[23]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[23]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[23]), .Y(n26825) );
  sky130_fd_sc_hd__o21ai_0 U16837 ( .A1(j202_soc_core_j22_cpu_memop_MEM__1_), 
        .A2(n24300), .B1(n24299), .Y(n24301) );
  sky130_fd_sc_hd__o21ai_0 U16838 ( .A1(n23896), .A2(n23895), .B1(
        j202_soc_core_uart_TOP_rx_valid), .Y(n23897) );
  sky130_fd_sc_hd__o21ai_0 U16839 ( .A1(n27484), .A2(n26099), .B1(n26097), .Y(
        n26102) );
  sky130_fd_sc_hd__clkinv_1 U16840 ( .A(n28532), .Y(n28534) );
  sky130_fd_sc_hd__o21ai_0 U16841 ( .A1(n24931), .A2(n22745), .B1(n22744), .Y(
        n22746) );
  sky130_fd_sc_hd__o21ai_0 U16842 ( .A1(n25810), .A2(n25815), .B1(n25809), .Y(
        n25811) );
  sky130_fd_sc_hd__nand3_1 U16843 ( .A(n14208), .B(n13062), .C(n14207), .Y(
        n26945) );
  sky130_fd_sc_hd__o21ai_0 U16844 ( .A1(n25933), .A2(n22705), .B1(n21178), .Y(
        n21179) );
  sky130_fd_sc_hd__clkinv_1 U16845 ( .A(n28537), .Y(n24859) );
  sky130_fd_sc_hd__o21ai_0 U16846 ( .A1(n27188), .A2(n27187), .B1(n27186), .Y(
        n27189) );
  sky130_fd_sc_hd__o21ai_0 U16847 ( .A1(n26587), .A2(n28882), .B1(n26586), .Y(
        n26590) );
  sky130_fd_sc_hd__o21ai_0 U16848 ( .A1(n11146), .A2(n12234), .B1(n25769), .Y(
        n25771) );
  sky130_fd_sc_hd__o21ai_0 U16849 ( .A1(n22980), .A2(n22655), .B1(n22654), .Y(
        n22656) );
  sky130_fd_sc_hd__o21ai_0 U16850 ( .A1(n27540), .A2(n27537), .B1(n28583), .Y(
        n27531) );
  sky130_fd_sc_hd__o21ai_0 U16851 ( .A1(n27540), .A2(
        j202_soc_core_cmt_core_00_cnt1[0]), .B1(n28583), .Y(n27521) );
  sky130_fd_sc_hd__clkinv_1 U16852 ( .A(n12046), .Y(n12259) );
  sky130_fd_sc_hd__clkinv_1 U16853 ( .A(n25378), .Y(n23544) );
  sky130_fd_sc_hd__o21ai_0 U16854 ( .A1(n23018), .A2(n25224), .B1(n22099), .Y(
        n22100) );
  sky130_fd_sc_hd__nand2_1 U16855 ( .A(n30105), .B(n26413), .Y(n27588) );
  sky130_fd_sc_hd__clkinv_1 U16856 ( .A(n26240), .Y(n28509) );
  sky130_fd_sc_hd__and2_0 U16857 ( .A(n28091), .B(n25901), .X(n25903) );
  sky130_fd_sc_hd__inv_2 U16858 ( .A(n23616), .Y(n23617) );
  sky130_fd_sc_hd__clkinv_1 U16859 ( .A(n25372), .Y(n12397) );
  sky130_fd_sc_hd__o21ai_0 U16860 ( .A1(n23356), .A2(n27336), .B1(n30171), .Y(
        n23359) );
  sky130_fd_sc_hd__clkinv_1 U16861 ( .A(n23270), .Y(n23280) );
  sky130_fd_sc_hd__o21ai_0 U16862 ( .A1(n26157), .A2(n26392), .B1(n28109), .Y(
        n26395) );
  sky130_fd_sc_hd__clkinv_1 U16863 ( .A(n29547), .Y(n23048) );
  sky130_fd_sc_hd__o21a_1 U16864 ( .A1(n23516), .A2(n12351), .B1(n26159), .X(
        n28498) );
  sky130_fd_sc_hd__clkinv_1 U16865 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .Y(n29257) );
  sky130_fd_sc_hd__o21ai_0 U16866 ( .A1(n27210), .A2(n27207), .B1(n27206), .Y(
        n27216) );
  sky130_fd_sc_hd__o21ai_0 U16867 ( .A1(n26490), .A2(n27288), .B1(n27289), .Y(
        n27250) );
  sky130_fd_sc_hd__o21ai_0 U16868 ( .A1(n26613), .A2(n26612), .B1(n27223), .Y(
        n26614) );
  sky130_fd_sc_hd__o21ai_0 U16869 ( .A1(n28865), .A2(n26549), .B1(n26548), .Y(
        n26550) );
  sky130_fd_sc_hd__clkinv_1 U16870 ( .A(n11666), .Y(n27991) );
  sky130_fd_sc_hd__clkinv_1 U16871 ( .A(n27915), .Y(n25479) );
  sky130_fd_sc_hd__o21ai_0 U16872 ( .A1(n26309), .A2(n22745), .B1(n19100), .Y(
        n19101) );
  sky130_fd_sc_hd__o21ai_0 U16873 ( .A1(n23557), .A2(n27990), .B1(n23556), .Y(
        n13043) );
  sky130_fd_sc_hd__o21ai_0 U16874 ( .A1(n23420), .A2(n28072), .B1(n24109), .Y(
        n28403) );
  sky130_fd_sc_hd__nand2_1 U16875 ( .A(n22560), .B(n22559), .Y(n24469) );
  sky130_fd_sc_hd__clkinv_1 U16876 ( .A(j202_soc_core_intc_core_00_rg_ipr[45]), 
        .Y(n25790) );
  sky130_fd_sc_hd__and2_0 U16877 ( .A(n27894), .B(n24604), .X(n30201) );
  sky130_fd_sc_hd__clkinv_1 U16878 ( .A(j202_soc_core_intc_core_00_rg_ipr[17]), 
        .Y(n25746) );
  sky130_fd_sc_hd__and2_0 U16879 ( .A(n29270), .B(n28726), .X(n29265) );
  sky130_fd_sc_hd__o21ai_0 U16880 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[7]), .A2(n28293), .B1(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_0_), .Y(
        n27552) );
  sky130_fd_sc_hd__nand2_1 U16881 ( .A(n30062), .B(n22739), .Y(n15268) );
  sky130_fd_sc_hd__o21ai_0 U16882 ( .A1(n28984), .A2(n29061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[12]), .Y(n28991) );
  sky130_fd_sc_hd__o21ai_0 U16883 ( .A1(j202_soc_core_cmt_core_00_cnt1[13]), 
        .A2(n26082), .B1(n26089), .Y(n26083) );
  sky130_fd_sc_hd__o21ai_0 U16884 ( .A1(n27540), .A2(n24971), .B1(n28583), .Y(
        n27545) );
  sky130_fd_sc_hd__o21ai_0 U16885 ( .A1(n28246), .A2(n29061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[0]), .Y(n28247) );
  sky130_fd_sc_hd__o21ai_0 U16886 ( .A1(n28931), .A2(n29061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[4]), .Y(n28932) );
  sky130_fd_sc_hd__o21ai_0 U16887 ( .A1(n28959), .A2(n29061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[8]), .Y(n28960) );
  sky130_fd_sc_hd__o21ai_0 U16888 ( .A1(n29016), .A2(n29061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[16]), .Y(n29017) );
  sky130_fd_sc_hd__o21ai_0 U16889 ( .A1(n29088), .A2(
        j202_soc_core_qspi_wb_wdat[18]), .B1(n29039), .Y(n29031) );
  sky130_fd_sc_hd__o21ai_0 U16890 ( .A1(n29088), .A2(
        j202_soc_core_qspi_wb_wdat[21]), .B1(n29039), .Y(n26844) );
  sky130_fd_sc_hd__o21ai_0 U16891 ( .A1(n29054), .A2(n29061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[24]), .Y(n29055) );
  sky130_fd_sc_hd__o21ai_0 U16892 ( .A1(n29088), .A2(
        j202_soc_core_qspi_wb_wdat[27]), .B1(n29039), .Y(n26806) );
  sky130_fd_sc_hd__o21ai_0 U16893 ( .A1(n29062), .A2(n29061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[28]), .Y(n29063) );
  sky130_fd_sc_hd__o21ai_0 U16894 ( .A1(n29088), .A2(
        j202_soc_core_qspi_wb_wdat[30]), .B1(n29039), .Y(n26792) );
  sky130_fd_sc_hd__nand3_2 U16895 ( .A(n23624), .B(n23623), .C(n23622), .Y(
        n24297) );
  sky130_fd_sc_hd__clkinv_1 U16896 ( .A(j202_soc_core_intc_core_00_rg_ipr[29]), 
        .Y(n25490) );
  sky130_fd_sc_hd__o21ai_0 U16897 ( .A1(n29095), .A2(n29093), .B1(
        j202_soc_core_uart_TOP_dpll_state[1]), .Y(n29094) );
  sky130_fd_sc_hd__o21ai_0 U16898 ( .A1(j202_soc_core_uart_BRG_br_cnt[7]), 
        .A2(n29180), .B1(n29178), .Y(n29179) );
  sky130_fd_sc_hd__o21ai_0 U16909 ( .A1(j202_soc_core_uart_BRG_br_cnt[3]), 
        .A2(n28631), .B1(n28625), .Y(n28622) );
  sky130_fd_sc_hd__o21ai_0 U16918 ( .A1(n28620), .A2(
        j202_soc_core_uart_BRG_ps[6]), .B1(n28619), .Y(n28621) );
  sky130_fd_sc_hd__clkinv_1 U16920 ( .A(j202_soc_core_intc_core_00_rg_ipr[9]), 
        .Y(n25163) );
  sky130_fd_sc_hd__o21ai_0 U16931 ( .A1(n26103), .A2(n26102), .B1(
        j202_soc_core_cmt_core_00_cnt0[15]), .Y(n26109) );
  sky130_fd_sc_hd__o21ai_0 U16938 ( .A1(n29169), .A2(n25005), .B1(n27480), .Y(
        n27438) );
  sky130_fd_sc_hd__o21ai_0 U16947 ( .A1(n29169), .A2(n27483), .B1(n27480), .Y(
        n27488) );
  sky130_fd_sc_hd__o21ai_0 U16958 ( .A1(n27484), .A2(n25015), .B1(n25014), .Y(
        n25016) );
  sky130_fd_sc_hd__clkinv_1 U16965 ( .A(j202_soc_core_intc_core_00_rg_ipr[16]), 
        .Y(n26686) );
  sky130_fd_sc_hd__o21ai_0 U16967 ( .A1(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_0_), .A2(
        n29585), .B1(n27701), .Y(n27698) );
  sky130_fd_sc_hd__clkinv_1 U16974 ( .A(j202_soc_core_intc_core_00_rg_ipr[34]), 
        .Y(n26711) );
  sky130_fd_sc_hd__or2_0 U16975 ( .A(n25079), .B(n25097), .X(n28316) );
  sky130_fd_sc_hd__clkinv_1 U16982 ( .A(j202_soc_core_intc_core_00_rg_ipr[65]), 
        .Y(n28552) );
  sky130_fd_sc_hd__clkinv_1 U16983 ( .A(j202_soc_core_intc_core_00_rg_ipr[31]), 
        .Y(n26709) );
  sky130_fd_sc_hd__nand2_2 U16986 ( .A(n23624), .B(n13056), .Y(n12534) );
  sky130_fd_sc_hd__o21ai_0 U16993 ( .A1(n27228), .A2(n27227), .B1(
        j202_soc_core_wbqspiflash_00_state[4]), .Y(n27244) );
  sky130_fd_sc_hd__o21ai_0 U16995 ( .A1(n28669), .A2(n26510), .B1(n26519), .Y(
        n25336) );
  sky130_fd_sc_hd__a21boi_0 U17009 ( .A1(n25768), .A2(n22732), .B1_N(n22473), 
        .Y(n22520) );
  sky130_fd_sc_hd__and2_0 U17021 ( .A(n27119), .B(n23583), .X(n13078) );
  sky130_fd_sc_hd__and2_0 U17022 ( .A(n27119), .B(n23568), .X(n13080) );
  sky130_fd_sc_hd__and2_0 U17023 ( .A(n27119), .B(n23585), .X(n13077) );
  sky130_fd_sc_hd__o21ai_0 U17035 ( .A1(j202_soc_core_cmt_core_00_str0), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[0]), .B1(n28554), .Y(
        n28555) );
  sky130_fd_sc_hd__o21ai_0 U17039 ( .A1(n28576), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[6]), .B1(n28579), .Y(
        n28577) );
  sky130_fd_sc_hd__o21ai_0 U17040 ( .A1(j202_soc_core_cmt_core_00_str1), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[0]), .B1(n28567), .Y(
        n28565) );
  sky130_fd_sc_hd__o21ai_0 U17043 ( .A1(n27848), .A2(n24181), .B1(n24180), .Y(
        n24182) );
  sky130_fd_sc_hd__o21ai_0 U17047 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[7]), .A2(n28287), .B1(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_0_), .Y(
        n24731) );
  sky130_fd_sc_hd__clkinv_1 U17049 ( .A(n11770), .Y(n27649) );
  sky130_fd_sc_hd__clkinv_1 U17050 ( .A(n12184), .Y(n24779) );
  sky130_fd_sc_hd__clkinv_1 U17055 ( .A(n12034), .Y(n12035) );
  sky130_fd_sc_hd__clkinv_1 U17056 ( .A(n25466), .Y(n27642) );
  sky130_fd_sc_hd__o21ai_0 U17058 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .A2(n21836), .B1(n21770), 
        .Y(n21780) );
  sky130_fd_sc_hd__clkinv_1 U17102 ( .A(n27644), .Y(n27856) );
  sky130_fd_sc_hd__inv_2 U17118 ( .A(n24447), .Y(n27721) );
  sky130_fd_sc_hd__nand3_1 U17125 ( .A(n29551), .B(n25027), .C(n30026), .Y(
        n27950) );
  sky130_fd_sc_hd__clkinv_1 U17139 ( .A(n29752), .Y(n23945) );
  sky130_fd_sc_hd__o21ai_0 U17140 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .A2(n21825), .B1(n20922), 
        .Y(n20928) );
  sky130_fd_sc_hd__o21ai_0 U17141 ( .A1(n29183), .A2(n24031), .B1(n23855), .Y(
        n28691) );
  sky130_fd_sc_hd__o21ai_0 U17148 ( .A1(j202_soc_core_wbqspiflash_00_spi_hold), 
        .A2(n26569), .B1(n26664), .Y(n26572) );
  sky130_fd_sc_hd__o21ai_0 U17149 ( .A1(n26625), .A2(n26624), .B1(n26623), .Y(
        n26626) );
  sky130_fd_sc_hd__nand3_1 U17156 ( .A(n11622), .B(n20716), .C(n21919), .Y(
        n12880) );
  sky130_fd_sc_hd__o21ai_0 U17159 ( .A1(n24693), .A2(n24692), .B1(n28417), .Y(
        n24694) );
  sky130_fd_sc_hd__buf_1 U17160 ( .A(n23999), .X(n25478) );
  sky130_fd_sc_hd__o21ai_0 U17164 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[4]), .A2(n24522), .B1(
        n24524), .Y(n24523) );
  sky130_fd_sc_hd__inv_2 U17170 ( .A(n12386), .Y(n11156) );
  sky130_fd_sc_hd__inv_2 U17188 ( .A(n10993), .Y(n30095) );
  sky130_fd_sc_hd__o21ai_0 U17192 ( .A1(n27828), .A2(n28052), .B1(n24679), .Y(
        j202_soc_core_j22_cpu_ml_N152) );
  sky130_fd_sc_hd__o21ai_0 U17198 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .A2(n29133), .B1(n29132), 
        .Y(j202_soc_core_wbqspiflash_00_lldriver_N422) );
  sky130_fd_sc_hd__o21ai_0 U17199 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .A2(n29256), .B1(n29137), 
        .Y(j202_soc_core_wbqspiflash_00_lldriver_N419) );
  sky130_fd_sc_hd__o21ai_0 U17207 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .A2(n29195), .B1(n29141), 
        .Y(j202_soc_core_wbqspiflash_00_lldriver_N395) );
  sky130_fd_sc_hd__o21ai_0 U17215 ( .A1(n26087), .A2(n26086), .B1(n26085), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[14]) );
  sky130_fd_sc_hd__o21ai_0 U17216 ( .A1(n26988), .A2(n26987), .B1(n26986), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[9]) );
  sky130_fd_sc_hd__o21ai_0 U17217 ( .A1(n25375), .A2(n27770), .B1(n25374), .Y(
        j202_soc_core_j22_cpu_ml_maclj[21]) );
  sky130_fd_sc_hd__o21ai_0 U17228 ( .A1(n28258), .A2(n28257), .B1(n28256), .Y(
        j202_soc_core_ahb2apb_02_N128) );
  sky130_fd_sc_hd__o21ai_0 U17235 ( .A1(n28927), .A2(n28926), .B1(n28925), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N43) );
  sky130_fd_sc_hd__o21ai_0 U17249 ( .A1(n29019), .A2(n29018), .B1(n29017), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N56) );
  sky130_fd_sc_hd__o21ai_0 U17251 ( .A1(n29057), .A2(n29056), .B1(n29055), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N64) );
  sky130_fd_sc_hd__o21ai_0 U17252 ( .A1(n29012), .A2(n29011), .B1(n29010), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N55) );
  sky130_fd_sc_hd__or2_1 U17260 ( .A(n12083), .B(n12084), .X(n12082) );
  sky130_fd_sc_hd__nand2_1 U17285 ( .A(n24297), .B(n29830), .Y(n30053) );
  sky130_fd_sc_hd__o21ai_0 U17302 ( .A1(n29099), .A2(n29098), .B1(n12069), .Y(
        j202_soc_core_uart_TOP_N43) );
  sky130_fd_sc_hd__o21ai_0 U17304 ( .A1(j202_soc_core_uart_TOP_tx_bit_cnt[0]), 
        .A2(n28595), .B1(n29827), .Y(j202_soc_core_uart_TOP_N58) );
  sky130_fd_sc_hd__o21ai_0 U17307 ( .A1(n29096), .A2(n29095), .B1(n29094), .Y(
        n24) );
  sky130_fd_sc_hd__o21ai_0 U17308 ( .A1(n27958), .A2(n27955), .B1(n27953), .Y(
        n26) );
  sky130_fd_sc_hd__o21ai_0 U17318 ( .A1(n27994), .A2(n25484), .B1(n25483), .Y(
        n28) );
  sky130_fd_sc_hd__o21ai_0 U17322 ( .A1(n26105), .A2(n26101), .B1(n26100), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[14]) );
  sky130_fd_sc_hd__o21ai_0 U17332 ( .A1(n27928), .A2(n28291), .B1(n27927), .Y(
        n29) );
  sky130_fd_sc_hd__o21ai_0 U17338 ( .A1(n27932), .A2(n28545), .B1(n27931), .Y(
        n32) );
  sky130_fd_sc_hd__o21ai_0 U17339 ( .A1(n25732), .A2(n27624), .B1(n25731), .Y(
        n33) );
  sky130_fd_sc_hd__o21ai_0 U17362 ( .A1(n25319), .A2(n27624), .B1(n25318), .Y(
        n35) );
  sky130_fd_sc_hd__and2_0 U17387 ( .A(n25662), .B(n27856), .X(n13105) );
  sky130_fd_sc_hd__and2_0 U17401 ( .A(n25893), .B(n27856), .X(n13104) );
  sky130_fd_sc_hd__o21ai_0 U17403 ( .A1(n25307), .A2(n27770), .B1(n25374), .Y(
        j202_soc_core_j22_cpu_ml_maclj[17]) );
  sky130_fd_sc_hd__o21ai_0 U17405 ( .A1(n27096), .A2(n27624), .B1(n27095), .Y(
        n37) );
  sky130_fd_sc_hd__o21ai_0 U17418 ( .A1(n24851), .A2(n27770), .B1(n25374), .Y(
        j202_soc_core_j22_cpu_ml_maclj[16]) );
  sky130_fd_sc_hd__o21ai_0 U17422 ( .A1(n28209), .A2(n28277), .B1(n28205), .Y(
        n45) );
  sky130_fd_sc_hd__o21ai_0 U17427 ( .A1(n26879), .A2(n28545), .B1(n26878), .Y(
        n60) );
  sky130_fd_sc_hd__o21ai_0 U17433 ( .A1(n27994), .A2(n27651), .B1(n27650), .Y(
        n66) );
  sky130_fd_sc_hd__o21ai_0 U17448 ( .A1(n27994), .A2(n27867), .B1(n27866), .Y(
        n67) );
  sky130_fd_sc_hd__clkinv_1 U17449 ( .A(n12533), .Y(n29866) );
  sky130_fd_sc_hd__o21ai_0 U17450 ( .A1(n27648), .A2(n25970), .B1(n25969), .Y(
        j202_soc_core_j22_cpu_rf_N3360) );
  sky130_fd_sc_hd__o21ai_0 U17461 ( .A1(n26981), .A2(n25937), .B1(n25936), .Y(
        j202_soc_core_j22_cpu_rf_N3357) );
  sky130_fd_sc_hd__o21ai_0 U17463 ( .A1(n26981), .A2(n26980), .B1(n26979), .Y(
        j202_soc_core_j22_cpu_rf_N3354) );
  sky130_fd_sc_hd__o21ai_0 U17466 ( .A1(n27648), .A2(n12256), .B1(n24860), .Y(
        j202_soc_core_j22_cpu_rf_N3363) );
  sky130_fd_sc_hd__o21ai_0 U17485 ( .A1(n26981), .A2(n25763), .B1(n25723), .Y(
        j202_soc_core_j22_cpu_rf_N3364) );
  sky130_fd_sc_hd__o21ai_0 U17496 ( .A1(n27614), .A2(n27613), .B1(n27612), .Y(
        j202_soc_core_wbqspiflash_00_N698) );
  sky130_fd_sc_hd__o21ai_0 U17497 ( .A1(n29087), .A2(n28829), .B1(n28833), .Y(
        j202_soc_core_wbqspiflash_00_N613) );
  sky130_fd_sc_hd__o21ai_0 U17501 ( .A1(n29087), .A2(n29084), .B1(n29083), .Y(
        j202_soc_core_wbqspiflash_00_N606) );
  sky130_fd_sc_hd__o21ai_0 U17540 ( .A1(n27309), .A2(n28685), .B1(n27308), .Y(
        j202_soc_core_wbqspiflash_00_N740) );
  sky130_fd_sc_hd__o21ai_0 U17545 ( .A1(n27184), .A2(n27183), .B1(n27182), .Y(
        j202_soc_core_wbqspiflash_00_N592) );
  sky130_fd_sc_hd__o21ai_0 U17556 ( .A1(n27994), .A2(n27593), .B1(n27592), .Y(
        n71) );
  sky130_fd_sc_hd__o21ai_0 U17563 ( .A1(n25144), .A2(n27770), .B1(n25143), .Y(
        j202_soc_core_j22_cpu_ml_maclj[30]) );
  sky130_fd_sc_hd__o21ai_0 U17565 ( .A1(n25262), .A2(n27770), .B1(n25254), .Y(
        j202_soc_core_j22_cpu_ml_maclj[25]) );
  sky130_fd_sc_hd__o21ai_0 U17566 ( .A1(n24741), .A2(n28293), .B1(n24740), .Y(
        n72) );
  sky130_fd_sc_hd__o21ai_0 U17576 ( .A1(n27674), .A2(n28293), .B1(n27673), .Y(
        n77) );
  sky130_fd_sc_hd__o21ai_0 U17583 ( .A1(n28171), .A2(n28287), .B1(n28167), .Y(
        n83) );
  sky130_fd_sc_hd__o21ai_0 U17596 ( .A1(n28213), .A2(n28284), .B1(n28212), .Y(
        n87) );
  sky130_fd_sc_hd__o21ai_0 U17623 ( .A1(n28218), .A2(n28287), .B1(n28214), .Y(
        n89) );
  sky130_fd_sc_hd__o21ai_0 U17645 ( .A1(n27128), .A2(n27624), .B1(n27127), .Y(
        n93) );
  sky130_fd_sc_hd__o21ai_0 U17652 ( .A1(n27367), .A2(n27624), .B1(n27366), .Y(
        n94) );
  sky130_fd_sc_hd__o21ai_0 U17655 ( .A1(n28902), .A2(n28910), .B1(n28901), .Y(
        n103) );
  sky130_fd_sc_hd__o21ai_0 U17656 ( .A1(n27550), .A2(n28291), .B1(n27549), .Y(
        n113) );
  sky130_fd_sc_hd__o21ai_0 U17669 ( .A1(n26981), .A2(n24909), .B1(n24908), .Y(
        j202_soc_core_j22_cpu_rf_N3355) );
  sky130_fd_sc_hd__o21ai_0 U17705 ( .A1(n28042), .A2(n28423), .B1(n28422), .Y(
        j202_soc_core_j22_cpu_ml_N194) );
  sky130_fd_sc_hd__o21ai_0 U17716 ( .A1(n23749), .A2(n25290), .B1(n25283), .Y(
        j202_soc_core_j22_cpu_rf_N3298) );
  sky130_fd_sc_hd__o21ai_0 U17727 ( .A1(n12333), .A2(n28379), .B1(n24611), .Y(
        n10618) );
  sky130_fd_sc_hd__o21ai_0 U17743 ( .A1(n28285), .A2(n28284), .B1(n28283), .Y(
        n115) );
  sky130_fd_sc_hd__and2_0 U17744 ( .A(n27093), .B(n29565), .X(n12142) );
  sky130_fd_sc_hd__o21ai_0 U17752 ( .A1(n28583), .A2(n27543), .B1(n27542), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[5]) );
  sky130_fd_sc_hd__and2_0 U17757 ( .A(n12181), .B(n27856), .X(n13097) );
  sky130_fd_sc_hd__o21ai_0 U17771 ( .A1(n26875), .A2(n28291), .B1(n26874), .Y(
        n133) );
  sky130_fd_sc_hd__and2_0 U17772 ( .A(n10966), .B(n29554), .X(n29638) );
  sky130_fd_sc_hd__clkinv_1 U17786 ( .A(n24074), .Y(n11185) );
  sky130_fd_sc_hd__o21ai_0 U17788 ( .A1(n28983), .A2(n28982), .B1(n28981), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N51) );
  sky130_fd_sc_hd__o21ai_0 U17869 ( .A1(n26570), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B1(n26463), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N314) );
  sky130_fd_sc_hd__o21ai_0 U17870 ( .A1(n27307), .A2(n26579), .B1(n26578), .Y(
        j202_soc_core_wbqspiflash_00_N708) );
  sky130_fd_sc_hd__o21ai_0 U17871 ( .A1(n27264), .A2(n26528), .B1(n26527), .Y(
        n10543) );
  sky130_fd_sc_hd__o21ai_0 U17873 ( .A1(n27763), .A2(n28423), .B1(n27758), .Y(
        j202_soc_core_j22_cpu_ml_N195) );
  sky130_fd_sc_hd__and2_0 U17874 ( .A(n27093), .B(n29556), .X(n12148) );
  sky130_fd_sc_hd__clkinv_1 U17888 ( .A(n12842), .Y(n29496) );
  sky130_fd_sc_hd__o21ai_0 U17897 ( .A1(n29599), .A2(n28207), .B1(n28206), .Y(
        n137) );
  sky130_fd_sc_hd__clkinv_1 U17898 ( .A(gpio_en_o[1]), .Y(io_oeb[1]) );
  sky130_fd_sc_hd__clkinv_1 U17927 ( .A(gpio_en_o[10]), .Y(io_oeb[30]) );
  sky130_fd_sc_hd__and2_0 U17934 ( .A(n12857), .B(n12856), .X(n29883) );
  sky130_fd_sc_hd__and2_0 U17954 ( .A(n12854), .B(n12853), .X(n29884) );
  sky130_fd_sc_hd__buf_1 U17955 ( .A(n12323), .X(n29560) );
  sky130_fd_sc_hd__conb_1 U17998 ( .LO(n29885), .HI(
        j202_soc_core_ahb2aqu_00_N127) );
  sky130_fd_sc_hd__clkinv_1 U18019 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        user_irq[0]) );
  sky130_fd_sc_hd__clkinv_1 U18053 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        user_irq[1]) );
  sky130_fd_sc_hd__clkinv_1 U18073 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        user_irq[2]) );
  sky130_fd_sc_hd__clkinv_1 U18075 ( .A(n29885), .Y(io_oeb[5]) );
  sky130_fd_sc_hd__clkinv_1 U18086 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[6]) );
  sky130_fd_sc_hd__clkinv_1 U18092 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[8]) );
  sky130_fd_sc_hd__clkinv_1 U18094 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[9]) );
  sky130_fd_sc_hd__clkinv_1 U18115 ( .A(n29885), .Y(io_oeb[14]) );
  sky130_fd_sc_hd__clkinv_1 U18132 ( .A(n29885), .Y(io_oeb[15]) );
  sky130_fd_sc_hd__clkinv_1 U18198 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[16]) );
  sky130_fd_sc_hd__clkinv_1 U18200 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[17]) );
  sky130_fd_sc_hd__clkinv_1 U18203 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[18]) );
  sky130_fd_sc_hd__clkinv_1 U18204 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[19]) );
  sky130_fd_sc_hd__clkinv_1 U18205 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[20]) );
  sky130_fd_sc_hd__clkinv_1 U18211 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[21]) );
  sky130_fd_sc_hd__clkinv_1 U18234 ( .A(n29885), .Y(io_oeb[22]) );
  sky130_fd_sc_hd__clkinv_1 U18274 ( .A(n29885), .Y(io_oeb[23]) );
  sky130_fd_sc_hd__clkinv_1 U18288 ( .A(n29885), .Y(io_oeb[24]) );
  sky130_fd_sc_hd__clkinv_1 U18290 ( .A(n29885), .Y(io_oeb[25]) );
  sky130_fd_sc_hd__clkinv_1 U18305 ( .A(n29885), .Y(io_oeb[37]) );
  sky130_fd_sc_hd__clkinv_1 U18306 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[5]) );
  sky130_fd_sc_hd__clkinv_1 U18342 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[14]) );
  sky130_fd_sc_hd__clkinv_1 U18343 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[15]) );
  sky130_fd_sc_hd__clkinv_1 U18393 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[22]) );
  sky130_fd_sc_hd__clkinv_1 U18397 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[23]) );
  sky130_fd_sc_hd__clkinv_1 U18414 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[24]) );
  sky130_fd_sc_hd__clkinv_1 U18427 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[25]) );
  sky130_fd_sc_hd__clkinv_1 U18451 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[37]) );
  sky130_fd_sc_hd__clkinv_1 U18455 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[32]) );
  sky130_fd_sc_hd__clkinv_1 U18476 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[33]) );
  sky130_fd_sc_hd__clkinv_1 U18486 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[34]) );
  sky130_fd_sc_hd__clkinv_1 U18492 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[35]) );
  sky130_fd_sc_hd__clkinv_1 U18496 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[36]) );
  sky130_fd_sc_hd__clkinv_1 U18519 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[37]) );
  sky130_fd_sc_hd__clkinv_1 U18522 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[38]) );
  sky130_fd_sc_hd__clkinv_1 U18531 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[39]) );
  sky130_fd_sc_hd__clkinv_1 U18535 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[40]) );
  sky130_fd_sc_hd__clkinv_1 U18539 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[41]) );
  sky130_fd_sc_hd__clkinv_1 U18656 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[42]) );
  sky130_fd_sc_hd__clkinv_1 U18657 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[43]) );
  sky130_fd_sc_hd__clkinv_1 U18660 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[44]) );
  sky130_fd_sc_hd__clkinv_1 U18667 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[45]) );
  sky130_fd_sc_hd__clkinv_1 U18673 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[46]) );
  sky130_fd_sc_hd__clkinv_1 U18678 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[47]) );
  sky130_fd_sc_hd__clkinv_1 U18687 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[48]) );
  sky130_fd_sc_hd__clkinv_1 U18777 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[49]) );
  sky130_fd_sc_hd__clkinv_1 U18820 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[50]) );
  sky130_fd_sc_hd__clkinv_1 U18825 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[51]) );
  sky130_fd_sc_hd__clkinv_1 U18833 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[52]) );
  sky130_fd_sc_hd__clkinv_1 U18835 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[53]) );
  sky130_fd_sc_hd__clkinv_1 U18837 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[54]) );
  sky130_fd_sc_hd__clkinv_1 U18838 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[55]) );
  sky130_fd_sc_hd__clkinv_1 U18852 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[56]) );
  sky130_fd_sc_hd__clkinv_1 U18873 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[57]) );
  sky130_fd_sc_hd__clkinv_1 U18905 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[58]) );
  sky130_fd_sc_hd__clkinv_1 U18909 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[59]) );
  sky130_fd_sc_hd__clkinv_1 U18913 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[60]) );
  sky130_fd_sc_hd__clkinv_1 U18916 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[61]) );
  sky130_fd_sc_hd__clkinv_1 U18932 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[62]) );
  sky130_fd_sc_hd__clkinv_1 U18948 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[63]) );
  sky130_fd_sc_hd__clkinv_1 U18954 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[64]) );
  sky130_fd_sc_hd__clkinv_1 U18956 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[65]) );
  sky130_fd_sc_hd__clkinv_1 U18961 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[66]) );
  sky130_fd_sc_hd__clkinv_1 U18962 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[67]) );
  sky130_fd_sc_hd__clkinv_1 U18963 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[68]) );
  sky130_fd_sc_hd__clkinv_1 U18969 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[69]) );
  sky130_fd_sc_hd__clkinv_1 U18981 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[70]) );
  sky130_fd_sc_hd__clkinv_1 U18982 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[71]) );
  sky130_fd_sc_hd__clkinv_1 U18986 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[72]) );
  sky130_fd_sc_hd__clkinv_1 U18990 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[73]) );
  sky130_fd_sc_hd__clkinv_1 U19005 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[74]) );
  sky130_fd_sc_hd__clkinv_1 U19006 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[75]) );
  sky130_fd_sc_hd__clkinv_1 U19007 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[76]) );
  sky130_fd_sc_hd__clkinv_1 U19015 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[77]) );
  sky130_fd_sc_hd__clkinv_1 U19020 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[78]) );
  sky130_fd_sc_hd__clkinv_1 U19028 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[79]) );
  sky130_fd_sc_hd__clkinv_1 U19032 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[80]) );
  sky130_fd_sc_hd__clkinv_1 U19033 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[81]) );
  sky130_fd_sc_hd__clkinv_1 U19044 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[82]) );
  sky130_fd_sc_hd__clkinv_1 U19052 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[83]) );
  sky130_fd_sc_hd__clkinv_1 U19066 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[84]) );
  sky130_fd_sc_hd__clkinv_1 U19075 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[85]) );
  sky130_fd_sc_hd__clkinv_1 U19086 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[86]) );
  sky130_fd_sc_hd__clkinv_1 U19101 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[87]) );
  sky130_fd_sc_hd__clkinv_1 U19114 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[88]) );
  sky130_fd_sc_hd__clkinv_1 U19121 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[89]) );
  sky130_fd_sc_hd__clkinv_1 U19143 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[90]) );
  sky130_fd_sc_hd__clkinv_1 U19164 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[91]) );
  sky130_fd_sc_hd__clkinv_1 U19165 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[92]) );
  sky130_fd_sc_hd__clkinv_1 U19172 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[93]) );
  sky130_fd_sc_hd__clkinv_1 U19176 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[94]) );
  sky130_fd_sc_hd__clkinv_1 U19179 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[95]) );
  sky130_fd_sc_hd__clkinv_1 U19203 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[96]) );
  sky130_fd_sc_hd__clkinv_1 U19205 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[97]) );
  sky130_fd_sc_hd__clkinv_1 U19211 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[98]) );
  sky130_fd_sc_hd__clkinv_1 U19225 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[99]) );
  sky130_fd_sc_hd__clkinv_1 U19295 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[100]) );
  sky130_fd_sc_hd__clkinv_1 U19310 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[101]) );
  sky130_fd_sc_hd__clkinv_1 U19354 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[102]) );
  sky130_fd_sc_hd__clkinv_1 U19378 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[103]) );
  sky130_fd_sc_hd__clkinv_1 U19434 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[104]) );
  sky130_fd_sc_hd__clkinv_1 U19435 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[105]) );
  sky130_fd_sc_hd__clkinv_1 U19552 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[106]) );
  sky130_fd_sc_hd__clkinv_1 U19555 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[107]) );
  sky130_fd_sc_hd__clkinv_1 U19577 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[108]) );
  sky130_fd_sc_hd__clkinv_1 U19609 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[109]) );
  sky130_fd_sc_hd__clkinv_1 U19645 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[110]) );
  sky130_fd_sc_hd__clkinv_1 U19649 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[111]) );
  sky130_fd_sc_hd__clkinv_1 U19650 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[112]) );
  sky130_fd_sc_hd__clkinv_1 U19700 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[113]) );
  sky130_fd_sc_hd__clkinv_1 U19725 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[114]) );
  sky130_fd_sc_hd__clkinv_1 U19743 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[115]) );
  sky130_fd_sc_hd__clkinv_1 U19748 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[116]) );
  sky130_fd_sc_hd__clkinv_1 U19775 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[117]) );
  sky130_fd_sc_hd__clkinv_1 U19794 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[118]) );
  sky130_fd_sc_hd__clkinv_1 U19830 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[119]) );
  sky130_fd_sc_hd__clkinv_1 U19858 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[120]) );
  sky130_fd_sc_hd__clkinv_1 U19872 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[121]) );
  sky130_fd_sc_hd__clkinv_1 U19913 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[122]) );
  sky130_fd_sc_hd__clkinv_1 U19934 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[123]) );
  sky130_fd_sc_hd__clkinv_1 U19962 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[124]) );
  sky130_fd_sc_hd__clkinv_1 U19999 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[125]) );
  sky130_fd_sc_hd__clkinv_1 U20004 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[126]) );
  sky130_fd_sc_hd__clkinv_1 U20005 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[127]) );
  sky130_fd_sc_hd__or2_0 U20014 ( .A(n23209), .B(n23218), .X(n30010) );
  sky130_fd_sc_hd__buf_1 U20217 ( .A(n12362), .X(n11550) );
  sky130_fd_sc_hd__clkinv_1 U20231 ( .A(n12362), .Y(n11728) );
  sky130_fd_sc_hd__and2_0 U20317 ( .A(n27344), .B(n27343), .X(n30013) );
  sky130_fd_sc_hd__inv_2 U20326 ( .A(n27739), .Y(n12820) );
  sky130_fd_sc_hd__o21a_1 U20359 ( .A1(n24448), .A2(n24447), .B1(n12213), .X(
        n30014) );
  sky130_fd_sc_hd__and3_1 U20386 ( .A(n19114), .B(n19113), .C(n19112), .X(
        n30015) );
  sky130_fd_sc_hd__or2_0 U20387 ( .A(n18168), .B(n18167), .X(n30016) );
  sky130_fd_sc_hd__and2_0 U20473 ( .A(n13361), .B(n13359), .X(n30019) );
  sky130_fd_sc_hd__and4_1 U20488 ( .A(n20728), .B(n20727), .C(n20726), .D(
        n20725), .X(n30020) );
  sky130_fd_sc_hd__inv_2 U20499 ( .A(n23947), .Y(n23392) );
  sky130_fd_sc_hd__o21a_1 U20528 ( .A1(n24125), .A2(n11903), .B1(n11900), .X(
        n30021) );
  sky130_fd_sc_hd__clkinv_1 U20665 ( .A(j202_soc_core_j22_cpu_ml_bufa[8]), .Y(
        n11116) );
  sky130_fd_sc_hd__xnor2_1 U20682 ( .A(j202_soc_core_j22_cpu_ml_bufa[6]), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .Y(n30022) );
  sky130_fd_sc_hd__and4_1 U20871 ( .A(n13771), .B(n13770), .C(n13769), .D(
        n13768), .X(n30023) );
  sky130_fd_sc_hd__and4_1 U20876 ( .A(n14279), .B(n14278), .C(n14277), .D(
        n14276), .X(n30024) );
  sky130_fd_sc_hd__inv_2 U21131 ( .A(n12862), .Y(n24281) );
  sky130_fd_sc_hd__and2_0 U21268 ( .A(n12365), .B(n12465), .X(n30025) );
  sky130_fd_sc_hd__nand3_1 U21340 ( .A(n25594), .B(n26916), .C(n26329), .Y(
        n25564) );
  sky130_fd_sc_hd__and2_0 U21403 ( .A(n25029), .B(n25028), .X(n30026) );
  sky130_fd_sc_hd__clkinv_1 U21452 ( .A(j202_soc_core_intc_core_00_rg_ipr[18]), 
        .Y(n30173) );
  sky130_fd_sc_hd__and3_1 U21529 ( .A(n15253), .B(n15246), .C(n15252), .X(
        n30028) );
  sky130_fd_sc_hd__nand2_1 U21623 ( .A(n12940), .B(n15256), .Y(n11981) );
  sky130_fd_sc_hd__clkinv_1 U21649 ( .A(n29594), .Y(n30132) );
  sky130_fd_sc_hd__and4_1 U21713 ( .A(n12574), .B(n21042), .C(n29440), .D(
        n29437), .X(n30029) );
  sky130_fd_sc_hd__nand3_1 U21716 ( .A(n19260), .B(n19258), .C(n19259), .Y(
        n19262) );
  sky130_fd_sc_hd__and2_4 U21804 ( .A(n28062), .B(n12107), .X(n30030) );
  sky130_fd_sc_hd__clkinv_2 U21810 ( .A(n23433), .Y(n23443) );
  sky130_fd_sc_hd__nand2_1 U21919 ( .A(n23432), .B(n23431), .Y(n23433) );
  sky130_fd_sc_hd__nor2_1 U22003 ( .A(n30032), .B(n30031), .Y(n23431) );
  sky130_fd_sc_hd__nor2_1 U22058 ( .A(n23994), .B(n23430), .Y(n30031) );
  sky130_fd_sc_hd__nand2_1 U22164 ( .A(n23429), .B(n23428), .Y(n30032) );
  sky130_fd_sc_hd__xnor2_1 U22194 ( .A(n30033), .B(n18508), .Y(n18561) );
  sky130_fd_sc_hd__xnor2_1 U22203 ( .A(n18511), .B(n18509), .Y(n30033) );
  sky130_fd_sc_hd__xnor2_1 U22206 ( .A(n18397), .B(n30034), .Y(n18423) );
  sky130_fd_sc_hd__xnor2_1 U22209 ( .A(n18395), .B(n18396), .Y(n30034) );
  sky130_fd_sc_hd__xnor2_1 U22264 ( .A(n18427), .B(n18426), .Y(n13031) );
  sky130_fd_sc_hd__nand2_1 U22335 ( .A(n30036), .B(n30035), .Y(n18427) );
  sky130_fd_sc_hd__nand2_1 U22354 ( .A(n18397), .B(n18396), .Y(n30035) );
  sky130_fd_sc_hd__nand2_1 U22378 ( .A(n30038), .B(n30037), .Y(n18505) );
  sky130_fd_sc_hd__nand2_1 U22392 ( .A(n18502), .B(n30040), .Y(n30037) );
  sky130_fd_sc_hd__o21ai_1 U22403 ( .A1(n30040), .A2(n18502), .B1(n18501), .Y(
        n30038) );
  sky130_fd_sc_hd__xnor2_1 U22413 ( .A(n18501), .B(n30039), .Y(n18543) );
  sky130_fd_sc_hd__xnor2_1 U22419 ( .A(n30040), .B(n18502), .Y(n30039) );
  sky130_fd_sc_hd__o22ai_1 U22432 ( .A1(n18533), .A2(n18365), .B1(n18532), 
        .B2(n18530), .Y(n30040) );
  sky130_fd_sc_hd__xnor2_1 U22456 ( .A(n18467), .B(n11876), .Y(n30041) );
  sky130_fd_sc_hd__nand3_2 U22461 ( .A(n11540), .B(n11538), .C(n11537), .Y(
        n22257) );
  sky130_fd_sc_hd__nand2_1 U22486 ( .A(n22220), .B(n22228), .Y(n30042) );
  sky130_fd_sc_hd__nand3_1 U22503 ( .A(n22264), .B(n22405), .C(n22404), .Y(
        n22267) );
  sky130_fd_sc_hd__a21boi_1 U22520 ( .A1(n13012), .A2(n13001), .B1_N(n15629), 
        .Y(n12292) );
  sky130_fd_sc_hd__nand3_1 U22585 ( .A(n12016), .B(n12014), .C(n12019), .Y(
        n22005) );
  sky130_fd_sc_hd__nand3_2 U22617 ( .A(n11725), .B(n24119), .C(n24118), .Y(
        n10611) );
  sky130_fd_sc_hd__nand2_1 U22630 ( .A(n11469), .B(n28417), .Y(n11725) );
  sky130_fd_sc_hd__inv_1 U22673 ( .A(n30043), .Y(n23449) );
  sky130_fd_sc_hd__nor2_1 U22691 ( .A(n27737), .B(n11377), .Y(n30043) );
  sky130_fd_sc_hd__inv_1 U22727 ( .A(n30044), .Y(n11573) );
  sky130_fd_sc_hd__nand2_1 U22893 ( .A(n23390), .B(n28116), .Y(n30044) );
  sky130_fd_sc_hd__nand3_2 U23024 ( .A(n11646), .B(n23406), .C(n28133), .Y(
        n11941) );
  sky130_fd_sc_hd__nand2_2 U23103 ( .A(n11667), .B(n12022), .Y(n12016) );
  sky130_fd_sc_hd__o21a_1 U23140 ( .A1(n25393), .A2(n25397), .B1(n26919), .X(
        n25395) );
  sky130_fd_sc_hd__buf_2 U23144 ( .A(n29492), .X(n10966) );
  sky130_fd_sc_hd__inv_1 U23147 ( .A(n20893), .Y(n30045) );
  sky130_fd_sc_hd__inv_2 U23202 ( .A(n30045), .Y(n30046) );
  sky130_fd_sc_hd__inv_1 U23206 ( .A(n17076), .Y(n20893) );
  sky130_fd_sc_hd__inv_2 U23230 ( .A(n30161), .Y(n24435) );
  sky130_fd_sc_hd__inv_2 U23236 ( .A(n30160), .Y(n24496) );
  sky130_fd_sc_hd__nand2_1 U23238 ( .A(n13037), .B(n30137), .Y(n30047) );
  sky130_fd_sc_hd__nand2_1 U23250 ( .A(n13037), .B(n30137), .Y(n30048) );
  sky130_fd_sc_hd__nand3_2 U23268 ( .A(n30165), .B(n11708), .C(n11707), .Y(
        n13037) );
  sky130_fd_sc_hd__nand2_1 U23274 ( .A(n13037), .B(n30137), .Y(n13036) );
  sky130_fd_sc_hd__inv_2 U23314 ( .A(n19262), .Y(n30127) );
  sky130_fd_sc_hd__inv_1 U23319 ( .A(n30203), .Y(n12359) );
  sky130_fd_sc_hd__clkinv_4 U23324 ( .A(n11158), .Y(n11029) );
  sky130_fd_sc_hd__inv_1 U23355 ( .A(n25209), .Y(n26456) );
  sky130_fd_sc_hd__nand2_1 U23409 ( .A(n22437), .B(n19277), .Y(n30128) );
  sky130_fd_sc_hd__nand3_1 U23526 ( .A(n12270), .B(n21047), .C(n21316), .Y(
        n12268) );
  sky130_fd_sc_hd__xnor2_1 U23535 ( .A(n30049), .B(n12887), .Y(n23484) );
  sky130_fd_sc_hd__nand2_1 U23544 ( .A(n21760), .B(n22919), .Y(n30049) );
  sky130_fd_sc_hd__buf_4 U23602 ( .A(n24957), .X(n30071) );
  sky130_fd_sc_hd__nand2_2 U23631 ( .A(n25970), .B(n25968), .Y(n30050) );
  sky130_fd_sc_hd__nand2_2 U23641 ( .A(n25970), .B(n25968), .Y(n30051) );
  sky130_fd_sc_hd__nand2_2 U23661 ( .A(n25970), .B(n25968), .Y(n26895) );
  sky130_fd_sc_hd__nand3_1 U23670 ( .A(n11371), .B(n11516), .C(n20091), .Y(
        n26168) );
  sky130_fd_sc_hd__o211ai_1 U23681 ( .A1(n26926), .A2(n24950), .B1(n24949), 
        .C1(n24948), .Y(n24951) );
  sky130_fd_sc_hd__inv_4 U23709 ( .A(n12372), .Y(n11158) );
  sky130_fd_sc_hd__nand4_1 U23762 ( .A(n12581), .B(n12576), .C(n16385), .D(
        n12577), .Y(n30054) );
  sky130_fd_sc_hd__nand2_2 U23768 ( .A(n12843), .B(n29827), .Y(n30055) );
  sky130_fd_sc_hd__nand2_2 U23800 ( .A(n12843), .B(n29830), .Y(n30056) );
  sky130_fd_sc_hd__nand2_2 U23801 ( .A(n12843), .B(n29830), .Y(n12277) );
  sky130_fd_sc_hd__nand4_1 U23804 ( .A(n12999), .B(n12998), .C(n12997), .D(
        n12996), .Y(n30057) );
  sky130_fd_sc_hd__nand2_1 U23884 ( .A(n20586), .B(n20588), .Y(n30059) );
  sky130_fd_sc_hd__nand2_1 U23950 ( .A(n20586), .B(n20588), .Y(n24357) );
  sky130_fd_sc_hd__and2_1 U24067 ( .A(n20091), .B(n20092), .X(n12129) );
  sky130_fd_sc_hd__inv_1 U24109 ( .A(n28092), .Y(n30060) );
  sky130_fd_sc_hd__inv_2 U24121 ( .A(n30060), .Y(n30061) );
  sky130_fd_sc_hd__inv_2 U24214 ( .A(n11981), .Y(n30062) );
  sky130_fd_sc_hd__a22o_1 U24240 ( .A1(n27810), .A2(n26941), .B1(n27808), .B2(
        n24879), .X(n24881) );
  sky130_fd_sc_hd__a21oi_1 U24249 ( .A1(n17040), .A2(n16729), .B1(n16728), .Y(
        n16734) );
  sky130_fd_sc_hd__a21oi_1 U24312 ( .A1(n17040), .A2(n15488), .B1(n15487), .Y(
        n15493) );
  sky130_fd_sc_hd__a22o_1 U24393 ( .A1(n27810), .A2(n26064), .B1(n27808), .B2(
        n26941), .X(n25402) );
  sky130_fd_sc_hd__nand2b_1 U24415 ( .A_N(n26941), .B(n27023), .Y(n26218) );
  sky130_fd_sc_hd__nand2b_1 U24428 ( .A_N(n27023), .B(n26941), .Y(n26301) );
  sky130_fd_sc_hd__nand3_2 U24459 ( .A(n15191), .B(n15190), .C(n15189), .Y(
        n30063) );
  sky130_fd_sc_hd__nand2_1 U24527 ( .A(n12064), .B(n28027), .Y(n24400) );
  sky130_fd_sc_hd__a2bb2o_1 U24569 ( .A1_N(n25940), .A2_N(n25939), .B1(n25938), 
        .B2(n26168), .X(n26194) );
  sky130_fd_sc_hd__nand2_4 U24572 ( .A(n17460), .B(n17459), .Y(n18036) );
  sky130_fd_sc_hd__nand2_1 U24603 ( .A(n15090), .B(n15091), .Y(n30064) );
  sky130_fd_sc_hd__nand2_1 U24726 ( .A(n30178), .B(n30065), .Y(n29442) );
  sky130_fd_sc_hd__inv_2 U24854 ( .A(n30064), .Y(n30065) );
  sky130_fd_sc_hd__nand2_2 U24904 ( .A(n24281), .B(n22739), .Y(n12729) );
  sky130_fd_sc_hd__inv_1 U24906 ( .A(n30063), .Y(n16100) );
  sky130_fd_sc_hd__nand3_1 U24909 ( .A(n24179), .B(n23511), .C(n23510), .Y(
        n23512) );
  sky130_fd_sc_hd__inv_1 U24910 ( .A(j202_soc_core_j22_cpu_ml_bufa[18]), .Y(
        n17408) );
  sky130_fd_sc_hd__and2_1 U24928 ( .A(n26191), .B(n26189), .X(n24156) );
  sky130_fd_sc_hd__nand3_1 U24960 ( .A(n10959), .B(n17089), .C(n17088), .Y(
        n17091) );
  sky130_fd_sc_hd__nand2_1 U25008 ( .A(n17091), .B(n13074), .Y(n30066) );
  sky130_fd_sc_hd__nand2_1 U25009 ( .A(n17091), .B(n13074), .Y(n20897) );
  sky130_fd_sc_hd__inv_2 U25023 ( .A(n12275), .Y(n30067) );
  sky130_fd_sc_hd__inv_2 U25024 ( .A(n12275), .Y(n30068) );
  sky130_fd_sc_hd__inv_2 U25027 ( .A(n12275), .Y(n13109) );
  sky130_fd_sc_hd__nand4_1 U25028 ( .A(n26945), .B(n12028), .C(n26175), .D(
        n11549), .Y(n24954) );
  sky130_fd_sc_hd__nor2_4 U25043 ( .A(n21048), .B(n12268), .Y(n29492) );
  sky130_fd_sc_hd__inv_1 U25089 ( .A(n12265), .Y(n30069) );
  sky130_fd_sc_hd__inv_2 U25192 ( .A(n30069), .Y(n30070) );
  sky130_fd_sc_hd__nand2_2 U25204 ( .A(n21187), .B(n21188), .Y(n12265) );
  sky130_fd_sc_hd__nand3_2 U25223 ( .A(n12846), .B(n12845), .C(n16887), .Y(
        n26158) );
  sky130_fd_sc_hd__nand3_1 U25305 ( .A(n30162), .B(n12724), .C(n17078), .Y(
        n30157) );
  sky130_fd_sc_hd__clkinv_1 U25326 ( .A(n17072), .Y(n10959) );
  sky130_fd_sc_hd__clkinv_1 U25424 ( .A(n29442), .Y(n12293) );
  sky130_fd_sc_hd__clkinv_2 U25428 ( .A(n12265), .Y(n12271) );
  sky130_fd_sc_hd__buf_2 U25455 ( .A(n12265), .X(n12466) );
  sky130_fd_sc_hd__nor2_1 U25486 ( .A(n23976), .B(n12272), .Y(n23977) );
  sky130_fd_sc_hd__nor2_1 U25498 ( .A(n23965), .B(n12272), .Y(n23966) );
  sky130_fd_sc_hd__nor2_2 U25587 ( .A(n23967), .B(n12272), .Y(n23968) );
  sky130_fd_sc_hd__nand2_1 U25638 ( .A(n21187), .B(n21188), .Y(n25024) );
  sky130_fd_sc_hd__inv_2 U25656 ( .A(n23968), .Y(n29822) );
  sky130_fd_sc_hd__nand3_4 U25675 ( .A(n13360), .B(n30019), .C(n13358), .Y(
        n24912) );
  sky130_fd_sc_hd__nand3_2 U25711 ( .A(n13429), .B(n11094), .C(n18860), .Y(
        n22983) );
  sky130_fd_sc_hd__buf_2 U25716 ( .A(n11388), .X(n26191) );
  sky130_fd_sc_hd__bufinv_8 U25737 ( .A(n11158), .Y(n30097) );
  sky130_fd_sc_hd__bufinv_8 U25742 ( .A(n11158), .Y(n30098) );
  sky130_fd_sc_hd__nand3_1 U25778 ( .A(n22008), .B(n10981), .C(n23421), .Y(
        n24547) );
  sky130_fd_sc_hd__a21oi_1 U25825 ( .A1(n11729), .A2(n11731), .B1(n11730), .Y(
        n11597) );
  sky130_fd_sc_hd__nand2_2 U25857 ( .A(n24606), .B(n23955), .Y(n30072) );
  sky130_fd_sc_hd__nand2_1 U25896 ( .A(n24606), .B(n23955), .Y(n23610) );
  sky130_fd_sc_hd__nand2_1 U25897 ( .A(n11175), .B(n11719), .Y(n30073) );
  sky130_fd_sc_hd__and2_1 U25905 ( .A(n23615), .B(n24406), .X(n24407) );
  sky130_fd_sc_hd__nand4_1 U25976 ( .A(n23515), .B(n23513), .C(n23512), .D(
        n23514), .Y(n30076) );
  sky130_fd_sc_hd__nand4_1 U26033 ( .A(n23515), .B(n23513), .C(n23512), .D(
        n23514), .Y(n30077) );
  sky130_fd_sc_hd__nand4_1 U26053 ( .A(n23515), .B(n23513), .C(n23512), .D(
        n23514), .Y(n26159) );
  sky130_fd_sc_hd__inv_1 U26063 ( .A(n27742), .Y(n30078) );
  sky130_fd_sc_hd__buf_2 U26121 ( .A(n24560), .X(n12228) );
  sky130_fd_sc_hd__dlygate4sd1_1 U26130 ( .A(n24612), .X(n12333) );
  sky130_fd_sc_hd__clkinv_1 U26164 ( .A(n25660), .Y(n28505) );
  sky130_fd_sc_hd__nand2_1 U26208 ( .A(n23408), .B(n24559), .Y(n30079) );
  sky130_fd_sc_hd__nand2_1 U26271 ( .A(n23408), .B(n24559), .Y(n24562) );
  sky130_fd_sc_hd__nand2_1 U26304 ( .A(n23402), .B(n11175), .Y(n12922) );
  sky130_fd_sc_hd__nand2_2 U26348 ( .A(n18338), .B(n18337), .Y(n30080) );
  sky130_fd_sc_hd__or2_1 U26357 ( .A(n18474), .B(n17586), .X(n30081) );
  sky130_fd_sc_hd__nand2_1 U26393 ( .A(n30081), .B(n30082), .Y(n17584) );
  sky130_fd_sc_hd__nand2_2 U26474 ( .A(n18338), .B(n18337), .Y(n11553) );
  sky130_fd_sc_hd__fah_1 U26494 ( .A(n17584), .B(n17585), .CI(n17583), .COUT(
        n17617), .SUM(n17591) );
  sky130_fd_sc_hd__nor2_1 U26576 ( .A(n12321), .B(n11579), .Y(n23427) );
  sky130_fd_sc_hd__nand2_1 U26618 ( .A(n12217), .B(n23955), .Y(n12874) );
  sky130_fd_sc_hd__nand2_1 U26623 ( .A(n28266), .B(n12942), .Y(n30083) );
  sky130_fd_sc_hd__nand2_1 U26646 ( .A(n28266), .B(n12942), .Y(n24684) );
  sky130_fd_sc_hd__o21ai_0 U26675 ( .A1(n27855), .A2(n28477), .B1(n25289), .Y(
        j202_soc_core_j22_cpu_rf_N323) );
  sky130_fd_sc_hd__clkbuf_1 U26717 ( .A(n25372), .X(n30084) );
  sky130_fd_sc_hd__nand3_2 U26881 ( .A(n11485), .B(n12398), .C(n25369), .Y(
        n25372) );
  sky130_fd_sc_hd__and3_1 U26913 ( .A(n21838), .B(n21839), .C(n21840), .X(
        n30085) );
  sky130_fd_sc_hd__buf_8 U26941 ( .A(n11137), .X(n10986) );
  sky130_fd_sc_hd__buf_8 U26960 ( .A(n11137), .X(n10985) );
  sky130_fd_sc_hd__buf_8 U27007 ( .A(n11137), .X(n10988) );
  sky130_fd_sc_hd__buf_8 U27048 ( .A(n11137), .X(n11121) );
  sky130_fd_sc_hd__buf_8 U27068 ( .A(n11137), .X(n11162) );
  sky130_fd_sc_hd__buf_8 U27206 ( .A(n11137), .X(n29820) );
  sky130_fd_sc_hd__clkinv_4 U27226 ( .A(n27584), .Y(n27583) );
  sky130_fd_sc_hd__inv_1 U27292 ( .A(n11358), .Y(n30086) );
  sky130_fd_sc_hd__nor2_2 U27308 ( .A(n28098), .B(n28393), .Y(n28345) );
  sky130_fd_sc_hd__o21ai_0 U27323 ( .A1(n24832), .A2(n25632), .B1(n25631), .Y(
        j202_soc_core_j22_cpu_rf_N3295) );
  sky130_fd_sc_hd__and2_1 U27348 ( .A(n25630), .B(n27856), .X(n12132) );
  sky130_fd_sc_hd__nand2_2 U27360 ( .A(n28151), .B(n28417), .Y(n28083) );
  sky130_fd_sc_hd__nand2_2 U27385 ( .A(n25932), .B(n25931), .Y(n25935) );
  sky130_fd_sc_hd__o21a_1 U27431 ( .A1(n27648), .A2(n25722), .B1(n25721), .X(
        n25723) );
  sky130_fd_sc_hd__nand4bb_1 U27447 ( .A_N(n28152), .B_N(n28151), .C(n28150), 
        .D(n28149), .Y(n28153) );
  sky130_fd_sc_hd__xnor2_1 U27487 ( .A(n18363), .B(n25761), .Y(n17795) );
  sky130_fd_sc_hd__buf_6 U27524 ( .A(j202_soc_core_j22_cpu_ml_bufa[17]), .X(
        n25761) );
  sky130_fd_sc_hd__inv_2 U27567 ( .A(n11569), .Y(n30087) );
  sky130_fd_sc_hd__nand2_2 U27577 ( .A(n30126), .B(n23411), .Y(n11569) );
  sky130_fd_sc_hd__nor2_1 U27636 ( .A(n12362), .B(n11579), .Y(n11578) );
  sky130_fd_sc_hd__nand2b_1 U27641 ( .A_N(n12238), .B(n11395), .Y(n11726) );
  sky130_fd_sc_hd__clkbuf_1 U27669 ( .A(n12318), .X(n11384) );
  sky130_fd_sc_hd__nand2_2 U27844 ( .A(n19542), .B(n19543), .Y(n30088) );
  sky130_fd_sc_hd__nand2_2 U27848 ( .A(n19542), .B(n19543), .Y(n29589) );
  sky130_fd_sc_hd__o22a_1 U27880 ( .A1(n30088), .A2(n23947), .B1(n23422), .B2(
        n24563), .X(n30089) );
  sky130_fd_sc_hd__inv_2 U27937 ( .A(n10990), .Y(n30090) );
  sky130_fd_sc_hd__clkinv_2 U27956 ( .A(n30090), .Y(n30091) );
  sky130_fd_sc_hd__inv_2 U28038 ( .A(n10991), .Y(n30092) );
  sky130_fd_sc_hd__clkinv_2 U28041 ( .A(n30092), .Y(n30093) );
  sky130_fd_sc_hd__inv_1 U28152 ( .A(n11133), .Y(n10991) );
  sky130_fd_sc_hd__clkinv_2 U28155 ( .A(n11135), .Y(n11075) );
  sky130_fd_sc_hd__clkinv_2 U28180 ( .A(n11135), .Y(n11032) );
  sky130_fd_sc_hd__clkinv_2 U28181 ( .A(n11135), .Y(n11026) );
  sky130_fd_sc_hd__clkinv_2 U28185 ( .A(n11135), .Y(n11078) );
  sky130_fd_sc_hd__clkinv_2 U28187 ( .A(n11135), .Y(n11077) );
  sky130_fd_sc_hd__clkinv_2 U28388 ( .A(n11135), .Y(n11076) );
  sky130_fd_sc_hd__buf_8 U28404 ( .A(n12370), .X(n11120) );
  sky130_fd_sc_hd__inv_4 U28405 ( .A(n11087), .Y(n30094) );
  sky130_fd_sc_hd__inv_4 U28428 ( .A(n11087), .Y(n11034) );
  sky130_fd_sc_hd__inv_12 U28445 ( .A(n23980), .Y(n11087) );
  sky130_fd_sc_hd__clkinv_4 U28456 ( .A(n30095), .Y(n30096) );
  sky130_fd_sc_hd__clkinv_2 U28461 ( .A(n11157), .Y(n11039) );
  sky130_fd_sc_hd__clkinv_2 U28486 ( .A(n11154), .Y(n11025) );
  sky130_fd_sc_hd__clkinv_4 U28496 ( .A(n30099), .Y(n30100) );
  sky130_fd_sc_hd__inv_1 U28504 ( .A(n30101), .Y(n17320) );
  sky130_fd_sc_hd__nand2_1 U28512 ( .A(n30103), .B(n30102), .Y(n30101) );
  sky130_fd_sc_hd__nand2_1 U28517 ( .A(j202_soc_core_memory0_ram_dout0[423]), 
        .B(n12156), .Y(n30102) );
  sky130_fd_sc_hd__nand2_1 U28522 ( .A(j202_soc_core_memory0_ram_dout0[359]), 
        .B(n21495), .Y(n30103) );
  sky130_fd_sc_hd__inv_2 U28543 ( .A(n30138), .Y(n30137) );
  sky130_fd_sc_hd__nand4_1 U28547 ( .A(n12005), .B(n12003), .C(n12004), .D(
        n30104), .Y(n12394) );
  sky130_fd_sc_hd__nand2_1 U28552 ( .A(j202_soc_core_memory0_ram_dout0[312]), 
        .B(n21503), .Y(n30104) );
  sky130_fd_sc_hd__nand2_1 U28575 ( .A(n11388), .B(n11205), .Y(n21694) );
  sky130_fd_sc_hd__nand3_2 U28586 ( .A(n12792), .B(n14727), .C(n12783), .Y(
        n11388) );
  sky130_fd_sc_hd__nand2_1 U28669 ( .A(n26412), .B(n26416), .Y(n30105) );
  sky130_fd_sc_hd__nor2_1 U28670 ( .A(n12422), .B(n12659), .Y(n12297) );
  sky130_fd_sc_hd__nand4_1 U28809 ( .A(n11791), .B(n11792), .C(n11793), .D(
        n16180), .Y(n12422) );
  sky130_fd_sc_hd__o21ai_2 U28873 ( .A1(n18670), .A2(n19106), .B1(n18669), .Y(
        n18671) );
  sky130_fd_sc_hd__nand3_2 U28926 ( .A(n20884), .B(n12969), .C(n12968), .Y(
        n23549) );
  sky130_fd_sc_hd__nand2_1 U28951 ( .A(n12967), .B(n12123), .Y(n12968) );
  sky130_fd_sc_hd__xnor2_1 U29002 ( .A(n18461), .B(n30106), .Y(n18450) );
  sky130_fd_sc_hd__xnor2_1 U29004 ( .A(n18462), .B(n18460), .Y(n30106) );
  sky130_fd_sc_hd__xnor2_1 U29036 ( .A(n18641), .B(n18642), .Y(n18463) );
  sky130_fd_sc_hd__nand2_1 U29058 ( .A(n30108), .B(n30107), .Y(n18641) );
  sky130_fd_sc_hd__nand2_1 U29060 ( .A(n18461), .B(n18462), .Y(n30107) );
  sky130_fd_sc_hd__o21ai_1 U29095 ( .A1(n18462), .A2(n18461), .B1(n18460), .Y(
        n30108) );
  sky130_fd_sc_hd__nand2_1 U29143 ( .A(n23408), .B(n12844), .Y(n28089) );
  sky130_fd_sc_hd__nand3_2 U29145 ( .A(n27122), .B(n30127), .C(n30015), .Y(
        n19263) );
  sky130_fd_sc_hd__xor2_1 U29195 ( .A(n17756), .B(n30109), .X(n17817) );
  sky130_fd_sc_hd__xor2_1 U29273 ( .A(n17757), .B(n17755), .X(n30109) );
  sky130_fd_sc_hd__xnor2_1 U29285 ( .A(n17753), .B(n30110), .Y(n17818) );
  sky130_fd_sc_hd__xnor2_1 U29292 ( .A(n17754), .B(n17752), .Y(n30110) );
  sky130_fd_sc_hd__nand2_1 U29444 ( .A(n30112), .B(n30111), .Y(n17835) );
  sky130_fd_sc_hd__nand2_1 U29543 ( .A(n30116), .B(n30119), .Y(n30111) );
  sky130_fd_sc_hd__nand2_1 U29586 ( .A(n17527), .B(n30113), .Y(n30112) );
  sky130_fd_sc_hd__nand2b_1 U29589 ( .A_N(n30116), .B(n30114), .Y(n30113) );
  sky130_fd_sc_hd__xnor2_1 U29621 ( .A(n30115), .B(n17527), .Y(n17813) );
  sky130_fd_sc_hd__xnor2_1 U29624 ( .A(n30119), .B(n30116), .Y(n30115) );
  sky130_fd_sc_hd__nand2_1 U29636 ( .A(n30118), .B(n30117), .Y(n30116) );
  sky130_fd_sc_hd__nand2_1 U29699 ( .A(n17756), .B(n17757), .Y(n30117) );
  sky130_fd_sc_hd__o21ai_1 U29744 ( .A1(n17757), .A2(n17756), .B1(n17755), .Y(
        n30118) );
  sky130_fd_sc_hd__nand2_1 U29750 ( .A(n30121), .B(n30120), .Y(n30119) );
  sky130_fd_sc_hd__nand2_1 U29777 ( .A(n17753), .B(n17754), .Y(n30120) );
  sky130_fd_sc_hd__o21ai_1 U29791 ( .A1(n17754), .A2(n17753), .B1(n17752), .Y(
        n30121) );
  sky130_fd_sc_hd__inv_1 U29950 ( .A(n30128), .Y(n22688) );
  sky130_fd_sc_hd__nand2_1 U29959 ( .A(n30123), .B(n30122), .Y(n18299) );
  sky130_fd_sc_hd__nand2_1 U29977 ( .A(n18069), .B(n18070), .Y(n30122) );
  sky130_fd_sc_hd__o21ai_1 U30002 ( .A1(n18070), .A2(n18069), .B1(n18068), .Y(
        n30123) );
  sky130_fd_sc_hd__xnor2_1 U30038 ( .A(n18068), .B(n30124), .Y(n18302) );
  sky130_fd_sc_hd__xnor2_1 U30061 ( .A(n18070), .B(n18069), .Y(n30124) );
  sky130_fd_sc_hd__nand4_1 U30069 ( .A(n24546), .B(n24660), .C(n12776), .D(
        n12583), .Y(n24408) );
  sky130_fd_sc_hd__nor2_4 U30070 ( .A(n28091), .B(n11706), .Y(n12583) );
  sky130_fd_sc_hd__nand3_1 U30071 ( .A(n12971), .B(n30194), .C(n30020), .Y(
        n12970) );
  sky130_fd_sc_hd__nor2_1 U30073 ( .A(n12977), .B(n11381), .Y(n12971) );
  sky130_fd_sc_hd__inv_2 U30136 ( .A(n30125), .Y(n12286) );
  sky130_fd_sc_hd__nand2_1 U30146 ( .A(n12205), .B(n29587), .Y(n30125) );
  sky130_fd_sc_hd__nand2_1 U30162 ( .A(n24615), .B(n24614), .Y(n12923) );
  sky130_fd_sc_hd__nand3_2 U30275 ( .A(n24405), .B(n29593), .C(n29587), .Y(
        n24615) );
  sky130_fd_sc_hd__nand4_1 U30424 ( .A(n10975), .B(n11571), .C(n11572), .D(
        n11573), .Y(n30126) );
  sky130_fd_sc_hd__nand4_1 U30454 ( .A(n11586), .B(n11584), .C(n11107), .D(
        n30129), .Y(n11583) );
  sky130_fd_sc_hd__inv_2 U30468 ( .A(n30130), .Y(n30129) );
  sky130_fd_sc_hd__nand2_1 U30509 ( .A(n20416), .B(n20424), .Y(n30130) );
  sky130_fd_sc_hd__nand2_1 U30600 ( .A(n30131), .B(n11807), .Y(n12742) );
  sky130_fd_sc_hd__nor2_1 U30629 ( .A(n11798), .B(n11803), .Y(n30131) );
  sky130_fd_sc_hd__nor2_1 U30633 ( .A(n23549), .B(n30132), .Y(n11535) );
  sky130_fd_sc_hd__xor2_1 U30640 ( .A(n12484), .B(n30133), .X(n17912) );
  sky130_fd_sc_hd__xnor2_1 U30670 ( .A(n17800), .B(n17801), .Y(n30133) );
  sky130_fd_sc_hd__xnor2_1 U30673 ( .A(n18305), .B(n30134), .Y(n18308) );
  sky130_fd_sc_hd__xnor2_1 U30697 ( .A(n18307), .B(n18306), .Y(n30134) );
  sky130_fd_sc_hd__xnor2_1 U30705 ( .A(n18312), .B(n18313), .Y(n30143) );
  sky130_fd_sc_hd__nand2_1 U30827 ( .A(n30136), .B(n30135), .Y(n18312) );
  sky130_fd_sc_hd__nand2_1 U30829 ( .A(n18306), .B(n18307), .Y(n30135) );
  sky130_fd_sc_hd__nand2_1 U30833 ( .A(n19692), .B(n21919), .Y(n30138) );
  sky130_fd_sc_hd__clkbuf_1 U30929 ( .A(n27899), .X(n30139) );
  sky130_fd_sc_hd__o22ai_1 U30930 ( .A1(n30142), .A2(n30141), .B1(n30140), 
        .B2(n30144), .Y(n18320) );
  sky130_fd_sc_hd__nor2_1 U30936 ( .A(n18313), .B(n18312), .Y(n30140) );
  sky130_fd_sc_hd__inv_1 U30974 ( .A(n18312), .Y(n30141) );
  sky130_fd_sc_hd__inv_2 U31012 ( .A(n18313), .Y(n30142) );
  sky130_fd_sc_hd__xor2_1 U31068 ( .A(n30144), .B(n30143), .X(n18317) );
  sky130_fd_sc_hd__xor2_1 U31120 ( .A(n17999), .B(n12166), .X(n30144) );
  sky130_fd_sc_hd__clkbuf_1 U31121 ( .A(j202_soc_core_j22_cpu_ml_bufa[10]), 
        .X(n30145) );
  sky130_fd_sc_hd__nand3_2 U31132 ( .A(n25564), .B(n11104), .C(n30146), .Y(
        n25383) );
  sky130_fd_sc_hd__inv_2 U31140 ( .A(n30147), .Y(n11098) );
  sky130_fd_sc_hd__nand2_1 U31154 ( .A(n27898), .B(n28089), .Y(n30147) );
  sky130_fd_sc_hd__inv_2 U31172 ( .A(n30148), .Y(n19542) );
  sky130_fd_sc_hd__nand3_2 U31180 ( .A(n12461), .B(n20893), .C(n11208), .Y(
        n30152) );
  sky130_fd_sc_hd__nand2_1 U31244 ( .A(n29546), .B(n12271), .Y(n29761) );
  sky130_fd_sc_hd__nand2_2 U31252 ( .A(n30150), .B(n11980), .Y(n21187) );
  sky130_fd_sc_hd__inv_1 U31283 ( .A(n30151), .Y(n11103) );
  sky130_fd_sc_hd__nand4_1 U31287 ( .A(n17065), .B(n17064), .C(n17063), .D(
        n17062), .Y(n30151) );
  sky130_fd_sc_hd__inv_2 U31296 ( .A(n30152), .Y(n11978) );
  sky130_fd_sc_hd__nand4_1 U31300 ( .A(n12579), .B(n11884), .C(n12578), .D(
        n30153), .Y(n11883) );
  sky130_fd_sc_hd__nand2_1 U31301 ( .A(j202_soc_core_memory0_ram_dout0[447]), 
        .B(n12156), .Y(n30153) );
  sky130_fd_sc_hd__nand2_1 U31350 ( .A(n30155), .B(n30154), .Y(n18217) );
  sky130_fd_sc_hd__nand2_1 U31442 ( .A(n18167), .B(n18168), .Y(n30154) );
  sky130_fd_sc_hd__nand2_1 U31472 ( .A(n18166), .B(n30016), .Y(n30155) );
  sky130_fd_sc_hd__xnor2_1 U31518 ( .A(n30156), .B(n18166), .Y(n18165) );
  sky130_fd_sc_hd__xnor2_1 U31553 ( .A(n18168), .B(n18167), .Y(n30156) );
  sky130_fd_sc_hd__inv_2 U31579 ( .A(n12293), .Y(n30163) );
  sky130_fd_sc_hd__xnor2_1 U31588 ( .A(n16092), .B(n30158), .Y(n25473) );
  sky130_fd_sc_hd__nand2_1 U31596 ( .A(n29514), .B(n12214), .Y(n30160) );
  sky130_fd_sc_hd__nand2_1 U31612 ( .A(n29499), .B(n12214), .Y(n30161) );
  sky130_fd_sc_hd__a21oi_2 U31618 ( .A1(n21029), .A2(n15071), .B1(n15070), .Y(
        n15381) );
  sky130_fd_sc_hd__nand2_1 U31624 ( .A(n12729), .B(n12727), .Y(n30164) );
  sky130_fd_sc_hd__nor2_1 U31625 ( .A(n11758), .B(n11753), .Y(n30165) );
  sky130_fd_sc_hd__inv_1 U31642 ( .A(n17236), .Y(n12769) );
  sky130_fd_sc_hd__nand4_1 U31645 ( .A(n17233), .B(n17234), .C(n17235), .D(
        n17232), .Y(n17236) );
  sky130_fd_sc_hd__inv_6 U31652 ( .A(n25135), .Y(n26897) );
  sky130_fd_sc_hd__nand2_2 U31798 ( .A(n25133), .B(n25132), .Y(n25135) );
  sky130_fd_sc_hd__nand4_1 U31813 ( .A(n20916), .B(n20915), .C(n20911), .D(
        n20910), .Y(n11915) );
  sky130_fd_sc_hd__nand2_1 U31834 ( .A(j202_soc_core_memory0_ram_dout0[396]), 
        .B(n21496), .Y(n20916) );
  sky130_fd_sc_hd__nand2_1 U31848 ( .A(n30166), .B(n28417), .Y(n27913) );
  sky130_fd_sc_hd__nand4_1 U31888 ( .A(n27908), .B(n12345), .C(n12251), .D(
        n27909), .Y(n30166) );
  sky130_fd_sc_hd__nand4_1 U31893 ( .A(n11739), .B(n11531), .C(n12801), .D(
        n12800), .Y(n11363) );
  sky130_fd_sc_hd__nand2_1 U31970 ( .A(j202_soc_core_memory0_ram_dout0[333]), 
        .B(n21490), .Y(n11739) );
  sky130_fd_sc_hd__nand2_1 U31976 ( .A(n11913), .B(n19934), .Y(n20886) );
  sky130_fd_sc_hd__nand2_1 U32035 ( .A(n30167), .B(n11400), .Y(n11399) );
  sky130_fd_sc_hd__nand4_1 U32080 ( .A(n22115), .B(n12210), .C(n22116), .D(
        n22117), .Y(n30167) );
  sky130_fd_sc_hd__a21oi_1 U32137 ( .A1(n22147), .A2(n26426), .B1(n22146), .Y(
        n25145) );
  sky130_fd_sc_hd__inv_2 U32188 ( .A(n30179), .Y(n30197) );
  sky130_fd_sc_hd__nand3_2 U32189 ( .A(n11661), .B(n20886), .C(n20888), .Y(
        n12273) );
  sky130_fd_sc_hd__a21oi_1 U32195 ( .A1(n27345), .A2(n30013), .B1(n29583), .Y(
        n27346) );
  sky130_fd_sc_hd__nand2_2 U32203 ( .A(n23377), .B(n23376), .Y(n27345) );
  sky130_fd_sc_hd__o21ai_1 U32219 ( .A1(n23352), .A2(n27322), .B1(n30168), .Y(
        n23257) );
  sky130_fd_sc_hd__nand2_1 U32228 ( .A(n27322), .B(n23357), .Y(n30168) );
  sky130_fd_sc_hd__buf_2 U32258 ( .A(n27319), .X(n30169) );
  sky130_fd_sc_hd__nand3_1 U32270 ( .A(n23363), .B(n23362), .C(n30170), .Y(
        n23371) );
  sky130_fd_sc_hd__inv_1 U32272 ( .A(n23364), .Y(n30170) );
  sky130_fd_sc_hd__nand2_1 U32299 ( .A(n27336), .B(n23353), .Y(n30171) );
  sky130_fd_sc_hd__clkinv_1 U32409 ( .A(n11666), .Y(n30188) );
  sky130_fd_sc_hd__o21ai_1 U32449 ( .A1(n30173), .A2(n27321), .B1(n30172), .Y(
        n23209) );
  sky130_fd_sc_hd__nand2_1 U32459 ( .A(n27321), .B(
        j202_soc_core_intc_core_00_rg_ipr[22]), .Y(n30172) );
  sky130_fd_sc_hd__o21ai_1 U32469 ( .A1(n11518), .A2(n17236), .B1(n12109), .Y(
        n12017) );
  sky130_fd_sc_hd__nor2_4 U32474 ( .A(n27743), .B(n24564), .Y(n28130) );
  sky130_fd_sc_hd__nand2_4 U32475 ( .A(n29589), .B(n12318), .Y(n27743) );
  sky130_fd_sc_hd__nor2_1 U32511 ( .A(n12252), .B(n12286), .Y(n11735) );
  sky130_fd_sc_hd__nor2_2 U32529 ( .A(n11724), .B(n24097), .Y(n12252) );
  sky130_fd_sc_hd__inv_1 U32602 ( .A(n30174), .Y(n20416) );
  sky130_fd_sc_hd__nand2_1 U32627 ( .A(n11602), .B(n11603), .Y(n30174) );
  sky130_fd_sc_hd__inv_2 U32655 ( .A(n27742), .Y(n24634) );
  sky130_fd_sc_hd__nand2_2 U32677 ( .A(n11621), .B(n23392), .Y(n27742) );
  sky130_fd_sc_hd__nor2_1 U32687 ( .A(n30177), .B(n30175), .Y(n30199) );
  sky130_fd_sc_hd__nor2b_1 U32704 ( .B_N(n30176), .A(n21933), .Y(n30175) );
  sky130_fd_sc_hd__inv_2 U32708 ( .A(n11203), .Y(n30176) );
  sky130_fd_sc_hd__nand2_1 U32743 ( .A(n11638), .B(n19540), .Y(n30177) );
  sky130_fd_sc_hd__nand3_1 U32772 ( .A(n16570), .B(n16572), .C(n16571), .Y(
        n17072) );
  sky130_fd_sc_hd__nand2_1 U32785 ( .A(n11388), .B(n22739), .Y(n30178) );
  sky130_fd_sc_hd__nand2_1 U32790 ( .A(n29519), .B(n12214), .Y(n30179) );
  sky130_fd_sc_hd__nand2_1 U32813 ( .A(n12214), .B(n29504), .Y(n30180) );
  sky130_fd_sc_hd__nand2_1 U32887 ( .A(n12214), .B(n29510), .Y(n30181) );
  sky130_fd_sc_hd__nand2_1 U32891 ( .A(n12214), .B(n29509), .Y(n30182) );
  sky130_fd_sc_hd__nand2_1 U32923 ( .A(n12214), .B(n29523), .Y(n30183) );
  sky130_fd_sc_hd__clkinv_2 U32938 ( .A(j202_soc_core_memory0_ram_dout0[497]), 
        .Y(n30184) );
  sky130_fd_sc_hd__inv_2 U32946 ( .A(n30185), .Y(n23624) );
  sky130_fd_sc_hd__nand2_1 U32985 ( .A(n11439), .B(n12269), .Y(n30185) );
  sky130_fd_sc_hd__xor2_1 U32987 ( .A(n16195), .B(n16196), .X(n27067) );
  sky130_fd_sc_hd__inv_2 U32992 ( .A(n14775), .Y(n16077) );
  sky130_fd_sc_hd__nand2_1 U32994 ( .A(n11853), .B(n29524), .Y(n30186) );
  sky130_fd_sc_hd__inv_2 U33025 ( .A(n12038), .Y(n24617) );
  sky130_fd_sc_hd__nand3_2 U33031 ( .A(n11741), .B(n28092), .C(n23597), .Y(
        n12038) );
  sky130_fd_sc_hd__nand4_2 U33045 ( .A(n25148), .B(n12323), .C(n30188), .D(
        n30187), .Y(n23396) );
  sky130_fd_sc_hd__inv_1 U33207 ( .A(n22005), .Y(n30187) );
  sky130_fd_sc_hd__o31a_1 U33213 ( .A1(n27717), .A2(n23969), .A3(n22452), .B1(
        n28109), .X(n30189) );
  sky130_fd_sc_hd__nor2_4 U33222 ( .A(n13393), .B(n13408), .Y(n13566) );
  sky130_fd_sc_hd__nand2_2 U33236 ( .A(n17409), .B(n17729), .Y(n17410) );
  sky130_fd_sc_hd__nor2_4 U33262 ( .A(n13401), .B(n13403), .Y(n13820) );
  sky130_fd_sc_hd__nand2_2 U33267 ( .A(n13477), .B(
        j202_soc_core_j22_cpu_regop_Ra__0_), .Y(n13294) );
  sky130_fd_sc_hd__clkinv_1 U33450 ( .A(n13836), .Y(n14052) );
  sky130_fd_sc_hd__or2_0 U33487 ( .A(n13415), .B(n13414), .X(n30190) );
  sky130_fd_sc_hd__clkinv_1 U33516 ( .A(n27786), .Y(n26411) );
  sky130_fd_sc_hd__and4_1 U33521 ( .A(n11736), .B(n11739), .C(n11738), .D(
        n11737), .X(n30198) );
  sky130_fd_sc_hd__clkinv_1 U33545 ( .A(n22232), .Y(n12557) );
  sky130_fd_sc_hd__clkinv_1 U33561 ( .A(n21917), .Y(n11203) );
  sky130_fd_sc_hd__clkinv_1 U33562 ( .A(n25397), .Y(n27785) );
  sky130_fd_sc_hd__clkinv_1 U33563 ( .A(j202_soc_core_j22_cpu_ma_M_address[1]), 
        .Y(n23511) );
  sky130_fd_sc_hd__inv_2 U33565 ( .A(n24593), .Y(n23384) );
  sky130_fd_sc_hd__buf_4 U33585 ( .A(n22003), .X(n11395) );
  sky130_fd_sc_hd__nand3_2 U33590 ( .A(n15268), .B(n15267), .C(n15266), .Y(
        n12299) );
  sky130_fd_sc_hd__o21ba_4 U33591 ( .A1(n12341), .A2(n27355), .B1_N(n27159), 
        .X(n24805) );
  sky130_fd_sc_hd__clkinv_2 U33602 ( .A(n25662), .Y(n27385) );
  sky130_fd_sc_hd__clkinv_2 U33604 ( .A(n25662), .Y(n12258) );
  sky130_fd_sc_hd__clkinv_2 U33623 ( .A(n25313), .Y(n12057) );
  sky130_fd_sc_hd__clkinv_2 U33624 ( .A(n25313), .Y(n12056) );
  sky130_fd_sc_hd__and3_1 U33628 ( .A(n27734), .B(n27733), .C(n27732), .X(
        n30202) );
  sky130_fd_sc_hd__clkinv_2 U33636 ( .A(n22007), .Y(n23387) );
  sky130_fd_sc_hd__buf_2 U33645 ( .A(n12278), .X(n24128) );
  sky130_fd_sc_hd__and2_2 U33646 ( .A(n23999), .B(n29828), .X(n30203) );
  sky130_fd_sc_hd__probe_p_8 U33649 ( .A(n12375), .X(n10987) );
  sky130_fd_sc_hd__inv_4 U33681 ( .A(n11085), .Y(n11060) );
  sky130_fd_sc_hd__clkinv_4 U33683 ( .A(n11060), .Y(n11022) );
  sky130_fd_sc_hd__inv_6 U33687 ( .A(n11060), .Y(n11063) );
endmodule

