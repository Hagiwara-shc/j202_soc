// SPDX-FileCopyrightText: 2022 SH CONSULTING K.K.
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

module j202_soc_core_wrapper ( wb_clk_i, wb_rst_i, wbs_stb_i, wbs_cyc_i, 
        wbs_we_i, wbs_sel_i, wbs_dat_i, wbs_adr_i, wbs_ack_o, wbs_dat_o, 
        la_data_in, la_data_out, la_oenb, io_in, io_out, io_oeb, analog_io, 
        user_clock2, user_irq );
  input [3:0] wbs_sel_i;
  input [31:0] wbs_dat_i;
  input [31:0] wbs_adr_i;
  output [31:0] wbs_dat_o;
  input [127:0] la_data_in;
  output [127:0] la_data_out;
  input [127:0] la_oenb;
  input [37:0] io_in;
  output [37:0] io_out;
  output [37:0] io_oeb;
  inout [28:0] analog_io;
  output [2:0] user_irq;
  input wb_clk_i, wb_rst_i, wbs_stb_i, wbs_cyc_i, wbs_we_i, user_clock2;
  output wbs_ack_o;
  wire   n3, n4, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n220, n230, n240, n250, n260, n270, n280, n290, n300, n310, n320,
         n330, n340, n350, n360, n370, n380, n390, n400, n410, n420, n430,
         n440, n450, n460, n470, j202_soc_core_qspi_wb_cyc,
         j202_soc_core_qspi_wb_ack, j202_soc_core_aquc_STB_,
         j202_soc_core_aquc_ADR__0_, j202_soc_core_aquc_ADR__2_,
         j202_soc_core_aquc_ADR__3_, j202_soc_core_aquc_ADR__4_,
         j202_soc_core_aquc_ADR__5_, j202_soc_core_aquc_ADR__6_,
         j202_soc_core_aquc_ADR__7_, j202_soc_core_aquc_SEL__0_,
         j202_soc_core_aquc_SEL__2_, j202_soc_core_aquc_SEL__3_,
         j202_soc_core_aquc_WE_, j202_soc_core_aquc_CE__0_,
         j202_soc_core_aquc_CE__1_, j202_soc_core_bldc_int,
         j202_soc_core_qspi_int, j202_soc_core_ahbcs_6__HREADY_,
         j202_soc_core_intr_vec__0_, j202_soc_core_intr_vec__1_,
         j202_soc_core_intr_vec__2_, j202_soc_core_intr_vec__3_,
         j202_soc_core_intr_vec__4_, j202_soc_core_intr_vec__6_,
         j202_soc_core_intr_level__0_, j202_soc_core_intr_level__1_,
         j202_soc_core_intr_level__2_, j202_soc_core_intr_level__3_,
         j202_soc_core_intr_level__4_, j202_soc_core_intr_req_,
         j202_soc_core_rst, j202_soc_core_rst1, j202_soc_core_rst0,
         j202_soc_core_j22_cpu_regop_M_Wm__0_,
         j202_soc_core_j22_cpu_regop_M_Wm__1_,
         j202_soc_core_j22_cpu_regop_M_Wm__2_,
         j202_soc_core_j22_cpu_regop_M_Wm__3_,
         j202_soc_core_j22_cpu_regop_M_Rn__0_,
         j202_soc_core_j22_cpu_regop_M_Rn__1_,
         j202_soc_core_j22_cpu_regop_M_Rn__2_,
         j202_soc_core_j22_cpu_regop_M_Rn__3_,
         j202_soc_core_j22_cpu_regop_Wm__0_,
         j202_soc_core_j22_cpu_regop_Wm__1_,
         j202_soc_core_j22_cpu_regop_Wm__2_,
         j202_soc_core_j22_cpu_regop_Wm__3_,
         j202_soc_core_j22_cpu_regop_We__1_,
         j202_soc_core_j22_cpu_regop_We__2_,
         j202_soc_core_j22_cpu_regop_We__3_,
         j202_soc_core_j22_cpu_regop_Rs__0_,
         j202_soc_core_j22_cpu_regop_Rs__1_,
         j202_soc_core_j22_cpu_regop_Rb__1_,
         j202_soc_core_j22_cpu_regop_Ra__0_,
         j202_soc_core_j22_cpu_regop_Ra__1_,
         j202_soc_core_j22_cpu_regop_imm__7_,
         j202_soc_core_j22_cpu_regop_Rn__0_,
         j202_soc_core_j22_cpu_regop_Rn__1_,
         j202_soc_core_j22_cpu_regop_Rn__2_,
         j202_soc_core_j22_cpu_regop_Rn__3_, j202_soc_core_j22_cpu_ifetch,
         j202_soc_core_j22_cpu_memop_Ma__0_,
         j202_soc_core_j22_cpu_memop_Ma__1_,
         j202_soc_core_j22_cpu_memop_MEM__0_,
         j202_soc_core_j22_cpu_memop_MEM__1_,
         j202_soc_core_j22_cpu_memop_MEM__2_,
         j202_soc_core_j22_cpu_memop_MEM__3_, j202_soc_core_j22_cpu_pc_hold,
         j202_soc_core_j22_cpu_istall, j202_soc_core_j22_cpu_intack,
         j202_soc_core_j22_cpu_N8, j202_soc_core_j22_cpu_rte4,
         j202_soc_core_j22_cpu_rfuo_sr__t_, j202_soc_core_j22_cpu_rfuo_sr__s_,
         j202_soc_core_j22_cpu_rfuo_sr__i__0_,
         j202_soc_core_j22_cpu_rfuo_sr__i__1_,
         j202_soc_core_j22_cpu_rfuo_sr__i__2_,
         j202_soc_core_j22_cpu_rfuo_sr__i__3_,
         j202_soc_core_j22_cpu_rfuo_sr__q_, j202_soc_core_j22_cpu_rfuo_sr__m_,
         j202_soc_core_j22_cpu_ifetchl, j202_soc_core_j22_cpu_id_opn_v_,
         j202_soc_core_j22_cpu_id_opn_inst__0_,
         j202_soc_core_j22_cpu_id_opn_inst__1_,
         j202_soc_core_j22_cpu_id_opn_inst__2_,
         j202_soc_core_j22_cpu_id_opn_inst__3_,
         j202_soc_core_j22_cpu_id_opn_inst__4_,
         j202_soc_core_j22_cpu_id_opn_inst__5_,
         j202_soc_core_j22_cpu_id_opn_inst__6_,
         j202_soc_core_j22_cpu_id_opn_inst__7_,
         j202_soc_core_j22_cpu_id_opn_inst__8_,
         j202_soc_core_j22_cpu_id_opn_inst__9_,
         j202_soc_core_j22_cpu_id_opn_inst__10_,
         j202_soc_core_j22_cpu_id_opn_inst__11_,
         j202_soc_core_j22_cpu_id_opn_inst__12_,
         j202_soc_core_j22_cpu_id_opn_inst__13_,
         j202_soc_core_j22_cpu_id_opn_inst__14_,
         j202_soc_core_j22_cpu_id_opn_inst__15_,
         j202_soc_core_j22_cpu_id_op2_v_,
         j202_soc_core_j22_cpu_id_op2_inst__0_,
         j202_soc_core_j22_cpu_id_op2_inst__1_,
         j202_soc_core_j22_cpu_id_op2_inst__2_,
         j202_soc_core_j22_cpu_id_op2_inst__3_,
         j202_soc_core_j22_cpu_id_op2_inst__4_,
         j202_soc_core_j22_cpu_id_op2_inst__5_,
         j202_soc_core_j22_cpu_id_op2_inst__6_,
         j202_soc_core_j22_cpu_id_op2_inst__7_,
         j202_soc_core_j22_cpu_id_op2_inst__8_,
         j202_soc_core_j22_cpu_id_op2_inst__9_,
         j202_soc_core_j22_cpu_id_op2_inst__10_,
         j202_soc_core_j22_cpu_id_op2_inst__11_,
         j202_soc_core_j22_cpu_id_op2_inst__12_,
         j202_soc_core_j22_cpu_id_op2_inst__13_,
         j202_soc_core_j22_cpu_id_op2_inst__14_,
         j202_soc_core_j22_cpu_id_op2_inst__15_,
         j202_soc_core_j22_cpu_id_idec_N959,
         j202_soc_core_j22_cpu_id_idec_N958,
         j202_soc_core_j22_cpu_id_idec_N957,
         j202_soc_core_j22_cpu_id_idec_N956,
         j202_soc_core_j22_cpu_id_idec_N937,
         j202_soc_core_j22_cpu_id_idec_N917,
         j202_soc_core_j22_cpu_id_idec_N900,
         j202_soc_core_j22_cpu_id_idec_N894,
         j202_soc_core_j22_cpu_id_idec_N857,
         j202_soc_core_j22_cpu_id_idec_N822, j202_soc_core_j22_cpu_rf_N3392,
         j202_soc_core_j22_cpu_rf_N3391, j202_soc_core_j22_cpu_rf_N3390,
         j202_soc_core_j22_cpu_rf_N3388, j202_soc_core_j22_cpu_rf_N3386,
         j202_soc_core_j22_cpu_rf_N3379, j202_soc_core_j22_cpu_rf_N3378,
         j202_soc_core_j22_cpu_rf_N3377, j202_soc_core_j22_cpu_rf_N3376,
         j202_soc_core_j22_cpu_rf_N3375, j202_soc_core_j22_cpu_rf_N3374,
         j202_soc_core_j22_cpu_rf_N3373, j202_soc_core_j22_cpu_rf_N3372,
         j202_soc_core_j22_cpu_rf_N3371, j202_soc_core_j22_cpu_rf_N3370,
         j202_soc_core_j22_cpu_rf_N3369, j202_soc_core_j22_cpu_rf_N3368,
         j202_soc_core_j22_cpu_rf_N3367, j202_soc_core_j22_cpu_rf_N3366,
         j202_soc_core_j22_cpu_rf_N3365, j202_soc_core_j22_cpu_rf_N3364,
         j202_soc_core_j22_cpu_rf_N3363, j202_soc_core_j22_cpu_rf_N3361,
         j202_soc_core_j22_cpu_rf_N3360, j202_soc_core_j22_cpu_rf_N3359,
         j202_soc_core_j22_cpu_rf_N3358, j202_soc_core_j22_cpu_rf_N3357,
         j202_soc_core_j22_cpu_rf_N3356, j202_soc_core_j22_cpu_rf_N3355,
         j202_soc_core_j22_cpu_rf_N3354, j202_soc_core_j22_cpu_rf_N3352,
         j202_soc_core_j22_cpu_rf_N3351, j202_soc_core_j22_cpu_rf_N3350,
         j202_soc_core_j22_cpu_rf_N3349, j202_soc_core_j22_cpu_rf_N3348,
         j202_soc_core_j22_cpu_rf_N3347, j202_soc_core_j22_cpu_rf_N3346,
         j202_soc_core_j22_cpu_rf_N3345, j202_soc_core_j22_cpu_rf_N3343,
         j202_soc_core_j22_cpu_rf_N3342, j202_soc_core_j22_cpu_rf_N3341,
         j202_soc_core_j22_cpu_rf_N3340, j202_soc_core_j22_cpu_rf_N3339,
         j202_soc_core_j22_cpu_rf_N3338, j202_soc_core_j22_cpu_rf_N3337,
         j202_soc_core_j22_cpu_rf_N3336, j202_soc_core_j22_cpu_rf_N3335,
         j202_soc_core_j22_cpu_rf_N3334, j202_soc_core_j22_cpu_rf_N3333,
         j202_soc_core_j22_cpu_rf_N3331, j202_soc_core_j22_cpu_rf_N3330,
         j202_soc_core_j22_cpu_rf_N3329, j202_soc_core_j22_cpu_rf_N3328,
         j202_soc_core_j22_cpu_rf_N3327, j202_soc_core_j22_cpu_rf_N3326,
         j202_soc_core_j22_cpu_rf_N3325, j202_soc_core_j22_cpu_rf_N3324,
         j202_soc_core_j22_cpu_rf_N3323, j202_soc_core_j22_cpu_rf_N3322,
         j202_soc_core_j22_cpu_rf_N3321, j202_soc_core_j22_cpu_rf_N3319,
         j202_soc_core_j22_cpu_rf_N3318, j202_soc_core_j22_cpu_rf_N3317,
         j202_soc_core_j22_cpu_rf_N3316, j202_soc_core_j22_cpu_rf_N3315,
         j202_soc_core_j22_cpu_rf_N3314, j202_soc_core_j22_cpu_rf_N3313,
         j202_soc_core_j22_cpu_rf_N3311, j202_soc_core_j22_cpu_rf_N3309,
         j202_soc_core_j22_cpu_rf_N3307, j202_soc_core_j22_cpu_rf_N3305,
         j202_soc_core_j22_cpu_rf_N3304, j202_soc_core_j22_cpu_rf_N3303,
         j202_soc_core_j22_cpu_rf_N3302, j202_soc_core_j22_cpu_rf_N3300,
         j202_soc_core_j22_cpu_rf_N3299, j202_soc_core_j22_cpu_rf_N3298,
         j202_soc_core_j22_cpu_rf_N3297, j202_soc_core_j22_cpu_rf_N3296,
         j202_soc_core_j22_cpu_rf_N3295, j202_soc_core_j22_cpu_rf_N3294,
         j202_soc_core_j22_cpu_rf_N3292, j202_soc_core_j22_cpu_rf_N3291,
         j202_soc_core_j22_cpu_rf_N3290, j202_soc_core_j22_cpu_rf_N3289,
         j202_soc_core_j22_cpu_rf_N3288, j202_soc_core_j22_cpu_rf_N3287,
         j202_soc_core_j22_cpu_rf_N3286, j202_soc_core_j22_cpu_rf_N3284,
         j202_soc_core_j22_cpu_rf_N3283, j202_soc_core_j22_cpu_rf_N3282,
         j202_soc_core_j22_cpu_rf_N3281, j202_soc_core_j22_cpu_rf_N3280,
         j202_soc_core_j22_cpu_rf_N3279, j202_soc_core_j22_cpu_rf_N3278,
         j202_soc_core_j22_cpu_rf_N3276, j202_soc_core_j22_cpu_rf_N3275,
         j202_soc_core_j22_cpu_rf_N3274, j202_soc_core_j22_cpu_rf_N3273,
         j202_soc_core_j22_cpu_rf_N3272, j202_soc_core_j22_cpu_rf_N3271,
         j202_soc_core_j22_cpu_rf_N3270, j202_soc_core_j22_cpu_rf_N3268,
         j202_soc_core_j22_cpu_rf_N3267, j202_soc_core_j22_cpu_rf_N3266,
         j202_soc_core_j22_cpu_rf_N3265, j202_soc_core_j22_cpu_rf_N3263,
         j202_soc_core_j22_cpu_rf_N3262, j202_soc_core_j22_cpu_rf_N3261,
         j202_soc_core_j22_cpu_rf_N3260, j202_soc_core_j22_cpu_rf_N3259,
         j202_soc_core_j22_cpu_rf_N3258, j202_soc_core_j22_cpu_rf_N3257,
         j202_soc_core_j22_cpu_rf_N3255, j202_soc_core_j22_cpu_rf_N3254,
         j202_soc_core_j22_cpu_rf_N3253, j202_soc_core_j22_cpu_rf_N3252,
         j202_soc_core_j22_cpu_rf_N3251, j202_soc_core_j22_cpu_rf_N3250,
         j202_soc_core_j22_cpu_rf_N3249, j202_soc_core_j22_cpu_rf_N3247,
         j202_soc_core_j22_cpu_rf_N3246, j202_soc_core_j22_cpu_rf_N3245,
         j202_soc_core_j22_cpu_rf_N3244, j202_soc_core_j22_cpu_rf_N3243,
         j202_soc_core_j22_cpu_rf_N3242, j202_soc_core_j22_cpu_rf_N3241,
         j202_soc_core_j22_cpu_rf_N3239, j202_soc_core_j22_cpu_rf_N3238,
         j202_soc_core_j22_cpu_rf_N3237, j202_soc_core_j22_cpu_rf_N3236,
         j202_soc_core_j22_cpu_rf_N3235, j202_soc_core_j22_cpu_rf_N3234,
         j202_soc_core_j22_cpu_rf_N3233, j202_soc_core_j22_cpu_rf_N3231,
         j202_soc_core_j22_cpu_rf_N3230, j202_soc_core_j22_cpu_rf_N3229,
         j202_soc_core_j22_cpu_rf_N3228, j202_soc_core_j22_cpu_rf_N3227,
         j202_soc_core_j22_cpu_rf_N3226, j202_soc_core_j22_cpu_rf_N3225,
         j202_soc_core_j22_cpu_rf_N3224, j202_soc_core_j22_cpu_rf_N3223,
         j202_soc_core_j22_cpu_rf_N3222, j202_soc_core_j22_cpu_rf_N3221,
         j202_soc_core_j22_cpu_rf_N3220, j202_soc_core_j22_cpu_rf_N3218,
         j202_soc_core_j22_cpu_rf_N3217, j202_soc_core_j22_cpu_rf_N3216,
         j202_soc_core_j22_cpu_rf_N3215, j202_soc_core_j22_cpu_rf_N3214,
         j202_soc_core_j22_cpu_rf_N3213, j202_soc_core_j22_cpu_rf_N3212,
         j202_soc_core_j22_cpu_rf_N3210, j202_soc_core_j22_cpu_rf_N3209,
         j202_soc_core_j22_cpu_rf_N3208, j202_soc_core_j22_cpu_rf_N3207,
         j202_soc_core_j22_cpu_rf_N3206, j202_soc_core_j22_cpu_rf_N3205,
         j202_soc_core_j22_cpu_rf_N3204, j202_soc_core_j22_cpu_rf_N3202,
         j202_soc_core_j22_cpu_rf_N3201, j202_soc_core_j22_cpu_rf_N3200,
         j202_soc_core_j22_cpu_rf_N3199, j202_soc_core_j22_cpu_rf_N3198,
         j202_soc_core_j22_cpu_rf_N3197, j202_soc_core_j22_cpu_rf_N3196,
         j202_soc_core_j22_cpu_rf_N3194, j202_soc_core_j22_cpu_rf_N3193,
         j202_soc_core_j22_cpu_rf_N3192, j202_soc_core_j22_cpu_rf_N3191,
         j202_soc_core_j22_cpu_rf_N3190, j202_soc_core_j22_cpu_rf_N3189,
         j202_soc_core_j22_cpu_rf_N3188, j202_soc_core_j22_cpu_rf_N3187,
         j202_soc_core_j22_cpu_rf_N3186, j202_soc_core_j22_cpu_rf_N3185,
         j202_soc_core_j22_cpu_rf_N3184, j202_soc_core_j22_cpu_rf_N3183,
         j202_soc_core_j22_cpu_rf_N3181, j202_soc_core_j22_cpu_rf_N3180,
         j202_soc_core_j22_cpu_rf_N3179, j202_soc_core_j22_cpu_rf_N3178,
         j202_soc_core_j22_cpu_rf_N3177, j202_soc_core_j22_cpu_rf_N3176,
         j202_soc_core_j22_cpu_rf_N3175, j202_soc_core_j22_cpu_rf_N3173,
         j202_soc_core_j22_cpu_rf_N3172, j202_soc_core_j22_cpu_rf_N3171,
         j202_soc_core_j22_cpu_rf_N3170, j202_soc_core_j22_cpu_rf_N3169,
         j202_soc_core_j22_cpu_rf_N3168, j202_soc_core_j22_cpu_rf_N3167,
         j202_soc_core_j22_cpu_rf_N3165, j202_soc_core_j22_cpu_rf_N3164,
         j202_soc_core_j22_cpu_rf_N3163, j202_soc_core_j22_cpu_rf_N3162,
         j202_soc_core_j22_cpu_rf_N3161, j202_soc_core_j22_cpu_rf_N3160,
         j202_soc_core_j22_cpu_rf_N3159, j202_soc_core_j22_cpu_rf_N3157,
         j202_soc_core_j22_cpu_rf_N3156, j202_soc_core_j22_cpu_rf_N3155,
         j202_soc_core_j22_cpu_rf_N3154, j202_soc_core_j22_cpu_rf_N3152,
         j202_soc_core_j22_cpu_rf_N3151, j202_soc_core_j22_cpu_rf_N3150,
         j202_soc_core_j22_cpu_rf_N3149, j202_soc_core_j22_cpu_rf_N3148,
         j202_soc_core_j22_cpu_rf_N3147, j202_soc_core_j22_cpu_rf_N3146,
         j202_soc_core_j22_cpu_rf_N3144, j202_soc_core_j22_cpu_rf_N3143,
         j202_soc_core_j22_cpu_rf_N3142, j202_soc_core_j22_cpu_rf_N3141,
         j202_soc_core_j22_cpu_rf_N3140, j202_soc_core_j22_cpu_rf_N3139,
         j202_soc_core_j22_cpu_rf_N3138, j202_soc_core_j22_cpu_rf_N3136,
         j202_soc_core_j22_cpu_rf_N3135, j202_soc_core_j22_cpu_rf_N3134,
         j202_soc_core_j22_cpu_rf_N3133, j202_soc_core_j22_cpu_rf_N3132,
         j202_soc_core_j22_cpu_rf_N3131, j202_soc_core_j22_cpu_rf_N3130,
         j202_soc_core_j22_cpu_rf_N3128, j202_soc_core_j22_cpu_rf_N3127,
         j202_soc_core_j22_cpu_rf_N3126, j202_soc_core_j22_cpu_rf_N3125,
         j202_soc_core_j22_cpu_rf_N3124, j202_soc_core_j22_cpu_rf_N3123,
         j202_soc_core_j22_cpu_rf_N3122, j202_soc_core_j22_cpu_rf_N3120,
         j202_soc_core_j22_cpu_rf_N3119, j202_soc_core_j22_cpu_rf_N3118,
         j202_soc_core_j22_cpu_rf_N3117, j202_soc_core_j22_cpu_rf_N3116,
         j202_soc_core_j22_cpu_rf_N3115, j202_soc_core_j22_cpu_rf_N3114,
         j202_soc_core_j22_cpu_rf_N3113, j202_soc_core_j22_cpu_rf_N3112,
         j202_soc_core_j22_cpu_rf_N3111, j202_soc_core_j22_cpu_rf_N3110,
         j202_soc_core_j22_cpu_rf_N3109, j202_soc_core_j22_cpu_rf_N3107,
         j202_soc_core_j22_cpu_rf_N3106, j202_soc_core_j22_cpu_rf_N3105,
         j202_soc_core_j22_cpu_rf_N3104, j202_soc_core_j22_cpu_rf_N3103,
         j202_soc_core_j22_cpu_rf_N3102, j202_soc_core_j22_cpu_rf_N3101,
         j202_soc_core_j22_cpu_rf_N3099, j202_soc_core_j22_cpu_rf_N3098,
         j202_soc_core_j22_cpu_rf_N3097, j202_soc_core_j22_cpu_rf_N3096,
         j202_soc_core_j22_cpu_rf_N3095, j202_soc_core_j22_cpu_rf_N3094,
         j202_soc_core_j22_cpu_rf_N3093, j202_soc_core_j22_cpu_rf_N3091,
         j202_soc_core_j22_cpu_rf_N3090, j202_soc_core_j22_cpu_rf_N3089,
         j202_soc_core_j22_cpu_rf_N3088, j202_soc_core_j22_cpu_rf_N3087,
         j202_soc_core_j22_cpu_rf_N3086, j202_soc_core_j22_cpu_rf_N3085,
         j202_soc_core_j22_cpu_rf_N3083, j202_soc_core_j22_cpu_rf_N3082,
         j202_soc_core_j22_cpu_rf_N3081, j202_soc_core_j22_cpu_rf_N3080,
         j202_soc_core_j22_cpu_rf_N3079, j202_soc_core_j22_cpu_rf_N3078,
         j202_soc_core_j22_cpu_rf_N3077, j202_soc_core_j22_cpu_rf_N3076,
         j202_soc_core_j22_cpu_rf_N3075, j202_soc_core_j22_cpu_rf_N3074,
         j202_soc_core_j22_cpu_rf_N3073, j202_soc_core_j22_cpu_rf_N3072,
         j202_soc_core_j22_cpu_rf_N3070, j202_soc_core_j22_cpu_rf_N3069,
         j202_soc_core_j22_cpu_rf_N3068, j202_soc_core_j22_cpu_rf_N3067,
         j202_soc_core_j22_cpu_rf_N3066, j202_soc_core_j22_cpu_rf_N3065,
         j202_soc_core_j22_cpu_rf_N3064, j202_soc_core_j22_cpu_rf_N3062,
         j202_soc_core_j22_cpu_rf_N3061, j202_soc_core_j22_cpu_rf_N3060,
         j202_soc_core_j22_cpu_rf_N3059, j202_soc_core_j22_cpu_rf_N3058,
         j202_soc_core_j22_cpu_rf_N3057, j202_soc_core_j22_cpu_rf_N3056,
         j202_soc_core_j22_cpu_rf_N3054, j202_soc_core_j22_cpu_rf_N3053,
         j202_soc_core_j22_cpu_rf_N3052, j202_soc_core_j22_cpu_rf_N3051,
         j202_soc_core_j22_cpu_rf_N3050, j202_soc_core_j22_cpu_rf_N3049,
         j202_soc_core_j22_cpu_rf_N3048, j202_soc_core_j22_cpu_rf_N3046,
         j202_soc_core_j22_cpu_rf_N3045, j202_soc_core_j22_cpu_rf_N3044,
         j202_soc_core_j22_cpu_rf_N3043, j202_soc_core_j22_cpu_rf_N3042,
         j202_soc_core_j22_cpu_rf_N3041, j202_soc_core_j22_cpu_rf_N3040,
         j202_soc_core_j22_cpu_rf_N3039, j202_soc_core_j22_cpu_rf_N3038,
         j202_soc_core_j22_cpu_rf_N3037, j202_soc_core_j22_cpu_rf_N3036,
         j202_soc_core_j22_cpu_rf_N3035, j202_soc_core_j22_cpu_rf_N3033,
         j202_soc_core_j22_cpu_rf_N3032, j202_soc_core_j22_cpu_rf_N3031,
         j202_soc_core_j22_cpu_rf_N3030, j202_soc_core_j22_cpu_rf_N3029,
         j202_soc_core_j22_cpu_rf_N3028, j202_soc_core_j22_cpu_rf_N3027,
         j202_soc_core_j22_cpu_rf_N3025, j202_soc_core_j22_cpu_rf_N3024,
         j202_soc_core_j22_cpu_rf_N3023, j202_soc_core_j22_cpu_rf_N3022,
         j202_soc_core_j22_cpu_rf_N3021, j202_soc_core_j22_cpu_rf_N3020,
         j202_soc_core_j22_cpu_rf_N3019, j202_soc_core_j22_cpu_rf_N3017,
         j202_soc_core_j22_cpu_rf_N3016, j202_soc_core_j22_cpu_rf_N3015,
         j202_soc_core_j22_cpu_rf_N3014, j202_soc_core_j22_cpu_rf_N3013,
         j202_soc_core_j22_cpu_rf_N3012, j202_soc_core_j22_cpu_rf_N3011,
         j202_soc_core_j22_cpu_rf_N3009, j202_soc_core_j22_cpu_rf_N3008,
         j202_soc_core_j22_cpu_rf_N3007, j202_soc_core_j22_cpu_rf_N3006,
         j202_soc_core_j22_cpu_rf_N3005, j202_soc_core_j22_cpu_rf_N3004,
         j202_soc_core_j22_cpu_rf_N3003, j202_soc_core_j22_cpu_rf_N3002,
         j202_soc_core_j22_cpu_rf_N3001, j202_soc_core_j22_cpu_rf_N3000,
         j202_soc_core_j22_cpu_rf_N2999, j202_soc_core_j22_cpu_rf_N2998,
         j202_soc_core_j22_cpu_rf_N2996, j202_soc_core_j22_cpu_rf_N2995,
         j202_soc_core_j22_cpu_rf_N2994, j202_soc_core_j22_cpu_rf_N2993,
         j202_soc_core_j22_cpu_rf_N2992, j202_soc_core_j22_cpu_rf_N2991,
         j202_soc_core_j22_cpu_rf_N2990, j202_soc_core_j22_cpu_rf_N2988,
         j202_soc_core_j22_cpu_rf_N2987, j202_soc_core_j22_cpu_rf_N2986,
         j202_soc_core_j22_cpu_rf_N2985, j202_soc_core_j22_cpu_rf_N2984,
         j202_soc_core_j22_cpu_rf_N2983, j202_soc_core_j22_cpu_rf_N2982,
         j202_soc_core_j22_cpu_rf_N2980, j202_soc_core_j22_cpu_rf_N2979,
         j202_soc_core_j22_cpu_rf_N2978, j202_soc_core_j22_cpu_rf_N2977,
         j202_soc_core_j22_cpu_rf_N2976, j202_soc_core_j22_cpu_rf_N2975,
         j202_soc_core_j22_cpu_rf_N2974, j202_soc_core_j22_cpu_rf_N2972,
         j202_soc_core_j22_cpu_rf_N2971, j202_soc_core_j22_cpu_rf_N2970,
         j202_soc_core_j22_cpu_rf_N2969, j202_soc_core_j22_cpu_rf_N2968,
         j202_soc_core_j22_cpu_rf_N2967, j202_soc_core_j22_cpu_rf_N2966,
         j202_soc_core_j22_cpu_rf_N2965, j202_soc_core_j22_cpu_rf_N2964,
         j202_soc_core_j22_cpu_rf_N2963, j202_soc_core_j22_cpu_rf_N2962,
         j202_soc_core_j22_cpu_rf_N2961, j202_soc_core_j22_cpu_rf_N2959,
         j202_soc_core_j22_cpu_rf_N2958, j202_soc_core_j22_cpu_rf_N2957,
         j202_soc_core_j22_cpu_rf_N2956, j202_soc_core_j22_cpu_rf_N2955,
         j202_soc_core_j22_cpu_rf_N2954, j202_soc_core_j22_cpu_rf_N2953,
         j202_soc_core_j22_cpu_rf_N2951, j202_soc_core_j22_cpu_rf_N2950,
         j202_soc_core_j22_cpu_rf_N2949, j202_soc_core_j22_cpu_rf_N2948,
         j202_soc_core_j22_cpu_rf_N2947, j202_soc_core_j22_cpu_rf_N2946,
         j202_soc_core_j22_cpu_rf_N2945, j202_soc_core_j22_cpu_rf_N2943,
         j202_soc_core_j22_cpu_rf_N2942, j202_soc_core_j22_cpu_rf_N2941,
         j202_soc_core_j22_cpu_rf_N2940, j202_soc_core_j22_cpu_rf_N2939,
         j202_soc_core_j22_cpu_rf_N2938, j202_soc_core_j22_cpu_rf_N2937,
         j202_soc_core_j22_cpu_rf_N2935, j202_soc_core_j22_cpu_rf_N2934,
         j202_soc_core_j22_cpu_rf_N2933, j202_soc_core_j22_cpu_rf_N2932,
         j202_soc_core_j22_cpu_rf_N2931, j202_soc_core_j22_cpu_rf_N2930,
         j202_soc_core_j22_cpu_rf_N2929, j202_soc_core_j22_cpu_rf_N2928,
         j202_soc_core_j22_cpu_rf_N2927, j202_soc_core_j22_cpu_rf_N2926,
         j202_soc_core_j22_cpu_rf_N2925, j202_soc_core_j22_cpu_rf_N2924,
         j202_soc_core_j22_cpu_rf_N2922, j202_soc_core_j22_cpu_rf_N2921,
         j202_soc_core_j22_cpu_rf_N2920, j202_soc_core_j22_cpu_rf_N2919,
         j202_soc_core_j22_cpu_rf_N2918, j202_soc_core_j22_cpu_rf_N2917,
         j202_soc_core_j22_cpu_rf_N2916, j202_soc_core_j22_cpu_rf_N2914,
         j202_soc_core_j22_cpu_rf_N2913, j202_soc_core_j22_cpu_rf_N2912,
         j202_soc_core_j22_cpu_rf_N2911, j202_soc_core_j22_cpu_rf_N2910,
         j202_soc_core_j22_cpu_rf_N2909, j202_soc_core_j22_cpu_rf_N2908,
         j202_soc_core_j22_cpu_rf_N2906, j202_soc_core_j22_cpu_rf_N2905,
         j202_soc_core_j22_cpu_rf_N2904, j202_soc_core_j22_cpu_rf_N2903,
         j202_soc_core_j22_cpu_rf_N2902, j202_soc_core_j22_cpu_rf_N2901,
         j202_soc_core_j22_cpu_rf_N2900, j202_soc_core_j22_cpu_rf_N2898,
         j202_soc_core_j22_cpu_rf_N2897, j202_soc_core_j22_cpu_rf_N2896,
         j202_soc_core_j22_cpu_rf_N2895, j202_soc_core_j22_cpu_rf_N2894,
         j202_soc_core_j22_cpu_rf_N2893, j202_soc_core_j22_cpu_rf_N2892,
         j202_soc_core_j22_cpu_rf_N2891, j202_soc_core_j22_cpu_rf_N2890,
         j202_soc_core_j22_cpu_rf_N2889, j202_soc_core_j22_cpu_rf_N2888,
         j202_soc_core_j22_cpu_rf_N2887, j202_soc_core_j22_cpu_rf_N2885,
         j202_soc_core_j22_cpu_rf_N2884, j202_soc_core_j22_cpu_rf_N2883,
         j202_soc_core_j22_cpu_rf_N2882, j202_soc_core_j22_cpu_rf_N2881,
         j202_soc_core_j22_cpu_rf_N2880, j202_soc_core_j22_cpu_rf_N2879,
         j202_soc_core_j22_cpu_rf_N2877, j202_soc_core_j22_cpu_rf_N2876,
         j202_soc_core_j22_cpu_rf_N2875, j202_soc_core_j22_cpu_rf_N2874,
         j202_soc_core_j22_cpu_rf_N2873, j202_soc_core_j22_cpu_rf_N2872,
         j202_soc_core_j22_cpu_rf_N2871, j202_soc_core_j22_cpu_rf_N2869,
         j202_soc_core_j22_cpu_rf_N2868, j202_soc_core_j22_cpu_rf_N2867,
         j202_soc_core_j22_cpu_rf_N2866, j202_soc_core_j22_cpu_rf_N2865,
         j202_soc_core_j22_cpu_rf_N2864, j202_soc_core_j22_cpu_rf_N2863,
         j202_soc_core_j22_cpu_rf_N2861, j202_soc_core_j22_cpu_rf_N2860,
         j202_soc_core_j22_cpu_rf_N2859, j202_soc_core_j22_cpu_rf_N2858,
         j202_soc_core_j22_cpu_rf_N2857, j202_soc_core_j22_cpu_rf_N2856,
         j202_soc_core_j22_cpu_rf_N2855, j202_soc_core_j22_cpu_rf_N2854,
         j202_soc_core_j22_cpu_rf_N2853, j202_soc_core_j22_cpu_rf_N2852,
         j202_soc_core_j22_cpu_rf_N2851, j202_soc_core_j22_cpu_rf_N2850,
         j202_soc_core_j22_cpu_rf_N2848, j202_soc_core_j22_cpu_rf_N2847,
         j202_soc_core_j22_cpu_rf_N2846, j202_soc_core_j22_cpu_rf_N2845,
         j202_soc_core_j22_cpu_rf_N2844, j202_soc_core_j22_cpu_rf_N2843,
         j202_soc_core_j22_cpu_rf_N2842, j202_soc_core_j22_cpu_rf_N2840,
         j202_soc_core_j22_cpu_rf_N2839, j202_soc_core_j22_cpu_rf_N2838,
         j202_soc_core_j22_cpu_rf_N2837, j202_soc_core_j22_cpu_rf_N2836,
         j202_soc_core_j22_cpu_rf_N2835, j202_soc_core_j22_cpu_rf_N2834,
         j202_soc_core_j22_cpu_rf_N2832, j202_soc_core_j22_cpu_rf_N2831,
         j202_soc_core_j22_cpu_rf_N2830, j202_soc_core_j22_cpu_rf_N2829,
         j202_soc_core_j22_cpu_rf_N2828, j202_soc_core_j22_cpu_rf_N2827,
         j202_soc_core_j22_cpu_rf_N2826, j202_soc_core_j22_cpu_rf_N2824,
         j202_soc_core_j22_cpu_rf_N2823, j202_soc_core_j22_cpu_rf_N2822,
         j202_soc_core_j22_cpu_rf_N2821, j202_soc_core_j22_cpu_rf_N2820,
         j202_soc_core_j22_cpu_rf_N2819, j202_soc_core_j22_cpu_rf_N2818,
         j202_soc_core_j22_cpu_rf_N2817, j202_soc_core_j22_cpu_rf_N2816,
         j202_soc_core_j22_cpu_rf_N2815, j202_soc_core_j22_cpu_rf_N2814,
         j202_soc_core_j22_cpu_rf_N2813, j202_soc_core_j22_cpu_rf_N2811,
         j202_soc_core_j22_cpu_rf_N2810, j202_soc_core_j22_cpu_rf_N2809,
         j202_soc_core_j22_cpu_rf_N2808, j202_soc_core_j22_cpu_rf_N2807,
         j202_soc_core_j22_cpu_rf_N2806, j202_soc_core_j22_cpu_rf_N2805,
         j202_soc_core_j22_cpu_rf_N2803, j202_soc_core_j22_cpu_rf_N2802,
         j202_soc_core_j22_cpu_rf_N2801, j202_soc_core_j22_cpu_rf_N2800,
         j202_soc_core_j22_cpu_rf_N2799, j202_soc_core_j22_cpu_rf_N2798,
         j202_soc_core_j22_cpu_rf_N2797, j202_soc_core_j22_cpu_rf_N2795,
         j202_soc_core_j22_cpu_rf_N2794, j202_soc_core_j22_cpu_rf_N2793,
         j202_soc_core_j22_cpu_rf_N2792, j202_soc_core_j22_cpu_rf_N2791,
         j202_soc_core_j22_cpu_rf_N2790, j202_soc_core_j22_cpu_rf_N2789,
         j202_soc_core_j22_cpu_rf_N2787, j202_soc_core_j22_cpu_rf_N2786,
         j202_soc_core_j22_cpu_rf_N2785, j202_soc_core_j22_cpu_rf_N2784,
         j202_soc_core_j22_cpu_rf_N2783, j202_soc_core_j22_cpu_rf_N2782,
         j202_soc_core_j22_cpu_rf_N2781, j202_soc_core_j22_cpu_rf_N2780,
         j202_soc_core_j22_cpu_rf_N2779, j202_soc_core_j22_cpu_rf_N2778,
         j202_soc_core_j22_cpu_rf_N2777, j202_soc_core_j22_cpu_rf_N2776,
         j202_soc_core_j22_cpu_rf_N2774, j202_soc_core_j22_cpu_rf_N2773,
         j202_soc_core_j22_cpu_rf_N2772, j202_soc_core_j22_cpu_rf_N2771,
         j202_soc_core_j22_cpu_rf_N2770, j202_soc_core_j22_cpu_rf_N2769,
         j202_soc_core_j22_cpu_rf_N2768, j202_soc_core_j22_cpu_rf_N2766,
         j202_soc_core_j22_cpu_rf_N2765, j202_soc_core_j22_cpu_rf_N2764,
         j202_soc_core_j22_cpu_rf_N2763, j202_soc_core_j22_cpu_rf_N2762,
         j202_soc_core_j22_cpu_rf_N2761, j202_soc_core_j22_cpu_rf_N2760,
         j202_soc_core_j22_cpu_rf_N2758, j202_soc_core_j22_cpu_rf_N2757,
         j202_soc_core_j22_cpu_rf_N2756, j202_soc_core_j22_cpu_rf_N2755,
         j202_soc_core_j22_cpu_rf_N2754, j202_soc_core_j22_cpu_rf_N2753,
         j202_soc_core_j22_cpu_rf_N2752, j202_soc_core_j22_cpu_rf_N2750,
         j202_soc_core_j22_cpu_rf_N2749, j202_soc_core_j22_cpu_rf_N2748,
         j202_soc_core_j22_cpu_rf_N2747, j202_soc_core_j22_cpu_rf_N2746,
         j202_soc_core_j22_cpu_rf_N2745, j202_soc_core_j22_cpu_rf_N2744,
         j202_soc_core_j22_cpu_rf_N2743, j202_soc_core_j22_cpu_rf_N2742,
         j202_soc_core_j22_cpu_rf_N2741, j202_soc_core_j22_cpu_rf_N2740,
         j202_soc_core_j22_cpu_rf_N2739, j202_soc_core_j22_cpu_rf_N2737,
         j202_soc_core_j22_cpu_rf_N2736, j202_soc_core_j22_cpu_rf_N2735,
         j202_soc_core_j22_cpu_rf_N2734, j202_soc_core_j22_cpu_rf_N2733,
         j202_soc_core_j22_cpu_rf_N2732, j202_soc_core_j22_cpu_rf_N2731,
         j202_soc_core_j22_cpu_rf_N2729, j202_soc_core_j22_cpu_rf_N2728,
         j202_soc_core_j22_cpu_rf_N2727, j202_soc_core_j22_cpu_rf_N2726,
         j202_soc_core_j22_cpu_rf_N2725, j202_soc_core_j22_cpu_rf_N2724,
         j202_soc_core_j22_cpu_rf_N2723, j202_soc_core_j22_cpu_rf_N2721,
         j202_soc_core_j22_cpu_rf_N2720, j202_soc_core_j22_cpu_rf_N2719,
         j202_soc_core_j22_cpu_rf_N2718, j202_soc_core_j22_cpu_rf_N2717,
         j202_soc_core_j22_cpu_rf_N2716, j202_soc_core_j22_cpu_rf_N2715,
         j202_soc_core_j22_cpu_rf_N2713, j202_soc_core_j22_cpu_rf_N2712,
         j202_soc_core_j22_cpu_rf_N2711, j202_soc_core_j22_cpu_rf_N2710,
         j202_soc_core_j22_cpu_rf_N2709, j202_soc_core_j22_cpu_rf_N2708,
         j202_soc_core_j22_cpu_rf_N2707, j202_soc_core_j22_cpu_rf_N2706,
         j202_soc_core_j22_cpu_rf_N2705, j202_soc_core_j22_cpu_rf_N2704,
         j202_soc_core_j22_cpu_rf_N2703, j202_soc_core_j22_cpu_rf_N2702,
         j202_soc_core_j22_cpu_rf_N2700, j202_soc_core_j22_cpu_rf_N2699,
         j202_soc_core_j22_cpu_rf_N2698, j202_soc_core_j22_cpu_rf_N2697,
         j202_soc_core_j22_cpu_rf_N2696, j202_soc_core_j22_cpu_rf_N2695,
         j202_soc_core_j22_cpu_rf_N2694, j202_soc_core_j22_cpu_rf_N2692,
         j202_soc_core_j22_cpu_rf_N2691, j202_soc_core_j22_cpu_rf_N2690,
         j202_soc_core_j22_cpu_rf_N2689, j202_soc_core_j22_cpu_rf_N2688,
         j202_soc_core_j22_cpu_rf_N2687, j202_soc_core_j22_cpu_rf_N2686,
         j202_soc_core_j22_cpu_rf_N2684, j202_soc_core_j22_cpu_rf_N2683,
         j202_soc_core_j22_cpu_rf_N2682, j202_soc_core_j22_cpu_rf_N2681,
         j202_soc_core_j22_cpu_rf_N2680, j202_soc_core_j22_cpu_rf_N2679,
         j202_soc_core_j22_cpu_rf_N2678, j202_soc_core_j22_cpu_rf_N2674,
         j202_soc_core_j22_cpu_rf_N2671, j202_soc_core_j22_cpu_rf_N2670,
         j202_soc_core_j22_cpu_rf_N2667, j202_soc_core_j22_cpu_rf_N2663,
         j202_soc_core_j22_cpu_rf_N2662, j202_soc_core_j22_cpu_rf_N2658,
         j202_soc_core_j22_cpu_rf_N2657, j202_soc_core_j22_cpu_rf_N2653,
         j202_soc_core_j22_cpu_rf_N2649, j202_soc_core_j22_cpu_rf_N2648,
         j202_soc_core_j22_cpu_rf_N2647, j202_soc_core_j22_cpu_rf_N2646,
         j202_soc_core_j22_cpu_rf_N2645, j202_soc_core_j22_cpu_rf_N2644,
         j202_soc_core_j22_cpu_rf_N2643, j202_soc_core_j22_cpu_rf_N2642,
         j202_soc_core_j22_cpu_rf_N2640, j202_soc_core_j22_cpu_rf_N2639,
         j202_soc_core_j22_cpu_rf_N2638, j202_soc_core_j22_cpu_rf_N2637,
         j202_soc_core_j22_cpu_rf_N2628, j202_soc_core_j22_cpu_rf_N2627,
         j202_soc_core_j22_cpu_rf_N2626, j202_soc_core_j22_cpu_rf_N2625,
         j202_soc_core_j22_cpu_rf_N329, j202_soc_core_j22_cpu_rf_N328,
         j202_soc_core_j22_cpu_rf_N327, j202_soc_core_j22_cpu_rf_N326,
         j202_soc_core_j22_cpu_rf_N325, j202_soc_core_j22_cpu_rf_N324,
         j202_soc_core_j22_cpu_rf_N323, j202_soc_core_j22_cpu_rf_N322,
         j202_soc_core_j22_cpu_rf_N321, j202_soc_core_j22_cpu_rf_N320,
         j202_soc_core_j22_cpu_rf_N319, j202_soc_core_j22_cpu_rf_N318,
         j202_soc_core_j22_cpu_rf_N317, j202_soc_core_j22_cpu_rf_N316,
         j202_soc_core_j22_cpu_rf_N315, j202_soc_core_j22_cpu_rf_N314,
         j202_soc_core_j22_cpu_rf_N313, j202_soc_core_j22_cpu_rf_N312,
         j202_soc_core_j22_cpu_rf_N311, j202_soc_core_j22_cpu_rf_N310,
         j202_soc_core_j22_cpu_rf_N309, j202_soc_core_j22_cpu_rf_N308,
         j202_soc_core_j22_cpu_rf_N307, j202_soc_core_j22_cpu_rf_N306,
         j202_soc_core_j22_cpu_rf_N305, j202_soc_core_j22_cpu_rf_N304,
         j202_soc_core_j22_cpu_rf_N303, j202_soc_core_j22_cpu_rf_N302,
         j202_soc_core_j22_cpu_rf_N301, j202_soc_core_j22_cpu_rf_N300,
         j202_soc_core_j22_cpu_rf_N299, j202_soc_core_j22_cpu_rf_N298,
         j202_soc_core_j22_cpu_ma_N56, j202_soc_core_j22_cpu_ma_N55,
         j202_soc_core_j22_cpu_ma_N54, j202_soc_core_j22_cpu_ma_N53,
         j202_soc_core_j22_cpu_ml_N429, j202_soc_core_j22_cpu_ml_N427,
         j202_soc_core_j22_cpu_ml_N426, j202_soc_core_j22_cpu_ml_N425,
         j202_soc_core_j22_cpu_ml_N424, j202_soc_core_j22_cpu_ml_N423,
         j202_soc_core_j22_cpu_ml_N422, j202_soc_core_j22_cpu_ml_N421,
         j202_soc_core_j22_cpu_ml_N420, j202_soc_core_j22_cpu_ml_N419,
         j202_soc_core_j22_cpu_ml_N418, j202_soc_core_j22_cpu_ml_N417,
         j202_soc_core_j22_cpu_ml_N416, j202_soc_core_j22_cpu_ml_N415,
         j202_soc_core_j22_cpu_ml_N414, j202_soc_core_j22_cpu_ml_N413,
         j202_soc_core_j22_cpu_ml_N412, j202_soc_core_j22_cpu_ml_N370,
         j202_soc_core_j22_cpu_ml_N369, j202_soc_core_j22_cpu_ml_N368,
         j202_soc_core_j22_cpu_ml_N367, j202_soc_core_j22_cpu_ml_N363,
         j202_soc_core_j22_cpu_ml_N362, j202_soc_core_j22_cpu_ml_N361,
         j202_soc_core_j22_cpu_ml_N360, j202_soc_core_j22_cpu_ml_N359,
         j202_soc_core_j22_cpu_ml_N357, j202_soc_core_j22_cpu_ml_N356,
         j202_soc_core_j22_cpu_ml_N354, j202_soc_core_j22_cpu_ml_N336,
         j202_soc_core_j22_cpu_ml_N335, j202_soc_core_j22_cpu_ml_N334,
         j202_soc_core_j22_cpu_ml_N333, j202_soc_core_j22_cpu_ml_N332,
         j202_soc_core_j22_cpu_ml_N331, j202_soc_core_j22_cpu_ml_N330,
         j202_soc_core_j22_cpu_ml_N329, j202_soc_core_j22_cpu_ml_N328,
         j202_soc_core_j22_cpu_ml_N327, j202_soc_core_j22_cpu_ml_N326,
         j202_soc_core_j22_cpu_ml_N325, j202_soc_core_j22_cpu_ml_N324,
         j202_soc_core_j22_cpu_ml_N323, j202_soc_core_j22_cpu_ml_N322,
         j202_soc_core_j22_cpu_ml_N321, j202_soc_core_j22_cpu_ml_N320,
         j202_soc_core_j22_cpu_ml_N319, j202_soc_core_j22_cpu_ml_N318,
         j202_soc_core_j22_cpu_ml_N317, j202_soc_core_j22_cpu_ml_N316,
         j202_soc_core_j22_cpu_ml_N315, j202_soc_core_j22_cpu_ml_N314,
         j202_soc_core_j22_cpu_ml_N313, j202_soc_core_j22_cpu_ml_N312,
         j202_soc_core_j22_cpu_ml_N311, j202_soc_core_j22_cpu_ml_N310,
         j202_soc_core_j22_cpu_ml_N309, j202_soc_core_j22_cpu_ml_N308,
         j202_soc_core_j22_cpu_ml_N307, j202_soc_core_j22_cpu_ml_N306,
         j202_soc_core_j22_cpu_ml_N305, j202_soc_core_j22_cpu_ml_N304,
         j202_soc_core_j22_cpu_ml_N303, j202_soc_core_j22_cpu_ml_N195,
         j202_soc_core_j22_cpu_ml_N194, j202_soc_core_j22_cpu_ml_N193,
         j202_soc_core_j22_cpu_ml_N192, j202_soc_core_j22_cpu_ml_N191,
         j202_soc_core_j22_cpu_ml_N156, j202_soc_core_j22_cpu_ml_N155,
         j202_soc_core_j22_cpu_ml_N154, j202_soc_core_j22_cpu_ml_N153,
         j202_soc_core_j22_cpu_ml_N152,
         j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_N497,
         j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_N487,
         j202_soc_core_ahb2apb_00_N143, j202_soc_core_ahb2apb_00_N142,
         j202_soc_core_ahb2apb_00_N141, j202_soc_core_ahb2apb_00_N140,
         j202_soc_core_ahb2apb_00_N139, j202_soc_core_ahb2apb_00_N138,
         j202_soc_core_ahb2apb_00_N137, j202_soc_core_ahb2apb_00_N136,
         j202_soc_core_ahb2apb_00_N135, j202_soc_core_ahb2apb_00_N134,
         j202_soc_core_ahb2apb_00_N133, j202_soc_core_ahb2apb_00_N132,
         j202_soc_core_ahb2apb_00_N131, j202_soc_core_ahb2apb_00_N130,
         j202_soc_core_ahb2apb_00_N129, j202_soc_core_ahb2apb_00_N128,
         j202_soc_core_ahb2apb_00_N127, j202_soc_core_ahb2apb_00_N90,
         j202_soc_core_ahb2apb_00_N89, j202_soc_core_ahb2apb_00_N55,
         j202_soc_core_ahb2apb_00_N30, j202_soc_core_ahb2apb_00_N29,
         j202_soc_core_ahb2apb_00_N28, j202_soc_core_ahb2apb_00_N27,
         j202_soc_core_ahb2apb_00_N26, j202_soc_core_ahb2apb_00_N25,
         j202_soc_core_ahb2apb_00_N24, j202_soc_core_ahb2apb_00_N23,
         j202_soc_core_ahb2apb_00_N22, j202_soc_core_cmt_core_00_cmf1,
         j202_soc_core_cmt_core_00_cmf0, j202_soc_core_cmt_core_00_str1,
         j202_soc_core_cmt_core_00_str0,
         j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_2,
         j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_1,
         j202_soc_core_cmt_core_00_cmt_apb_00_nxt_state_0_,
         j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen,
         j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_nxt_latch_status_0_,
         j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_0_,
         j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_nxt_latch_status_0_,
         j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_0_,
         j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt1_to1,
         j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt0_to1,
         j202_soc_core_ahb2apb_01_N159, j202_soc_core_ahb2apb_01_N158,
         j202_soc_core_ahb2apb_01_N157, j202_soc_core_ahb2apb_01_N156,
         j202_soc_core_ahb2apb_01_N155, j202_soc_core_ahb2apb_01_N154,
         j202_soc_core_ahb2apb_01_N153, j202_soc_core_ahb2apb_01_N152,
         j202_soc_core_ahb2apb_01_N151, j202_soc_core_ahb2apb_01_N150,
         j202_soc_core_ahb2apb_01_N149, j202_soc_core_ahb2apb_01_N148,
         j202_soc_core_ahb2apb_01_N147, j202_soc_core_ahb2apb_01_N146,
         j202_soc_core_ahb2apb_01_N145, j202_soc_core_ahb2apb_01_N144,
         j202_soc_core_ahb2apb_01_N143, j202_soc_core_ahb2apb_01_N142,
         j202_soc_core_ahb2apb_01_N141, j202_soc_core_ahb2apb_01_N140,
         j202_soc_core_ahb2apb_01_N139, j202_soc_core_ahb2apb_01_N138,
         j202_soc_core_ahb2apb_01_N137, j202_soc_core_ahb2apb_01_N136,
         j202_soc_core_ahb2apb_01_N135, j202_soc_core_ahb2apb_01_N134,
         j202_soc_core_ahb2apb_01_N133, j202_soc_core_ahb2apb_01_N132,
         j202_soc_core_ahb2apb_01_N131, j202_soc_core_ahb2apb_01_N130,
         j202_soc_core_ahb2apb_01_N129, j202_soc_core_ahb2apb_01_N128,
         j202_soc_core_ahb2apb_01_N123, j202_soc_core_ahb2apb_01_N91,
         j202_soc_core_ahb2apb_01_N90, j202_soc_core_ahb2apb_01_N22,
         j202_soc_core_intc_core_00_cp_intack_all_0_,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_0__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_1__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_2__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_3__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_4__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_5__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_6__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_7__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_8__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_9__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_10__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_11__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_12__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_13__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_14__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_15__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N23,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N22,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N21,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N20,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N19,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N18,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N17,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N16,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N15,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N14,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N13,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N12,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N11,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N10,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N9,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N8,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N7,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N6,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N5,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N4,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N23,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N22,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N21,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N20,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N19,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N18,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N17,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N16,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N15,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N14,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N13,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N12,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N11,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N10,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N9,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N8,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N7,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N6,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N5,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N4,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N3,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_req_N3,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N6,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N5,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N4,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N3,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N6,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N5,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N4,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N3,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N9,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N7,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N6,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N5,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N4,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N3,
         j202_soc_core_ahb2apb_02_N159, j202_soc_core_ahb2apb_02_N158,
         j202_soc_core_ahb2apb_02_N157, j202_soc_core_ahb2apb_02_N156,
         j202_soc_core_ahb2apb_02_N155, j202_soc_core_ahb2apb_02_N154,
         j202_soc_core_ahb2apb_02_N153, j202_soc_core_ahb2apb_02_N152,
         j202_soc_core_ahb2apb_02_N151, j202_soc_core_ahb2apb_02_N150,
         j202_soc_core_ahb2apb_02_N149, j202_soc_core_ahb2apb_02_N148,
         j202_soc_core_ahb2apb_02_N147, j202_soc_core_ahb2apb_02_N146,
         j202_soc_core_ahb2apb_02_N145, j202_soc_core_ahb2apb_02_N144,
         j202_soc_core_ahb2apb_02_N143, j202_soc_core_ahb2apb_02_N142,
         j202_soc_core_ahb2apb_02_N141, j202_soc_core_ahb2apb_02_N140,
         j202_soc_core_ahb2apb_02_N139, j202_soc_core_ahb2apb_02_N138,
         j202_soc_core_ahb2apb_02_N137, j202_soc_core_ahb2apb_02_N136,
         j202_soc_core_ahb2apb_02_N135, j202_soc_core_ahb2apb_02_N134,
         j202_soc_core_ahb2apb_02_N133, j202_soc_core_ahb2apb_02_N132,
         j202_soc_core_ahb2apb_02_N131, j202_soc_core_ahb2apb_02_N130,
         j202_soc_core_ahb2apb_02_N129, j202_soc_core_ahb2apb_02_N128,
         j202_soc_core_ahb2apb_02_N123, j202_soc_core_ahb2apb_02_N91,
         j202_soc_core_ahb2apb_02_N90, j202_soc_core_ahb2apb_02_N22,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N34,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N33,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N32,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N31,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N30,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N29,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N28,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N27,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N26,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N25,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N24,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N23,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N22,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N21,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N20,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N19,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N18,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N17,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N16,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N15,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N14,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N13,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N12,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N11,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N10,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N9,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N8,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N7,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N6,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N5,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N4,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N3,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N71,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N70,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N69,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N68,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N67,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N66,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N65,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N64,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N63,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N62,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N61,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N60,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N59,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N58,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N57,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N56,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N55,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N54,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N53,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N52,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N51,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N50,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N49,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N48,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N47,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N46,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N45,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N44,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N43,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N42,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N41,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N40,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N34,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N33,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N32,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N31,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N30,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N29,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N28,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N27,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N25,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N24,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N23,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N22,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N21,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N20,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N19,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N16,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N11,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N6,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N4,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N3,
         j202_soc_core_ahb2aqu_00_N164, j202_soc_core_ahb2aqu_00_N163,
         j202_soc_core_ahb2aqu_00_N161, j202_soc_core_ahb2aqu_00_N136,
         j202_soc_core_ahb2aqu_00_N135, j202_soc_core_ahb2aqu_00_N134,
         j202_soc_core_ahb2aqu_00_N133, j202_soc_core_ahb2aqu_00_N132,
         j202_soc_core_ahb2aqu_00_N131, j202_soc_core_ahb2aqu_00_N127,
         j202_soc_core_ahb2aqu_00_N98, j202_soc_core_ahb2aqu_00_N95,
         j202_soc_core_ahb2aqu_00_aqu_st_0_, j202_soc_core_uart_sio_ce_x4,
         j202_soc_core_uart_sio_ce, j202_soc_core_uart_RDRXD1,
         j202_soc_core_uart_WRTXD1, j202_soc_core_uart_TOP_N137,
         j202_soc_core_uart_TOP_N128, j202_soc_core_uart_TOP_N123,
         j202_soc_core_uart_TOP_N118, j202_soc_core_uart_TOP_rx_sio_ce_r2,
         j202_soc_core_uart_TOP_rx_sio_ce_r1, j202_soc_core_uart_TOP_N102,
         j202_soc_core_uart_TOP_N101, j202_soc_core_uart_TOP_change,
         j202_soc_core_uart_TOP_N95, j202_soc_core_uart_TOP_rx_valid_r,
         j202_soc_core_uart_TOP_rx_valid, j202_soc_core_uart_TOP_N89,
         j202_soc_core_uart_TOP_N88, j202_soc_core_uart_TOP_N87,
         j202_soc_core_uart_TOP_N85, j202_soc_core_uart_TOP_rx_sio_ce,
         j202_soc_core_uart_TOP_rx_go, j202_soc_core_uart_TOP_rxd_r,
         j202_soc_core_uart_TOP_rxd_s, j202_soc_core_uart_TOP_N61,
         j202_soc_core_uart_TOP_N60, j202_soc_core_uart_TOP_N59,
         j202_soc_core_uart_TOP_N58, j202_soc_core_uart_TOP_N57,
         j202_soc_core_uart_TOP_N43, j202_soc_core_uart_TOP_shift_en_r,
         j202_soc_core_uart_TOP_N33, j202_soc_core_uart_TOP_N32,
         j202_soc_core_uart_TOP_N31, j202_soc_core_uart_TOP_N30,
         j202_soc_core_uart_TOP_N29, j202_soc_core_uart_TOP_N28,
         j202_soc_core_uart_TOP_N27, j202_soc_core_uart_TOP_N26,
         j202_soc_core_uart_TOP_N25, j202_soc_core_uart_TOP_N24,
         j202_soc_core_uart_TOP_load, j202_soc_core_uart_TOP_shift_en,
         j202_soc_core_uart_TOP_N16, j202_soc_core_uart_TOP_txf_empty_r,
         j202_soc_core_uart_TOP_tx_fifo_N42,
         j202_soc_core_uart_TOP_tx_fifo_N41, j202_soc_core_uart_TOP_tx_fifo_gb,
         j202_soc_core_uart_TOP_rx_fifo_N42,
         j202_soc_core_uart_TOP_rx_fifo_N41, j202_soc_core_uart_TOP_rx_fifo_gb,
         j202_soc_core_uart_BRG_N59, j202_soc_core_uart_BRG_sio_ce_r,
         j202_soc_core_uart_BRG_N57, j202_soc_core_uart_BRG_N55,
         j202_soc_core_uart_BRG_sio_ce_x4_t,
         j202_soc_core_uart_BRG_sio_ce_x4_r, j202_soc_core_uart_BRG_N47,
         j202_soc_core_uart_BRG_N42, j202_soc_core_uart_BRG_N41,
         j202_soc_core_uart_BRG_N40, j202_soc_core_uart_BRG_N39,
         j202_soc_core_uart_BRG_N38, j202_soc_core_uart_BRG_N37,
         j202_soc_core_uart_BRG_N36, j202_soc_core_uart_BRG_N35,
         j202_soc_core_uart_BRG_br_clr, j202_soc_core_uart_BRG_N21,
         j202_soc_core_uart_BRG_N19, j202_soc_core_uart_BRG_N18,
         j202_soc_core_uart_BRG_N17, j202_soc_core_uart_BRG_N16,
         j202_soc_core_uart_BRG_N15, j202_soc_core_uart_BRG_N14,
         j202_soc_core_uart_BRG_N13, j202_soc_core_uart_BRG_N12,
         j202_soc_core_uart_BRG_ps_clr, j202_soc_core_bldc_core_00_adc_en,
         j202_soc_core_bldc_core_00_pwm_en,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_nxt_bldc_int,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_0_,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_wen,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_nxt_latch_status_0_,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_0_,
         j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_2,
         j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1,
         j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posc,
         j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_negb,
         j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posb,
         j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posa,
         j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld,
         j202_soc_core_ahb2wbqspi_00_stb_o, j202_soc_core_wbqspiflash_00_N755,
         j202_soc_core_wbqspiflash_00_N750, j202_soc_core_wbqspiflash_00_N747,
         j202_soc_core_wbqspiflash_00_N746, j202_soc_core_wbqspiflash_00_N745,
         j202_soc_core_wbqspiflash_00_N743, j202_soc_core_wbqspiflash_00_N742,
         j202_soc_core_wbqspiflash_00_N741, j202_soc_core_wbqspiflash_00_N740,
         j202_soc_core_wbqspiflash_00_N739, j202_soc_core_wbqspiflash_00_N738,
         j202_soc_core_wbqspiflash_00_N737, j202_soc_core_wbqspiflash_00_N736,
         j202_soc_core_wbqspiflash_00_N735, j202_soc_core_wbqspiflash_00_N734,
         j202_soc_core_wbqspiflash_00_N733, j202_soc_core_wbqspiflash_00_N730,
         j202_soc_core_wbqspiflash_00_N729, j202_soc_core_wbqspiflash_00_N728,
         j202_soc_core_wbqspiflash_00_N727, j202_soc_core_wbqspiflash_00_N726,
         j202_soc_core_wbqspiflash_00_N725, j202_soc_core_wbqspiflash_00_N724,
         j202_soc_core_wbqspiflash_00_N723, j202_soc_core_wbqspiflash_00_N722,
         j202_soc_core_wbqspiflash_00_N721, j202_soc_core_wbqspiflash_00_N719,
         j202_soc_core_wbqspiflash_00_N718, j202_soc_core_wbqspiflash_00_N717,
         j202_soc_core_wbqspiflash_00_N716, j202_soc_core_wbqspiflash_00_N715,
         j202_soc_core_wbqspiflash_00_N714, j202_soc_core_wbqspiflash_00_N713,
         j202_soc_core_wbqspiflash_00_N712, j202_soc_core_wbqspiflash_00_N711,
         j202_soc_core_wbqspiflash_00_N710, j202_soc_core_wbqspiflash_00_N709,
         j202_soc_core_wbqspiflash_00_N708, j202_soc_core_wbqspiflash_00_N698,
         j202_soc_core_wbqspiflash_00_N697, j202_soc_core_wbqspiflash_00_N696,
         j202_soc_core_wbqspiflash_00_N695, j202_soc_core_wbqspiflash_00_N694,
         j202_soc_core_wbqspiflash_00_N688, j202_soc_core_wbqspiflash_00_N687,
         j202_soc_core_wbqspiflash_00_N686, j202_soc_core_wbqspiflash_00_N685,
         j202_soc_core_wbqspiflash_00_N684, j202_soc_core_wbqspiflash_00_N683,
         j202_soc_core_wbqspiflash_00_N682, j202_soc_core_wbqspiflash_00_N681,
         j202_soc_core_wbqspiflash_00_N674, j202_soc_core_wbqspiflash_00_N673,
         j202_soc_core_wbqspiflash_00_N672, j202_soc_core_wbqspiflash_00_N671,
         j202_soc_core_wbqspiflash_00_N670, j202_soc_core_wbqspiflash_00_N669,
         j202_soc_core_wbqspiflash_00_N668, j202_soc_core_wbqspiflash_00_N667,
         j202_soc_core_wbqspiflash_00_N663, j202_soc_core_wbqspiflash_00_N629,
         j202_soc_core_wbqspiflash_00_N628, j202_soc_core_wbqspiflash_00_N623,
         j202_soc_core_wbqspiflash_00_N622, j202_soc_core_wbqspiflash_00_N621,
         j202_soc_core_wbqspiflash_00_N620, j202_soc_core_wbqspiflash_00_N619,
         j202_soc_core_wbqspiflash_00_N618, j202_soc_core_wbqspiflash_00_N617,
         j202_soc_core_wbqspiflash_00_N616, j202_soc_core_wbqspiflash_00_N615,
         j202_soc_core_wbqspiflash_00_N614, j202_soc_core_wbqspiflash_00_N613,
         j202_soc_core_wbqspiflash_00_N612, j202_soc_core_wbqspiflash_00_N611,
         j202_soc_core_wbqspiflash_00_N609, j202_soc_core_wbqspiflash_00_N608,
         j202_soc_core_wbqspiflash_00_N607, j202_soc_core_wbqspiflash_00_N606,
         j202_soc_core_wbqspiflash_00_N605, j202_soc_core_wbqspiflash_00_N594,
         j202_soc_core_wbqspiflash_00_N592, j202_soc_core_wbqspiflash_00_N590,
         j202_soc_core_wbqspiflash_00_spif_cmd,
         j202_soc_core_wbqspiflash_00_spif_req,
         j202_soc_core_wbqspiflash_00_N86,
         j202_soc_core_wbqspiflash_00_alt_ctrl,
         j202_soc_core_wbqspiflash_00_N85,
         j202_soc_core_wbqspiflash_00_alt_cmd,
         j202_soc_core_wbqspiflash_00_spif_ctrl,
         j202_soc_core_wbqspiflash_00_spif_override,
         j202_soc_core_wbqspiflash_00_quad_mode_enabled,
         j202_soc_core_wbqspiflash_00_write_protect,
         j202_soc_core_wbqspiflash_00_dirty_sector,
         j202_soc_core_wbqspiflash_00_write_in_progress,
         j202_soc_core_wbqspiflash_00_w_qspi_cs_n,
         j202_soc_core_wbqspiflash_00_w_qspi_sck,
         j202_soc_core_wbqspiflash_00_spi_busy,
         j202_soc_core_wbqspiflash_00_spi_valid,
         j202_soc_core_wbqspiflash_00_spi_dir,
         j202_soc_core_wbqspiflash_00_spi_spd,
         j202_soc_core_wbqspiflash_00_spi_hold,
         j202_soc_core_wbqspiflash_00_spi_wr,
         j202_soc_core_wbqspiflash_00_lldriver_N430,
         j202_soc_core_wbqspiflash_00_lldriver_N429,
         j202_soc_core_wbqspiflash_00_lldriver_N428,
         j202_soc_core_wbqspiflash_00_lldriver_N427,
         j202_soc_core_wbqspiflash_00_lldriver_N426,
         j202_soc_core_wbqspiflash_00_lldriver_N425,
         j202_soc_core_wbqspiflash_00_lldriver_N424,
         j202_soc_core_wbqspiflash_00_lldriver_N423,
         j202_soc_core_wbqspiflash_00_lldriver_N422,
         j202_soc_core_wbqspiflash_00_lldriver_N421,
         j202_soc_core_wbqspiflash_00_lldriver_N420,
         j202_soc_core_wbqspiflash_00_lldriver_N419,
         j202_soc_core_wbqspiflash_00_lldriver_N418,
         j202_soc_core_wbqspiflash_00_lldriver_N417,
         j202_soc_core_wbqspiflash_00_lldriver_N416,
         j202_soc_core_wbqspiflash_00_lldriver_N415,
         j202_soc_core_wbqspiflash_00_lldriver_N414,
         j202_soc_core_wbqspiflash_00_lldriver_N413,
         j202_soc_core_wbqspiflash_00_lldriver_N412,
         j202_soc_core_wbqspiflash_00_lldriver_N411,
         j202_soc_core_wbqspiflash_00_lldriver_N410,
         j202_soc_core_wbqspiflash_00_lldriver_N409,
         j202_soc_core_wbqspiflash_00_lldriver_N408,
         j202_soc_core_wbqspiflash_00_lldriver_N407,
         j202_soc_core_wbqspiflash_00_lldriver_N406,
         j202_soc_core_wbqspiflash_00_lldriver_N405,
         j202_soc_core_wbqspiflash_00_lldriver_N404,
         j202_soc_core_wbqspiflash_00_lldriver_N403,
         j202_soc_core_wbqspiflash_00_lldriver_N402,
         j202_soc_core_wbqspiflash_00_lldriver_N401,
         j202_soc_core_wbqspiflash_00_lldriver_N400,
         j202_soc_core_wbqspiflash_00_lldriver_N399,
         j202_soc_core_wbqspiflash_00_lldriver_N398,
         j202_soc_core_wbqspiflash_00_lldriver_N397,
         j202_soc_core_wbqspiflash_00_lldriver_N396,
         j202_soc_core_wbqspiflash_00_lldriver_N395,
         j202_soc_core_wbqspiflash_00_lldriver_N394,
         j202_soc_core_wbqspiflash_00_lldriver_N393,
         j202_soc_core_wbqspiflash_00_lldriver_N392,
         j202_soc_core_wbqspiflash_00_lldriver_N391,
         j202_soc_core_wbqspiflash_00_lldriver_N389,
         j202_soc_core_wbqspiflash_00_lldriver_N361,
         j202_soc_core_wbqspiflash_00_lldriver_N360,
         j202_soc_core_wbqspiflash_00_lldriver_N359,
         j202_soc_core_wbqspiflash_00_lldriver_N358,
         j202_soc_core_wbqspiflash_00_lldriver_N356,
         j202_soc_core_wbqspiflash_00_lldriver_N355,
         j202_soc_core_wbqspiflash_00_lldriver_N354,
         j202_soc_core_wbqspiflash_00_lldriver_N326,
         j202_soc_core_wbqspiflash_00_lldriver_N325,
         j202_soc_core_wbqspiflash_00_lldriver_N324,
         j202_soc_core_wbqspiflash_00_lldriver_N323,
         j202_soc_core_wbqspiflash_00_lldriver_N321,
         j202_soc_core_wbqspiflash_00_lldriver_N319,
         j202_soc_core_wbqspiflash_00_lldriver_N318,
         j202_soc_core_wbqspiflash_00_lldriver_N317,
         j202_soc_core_wbqspiflash_00_lldriver_N316,
         j202_soc_core_wbqspiflash_00_lldriver_N315,
         j202_soc_core_wbqspiflash_00_lldriver_N314,
         j202_soc_core_wbqspiflash_00_lldriver_N313,
         j202_soc_core_wbqspiflash_00_lldriver_N312,
         j202_soc_core_wbqspiflash_00_lldriver_N311,
         j202_soc_core_wbqspiflash_00_lldriver_N310,
         j202_soc_core_wbqspiflash_00_lldriver_N308,
         j202_soc_core_wbqspiflash_00_lldriver_N307,
         j202_soc_core_wbqspiflash_00_lldriver_r_dir,
         j202_soc_core_wbqspiflash_00_lldriver_r_spd,
         j202_soc_core_bootrom_00_sel_w, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10539, n10540,
         n10541, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10561, n10562, n10563, n10565, n10566, n10567,
         n10568, n10569, n10570, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10605, n10606, n10607, n10608, n10674, n10675, n10676,
         n10678, n10679, n10745, n10746, n10747, n10748, n10904, n10905,
         n10906, n10907, n10911, DP_OP_1508J1_126_2326_n3,
         DP_OP_1508J1_126_2326_n4, DP_OP_1508J1_126_2326_n6,
         U7_RSOP_1495_C3_DATA3_2, n10920, n10921, n10922, n10923, n10926,
         n10929, n10930, n10931, n10932, n10933, n10934, n10938, n10939,
         n10940, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10957, n10958,
         n10959, n10960, n10961, n10963, n10964, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11316, n11317, n11318, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11348, n11349, n11350, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11611, n11612, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11726, n11727,
         n11728, n11729, n11730, n11732, n11733, n11734, n11735, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11864, n11865, n11866, n11867,
         n11868, n11869, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11989, n11990, n11991,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12040, n12041, n12042,
         n12045, n12046, n12047, n12048, n12049, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12060, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12109, n12110, n12111, n12112,
         n12114, n12115, n12116, n12117, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12146, n12147, n12148, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12180, n12181, n12182, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12520, n12521, n12522, n12523, n12524,
         n12526, n12527, n12528, n12529, n12530, n12531, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12581, n12582, n12583,
         n12584, n12585, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12902, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12974, n12975, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13100, n13101,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13183, n13184, n13185, n13186,
         n13187, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16358, n16359, n16360,
         n16361, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198,
         n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
         n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
         n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222,
         n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
         n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238,
         n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246,
         n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
         n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
         n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270,
         n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278,
         n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286,
         n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
         n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
         n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310,
         n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318,
         n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326,
         n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
         n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342,
         n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350,
         n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
         n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
         n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374,
         n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382,
         n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390,
         n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398,
         n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406,
         n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414,
         n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422,
         n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430,
         n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438,
         n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446,
         n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454,
         n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462,
         n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470,
         n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478,
         n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486,
         n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494,
         n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502,
         n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510,
         n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518,
         n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526,
         n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534,
         n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542,
         n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550,
         n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558,
         n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566,
         n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574,
         n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582,
         n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590,
         n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598,
         n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606,
         n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614,
         n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622,
         n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630,
         n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638,
         n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646,
         n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654,
         n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662,
         n21663, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
         n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
         n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
         n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
         n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
         n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711,
         n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719,
         n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
         n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
         n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
         n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
         n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759,
         n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
         n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
         n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
         n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
         n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
         n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807,
         n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
         n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
         n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831,
         n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
         n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
         n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855,
         n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863,
         n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
         n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879,
         n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
         n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
         n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
         n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
         n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
         n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
         n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
         n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
         n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
         n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
         n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999,
         n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
         n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
         n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
         n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
         n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
         n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
         n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
         n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
         n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071,
         n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
         n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
         n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095,
         n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
         n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111,
         n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119,
         n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
         n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
         n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143,
         n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151,
         n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
         n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167,
         n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
         n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183,
         n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
         n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
         n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
         n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215,
         n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223,
         n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
         n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239,
         n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247,
         n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255,
         n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263,
         n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271,
         n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
         n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287,
         n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295,
         n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
         n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311,
         n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
         n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
         n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
         n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343,
         n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
         n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359,
         n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367,
         n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375,
         n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383,
         n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391,
         n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399,
         n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
         n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415,
         n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423,
         n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431,
         n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439,
         n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
         n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455,
         n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463,
         n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
         n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479,
         n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487,
         n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495,
         n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503,
         n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511,
         n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519,
         n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527,
         n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535,
         n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543,
         n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551,
         n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559,
         n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567,
         n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575,
         n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583,
         n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591,
         n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599,
         n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607,
         n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615,
         n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623,
         n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631,
         n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639,
         n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647,
         n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655,
         n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663,
         n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671,
         n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679,
         n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687,
         n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695,
         n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703,
         n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711,
         n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719,
         n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727,
         n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735,
         n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743,
         n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751,
         n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759,
         n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767,
         n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775,
         n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783,
         n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791,
         n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799,
         n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807,
         n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815,
         n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823,
         n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831,
         n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839,
         n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847,
         n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855,
         n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863,
         n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871,
         n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879,
         n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887,
         n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895,
         n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903,
         n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911,
         n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919,
         n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927,
         n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935,
         n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943,
         n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951,
         n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959,
         n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967,
         n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975,
         n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983,
         n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991,
         n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999,
         n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007,
         n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015,
         n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023,
         n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031,
         n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039,
         n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047,
         n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055,
         n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063,
         n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071,
         n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079,
         n23080, n23081, n23082, n23083, n23084, n23086, n23087, n23088,
         n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096,
         n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104,
         n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112,
         n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120,
         n23121, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23208, n23209, n23210,
         n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218,
         n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226,
         n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234,
         n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242,
         n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250,
         n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258,
         n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266,
         n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274,
         n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282,
         n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290,
         n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298,
         n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306,
         n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314,
         n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322,
         n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330,
         n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338,
         n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346,
         n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354,
         n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362,
         n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370,
         n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378,
         n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386,
         n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394,
         n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402,
         n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410,
         n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418,
         n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426,
         n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434,
         n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442,
         n23443, n23444, n23445, n23446, n23447, n23449, n23450, n23451,
         n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459,
         n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
         n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
         n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483,
         n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
         n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499,
         n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
         n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515,
         n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
         n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531,
         n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
         n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
         n23548, n23549, n23552, n23553, n23554, n23555, n23556, n23557,
         n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565,
         n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573,
         n23574, n23575, n23576, n23577, n23578, n23580, n23581, n23582,
         n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590,
         n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598,
         n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606,
         n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614,
         n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622,
         n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630,
         n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638,
         n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646,
         n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654,
         n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662,
         n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670,
         n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678,
         n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686,
         n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694,
         n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702,
         n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710,
         n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718,
         n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726,
         n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734,
         n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742,
         n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750,
         n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758,
         n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766,
         n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774,
         n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782,
         n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790,
         n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798,
         n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806,
         n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
         n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
         n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835,
         n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
         n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851,
         n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859,
         n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867,
         n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
         n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
         n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891,
         n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
         n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907,
         n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
         n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
         n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
         n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
         n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964,
         n23965, n23966, n23967, n23968, n23970, n23971, n23972, n23973,
         n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981,
         n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989,
         n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997,
         n23998, n23999, n24000, n24001, n24002, n24003, n24005, n24006,
         n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014,
         n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022,
         n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030,
         n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038,
         n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046,
         n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054,
         n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062,
         n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070,
         n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078,
         n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086,
         n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094,
         n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102,
         n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110,
         n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118,
         n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126,
         n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134,
         n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142,
         n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150,
         n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158,
         n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166,
         n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174,
         n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182,
         n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190,
         n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200,
         n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208,
         n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216,
         n24217, n24218, n24219, n24220, n24221, n24222, n24225, n24226,
         n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234,
         n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242,
         n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250,
         n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258,
         n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266,
         n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274,
         n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282,
         n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290,
         n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298,
         n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306,
         n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314,
         n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322,
         n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330,
         n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338,
         n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346,
         n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354,
         n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362,
         n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370,
         n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378,
         n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386,
         n24387, n24388, n24389, n24390, n24392, n24393, n24394, n24395,
         n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
         n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411,
         n24412, n24413, n24414, n24415, n24417, n24418, n24419, n24420,
         n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428,
         n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436,
         n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444,
         n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452,
         n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460,
         n24461, n24462, n24463, n24464, n24465, n24466, n24468, n24469,
         n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477,
         n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485,
         n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493,
         n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501,
         n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509,
         n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517,
         n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525,
         n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533,
         n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541,
         n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549,
         n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557,
         n24558, n24559, n24560, n24561, n24562, n24564, n24565, n24566,
         n24567, n24569, n24570, n24571, n24572, n24573, n24574, n24575,
         n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583,
         n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591,
         n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599,
         n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607,
         n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615,
         n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623,
         n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631,
         n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639,
         n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647,
         n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655,
         n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663,
         n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671,
         n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679,
         n24680, n24681, n24682, n24684, n24685, n24686, n24687, n24688,
         n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696,
         n24697, n24698, n24699, n24700, n24702, n24703, n24704, n24705,
         n24706, n24707, n24709, n24710, n24711, n24712, n24713, n24714,
         n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722,
         n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730,
         n24731, n24732, n24733, n24734, n24736, n24737, n24738, n24739,
         n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748,
         n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756,
         n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764,
         n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772,
         n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780,
         n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788,
         n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796,
         n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804,
         n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812,
         n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820,
         n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828,
         n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836,
         n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844,
         n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852,
         n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860,
         n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868,
         n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876,
         n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884,
         n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892,
         n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900,
         n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908,
         n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916,
         n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924,
         n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932,
         n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940,
         n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948,
         n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956,
         n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964,
         n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972,
         n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980,
         n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988,
         n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996,
         n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004,
         n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012,
         n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020,
         n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028,
         n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036,
         n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044,
         n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052,
         n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060,
         n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068,
         n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076,
         n25077, n25078, n25080, n25081, n25082, n25083, n25084, n25085,
         n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093,
         n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101,
         n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109,
         n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117,
         n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125,
         n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133,
         n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141,
         n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149,
         n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157,
         n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165,
         n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173,
         n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181,
         n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189,
         n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197,
         n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205,
         n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213,
         n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221,
         n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229,
         n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237,
         n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245,
         n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253,
         n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261,
         n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269,
         n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277,
         n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285,
         n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293,
         n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301,
         n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309,
         n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317,
         n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325,
         n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333,
         n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341,
         n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349,
         n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357,
         n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365,
         n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373,
         n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381,
         n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389,
         n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397,
         n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405,
         n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413,
         n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421,
         n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429,
         n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437,
         n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445,
         n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453,
         n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461,
         n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469,
         n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477,
         n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485,
         n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493,
         n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501,
         n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509,
         n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517,
         n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525,
         n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533,
         n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541,
         n25542, n25544, n25545, n25546, n25547, n25548, n25549, n25550,
         n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558,
         n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566,
         n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574,
         n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582,
         n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590,
         n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598,
         n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606,
         n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614,
         n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622,
         n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630,
         n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638,
         n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646,
         n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654,
         n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662,
         n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670,
         n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678,
         n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686,
         n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694,
         n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702,
         n25703, n25704, n25705, n25706, n25707, n25708, n25709, n25710,
         n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718,
         n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726,
         n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734,
         n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742,
         n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750,
         n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758,
         n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766,
         n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774,
         n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782,
         n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790,
         n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798,
         n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806,
         n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814,
         n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822,
         n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830,
         n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838,
         n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846,
         n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854,
         n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862,
         n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870,
         n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878,
         n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886,
         n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894,
         n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902,
         n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910,
         n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918,
         n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926,
         n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934,
         n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942,
         n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950,
         n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958,
         n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966,
         n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974,
         n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982,
         n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990,
         n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998,
         n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006,
         n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014,
         n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022,
         n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030,
         n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038,
         n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046,
         n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054,
         n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062,
         n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070,
         n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078,
         n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086,
         n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094,
         n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102,
         n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110,
         n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118,
         n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126,
         n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134,
         n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142,
         n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150,
         n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158,
         n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166,
         n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174,
         n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182,
         n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190,
         n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198,
         n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206,
         n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214,
         n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222,
         n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230,
         n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238,
         n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246,
         n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254,
         n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262,
         n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270,
         n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278,
         n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286,
         n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294,
         n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302,
         n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310,
         n26311, n26312, n26313, n26314, n26315, n26317, n26318, n26319,
         n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327,
         n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335,
         n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343,
         n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351,
         n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359,
         n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367,
         n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375,
         n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383,
         n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391,
         n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399,
         n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407,
         n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415,
         n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423,
         n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431,
         n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439,
         n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26447,
         n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455,
         n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463,
         n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471,
         n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479,
         n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487,
         n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495,
         n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503,
         n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511,
         n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519,
         n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527,
         n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535,
         n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543,
         n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551,
         n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559,
         n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567,
         n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575,
         n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26584,
         n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592,
         n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600,
         n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608,
         n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616,
         n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624,
         n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632,
         n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640,
         n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648,
         n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656,
         n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664,
         n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672,
         n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680,
         n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688,
         n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696,
         n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704,
         n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712,
         n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720,
         n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728,
         n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736,
         n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744,
         n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752,
         n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760,
         n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768,
         n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776,
         n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784,
         n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792,
         n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800,
         n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808,
         n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816,
         n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824,
         n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832,
         n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840,
         n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848,
         n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856,
         n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864,
         n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872,
         n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880,
         n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888,
         n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896,
         n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904,
         n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912,
         n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920,
         n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928,
         n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936,
         n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944,
         n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952,
         n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960,
         n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968,
         n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976,
         n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984,
         n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992,
         n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000,
         n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008,
         n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016,
         n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024,
         n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032,
         n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040,
         n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048,
         n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056,
         n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064,
         n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072,
         n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080,
         n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088,
         n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096,
         n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104,
         n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112,
         n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120,
         n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128,
         n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136,
         n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144,
         n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152,
         n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160,
         n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168,
         n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176,
         n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184,
         n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192,
         n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200,
         n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208,
         n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216,
         n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224,
         n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232,
         n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240,
         n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248,
         n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256,
         n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264,
         n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272,
         n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280,
         n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288,
         n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296,
         n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304,
         n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312,
         n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320,
         n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328,
         n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336,
         n27337, n27338, n27339, n27340, n27341, n27342, n27343, n27344,
         n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352,
         n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360,
         n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368,
         n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376,
         n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384,
         n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392,
         n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400,
         n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408,
         n27409, n27410, n27411, n27412, n27413, n27414, n27415, n27416,
         n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424,
         n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432,
         n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440,
         n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448,
         n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456,
         n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464,
         n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472,
         n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480,
         n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488,
         n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496,
         n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504,
         n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512,
         n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520,
         n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528,
         n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536,
         n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544,
         n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552,
         n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560,
         n27561, n27562, n27563, n27564, n27565, n27566, n27567, n27568,
         n27569, n27570, n27571, n27572, n27573, n27574, n27575, n27576,
         n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584,
         n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592,
         n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600,
         n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608,
         n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616,
         n27617, n27618, n27619, n27620, n27621, n27622, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27778,
         n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786,
         n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794,
         n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802,
         n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810,
         n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818,
         n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826,
         n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834,
         n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842,
         n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850,
         n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858,
         n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866,
         n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874,
         n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882,
         n27883, n27884, n27885, n27887, n27888, n27889, n27890, n27891,
         n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899,
         n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907,
         n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915,
         n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923,
         n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931,
         n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939,
         n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947,
         n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955,
         n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963,
         n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971,
         n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979,
         n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987,
         n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995,
         n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003,
         n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011,
         n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019,
         n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027,
         n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035,
         n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043,
         n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051,
         n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059,
         n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067,
         n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075,
         n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083,
         n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091,
         n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099,
         n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107,
         n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115,
         n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123,
         n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131,
         n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139,
         n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147,
         n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155,
         n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163,
         n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171,
         n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179,
         n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187,
         n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195,
         n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203,
         n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211,
         n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219,
         n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227,
         n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235,
         n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243,
         n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251,
         n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259,
         n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267,
         n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275,
         n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283,
         n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291,
         n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299,
         n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307,
         n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315,
         n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323,
         n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331,
         n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339,
         n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347,
         n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355,
         n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363,
         n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371,
         n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379,
         n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387,
         n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395,
         n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403,
         n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411,
         n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419,
         n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427,
         n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435,
         n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443,
         n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451,
         n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459,
         n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467,
         n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475,
         n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483,
         n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491,
         n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499,
         n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507,
         n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515,
         n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523,
         n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531,
         n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539,
         n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
         n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555,
         n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563,
         n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571,
         n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579,
         n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587,
         n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595,
         n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603,
         n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611,
         n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
         n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627,
         n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635,
         n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643,
         n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651,
         n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659,
         n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667,
         n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675,
         n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683,
         n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691,
         n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699,
         n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707,
         n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715,
         n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723,
         n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731,
         n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739,
         n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747,
         n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755,
         n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763,
         n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771,
         n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779,
         n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787,
         n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795,
         n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803,
         n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811,
         n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819,
         n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827,
         n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835,
         n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843,
         n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851,
         n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859,
         n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867,
         n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875,
         n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883,
         n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891,
         n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899,
         n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907,
         n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915,
         n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923,
         n28924, n28926, n28927, n28928, n28929, n28930, n28931, n28932,
         n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940,
         n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948,
         n28949, n28950, n28951, n28952, n28953, n28954, n28955, n28956,
         n28957, n28958, n28959, n28960, n28961, n28962, n28963, n28964,
         n28965, n28966, n28967, n28968, n28969, n28970, n28971, n28972,
         n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980,
         n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988,
         n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996,
         n28997, n28998, n28999, n29000, n29001, n29002, n29003, n29004,
         n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012,
         n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020,
         n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028,
         n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036,
         n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044,
         n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052,
         n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060,
         n29061, n29062, n29063, n29064, n29065, n29066, n29067, n29068,
         n29069, n29070, n29071, n29072, n29073, n29074, n29075, n29076,
         n29077, n29078, n29079, n29080, n29081, n29082, n29083, n29084,
         n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092,
         n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119,
         n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127,
         n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135,
         n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143,
         n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151,
         n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159,
         n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167,
         n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175,
         n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183,
         n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191,
         n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199,
         n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207,
         n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215,
         n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223,
         n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231,
         n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239,
         n29240, n29242, n29243, n29244, n29245, n29246, n29247, n29248,
         n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29256,
         n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264,
         n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272,
         n29273, n29274, n29275, n29276, n29277, n29278, n29279, n29280,
         n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288,
         n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296,
         n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304,
         n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312,
         n29313, n29315, n29316, n29317, n29321, n29322, n29323, n29324,
         n29325, n29326, n29327, n29328, n29329, n29344, n29345, n29346,
         n29347, n29349, n29350, n29351, n29352, n29354, n29355, n29356,
         n29357, n29358, n29359, n29360, n29361, n29362, n29363, n29488,
         n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496,
         n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504,
         n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512,
         n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520,
         n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528,
         n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536,
         n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544,
         n29545, n29546, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412,
         SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414,
         SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416,
         SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418,
         SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420,
         SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422,
         SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424,
         SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426,
         SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428,
         SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430,
         SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432,
         SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434,
         SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436,
         SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438,
         SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440,
         SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442,
         SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444,
         SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446,
         SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448,
         SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450,
         SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452,
         SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454,
         SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456,
         SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458,
         SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460,
         SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_462,
         SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_464,
         SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_466,
         SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_468,
         SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_470,
         SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_472,
         SYNOPSYS_UNCONNECTED_473, SYNOPSYS_UNCONNECTED_474,
         SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_476,
         SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_478,
         SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_480,
         SYNOPSYS_UNCONNECTED_481, SYNOPSYS_UNCONNECTED_482,
         SYNOPSYS_UNCONNECTED_483, SYNOPSYS_UNCONNECTED_484,
         SYNOPSYS_UNCONNECTED_485, SYNOPSYS_UNCONNECTED_486,
         SYNOPSYS_UNCONNECTED_487, SYNOPSYS_UNCONNECTED_488,
         SYNOPSYS_UNCONNECTED_489, SYNOPSYS_UNCONNECTED_490,
         SYNOPSYS_UNCONNECTED_491, SYNOPSYS_UNCONNECTED_492,
         SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_494,
         SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_496,
         SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_498,
         SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_500,
         SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_502,
         SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_504,
         SYNOPSYS_UNCONNECTED_505, SYNOPSYS_UNCONNECTED_506,
         SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_508,
         SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_510,
         SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_512;
  wire   [31:0] gpio_en_o;
  wire   [1:0] start_n_reg;
  wire   [31:0] j202_soc_core_qspi_wb_wdat;
  wire   [24:2] j202_soc_core_qspi_wb_addr;
  wire   [15:0] j202_soc_core_prdata;
  wire   [6:0] j202_soc_core_paddr;
  wire   [7:0] j202_soc_core_pstrb;
  wire   [0:2] j202_soc_core_pwrite;
  wire   [5:0] j202_soc_core_j22_cpu_exuop_EXU_;
  wire   [4:0] j202_soc_core_j22_cpu_macop_MAC_;
  wire   [31:0] j202_soc_core_j22_cpu_pc;
  wire   [4:0] j202_soc_core_j22_cpu_opst;
  wire   [31:0] j202_soc_core_j22_cpu_rf_tmp;
  wire   [31:0] j202_soc_core_j22_cpu_rf_vbr;
  wire   [31:0] j202_soc_core_j22_cpu_rf_gbr;
  wire   [31:0] j202_soc_core_j22_cpu_rf_pr;
  wire   [511:0] j202_soc_core_j22_cpu_rf_gpr;
  wire   [1:0] j202_soc_core_j22_cpu_ma_M_address;
  wire   [1:0] j202_soc_core_j22_cpu_ma_M_area;
  wire   [3:0] j202_soc_core_j22_cpu_ma_M_MEM;
  wire   [31:0] j202_soc_core_j22_cpu_ml_maclj;
  wire   [31:0] j202_soc_core_j22_cpu_ml_machj;
  wire   [31:0] j202_soc_core_j22_cpu_ml_mach;
  wire   [31:0] j202_soc_core_j22_cpu_ml_macl;
  wire   [32:0] j202_soc_core_j22_cpu_ml_bufb;
  wire   [32:0] j202_soc_core_j22_cpu_ml_bufa;
  wire   [4:0] j202_soc_core_j22_cpu_ml_X_macop_MAC_;
  wire   [4:0] j202_soc_core_j22_cpu_ml_M_macop_MAC_;
  wire   [511:0] j202_soc_core_memory0_ram_dout0;
  wire   [15:0] j202_soc_core_memory0_ram_dout0_sel;
  wire   [111:0] j202_soc_core_ahblite_interconnect_s_hrdata;
  wire  
         [0:6] j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel
;
  wire   [2:0] j202_soc_core_ahb2apb_00_state;
  wire   [15:0] j202_soc_core_cmt_core_00_cnt1;
  wire   [15:0] j202_soc_core_cmt_core_00_cnt0;
  wire   [15:0] j202_soc_core_cmt_core_00_const1;
  wire   [15:0] j202_soc_core_cmt_core_00_const0;
  wire   [15:0] j202_soc_core_cmt_core_00_wdata_cnt0;
  wire   [1:0] j202_soc_core_cmt_core_00_cks1;
  wire   [1:0] j202_soc_core_cmt_core_00_cks0;
  wire   [7:0] j202_soc_core_cmt_core_00_reg_addr;
  wire   [1:0] j202_soc_core_cmt_core_00_cmt_apb_00_state;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata;
  wire   [6:2] j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1;
  wire   [6:2] j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1;
  wire   [9:0] j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1;
  wire   [9:0] j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0;
  wire   [9:0] j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0;
  wire   [9:0] j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0;
  wire   [2:0] j202_soc_core_ahb2apb_01_state;
  wire   [1:0] j202_soc_core_ahb2apb_01_hsize_buf;
  wire   [20:0] j202_soc_core_intc_core_00_in_intreq;
  wire   [127:0] j202_soc_core_intc_core_00_rg_ipr;
  wire   [127:0] j202_soc_core_intc_core_00_rg_itgt;
  wire   [20:0] j202_soc_core_intc_core_00_rg_irqc;
  wire   [31:0] j202_soc_core_intc_core_00_rg_ie;
  wire   [7:0] j202_soc_core_intc_core_00_rg_eimk;
  wire   [15:0] j202_soc_core_intc_core_00_rg_sint;
  wire   [11:0] j202_soc_core_intc_core_00_bs_addr;
  wire  
         [20:0] j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int
;
  wire  
         [6:0] j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch
;
  wire   [2:0] j202_soc_core_ahb2apb_02_state;
  wire   [1:0] j202_soc_core_ahb2apb_02_hsize_buf;
  wire   [7:0] j202_soc_core_gpio_core_00_reg_addr;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_dtr;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_isr;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_ier;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1;
  wire   [7:0] j202_soc_core_uart_din_i;
  wire   [7:0] j202_soc_core_uart_div1;
  wire   [7:0] j202_soc_core_uart_div0;
  wire   [1:0] j202_soc_core_uart_TOP_dpll_state;
  wire   [3:0] j202_soc_core_uart_TOP_rx_bit_cnt;
  wire   [3:0] j202_soc_core_uart_TOP_tx_bit_cnt;
  wire   [8:0] j202_soc_core_uart_TOP_hold_reg;
  wire   [9:2] j202_soc_core_uart_TOP_rxr;
  wire   [31:0] j202_soc_core_uart_TOP_tx_fifo_mem;
  wire   [1:0] j202_soc_core_uart_TOP_tx_fifo_rp;
  wire   [1:0] j202_soc_core_uart_TOP_tx_fifo_wp;
  wire   [31:0] j202_soc_core_uart_TOP_rx_fifo_mem;
  wire   [1:0] j202_soc_core_uart_TOP_rx_fifo_rp;
  wire   [1:0] j202_soc_core_uart_TOP_rx_fifo_wp;
  wire   [1:0] j202_soc_core_uart_BRG_cnt;
  wire   [7:0] j202_soc_core_uart_BRG_br_cnt;
  wire   [7:0] j202_soc_core_uart_BRG_ps;
  wire   [2:0] j202_soc_core_bldc_core_00_hall_value;
  wire   [2:0] j202_soc_core_bldc_core_00_comm;
  wire   [11:0] j202_soc_core_bldc_core_00_pwm_period;
  wire   [11:0] j202_soc_core_bldc_core_00_pwm_duty;
  wire   [23:0] j202_soc_core_bldc_core_00_wdata;
  wire   [7:0] j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1;
  wire   [1:0] j202_soc_core_bldc_core_00_bldc_wb_slave_00_state;
  wire  
         [2:0] j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status
;
  wire   [2:0] j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3;
  wire   [2:0] j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2;
  wire   [2:0] j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1;
  wire   [11:1] j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt;
  wire   [11:0] j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt;
  wire   [31:0] j202_soc_core_wbqspiflash_00_spif_data;
  wire   [7:0] j202_soc_core_wbqspiflash_00_last_status;
  wire   [9:0] j202_soc_core_wbqspiflash_00_reset_counter;
  wire   [4:0] j202_soc_core_wbqspiflash_00_state;
  wire   [7:0] j202_soc_core_wbqspiflash_00_erased_sector;
  wire   [23:2] j202_soc_core_wbqspiflash_00_w_spif_addr;
  wire   [3:0] j202_soc_core_wbqspiflash_00_w_qspi_dat;
  wire   [1:0] j202_soc_core_wbqspiflash_00_w_qspi_mod;
  wire   [31:0] j202_soc_core_wbqspiflash_00_spi_out;
  wire   [1:0] j202_soc_core_wbqspiflash_00_spi_len;
  wire   [31:0] j202_soc_core_wbqspiflash_00_spi_in;
  wire   [5:0] j202_soc_core_wbqspiflash_00_lldriver_spi_len;
  wire   [31:0] j202_soc_core_wbqspiflash_00_lldriver_r_word;
  wire   [30:0] j202_soc_core_wbqspiflash_00_lldriver_r_input;
  wire   [2:0] j202_soc_core_wbqspiflash_00_lldriver_state;
  wire   [17:2] j202_soc_core_bootrom_00_address_w;

  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_15__ram ( 
        .din0({n29299, n29297, n29293, n29291, n29289, n29287, n29285, n29283, 
        n29281, n29279, n29277, n29275, n29271, n29269, n29267, n29265, n29263, 
        n29261, n29259, n29257, n29255, n29253, n29312, n29310, n29308, n29306, 
        n29304, n29302, n29301, n29295, n29273, n29251}), .dout0(
        j202_soc_core_memory0_ram_dout0[511:480]), .addr0({n11090, n12528, 
        n12537, n11034, n10952, n12523, n10999, n12401, n29246}), .wmask0({
        n11023, n11097, n11009, n12539}), .dout1({SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_1}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10558), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_14__ram ( 
        .din0({n29300, n29298, n29294, n29292, n29290, n29288, n29286, n29284, 
        n29282, n29280, n29278, n29276, n29272, n29270, n29268, n29266, n29264, 
        n29262, n29260, n29258, n29256, n29254, n29313, n29311, n29309, n29307, 
        n29305, n29303, n12121, n29296, n29274, n29252}), .dout0(
        j202_soc_core_memory0_ram_dout0[479:448]), .addr0({n12407, n10992, 
        n12536, n11032, n10955, n12530, n10997, n11006, n12541}), .wmask0({
        n11013, n12413, n11002, n12539}), .dout1({SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_33}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10557), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_13__ram ( 
        .din0({n29299, n29297, n29293, n29291, n29289, n29287, n29285, n29283, 
        n29281, n29279, n29277, n29275, n29271, n29269, n29267, n29265, n29263, 
        n29261, n29259, n29257, n29255, n29253, n29312, n29310, n29308, n29306, 
        n29304, n29302, n12121, n29295, n29273, n29251}), .dout0(
        j202_soc_core_memory0_ram_dout0[447:416]), .addr0({n12407, n12527, 
        n12535, n11027, n10947, n12524, n10997, n11006, n29245}), .wmask0({
        n11022, n11018, n11021, n11017}), .dout1({SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_96, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_90, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_65}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10556), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_12__ram ( 
        .din0({n29300, n29298, n29294, n29292, n29290, n29288, n29286, n29284, 
        n29282, n29280, n29278, n29276, n29272, n29270, n29268, n29266, n29264, 
        n29262, n29260, n29258, n29256, n29254, n29313, n29311, n29309, n29307, 
        n29305, n29303, n12121, n29296, n29274, n29252}), .dout0(
        j202_soc_core_memory0_ram_dout0[415:384]), .addr0({n11014, n10996, 
        n29512, n11035, n10949, n12531, n12409, n11087, n10951}), .wmask0({
        n11025, n11019, n11021, n12540}), .dout1({SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_118, 
        SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_116, 
        SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_114, 
        SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_112, 
        SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_110, 
        SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_128, 
        SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_126, 
        SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_124, 
        SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_122, 
        SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_108, 
        SYNOPSYS_UNCONNECTED_97}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10555), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_11__ram ( 
        .din0({n29299, n29297, n29293, n29291, n29289, n29287, n29285, n29283, 
        n29281, n29279, n29277, n29275, n29271, n29269, n29267, n29265, n29263, 
        n29261, n29259, n29257, n29255, n29253, n29312, n29310, n29308, n29306, 
        n29304, n29302, n29301, n29295, n29273, n29251}), .dout0(
        j202_soc_core_memory0_ram_dout0[383:352]), .addr0({n11014, n10993, 
        n12518, n11033, n10948, n29525, n10998, n12406, n10945}), .wmask0({
        n11024, n12412, n11009, n11003}), .dout1({SYNOPSYS_UNCONNECTED_153, 
        SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_140, 
        SYNOPSYS_UNCONNECTED_129}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10554), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_10__ram ( 
        .din0({n29300, n29298, n29294, n29292, n29290, n29288, n29286, n29284, 
        n29282, n29280, n29278, n29276, n29272, n29270, n29268, n29266, n29264, 
        n29262, n29260, n29258, n29256, n29254, n29313, n29311, n29309, n29307, 
        n29305, n29303, n29301, n29296, n29274, n29252}), .dout0(
        j202_soc_core_memory0_ram_dout0[351:320]), .addr0({n11101, n12527, 
        n12537, n11029, n10948, n29526, n12403, n11007, n29246}), .wmask0({
        n11025, n11097, n11002, n11003}), .dout1({SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_178, 
        SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_176, 
        SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_174, 
        SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_171, 
        SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_169, 
        SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_167, 
        SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_165, 
        SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_163, 
        SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_192, 
        SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_190, 
        SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_188, 
        SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_186, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_172, 
        SYNOPSYS_UNCONNECTED_161}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10553), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_9__ram ( 
        .din0({n29299, n29297, n29293, n29291, n29289, n29287, n29285, n29283, 
        n29281, n29279, n29277, n29275, n29271, n29269, n29267, n29265, n29263, 
        n29261, n29259, n29257, n29255, n29253, n29312, n29310, n29308, n29306, 
        n29304, n29302, n29301, n29295, n29273, n29251}), .dout0(
        j202_soc_core_memory0_ram_dout0[319:288]), .addr0({n11090, n12526, 
        n12521, n11035, n10954, n12523, n12409, n29247, n11091}), .wmask0({
        n11024, n11000, n11099, n11088}), .dout1({SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_214, 
        SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_212, 
        SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_210, 
        SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_208, 
        SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_206, 
        SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_224, 
        SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_222, 
        SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_220, 
        SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_218, 
        SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_204, 
        SYNOPSYS_UNCONNECTED_193}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10552), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_8__ram ( 
        .din0({n29300, n29298, n29294, n29292, n29290, n29288, n29286, n29284, 
        n29282, n29280, n29278, n29276, n29272, n29270, n29268, n29266, n29264, 
        n29262, n29260, n29258, n29256, n29254, n29313, n29311, n29309, n29307, 
        n29305, n29303, n12121, n29296, n29274, n29252}), .dout0(
        j202_soc_core_memory0_ram_dout0[287:256]), .addr0({n12402, n10994, 
        n12535, n11028, n10949, n12530, n10991, n12401, n12541}), .wmask0({
        n11023, n12404, n11020, n11121}), .dout1({SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_246, 
        SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_244, 
        SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_242, 
        SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_240, 
        SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_238, 
        SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_256, 
        SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_254, 
        SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_252, 
        SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_250, 
        SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_236, 
        SYNOPSYS_UNCONNECTED_225}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10551), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_7__ram ( 
        .din0({n29299, n29297, n29293, n29291, n29289, n29287, n29285, n29283, 
        n29281, n29279, n29277, n29275, n29271, n29269, n29267, n29265, n29263, 
        n29261, n29259, n29257, n29255, n29253, n29312, n29310, n29308, n29306, 
        n29304, n29302, n29301, n29295, n29273, n29251}), .dout0(
        j202_soc_core_memory0_ram_dout0[255:224]), .addr0({n10943, n10994, 
        n29528, n11033, n10950, n12524, n10998, n11007, n10946}), .wmask0({
        n11013, n11000, n11123, n11004}), .dout1({SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_278, 
        SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_276, 
        SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_274, 
        SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_272, 
        SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_270, 
        SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_288, 
        SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_286, 
        SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_284, 
        SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_282, 
        SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_268, 
        SYNOPSYS_UNCONNECTED_257}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10550), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_6__ram ( 
        .din0({n29300, n29298, n29294, n29292, n29290, n29288, n29286, n29284, 
        n29282, n29280, n29278, n29276, n29272, n29270, n29268, n29266, n29264, 
        n29262, n29260, n29258, n29256, n29254, n29313, n29311, n29309, n29307, 
        n29305, n29303, n12121, n29296, n29274, n29252}), .dout0(
        j202_soc_core_memory0_ram_dout0[223:192]), .addr0({n11101, n10992, 
        n29509, n11032, n10953, n12531, n11092, n11031, n12408}), .wmask0({
        n11119, n12404, n11099, n11017}), .dout1({SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_299, 
        SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_297, 
        SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_295, 
        SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_293, 
        SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_291, 
        SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_320, 
        SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_318, 
        SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_316, 
        SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_314, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_289}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10549), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_5__ram ( 
        .din0({n29299, n29297, n29293, n29291, n29289, n29287, n29285, n29283, 
        n29281, n29279, n29277, n29275, n29271, n29269, n29267, n29265, n29263, 
        n29261, n29259, n29257, n29255, n29253, n29312, n29310, n29308, n29306, 
        n29304, n29302, n29301, n29295, n29273, n29251}), .dout0(
        j202_soc_core_memory0_ram_dout0[191:160]), .addr0({n10943, n10995, 
        n12536, n11030, n10950, n29527, n10999, n11031, n10946}), .wmask0({
        n11012, n12412, n11011, n11016}), .dout1({SYNOPSYS_UNCONNECTED_345, 
        SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_338, 
        SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_336, 
        SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_334, 
        SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_331, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_352, 
        SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_350, 
        SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_348, 
        SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_346, 
        SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_332, 
        SYNOPSYS_UNCONNECTED_321}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10548), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_4__ram ( 
        .din0({n29300, n29298, n29294, n29292, n29290, n29288, n29286, n29284, 
        n29282, n29280, n29278, n29276, n29272, n29270, n29268, n29266, n29264, 
        n29262, n29260, n29258, n29256, n29254, n29313, n29311, n29309, n29307, 
        n29305, n29303, n12121, n29296, n29274, n29252}), .dout0(
        j202_soc_core_memory0_ram_dout0[159:128]), .addr0({n10944, n10996, 
        n29511, n11034, n10953, n29527, n12403, n11005, n10951}), .wmask0({
        n11013, n12405, n11001, n12540}), .dout1({SYNOPSYS_UNCONNECTED_377, 
        SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_374, 
        SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_372, 
        SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_370, 
        SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_368, 
        SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_366, 
        SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_363, 
        SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_361, 
        SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_359, 
        SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_357, 
        SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_355, 
        SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_384, 
        SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_382, 
        SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_380, 
        SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_378, 
        SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_364, 
        SYNOPSYS_UNCONNECTED_353}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10547), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_3__ram ( 
        .din0({n29299, n29297, n29293, n29291, n29289, n29287, n29285, n29283, 
        n29281, n29279, n29277, n29275, n29271, n29269, n29267, n29265, n29263, 
        n29261, n29259, n29257, n29255, n29253, n29312, n29310, n29308, n29306, 
        n29304, n29302, n29301, n29295, n29273, n29251}), .dout0(
        j202_soc_core_memory0_ram_dout0[127:96]), .addr0({n11015, n10995, 
        n12517, n11030, n10947, n12522, n12410, n29247, n10945}), .wmask0({
        n11119, n11019, n11020, n11004}), .dout1({SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_406, 
        SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_404, 
        SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_402, 
        SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_400, 
        SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_398, 
        SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_389, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_416, 
        SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_414, 
        SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_412, 
        SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_410, 
        SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_396, 
        SYNOPSYS_UNCONNECTED_385}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10546), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_2__ram ( 
        .din0({n29300, n29298, n29294, n29292, n29290, n29288, n29286, n29284, 
        n29282, n29280, n29278, n29276, n29272, n29270, n29268, n29266, n29264, 
        n29262, n29260, n29258, n29256, n29254, n29313, n29311, n29309, n29307, 
        n29305, n29303, n12121, n29296, n29274, n29252}), .dout0(
        j202_soc_core_memory0_ram_dout0[95:64]), .addr0({n12402, n12528, 
        n12517, n11027, n10955, n12529, n11092, n11005, n11091}), .wmask0({
        n11013, n11018, n11123, n11121}), .dout1({SYNOPSYS_UNCONNECTED_441, 
        SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_438, 
        SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_436, 
        SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_434, 
        SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_432, 
        SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_430, 
        SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_427, 
        SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_425, 
        SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_423, 
        SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_421, 
        SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_419, 
        SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_448, 
        SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_446, 
        SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_444, 
        SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_442, 
        SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_428, 
        SYNOPSYS_UNCONNECTED_417}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10545), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_1__ram ( 
        .din0({n29299, n29297, n29293, n29291, n29289, n29287, n29285, n29283, 
        n29281, n29279, n29277, n29275, n29271, n29269, n29267, n29265, n29263, 
        n29261, n29259, n29257, n29255, n29253, n29312, n29310, n29308, n29306, 
        n29304, n29302, n29301, n29295, n29273, n29251}), .dout0(
        j202_soc_core_memory0_ram_dout0[63:32]), .addr0({n11015, n10993, 
        n12520, n11028, n10954, n12522, n10991, n12406, n29245}), .wmask0({
        n11119, n12405, n11001, n11016}), .dout1({SYNOPSYS_UNCONNECTED_473, 
        SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_470, 
        SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_468, 
        SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_466, 
        SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_464, 
        SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_462, 
        SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_459, 
        SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_457, 
        SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_455, 
        SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_453, 
        SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_451, 
        SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_480, 
        SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_478, 
        SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_476, 
        SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_474, 
        SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_460, 
        SYNOPSYS_UNCONNECTED_449}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10544), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_0__ram ( 
        .din0({n29300, n29298, n29294, n29292, n29290, n29288, n29286, n29284, 
        n29282, n29280, n29278, n29276, n29272, n29270, n29268, n29266, n29264, 
        n29262, n29260, n29258, n29256, n29254, n29313, n29311, n29309, n29307, 
        n29305, n29303, n12121, n29296, n29274, n29252}), .dout0(
        j202_soc_core_memory0_ram_dout0[31:0]), .addr0({n10944, n12526, n29510, 
        n11029, n10952, n12529, n12410, n11087, n10932}), .wmask0({n11119, 
        n12413, n11011, n11088}), .dout1({SYNOPSYS_UNCONNECTED_505, 
        SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_502, 
        SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_500, 
        SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_498, 
        SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_496, 
        SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_494, 
        SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_491, 
        SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_489, 
        SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_487, 
        SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_485, 
        SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_483, 
        SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_512, 
        SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_510, 
        SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_508, 
        SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_506, 
        SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_492, 
        SYNOPSYS_UNCONNECTED_481}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10543), .web0(n23581), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_fd_sc_hd__dfxtp_1 start_n_reg_reg_0_ ( .D(n3), .CLK(wb_clk_i), .Q(
        start_n_reg[0]) );
  sky130_fd_sc_hd__dfxtp_1 start_n_reg_reg_1_ ( .D(n4), .CLK(wb_clk_i), .Q(
        start_n_reg[1]) );
  sky130_fd_sc_hd__edfxtp_1 ready_reg ( .D(n29092), .DE(n470), .CLK(wb_clk_i), 
        .Q(wbs_ack_o) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_31_ ( .D(n460), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[31]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_30_ ( .D(n450), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[30]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_29_ ( .D(n440), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[29]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_28_ ( .D(n430), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[28]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_27_ ( .D(n420), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[27]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_26_ ( .D(n410), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[26]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_25_ ( .D(n400), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[25]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_24_ ( .D(n390), .DE(n380), .CLK(
        wb_clk_i), .Q(wbs_dat_o[24]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_23_ ( .D(n370), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[23]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_22_ ( .D(n360), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[22]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_21_ ( .D(n350), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[21]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_20_ ( .D(n340), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[20]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_19_ ( .D(n330), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[19]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_18_ ( .D(n320), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[18]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_17_ ( .D(n310), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[17]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_16_ ( .D(n300), .DE(n290), .CLK(
        wb_clk_i), .Q(wbs_dat_o[16]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_15_ ( .D(n280), .DE(n20), .CLK(
        wb_clk_i), .Q(wbs_dat_o[15]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_14_ ( .D(n270), .DE(n20), .CLK(
        wb_clk_i), .Q(wbs_dat_o[14]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_13_ ( .D(n260), .DE(n20), .CLK(
        wb_clk_i), .Q(wbs_dat_o[13]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_12_ ( .D(n250), .DE(n20), .CLK(
        wb_clk_i), .Q(wbs_dat_o[12]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_11_ ( .D(n240), .DE(n20), .CLK(
        wb_clk_i), .Q(wbs_dat_o[11]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_10_ ( .D(n230), .DE(n20), .CLK(
        wb_clk_i), .Q(wbs_dat_o[10]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_9_ ( .D(n220), .DE(n20), .CLK(wb_clk_i), .Q(wbs_dat_o[9]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_8_ ( .D(n21), .DE(n20), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[8]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_7_ ( .D(n19), .DE(n12), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[7]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_6_ ( .D(n18), .DE(n12), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[6]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_5_ ( .D(n17), .DE(n12), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[5]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_4_ ( .D(n16), .DE(n12), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[4]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_3_ ( .D(n15), .DE(n12), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[3]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_2_ ( .D(n14), .DE(n12), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[2]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_1_ ( .D(n13), .DE(n12), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[1]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_0_ ( .D(n11), .DE(n10), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_rst0_reg ( .D(n10487), .CLK(wb_clk_i), 
        .Q(j202_soc_core_rst0) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_rst1_reg ( .D(j202_soc_core_rst0), 
        .CLK(wb_clk_i), .Q(j202_soc_core_rst1) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_0_ ( 
        .D(n29152), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_1_ ( 
        .D(n29151), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_2_ ( 
        .D(n29150), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_3_ ( 
        .D(n29149), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_4_ ( 
        .D(n29148), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_5_ ( 
        .D(n29147), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_6_ ( 
        .D(n29146), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_7_ ( 
        .D(n29145), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_8_ ( 
        .D(n29144), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_9_ ( 
        .D(n29143), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_10_ ( 
        .D(n29142), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_11_ ( 
        .D(n29141), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_12_ ( 
        .D(n29140), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_13_ ( 
        .D(n29139), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_14_ ( 
        .D(n29138), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_15_ ( 
        .D(n29137), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_16_ ( 
        .D(n29136), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_17_ ( 
        .D(n29135), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_18_ ( 
        .D(n29134), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_19_ ( 
        .D(n29133), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_20_ ( 
        .D(n29132), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_21_ ( 
        .D(n29131), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_22_ ( 
        .D(n29130), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_23_ ( 
        .D(n29129), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_24_ ( 
        .D(n29128), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_25_ ( 
        .D(n29127), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_26_ ( 
        .D(n29126), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_27_ ( 
        .D(n29125), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_28_ ( 
        .D(n29124), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_29_ ( 
        .D(n29123), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_30_ ( 
        .D(n29122), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_31_ ( 
        .D(n29121), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_0_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N3), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_1_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N4), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_2_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N5), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_3_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N6), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_4_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N7), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_5_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N8), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_6_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N9), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_7_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N10), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_8_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N11), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_9_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N12), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_10_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N13), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[10])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_11_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N14), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[11])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_12_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N15), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[12])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_13_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N16), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_14_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N17), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_15_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N18), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_16_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N19), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_17_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N20), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[17])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_18_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N21), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[18])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_19_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N22), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[19])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_20_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N23), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[20])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_21_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[21])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_22_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N25), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[22])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_23_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N26), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[23])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_24_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N27), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[24])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_25_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N28), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[25])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_26_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N29), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[26])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_27_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N30), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[27])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_28_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N31), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[28])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_29_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N32), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[29])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_30_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N33), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[30])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_31_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N34), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[31])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_0_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N3), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_1_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N4), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_2_ ( 
        .D(n29225), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_3_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N6), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_4_ ( 
        .D(n29083), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_5_ ( 
        .D(n29224), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_6_ ( 
        .D(n29230), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_7_ ( 
        .D(n29223), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_8_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N11), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_9_ ( 
        .D(n29229), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_10_ ( 
        .D(n29228), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_11_ ( 
        .D(n29222), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_12_ ( 
        .D(n29084), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_13_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N16), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[13])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_14_ ( 
        .D(n29227), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_15_ ( 
        .D(n29226), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_16_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N19), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[16])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_17_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N20), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[17])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_18_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N21), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[18])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_19_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N22), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[19])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_20_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N23), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[20])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_21_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[21])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_22_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N25), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[22])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_23_ ( 
        .D(n29085), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_24_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N27), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[24])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_25_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N28), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[25])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_26_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N29), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[26])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_27_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N30), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[27])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_28_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N31), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[28])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_29_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N32), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[29])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_30_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N33), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[30])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_31_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N34), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[31])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rxd_s_reg ( .D(io_in[5]), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rxd_s) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rxd_r_reg ( .D(
        j202_soc_core_uart_TOP_rxd_s), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rxd_r) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1_reg_0_ ( 
        .D(io_in[22]), .CLK(wb_clk_i), .RESET_B(n29594), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2_reg_0_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[0]), .CLK(
        wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3_reg_0_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[0]), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1_reg_1_ ( 
        .D(io_in[23]), .CLK(wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2_reg_1_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[1]), .CLK(
        wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3_reg_1_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[1]), .CLK(
        wb_clk_i), .RESET_B(n12142), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1_reg_2_ ( 
        .D(io_in[24]), .CLK(wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2_reg_2_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[2]), .CLK(
        wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3_reg_2_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[2]), .CLK(
        wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1_reg ( 
        .D(n29076), .CLK(wb_clk_i), .RESET_B(n12142), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_2_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1), .CLK(
        wb_clk_i), .RESET_B(n12142), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_2) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_o_reg_2_ ( 
        .D(n138), .CLK(wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_bldc_core_00_hall_value[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status_reg_2_ ( 
        .D(j202_soc_core_bldc_core_00_hall_value[2]), .CLK(wb_clk_i), 
        .RESET_B(n29595), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_o_reg_0_ ( 
        .D(n137), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_hall_value[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status_reg_0_ ( 
        .D(j202_soc_core_bldc_core_00_hall_value[0]), .CLK(wb_clk_i), 
        .RESET_B(n29591), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_o_reg_1_ ( 
        .D(n136), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_bldc_core_00_hall_value[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status_reg_1_ ( 
        .D(j202_soc_core_bldc_core_00_hall_value[1]), .CLK(wb_clk_i), 
        .RESET_B(n29591), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_0_ ( 
        .D(n29008), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_1_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[1]), .CLK(
        wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_2_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[2]), .CLK(
        wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_3_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[3]), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_4_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[4]), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_5_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[5]), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_6_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[6]), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_7_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[7]), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_8_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[8]), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_9_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[9]), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_10_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[10]), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_11_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[11]), .CLK(
        wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_bootrom_00_sel_w_reg ( .D(n29505), 
        .CLK(wb_clk_i), .Q(j202_soc_core_bootrom_00_sel_w) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_ifetchl_reg ( .D(
        j202_soc_core_j22_cpu_ifetch), .DE(j202_soc_core_ahbcs_6__HREADY_), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ifetchl) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_area_reg_0_ ( .D(n10541), .DE(n10562), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ma_M_area[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aqu_st_reg_0_ ( .D(n29589), .DE(j202_soc_core_ahb2aqu_00_N95), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2aqu_00_aqu_st_0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_STB_ ( .D(
        n29114), .DE(j202_soc_core_ahb2aqu_00_N127), .CLK(wb_clk_i), .Q(
        j202_soc_core_aquc_STB_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_area_reg_1_ ( .D(n10540), .DE(n10562), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ma_M_area[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_WE_ ( .D(n12902), .DE(j202_soc_core_ahb2aqu_00_N95), .CLK(wb_clk_i), .Q(j202_soc_core_aquc_WE_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_state_reg_0_ ( 
        .D(n28915), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_1_ ( .D(
        n10567), .DE(n10563), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_opst[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rb__1_ ( 
        .D(n10582), .DE(n29117), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rb__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__2_ ( .D(
        j202_soc_core_ahb2aqu_00_N131), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_ADR__2_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_2_ ( 
        .D(j202_soc_core_aquc_ADR__2_), .CLK(wb_clk_i), .RESET_B(n29594), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_2_ ( .D(
        n29012), .DE(n29505), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__15_ ( 
        .D(n28983), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_15_ ( 
        .D(j202_soc_core_qspi_wb_wdat[15]), .CLK(wb_clk_i), .RESET_B(n29591), 
        .Q(j202_soc_core_bldc_core_00_wdata[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_15_ ( 
        .D(j202_soc_core_qspi_wb_wdat[15]), .CLK(wb_clk_i), .RESET_B(n29592), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_15_ ( 
        .D(n28927), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_15_ ( .D(
        j202_soc_core_ahb2apb_02_N143), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[47]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__7_ ( 
        .D(n10496), .DE(n10585), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__7_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__7_ ( .D(
        j202_soc_core_ahb2aqu_00_N136), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_ADR__7_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_7_ ( 
        .D(j202_soc_core_aquc_ADR__7_), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_7_ ( .D(
        n29010), .DE(n29506), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rn__3_ ( 
        .D(n10577), .DE(n29322), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rn__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__10_ ( 
        .D(n28978), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_10_ ( 
        .D(j202_soc_core_qspi_wb_wdat[10]), .CLK(wb_clk_i), .RESET_B(n29591), 
        .Q(j202_soc_core_bldc_core_00_wdata[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_10_ ( 
        .D(j202_soc_core_qspi_wb_wdat[10]), .CLK(wb_clk_i), .RESET_B(n29595), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_10_ ( 
        .D(n28928), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_10_ ( .D(
        j202_soc_core_ahb2apb_02_N138), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[42]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__0_ ( 
        .D(n10586), .DE(n10563), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__4_ ( .D(
        j202_soc_core_j22_cpu_ml_N195), .DE(j202_soc_core_ahbcs_6__HREADY_), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_M_macop_MAC_[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_Ma__1_ ( 
        .D(n10503), .DE(n10573), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_memop_Ma__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_4_ ( 
        .D(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_N487), .DE(n10562), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_20_ ( .D(
        j202_soc_core_j22_cpu_rf_N318), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__12_ ( 
        .D(n28980), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_12_ ( 
        .D(j202_soc_core_qspi_wb_wdat[12]), .CLK(wb_clk_i), .RESET_B(n12142), 
        .Q(j202_soc_core_bldc_core_00_wdata[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_12_ ( 
        .D(j202_soc_core_qspi_wb_wdat[12]), .CLK(wb_clk_i), .RESET_B(n29593), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__0_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__3_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_4_ ( 
        .D(n29059), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__4_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_6_ ( 
        .D(n29354), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__6_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__2_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_4_ ( 
        .D(n29069), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__4_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__1_ ( .D(
        n28950), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__2_ ( .D(
        n29326), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__3_ ( .D(
        n28921), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__7_ ( .D(
        n12727), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__7_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__10_ ( .D(
        n28971), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__10_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__11_ ( .D(
        n12175), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__11_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__12_ ( .D(
        n29328), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__12_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__15_ ( .D(
        n28917), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__15_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__0_ ( .D(
        n28926), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_v_ ( .D(n29357), 
        .DE(n10536), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_id_opn_v_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Wm__3_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N900), .DE(n10607), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_Wm__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_2_ ( .D(
        n10566), .DE(n10563), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_opst[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__4_ ( 
        .D(n10590), .DE(n10563), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_address_reg_1_ ( .D(
        n29033), .DE(n29347), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_address[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_1_ ( 
        .D(n10960), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_SEL__3_ ( .D(
        j202_soc_core_ahb2aqu_00_N164), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_SEL__3_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_1_ ( .D(n135), .CLK(
        wb_clk_i), .RESET_B(n29594), .Q(j202_soc_core_uart_div0[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__3_ ( .D(
        j202_soc_core_ahb2aqu_00_N132), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_ADR__3_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_3_ ( 
        .D(j202_soc_core_aquc_ADR__3_), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_3_ ( .D(
        n29013), .DE(n29506), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__8_ ( .D(
        n21914), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__8_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__0_ ( 
        .D(n10594), .DE(n29117), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_istall_reg ( .D(n10559), 
        .DE(n10608), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_istall) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_v_ ( .D(n28965), 
        .DE(j202_soc_core_ahbcs_6__HREADY_), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_v_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__0_ ( .D(
        n29036), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__1_ ( .D(
        n29071), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__2_ ( .D(
        n13272), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__3_ ( .D(
        n11767), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__6_ ( .D(
        n12617), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__6_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__7_ ( .D(
        n12472), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__7_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__8_ ( .D(
        n29015), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__8_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__9_ ( .D(
        n12376), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__9_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__10_ ( .D(
        n29077), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__10_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__11_ ( .D(
        n29009), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__11_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__12_ ( .D(
        n29524), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__12_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__15_ ( .D(
        n12757), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__15_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_30_ ( .D(
        j202_soc_core_j22_cpu_rf_N328), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_5_ ( 
        .D(n29323), .DE(n10562), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_2_ ( .D(
        n29012), .DE(n11125), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_3_ ( .D(
        n29013), .DE(n11125), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_7_ ( .D(
        n29010), .DE(n11125), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_18_ ( 
        .D(n28919), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_20_ ( 
        .D(n28918), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_req_reg ( .D(
        n10505), .DE(n29220), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_req) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_ack_reg ( .D(
        j202_soc_core_wbqspiflash_00_N730), .DE(
        j202_soc_core_wbqspiflash_00_N729), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_ack) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_stb_o_reg ( .D(n11125), 
        .DE(n10539), .CLK(wb_clk_i), .Q(j202_soc_core_ahb2wbqspi_00_stb_o) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_cyc_o_reg ( .D(n11125), 
        .DE(n10539), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_cyc) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_1_ ( .D(
        j202_soc_core_wbqspiflash_00_N725), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_hold_reg ( .D(
        j202_soc_core_wbqspiflash_00_N590), .DE(
        j202_soc_core_wbqspiflash_00_N745), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_hold) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_state_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N308), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N307), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_state[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_busy_reg ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N321), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_busy) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_write_in_progress_reg ( 
        .D(j202_soc_core_wbqspiflash_00_N709), .DE(
        j202_soc_core_wbqspiflash_00_N708), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_write_in_progress) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_31_ ( .D(
        n10506), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_2_ ( .D(
        j202_soc_core_wbqspiflash_00_N726), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_0_ ( .D(
        j202_soc_core_wbqspiflash_00_N724), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_len_reg_1_ ( .D(
        j202_soc_core_wbqspiflash_00_N737), .DE(
        j202_soc_core_wbqspiflash_00_N735), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_len[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N429), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_state_reg_1_ ( 
        .D(n29091), .DE(j202_soc_core_wbqspiflash_00_lldriver_N307), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_state_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N310), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N307), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_state[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_valid_reg ( 
        .D(n29056), .CLK(wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_valid)
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_sck_reg ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N312), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_sck) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_cs_n_reg ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N314), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N313), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_cs_n) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_write_protect_reg ( 
        .D(j202_soc_core_wbqspiflash_00_N722), .DE(
        j202_soc_core_wbqspiflash_00_N721), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_write_protect) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_28_ ( 
        .D(j202_soc_core_wbqspiflash_00_N695), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_0_ ( 
        .D(n11892), .DE(n10562), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_00_state_reg_0_ ( .D(
        j202_soc_core_ahb2apb_00_N89), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_00_state[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_00_state_reg_2_ ( .D(n29221), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2apb_00_state[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_00_state_reg_1_ ( .D(
        j202_soc_core_ahb2apb_00_N90), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_00_state[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_state_reg_1_ ( 
        .D(n28969), .CLK(wb_clk_i), .RESET_B(n12142), .Q(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_state_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_apb_00_nxt_state_0_), .CLK(wb_clk_i), 
        .RESET_B(n12142), .Q(j202_soc_core_cmt_core_00_cmt_apb_00_state[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_hwrite_buf_reg ( .D(
        j202_soc_core_ahb2apb_00_N55), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_pwrite[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_1_reg ( 
        .D(j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen), .CLK(wb_clk_i), 
        .RESET_B(n12142), .Q(j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_1)
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_2_reg ( 
        .D(j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_1), .CLK(wb_clk_i), 
        .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_2)
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_7_ ( .D(
        j202_soc_core_ahb2apb_00_N30), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_7_ ( 
        .D(j202_soc_core_paddr[6]), .CLK(wb_clk_i), .RESET_B(n12142), .Q(
        j202_soc_core_cmt_core_00_reg_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_3_ ( .D(
        j202_soc_core_ahb2apb_00_N26), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_3_ ( 
        .D(j202_soc_core_paddr[2]), .CLK(wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_cmt_core_00_reg_addr[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_2_ ( 
        .D(n10961), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_cmt_core_00_reg_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_00_N24), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_1_ ( 
        .D(j202_soc_core_paddr[1]), .CLK(wb_clk_i), .RESET_B(n12142), .Q(
        j202_soc_core_cmt_core_00_reg_addr[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_6_ ( 
        .D(n134), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_16_ ( 
        .D(n29359), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[16])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_16_ ( .D(
        j202_soc_core_ahb2apb_01_N144), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[80]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_16_ ( 
        .D(n28946), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_3_ ( 
        .D(n29065), .DE(n10562), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_CE__1_ ( .D(
        j202_soc_core_ahb2aqu_00_N98), .DE(j202_soc_core_ahb2aqu_00_N95), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_CE__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_19_ ( 
        .D(n28920), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_17_ ( 
        .D(j202_soc_core_qspi_wb_addr[19]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_dirty_sector_reg ( 
        .D(n28968), .DE(j202_soc_core_wbqspiflash_00_N719), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_dirty_sector) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_30_ ( 
        .D(j202_soc_core_wbqspiflash_00_N697), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__14_ ( .D(
        n12735), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__14_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_21_ ( .D(
        j202_soc_core_j22_cpu_rf_N319), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__13_ ( .D(
        n29329), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__13_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__13_ ( .D(
        n11646), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__13_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__14_ ( .D(
        n29327), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__14_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_14_ ( 
        .D(n29030), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_0_ ( .D(
        n29027), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__t_ ( .D(
        j202_soc_core_j22_cpu_rf_N2626), .DE(j202_soc_core_j22_cpu_rf_N2625), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__t_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_19_ ( .D(
        j202_soc_core_j22_cpu_rf_N317), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__11_ ( 
        .D(n28979), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_11_ ( 
        .D(j202_soc_core_qspi_wb_wdat[11]), .CLK(wb_clk_i), .RESET_B(n29592), 
        .Q(j202_soc_core_bldc_core_00_wdata[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_11_ ( 
        .D(j202_soc_core_qspi_wb_wdat[11]), .CLK(wb_clk_i), .RESET_B(n29593), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[11]), .CLK(
        wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cnt1[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[11]), .CLK(wb_clk_i), .RESET_B(
        n29592), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmf1_o_reg ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt1_to1), .CLK(
        wb_clk_i), .RESET_B(n12142), .Q(j202_soc_core_cmt_core_00_cmf1) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[9]), .CLK(wb_clk_i), .RESET_B(n29595), .Q(j202_soc_core_cmt_core_00_cnt1[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[9]), .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[9]), .CLK(wb_clk_i), 
        .RESET_B(n29592), .Q(j202_soc_core_prdata[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_9_ ( .D(
        j202_soc_core_ahb2apb_00_N137), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[105])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__9_ ( .D(
        n12771), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__9_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_9_ ( .D(
        n29032), .DE(n11125), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_9_ ( .D(
        n29032), .DE(n17160), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3204), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[455]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__14_ ( 
        .D(n28982), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_14_ ( 
        .D(j202_soc_core_qspi_wb_wdat[14]), .CLK(wb_clk_i), .RESET_B(n29592), 
        .Q(j202_soc_core_bldc_core_00_wdata[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_14_ ( 
        .D(j202_soc_core_qspi_wb_wdat[14]), .CLK(wb_clk_i), .RESET_B(n12142), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__i__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3390), .DE(j202_soc_core_j22_cpu_rf_N3391), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__i__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_6_ ( .D(
        j202_soc_core_ahb2apb_00_N29), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_6_ ( 
        .D(j202_soc_core_paddr[5]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_cmt_core_00_reg_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__6_ ( .D(
        j202_soc_core_ahb2aqu_00_N135), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_ADR__6_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_6_ ( 
        .D(j202_soc_core_aquc_ADR__6_), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_6_ ( .D(
        n29011), .DE(n11125), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_6_ ( .D(
        n29011), .DE(n17160), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_17_ ( 
        .D(n28922), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_17_ ( .D(
        n28922), .DE(n17160), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__5_ ( .D(
        n29072), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__5_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_5_ ( .D(
        j202_soc_core_ahb2apb_00_N28), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_5_ ( 
        .D(j202_soc_core_paddr[4]), .CLK(wb_clk_i), .RESET_B(n12142), .Q(
        j202_soc_core_cmt_core_00_reg_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__5_ ( .D(
        j202_soc_core_ahb2aqu_00_N134), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_ADR__5_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_5_ ( 
        .D(j202_soc_core_aquc_ADR__5_), .CLK(wb_clk_i), .RESET_B(n29594), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_5_ ( .D(
        n29035), .DE(n11125), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_5_ ( .D(
        n29035), .DE(n29506), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__4_ ( .D(
        n28923), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__4_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__4_ ( .D(
        n29075), .DE(n29116), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__4_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_MEM__1_ ( 
        .D(n10591), .DE(n10563), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_memop_MEM__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_MEM_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ma_N54), .DE(n10562), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_MEM[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_SEL__2_ ( .D(
        j202_soc_core_ahb2aqu_00_N163), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_SEL__2_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_1_ ( .D(n133), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_uart_div1[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_br_clr_reg ( .D(
        j202_soc_core_uart_BRG_N47), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_clr) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_x4_r_reg ( .D(
        j202_soc_core_uart_BRG_br_clr), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_sio_ce_x4_r) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_x4_t_reg ( .D(n29081), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_BRG_sio_ce_x4_t) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_x4_reg ( .D(
        j202_soc_core_uart_BRG_sio_ce_x4_t), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_sio_ce_x4) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_change_reg ( .D(
        j202_soc_core_uart_TOP_N102), .DE(j202_soc_core_uart_TOP_N101), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_change) );
  sky130_fd_sc_hd__dfstp_1 j202_soc_core_uart_TOP_dpll_state_reg_0_ ( .D(n132), 
        .CLK(wb_clk_i), .SET_B(n29593), .Q(
        j202_soc_core_uart_TOP_dpll_state[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_sio_ce_r1_reg ( .D(n29087), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_sio_ce_r1) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_sio_ce_r2_reg ( .D(
        j202_soc_core_uart_TOP_rx_sio_ce_r1), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_sio_ce_r2) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_sio_ce_reg ( .D(
        j202_soc_core_uart_TOP_N118), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_sio_ce) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_9_ ( .D(
        j202_soc_core_uart_TOP_rxd_s), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_8_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_7_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_6_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_5_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_4_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_3_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_2_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_bit_cnt_reg_0_ ( .D(
        n29232), .DE(j202_soc_core_uart_TOP_N85), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_bit_cnt[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_bit_cnt_reg_1_ ( .D(
        j202_soc_core_uart_TOP_N87), .DE(j202_soc_core_uart_TOP_N85), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_bit_cnt[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_bit_cnt_reg_2_ ( .D(
        j202_soc_core_uart_TOP_N88), .DE(j202_soc_core_uart_TOP_N85), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_bit_cnt[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_bit_cnt_reg_3_ ( .D(
        j202_soc_core_uart_TOP_N89), .DE(j202_soc_core_uart_TOP_N85), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_bit_cnt[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_go_reg ( .D(
        j202_soc_core_uart_TOP_N128), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_go) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_valid_reg ( .D(n10911), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_valid) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_valid_r_reg ( .D(
        j202_soc_core_uart_TOP_rx_valid), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_valid_r) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_rx_fifo_wp_reg_0_ ( .D(n131), 
        .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_uart_TOP_rx_fifo_wp[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_rx_fifo_wp_reg_1_ ( .D(n130), 
        .CLK(wb_clk_i), .RESET_B(n29594), .Q(
        j202_soc_core_uart_TOP_rx_fifo_wp[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__0_ ( .D(
        j202_soc_core_uart_TOP_rxr[2]), .DE(n29355), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__7_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(n29355), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__6_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(n29355), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__5_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(n29355), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__4_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(n29355), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__3_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(n29355), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__2_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(n29355), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__1_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(n29355), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__0_ ( .D(
        j202_soc_core_uart_TOP_rxr[2]), .DE(n29349), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__7_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(n29349), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__6_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(n29349), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__5_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(n29349), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__4_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(n29349), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__3_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(n29349), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__2_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(n29349), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__1_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(n29349), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__0_ ( .D(
        j202_soc_core_uart_TOP_rxr[2]), .DE(n29351), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__7_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(n29351), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__6_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(n29351), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__5_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(n29351), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__4_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(n29351), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__3_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(n29351), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__2_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(n29351), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__1_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(n29351), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__0_ ( .D(
        j202_soc_core_uart_TOP_rxr[2]), .DE(n29350), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__7_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(n29350), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__6_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(n29350), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__5_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(n29350), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__5_ ( .D(
        n29325), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__5_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__13_ ( 
        .D(n28981), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_13_ ( 
        .D(j202_soc_core_qspi_wb_wdat[13]), .CLK(wb_clk_i), .RESET_B(n29592), 
        .Q(j202_soc_core_bldc_core_00_wdata[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_13_ ( 
        .D(j202_soc_core_qspi_wb_wdat[13]), .CLK(wb_clk_i), .RESET_B(n29592), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__i__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3388), .DE(j202_soc_core_j22_cpu_rf_N3391), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__i__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N302), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_4_ ( .D(
        j202_soc_core_ahb2apb_00_N27), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_4_ ( 
        .D(j202_soc_core_paddr[3]), .CLK(wb_clk_i), .RESET_B(n12142), .Q(
        j202_soc_core_cmt_core_00_reg_addr[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_14_ ( 
        .D(n129), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_cmt_core_00_const0[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_13_ ( 
        .D(n128), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_const0[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_12_ ( 
        .D(n127), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_cmt_core_00_const0[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_11_ ( 
        .D(n126), .CLK(wb_clk_i), .RESET_B(n12142), .Q(
        j202_soc_core_cmt_core_00_const0[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_10_ ( 
        .D(n125), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_const0[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_15_ ( 
        .D(n124), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_const0[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_14_ ( 
        .D(n123), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_const1[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_13_ ( 
        .D(n122), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_const1[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_12_ ( 
        .D(n121), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_cmt_core_00_const1[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_11_ ( 
        .D(n120), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_const1[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_10_ ( 
        .D(n119), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_const1[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_15_ ( 
        .D(n118), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_cmt_core_00_const1[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__4_ ( .D(
        j202_soc_core_ahb2aqu_00_N133), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_ADR__4_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_4_ ( 
        .D(j202_soc_core_aquc_ADR__4_), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_4_ ( .D(
        n29034), .DE(n11125), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_4_ ( .D(
        n29034), .DE(n29506), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_31_ ( .D(
        j202_soc_core_j22_cpu_rf_N329), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_31_ ( .D(n12272), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__8_ ( .D(
        n29007), .DE(n29356), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_8_ ( 
        .D(j202_soc_core_qspi_wb_wdat[8]), .CLK(wb_clk_i), .RESET_B(n12142), 
        .Q(j202_soc_core_bldc_core_00_wdata[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_8_ ( 
        .D(j202_soc_core_qspi_wb_wdat[8]), .CLK(wb_clk_i), .RESET_B(n12142), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_8_ ( 
        .D(n117), .CLK(wb_clk_i), .RESET_B(n29594), .Q(
        j202_soc_core_cmt_core_00_const1[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_8_ ( 
        .D(n116), .CLK(wb_clk_i), .RESET_B(n29594), .Q(
        j202_soc_core_cmt_core_00_const0[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__i__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3386), .DE(j202_soc_core_j22_cpu_rf_N3391), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__i__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_6_ ( .D(
        j202_soc_core_j22_cpu_ml_N309), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_24_ ( 
        .D(n28924), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_len_reg_0_ ( .D(
        j202_soc_core_wbqspiflash_00_N736), .DE(
        j202_soc_core_wbqspiflash_00_N735), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_len[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_26_ ( 
        .D(n29165), .DE(j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_26_ ( .D(
        j202_soc_core_j22_cpu_rf_N324), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2671), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_28_ ( .D(n12271), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_30_ ( .D(n13336), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2674), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_16_ ( .D(
        n28946), .DE(n17160), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_14_ ( .D(
        n29030), .DE(n17160), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_6_ ( 
        .D(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_N497), .DE(n10562), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_29_ ( .D(
        j202_soc_core_j22_cpu_rf_N327), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_13_ ( .D(n24561), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_13_ ( 
        .D(n28947), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_13_ ( .D(
        n28947), .DE(n17160), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_1_ ( .D(
        n29028), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N301), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__3_ ( .D(
        n29002), .DE(n29356), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_3_ ( 
        .D(j202_soc_core_qspi_wb_wdat[3]), .CLK(wb_clk_i), .RESET_B(n29591), 
        .Q(j202_soc_core_bldc_core_00_wdata[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_3_ ( 
        .D(j202_soc_core_qspi_wb_wdat[3]), .CLK(wb_clk_i), .RESET_B(n29595), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_3_ ( 
        .D(n115), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_cmt_core_00_const1[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_3_ ( 
        .D(n114), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_const0[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_3_ ( 
        .D(n113), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_3_ ( 
        .D(n112), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_3_ ( .D(
        j202_soc_core_j22_cpu_id_idec_N894), .DE(n10563), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_opst[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_MEM__2_ ( 
        .D(n10592), .DE(n10563), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_memop_MEM__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_MEM_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ma_N55), .DE(n10562), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_MEM[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__5_ ( 
        .D(n10599), .DE(n29117), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_4_ ( .D(
        n10568), .DE(n10563), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_opst[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rs__0_ ( 
        .D(n29079), .DE(n29117), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rs__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_We__1_ ( 
        .D(n10603), .DE(n10607), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_We__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Wm__1_ ( 
        .D(n10601), .DE(n10607), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Wm__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_0_ ( .D(
        n10570), .DE(n10563), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_opst[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_MEM__3_ ( 
        .D(n10593), .DE(n10563), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_memop_MEM__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_MEM_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ma_N56), .DE(n10562), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_MEM[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_intack_reg ( .D(
        j202_soc_core_j22_cpu_id_idec_N822), .DE(n10565), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_intack) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intack_all_dout_reg_0_ ( 
        .D(n12071), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_cp_intack_all_0_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N3), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N4), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N5), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N6), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N9), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rte4_reg ( .D(
        j202_soc_core_j22_cpu_N8), .DE(n10565), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rte4) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Wm__2_ ( 
        .D(n10602), .DE(n10607), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Wm__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Wm__0_ ( 
        .D(n10600), .DE(n10607), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Wm__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_MEM__0_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N937), .DE(n10563), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_memop_MEM__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_MEM_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ma_N53), .DE(n10562), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_MEM[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Rn__3_ ( 
        .D(j202_soc_core_j22_cpu_regop_Rn__3_), .DE(n29362), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Rn__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Wm__0_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N956), .DE(n10561), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Wm__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Wm__3_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N959), .DE(n10561), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Wm__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Wm__2_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N958), .DE(n10561), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Wm__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Wm__1_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N957), .DE(n10561), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Wm__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__23_ ( 
        .D(n28992), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[23]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_23_ ( 
        .D(j202_soc_core_qspi_wb_wdat[23]), .CLK(wb_clk_i), .RESET_B(n29592), 
        .Q(j202_soc_core_bldc_core_00_wdata[23]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_7_ ( .D(n111), .CLK(
        wb_clk_i), .RESET_B(n29595), .Q(j202_soc_core_uart_div1[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__21_ ( 
        .D(n28990), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[21]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_21_ ( 
        .D(j202_soc_core_qspi_wb_wdat[21]), .CLK(wb_clk_i), .RESET_B(n29594), 
        .Q(j202_soc_core_bldc_core_00_wdata[21]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_5_ ( .D(n110), .CLK(
        wb_clk_i), .RESET_B(n29594), .Q(j202_soc_core_uart_div1[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__20_ ( 
        .D(n28989), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[20]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_20_ ( 
        .D(j202_soc_core_qspi_wb_wdat[20]), .CLK(wb_clk_i), .RESET_B(n29591), 
        .Q(j202_soc_core_bldc_core_00_wdata[20]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_4_ ( .D(n109), .CLK(
        wb_clk_i), .RESET_B(n29591), .Q(j202_soc_core_uart_div1[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__18_ ( 
        .D(n28986), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[18]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_18_ ( 
        .D(j202_soc_core_qspi_wb_wdat[18]), .CLK(wb_clk_i), .RESET_B(n29594), 
        .Q(j202_soc_core_bldc_core_00_wdata[18]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_2_ ( .D(n108), .CLK(
        wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_uart_div1[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__7_ ( .D(
        n29006), .DE(n29356), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_7_ ( 
        .D(j202_soc_core_qspi_wb_wdat[7]), .CLK(wb_clk_i), .RESET_B(n29592), 
        .Q(j202_soc_core_bldc_core_00_wdata[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_7_ ( 
        .D(j202_soc_core_qspi_wb_wdat[7]), .CLK(wb_clk_i), .RESET_B(n29595), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_7_ ( 
        .D(n107), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_cmt_core_00_const1[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_7_ ( 
        .D(n106), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_const0[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_nxt_latch_status_0_), 
        .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__6_ ( .D(
        n29005), .DE(n29356), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_6_ ( 
        .D(j202_soc_core_qspi_wb_wdat[6]), .CLK(wb_clk_i), .RESET_B(n29591), 
        .Q(j202_soc_core_bldc_core_00_wdata[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_6_ ( 
        .D(j202_soc_core_qspi_wb_wdat[6]), .CLK(wb_clk_i), .RESET_B(n29595), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_6_ ( 
        .D(n105), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_cmt_core_00_const1[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_6_ ( 
        .D(n104), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_cmt_core_00_const0[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_6_ ( 
        .D(n103), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_17_ ( 
        .D(n29360), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[17])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__5_ ( .D(
        n29004), .DE(n29356), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_5_ ( 
        .D(j202_soc_core_qspi_wb_wdat[5]), .CLK(wb_clk_i), .RESET_B(n29595), 
        .Q(j202_soc_core_bldc_core_00_wdata[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_5_ ( 
        .D(j202_soc_core_qspi_wb_wdat[5]), .CLK(wb_clk_i), .RESET_B(n29592), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_5_ ( 
        .D(n102), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_cmt_core_00_const1[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_5_ ( 
        .D(n101), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_cmt_core_00_const0[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_5_ ( 
        .D(n100), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_5_ ( 
        .D(n99), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__4_ ( .D(
        n29003), .DE(n29356), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_4_ ( 
        .D(j202_soc_core_qspi_wb_wdat[4]), .CLK(wb_clk_i), .RESET_B(n29593), 
        .Q(j202_soc_core_bldc_core_00_wdata[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_4_ ( 
        .D(j202_soc_core_qspi_wb_wdat[4]), .CLK(wb_clk_i), .RESET_B(n29593), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_4_ ( 
        .D(n98), .CLK(wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_cmt_core_00_const1[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_4_ ( 
        .D(n97), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_const0[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_4_ ( 
        .D(n96), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_4_ ( 
        .D(n95), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_pc_hold_reg ( .D(
        n10569), .DE(n10563), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_pc_hold) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_Ma__0_ ( 
        .D(n10504), .DE(n10573), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_memop_Ma__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_We__2_ ( 
        .D(n10579), .DE(n10607), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_We__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rn__2_ ( 
        .D(n10576), .DE(n29322), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rn__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Rn__2_ ( 
        .D(j202_soc_core_j22_cpu_regop_Rn__2_), .DE(n29362), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Rn__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rn__1_ ( 
        .D(n10575), .DE(n29322), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rn__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Rn__1_ ( 
        .D(j202_soc_core_j22_cpu_regop_Rn__1_), .DE(n29362), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Rn__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rn__0_ ( 
        .D(n10574), .DE(n29322), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rn__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Rn__0_ ( 
        .D(j202_soc_core_j22_cpu_regop_Rn__0_), .DE(n29362), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Rn__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__4_ ( 
        .D(n10598), .DE(n29117), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__3_ ( 
        .D(n10597), .DE(n29117), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__2_ ( 
        .D(n10596), .DE(n29117), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_We__3_ ( 
        .D(n12494), .DE(n10607), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_We__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3324), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3313), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3314), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3315), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3316), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3317), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3311), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3338), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3340), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3341), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3342), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3343), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2644), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2645), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2646), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2647), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2648), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2649), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2642), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3302), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3303), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3304), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3305), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3299), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3284), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3278), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3276), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3275), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3274), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3273), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3272), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3347), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3348), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3349), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3350), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3351), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3352), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3359), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3374), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3376), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3377), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3378), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3379), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2710), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2713), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2712), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2711), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2707), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2692), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2686), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2680), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2681), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2682), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2683), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2684), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2747), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[60]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2750), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[63]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2749), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[62]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2748), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[61]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2744), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[58]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2729), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[45]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2723), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[39]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2717), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[34]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2718), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[35]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2719), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[36]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2720), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[37]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2721), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[38]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2784), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[92]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2787), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[95]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2786), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[94]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2785), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[93]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2781), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[90]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2766), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[77]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2760), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[71]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2754), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[66]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2755), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[67]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2756), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[68]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2757), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[69]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2758), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[70]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2821), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[124]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2824), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[127]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2823), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[126]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2822), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[125]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2818), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[122]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2803), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[109]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2797), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[103]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2791), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[98]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2792), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[99]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2793), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[100]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2794), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[101]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2795), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[102]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2858), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[156]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2861), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[159]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2860), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[158]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2859), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[157]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2855), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[154]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2840), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[141]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2834), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[135]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2828), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[130]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2829), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[131]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2830), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[132]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2831), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[133]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2832), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[134]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2895), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[188]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2898), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[191]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2897), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[190]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2896), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[189]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2892), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[186]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2877), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[173]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2871), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[167]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2865), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[162]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2866), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[163]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2867), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[164]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2868), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[165]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2869), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[166]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2932), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[220]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2935), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[223]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2934), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[222]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2933), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[221]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2929), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[218]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2914), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[205]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2908), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[199]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2902), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[194]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2903), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[195]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2904), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[196]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2905), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[197]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2906), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[198]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2969), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[252]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2972), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[255]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2971), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[254]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2970), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[253]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2966), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[250]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2951), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[237]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2945), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[231]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2939), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[226]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2940), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[227]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2941), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[228]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2942), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[229]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2943), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[230]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3006), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[284]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3009), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[287]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3008), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[286]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3007), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[285]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3003), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[282]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2988), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[269]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2982), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[263]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2976), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[258]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2977), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[259]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2978), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[260]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2979), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[261]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2980), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[262]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3043), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[316]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3046), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[319]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3045), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[318]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3044), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[317]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3040), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[314]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3025), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[301]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3019), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[295]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3013), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[290]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3014), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[291]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3015), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[292]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3016), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[293]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3017), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[294]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3080), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[348]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3083), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[351]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3082), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[350]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3081), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[349]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3077), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[346]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3062), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[333]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3056), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[327]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3050), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[322]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3051), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[323]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3052), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[324]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3053), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[325]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3054), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[326]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3117), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[380]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3120), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[383]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3119), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[382]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3118), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[381]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3114), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[378]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3099), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[365]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3093), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[359]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3087), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[354]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3088), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[355]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3089), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[356]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3090), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[357]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3091), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[358]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3154), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[412]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3157), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[415]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3156), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[414]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3155), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[413]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3151), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[410]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3136), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[397]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3130), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[391]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3124), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[386]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3125), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[387]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3126), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[388]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3127), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[389]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3128), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[390]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3191), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[444]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3194), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[447]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3193), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[446]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3192), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[445]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3188), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[442]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3173), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[429]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3167), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[423]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3161), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[418]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3162), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[419]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3163), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[420]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3164), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[421]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3165), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[422]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3228), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[476]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3231), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[479]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3230), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[478]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3229), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[477]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3225), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[474]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3210), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[461]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3198), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[450]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3199), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[451]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3200), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[452]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3201), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[453]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3202), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[454]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3265), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[508]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3268), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[511]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3267), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[510]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3266), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[509]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3262), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[506]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3247), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[493]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3241), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[487]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3235), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[482]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3236), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[483]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3237), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[484]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3238), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[485]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3239), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[486]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__3_ ( 
        .D(n10589), .DE(n10563), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__2_ ( 
        .D(n10588), .DE(n10563), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__1_ ( 
        .D(n10587), .DE(n10563), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_2_ ( .D(
        j202_soc_core_j22_cpu_rf_N300), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_5_ ( .D(
        j202_soc_core_j22_cpu_rf_N303), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_6_ ( .D(
        j202_soc_core_j22_cpu_rf_N304), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_13_ ( .D(
        j202_soc_core_j22_cpu_rf_N311), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_28_ ( .D(
        j202_soc_core_j22_cpu_rf_N326), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Ra__1_ ( 
        .D(n10583), .DE(n29117), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Ra__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Ra__0_ ( 
        .D(n10606), .DE(n29117), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Ra__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rs__1_ ( 
        .D(n10605), .DE(n29117), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rs__1_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_req_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_req_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intr_req_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_00_N23), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_0_ ( 
        .D(j202_soc_core_paddr[0]), .CLK(wb_clk_i), .RESET_B(n12142), .Q(
        j202_soc_core_cmt_core_00_reg_addr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__0_ ( .D(
        n28964), .DE(j202_soc_core_ahb2aqu_00_N127), .CLK(wb_clk_i), .Q(
        j202_soc_core_aquc_ADR__0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_0_ ( 
        .D(j202_soc_core_aquc_ADR__0_), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_SEL__0_ ( .D(
        j202_soc_core_ahb2aqu_00_N161), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_SEL__0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_RDRXD1_reg ( .D(n29029), .CLK(
        wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_uart_RDRXD1) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_rx_fifo_rp_reg_0_ ( .D(n94), 
        .CLK(wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_uart_TOP_rx_fifo_rp[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_rx_fifo_rp_reg_1_ ( .D(n93), 
        .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_uart_TOP_rx_fifo_rp[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_gb_reg ( .D(
        j202_soc_core_uart_TOP_rx_fifo_N42), .DE(
        j202_soc_core_uart_TOP_rx_fifo_N41), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_gb) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_3_ ( .D(n92), .CLK(
        wb_clk_i), .RESET_B(n29591), .Q(j202_soc_core_uart_din_i[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_4_ ( .D(n91), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_uart_din_i[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_5_ ( .D(n90), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_uart_din_i[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_6_ ( .D(n89), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_uart_din_i[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_7_ ( .D(n88), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_uart_din_i[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_WRTXD1_reg ( .D(n28967), .CLK(
        wb_clk_i), .RESET_B(n29595), .Q(j202_soc_core_uart_WRTXD1) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_tx_fifo_wp_reg_0_ ( .D(n87), 
        .CLK(wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_uart_TOP_tx_fifo_wp[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_tx_fifo_wp_reg_1_ ( .D(n86), 
        .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_uart_TOP_tx_fifo_wp[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__7_ ( .D(
        j202_soc_core_uart_din_i[7]), .DE(n29346), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__6_ ( .D(
        j202_soc_core_uart_din_i[6]), .DE(n29346), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__5_ ( .D(
        j202_soc_core_uart_din_i[5]), .DE(n29346), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__4_ ( .D(
        j202_soc_core_uart_din_i[4]), .DE(n29346), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__3_ ( .D(
        j202_soc_core_uart_din_i[3]), .DE(n29346), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__7_ ( .D(
        j202_soc_core_uart_din_i[7]), .DE(n29344), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__6_ ( .D(
        j202_soc_core_uart_din_i[6]), .DE(n29344), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__5_ ( .D(
        j202_soc_core_uart_din_i[5]), .DE(n29344), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__4_ ( .D(
        j202_soc_core_uart_din_i[4]), .DE(n29344), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__3_ ( .D(
        j202_soc_core_uart_din_i[3]), .DE(n29344), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__7_ ( .D(
        j202_soc_core_uart_din_i[7]), .DE(n29352), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__6_ ( .D(
        j202_soc_core_uart_din_i[6]), .DE(n29352), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__5_ ( .D(
        j202_soc_core_uart_din_i[5]), .DE(n29352), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__4_ ( .D(
        j202_soc_core_uart_din_i[4]), .DE(n29352), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__3_ ( .D(
        j202_soc_core_uart_din_i[3]), .DE(n29352), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__7_ ( .D(
        j202_soc_core_uart_din_i[7]), .DE(n29345), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__6_ ( .D(
        j202_soc_core_uart_din_i[6]), .DE(n29345), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__5_ ( .D(
        j202_soc_core_uart_din_i[5]), .DE(n29345), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__4_ ( .D(
        j202_soc_core_uart_din_i[4]), .DE(n29345), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__3_ ( .D(
        j202_soc_core_uart_din_i[3]), .DE(n29345), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_address_reg_0_ ( .D(
        n29061), .DE(n29347), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_address[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3307), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3270), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2678), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3233), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[480]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2715), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[32]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2752), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[64]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2789), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[96]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2826), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[128]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2863), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[160]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2900), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[192]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2937), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[224]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2974), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[256]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3011), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[288]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3048), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[320]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3085), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[352]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3122), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[384]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3159), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[416]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3196), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[448]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_0_ ( .D(
        j202_soc_core_j22_cpu_rf_N298), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3345), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3370), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3335), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3296), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2704), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2741), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[55]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2778), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[87]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2815), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[119]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2852), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[151]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2889), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[183]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2926), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[215]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2963), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[247]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3000), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[279]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3037), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[311]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3074), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[343]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3111), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[375]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3148), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[407]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3185), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[439]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3222), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[471]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3259), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[503]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2667), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_23_ ( .D(
        j202_soc_core_j22_cpu_rf_N321), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3373), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3337), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3298), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2706), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2743), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[57]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2780), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[89]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2817), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[121]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2854), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[153]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2891), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[185]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2928), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[217]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2965), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[249]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3002), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[281]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3039), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[313]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3076), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[345]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3113), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[377]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3150), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[409]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3187), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[441]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3224), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[473]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3261), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[505]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2670), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_25_ ( .D(
        j202_soc_core_j22_cpu_rf_N323), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3355), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3319), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3280), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2688), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2725), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[41]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2762), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[73]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2799), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[105]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2836), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[137]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2873), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[169]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2910), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[201]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2947), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[233]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2984), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[265]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3021), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[297]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3058), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[329]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3095), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[361]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3132), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[393]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3169), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[425]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3206), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[457]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3243), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[489]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_9_ ( .D(n13329), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__m_ ( .D(
        j202_soc_core_j22_cpu_rf_N2640), .DE(j202_soc_core_j22_cpu_rf_N2639), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__m_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3309), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3271), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2679), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2716), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[33]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2753), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[65]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2790), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[97]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2827), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[129]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2864), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[161]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2901), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[193]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2938), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[225]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2975), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[257]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3012), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[289]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3049), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[321]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3086), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[353]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3123), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[385]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3160), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[417]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3197), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[449]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3234), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[481]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2643), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__s_ ( .D(
        j202_soc_core_j22_cpu_rf_N2628), .DE(j202_soc_core_j22_cpu_rf_N2627), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__s_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__0_ ( .D(
        j202_soc_core_j22_cpu_ml_N191), .DE(j202_soc_core_ahbcs_6__HREADY_), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__2_ ( .D(
        j202_soc_core_j22_cpu_ml_N193), .DE(j202_soc_core_ahbcs_6__HREADY_), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_M_macop_MAC_[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__3_ ( .D(
        j202_soc_core_j22_cpu_ml_N194), .DE(j202_soc_core_ahbcs_6__HREADY_), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_M_macop_MAC_[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__1_ ( .D(
        j202_soc_core_j22_cpu_ml_N192), .DE(j202_soc_core_ahbcs_6__HREADY_), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_6_ ( .D(n29321), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_mach[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_7_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[7]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_6_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[6]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ml_N303), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[0]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[0]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__0_ ( .D(
        n28977), .DE(n29356), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_0_ ( 
        .D(j202_soc_core_qspi_wb_wdat[0]), .CLK(wb_clk_i), .RESET_B(n12142), 
        .Q(j202_soc_core_bldc_core_00_wdata[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_0_ ( .D(n85), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_uart_din_i[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__0_ ( .D(
        j202_soc_core_uart_din_i[0]), .DE(n29345), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__0_ ( .D(
        j202_soc_core_uart_din_i[0]), .DE(n29352), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__0_ ( .D(
        j202_soc_core_uart_din_i[0]), .DE(n29344), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__0_ ( .D(
        j202_soc_core_uart_din_i[0]), .DE(n29346), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_0_ ( 
        .D(j202_soc_core_qspi_wb_wdat[0]), .CLK(wb_clk_i), .RESET_B(n29593), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_0_ ( 
        .D(n84), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_cmt_core_00_const1[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_0_ ( 
        .D(n83), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_cmt_core_00_const0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_0_ ( 
        .D(n82), .CLK(wb_clk_i), .RESET_B(n29594), .Q(
        j202_soc_core_cmt_core_00_cks1[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_0_ ( 
        .D(n81), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_cmt_core_00_cks0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmstr_reg_reg_o_reg_0_ ( 
        .D(n80), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_cmt_core_00_str0) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ml_N304), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[1]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[1]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ml_N305), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[2]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[2]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__2_ ( .D(
        n28999), .DE(n29356), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_2_ ( 
        .D(j202_soc_core_qspi_wb_wdat[2]), .CLK(wb_clk_i), .RESET_B(n29595), 
        .Q(j202_soc_core_bldc_core_00_wdata[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_2_ ( .D(n79), .CLK(
        wb_clk_i), .RESET_B(n29591), .Q(j202_soc_core_uart_din_i[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__2_ ( .D(
        j202_soc_core_uart_din_i[2]), .DE(n29345), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__2_ ( .D(
        j202_soc_core_uart_din_i[2]), .DE(n29352), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__2_ ( .D(
        j202_soc_core_uart_din_i[2]), .DE(n29344), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__2_ ( .D(
        j202_soc_core_uart_din_i[2]), .DE(n29346), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_2_ ( 
        .D(j202_soc_core_qspi_wb_wdat[2]), .CLK(wb_clk_i), .RESET_B(n29595), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_2_ ( 
        .D(n78), .CLK(wb_clk_i), .RESET_B(n29594), .Q(
        j202_soc_core_cmt_core_00_const1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_2_ ( 
        .D(n77), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_cmt_core_00_const0[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_2_ ( 
        .D(n76), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_2_ ( 
        .D(n75), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ml_N306), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[3]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[3]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_4_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[4]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_4_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[4]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_5_ ( .D(
        j202_soc_core_j22_cpu_ml_N308), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_5_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[5]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_5_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[5]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_7_ ( .D(
        j202_soc_core_j22_cpu_ml_N310), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_7_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[7]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_9_ ( .D(
        j202_soc_core_j22_cpu_ml_N312), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_9_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[9]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_9_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[9]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_13_ ( .D(
        j202_soc_core_j22_cpu_ml_N316), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_13_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[13]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_13_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[13]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_20_ ( .D(
        j202_soc_core_j22_cpu_ml_N359), .DE(n29119), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_4_ ( .D(
        j202_soc_core_j22_cpu_ml_N416), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_21_ ( .D(
        j202_soc_core_j22_cpu_ml_N360), .DE(n29119), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_5_ ( .D(
        j202_soc_core_j22_cpu_ml_N417), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_23_ ( .D(
        j202_soc_core_j22_cpu_ml_N362), .DE(n29119), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_7_ ( .D(
        j202_soc_core_j22_cpu_ml_N419), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_25_ ( .D(n12253), 
        .DE(n29119), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_9_ ( .D(
        j202_soc_core_j22_cpu_ml_N421), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_26_ ( .D(n12252), 
        .DE(n29119), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_28_ ( .D(
        j202_soc_core_j22_cpu_ml_N367), .DE(n29119), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_30_ ( .D(
        j202_soc_core_j22_cpu_ml_N369), .DE(n29119), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_19_ ( .D(
        j202_soc_core_j22_cpu_ml_N357), .DE(n29119), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ml_N415), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_18_ ( .D(
        j202_soc_core_j22_cpu_ml_N356), .DE(n29119), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ml_N414), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3364), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3328), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3289), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2697), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2734), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[49]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2771), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[81]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2808), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[113]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2845), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[145]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2882), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[177]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2919), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[209]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2956), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[241]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2993), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[273]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3030), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[305]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3067), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[337]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3104), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[369]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3141), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[401]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3178), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[433]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3215), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[465]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3252), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[497]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_17_ ( .D(n13334), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3366), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3330), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3291), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2699), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2736), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[51]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2773), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[83]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2810), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[115]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2847), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[147]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2884), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[179]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2921), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[211]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2958), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[243]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2995), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[275]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3032), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[307]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3069), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[339]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3106), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[371]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3143), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[403]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3180), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[435]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3217), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[467]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3254), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[499]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2663), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3375), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3339), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3300), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2708), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2745), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[59]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2782), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[91]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2819), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[123]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2856), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[155]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2893), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[187]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2930), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[219]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2967), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[251]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3004), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[283]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3041), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[315]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3078), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[347]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3115), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[379]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3152), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[411]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3189), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[443]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3226), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[475]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3263), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[507]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_27_ ( .D(n12270), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_27_ ( .D(n13277), 
        .DE(n29119), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_27_ ( .D(
        j202_soc_core_j22_cpu_rf_N325), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3357), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3322), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3282), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2690), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2727), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[43]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2764), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[75]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2801), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[107]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2838), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[139]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2875), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[171]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2912), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[203]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2949), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[235]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2986), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[267]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3023), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[299]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3060), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[331]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3097), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[363]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3134), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[395]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3171), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[427]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3208), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[459]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3245), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[491]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_11_ ( .D(n12267), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3358), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3323), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3283), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2691), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2728), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[44]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2765), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[76]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2802), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[108]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2839), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[140]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2876), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[172]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2913), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[204]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2950), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[236]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2987), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[268]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3024), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[300]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3061), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[332]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3098), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[364]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3135), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[396]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3172), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[428]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3209), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[460]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3246), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[492]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_12_ ( .D(n12256), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3360), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3325), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3286), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2694), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2731), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[46]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2768), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[78]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2805), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[110]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2842), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[142]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2879), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[174]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2916), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[206]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2953), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[238]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2990), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[270]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3027), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[302]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3064), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[334]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3101), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[366]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3138), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[398]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3175), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[430]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3212), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[462]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3249), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[494]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2657), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3369), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3334), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3295), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2703), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2740), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[54]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2777), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[86]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2814), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[118]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2851), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[150]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2888), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[182]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2925), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[214]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2962), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[246]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2999), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[278]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3036), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[310]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3073), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[342]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3110), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[374]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3147), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[406]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3184), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[438]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3221), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[470]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3258), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[502]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_22_ ( .D(n13322), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_22_ ( .D(
        j202_soc_core_j22_cpu_ml_N361), .DE(n29119), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_22_ ( .D(
        j202_soc_core_j22_cpu_rf_N320), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3372), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3336), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3297), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2705), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2742), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[56]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2779), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[88]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2816), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[120]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2853), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[152]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2890), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[184]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2927), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[216]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2964), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[248]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3001), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[280]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3038), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[312]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3075), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[344]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3112), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[376]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3149), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[408]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3186), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[440]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3223), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[472]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3260), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[504]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_24_ ( .D(n29115), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_24_ ( .D(
        j202_soc_core_j22_cpu_ml_N363), .DE(n29119), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_24_ ( .D(
        j202_soc_core_j22_cpu_rf_N322), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3354), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3318), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3279), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2687), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2724), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[40]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2761), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[72]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2798), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[104]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2835), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[136]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2872), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[168]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2909), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[200]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2946), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[232]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2983), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[264]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3020), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[296]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3057), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[328]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3094), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[360]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3131), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[392]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3168), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[424]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3205), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[456]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3242), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[488]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_8_ ( .D(n12268), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3356), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3321), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3281), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2689), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2726), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[42]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2763), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[74]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2800), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[106]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2837), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[138]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2874), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[170]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2911), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[202]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2948), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[234]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2985), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[266]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3022), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[298]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3059), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[330]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3096), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[362]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3133), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[394]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3170), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[426]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3207), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[458]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3244), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[490]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2653), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_10_ ( .D(
        j202_soc_core_j22_cpu_ml_N313), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_10_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[10]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_10_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[10]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_10_ ( .D(
        j202_soc_core_j22_cpu_ml_N422), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N308), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_10_ ( 
        .D(n29063), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_10_ ( .D(
        n29063), .DE(n29505), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3363), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3327), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3288), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2696), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2733), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[48]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2770), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[80]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2807), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[112]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2844), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[144]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2881), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[176]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2918), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[208]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2955), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[240]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2992), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[272]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3029), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[304]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3066), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[336]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3103), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[368]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3140), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[400]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3177), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[432]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3214), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[464]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3251), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[496]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_16_ ( .D(n13331), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3361), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3326), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3287), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2695), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2732), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[47]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2769), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[79]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2806), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[111]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2843), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[143]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2880), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[175]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2917), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[207]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2954), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[239]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2991), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[271]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3028), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[303]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3065), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[335]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3102), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[367]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3139), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[399]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3176), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[431]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3213), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[463]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3250), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[495]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2658), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_15_ ( .D(
        j202_soc_core_j22_cpu_ml_N318), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_15_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[15]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_15_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[15]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_18_ ( .D(
        j202_soc_core_j22_cpu_ml_N321), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_18_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[18]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_18_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[18]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_19_ ( .D(
        j202_soc_core_j22_cpu_ml_N322), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_19_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[19]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_19_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[19]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_20_ ( .D(
        j202_soc_core_j22_cpu_ml_N324), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_20_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[20]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_20_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[20]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_21_ ( .D(
        j202_soc_core_j22_cpu_ml_N325), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_21_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[21]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_21_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[21]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_22_ ( .D(
        j202_soc_core_j22_cpu_ml_N326), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_22_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[22]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_22_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[22]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__22_ ( 
        .D(n28991), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[22]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_22_ ( 
        .D(j202_soc_core_qspi_wb_wdat[22]), .CLK(wb_clk_i), .RESET_B(n29592), 
        .Q(j202_soc_core_bldc_core_00_wdata[22]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_6_ ( .D(n74), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_uart_div1[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_23_ ( .D(
        j202_soc_core_j22_cpu_ml_N327), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_23_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[23]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_23_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[23]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_24_ ( .D(
        j202_soc_core_j22_cpu_ml_N328), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_24_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[24]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_24_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[24]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_25_ ( .D(
        j202_soc_core_j22_cpu_ml_N329), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_25_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[25]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_25_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[25]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_26_ ( .D(
        j202_soc_core_j22_cpu_ml_N330), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_26_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[26]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_26_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[26]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__26_ ( 
        .D(n28995), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[26]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_2_ ( .D(n73), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_uart_div0[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_27_ ( .D(
        j202_soc_core_j22_cpu_ml_N331), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_27_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[27]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_27_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[27]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_28_ ( .D(
        j202_soc_core_j22_cpu_ml_N332), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_28_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[28]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_28_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[28]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_29_ ( .D(
        j202_soc_core_j22_cpu_ml_N333), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_29_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[29]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_29_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[29]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__29_ ( 
        .D(n28998), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[29]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_5_ ( .D(n72), .CLK(
        wb_clk_i), .RESET_B(n29595), .Q(j202_soc_core_uart_div0[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_30_ ( .D(
        j202_soc_core_j22_cpu_ml_N334), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_30_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[30]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_30_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[30]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_31_ ( .D(
        j202_soc_core_j22_cpu_ml_N335), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_31_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[31]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_31_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[31]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_32_ ( .D(
        j202_soc_core_j22_cpu_ml_N336), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[32]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_15_ ( .D(
        j202_soc_core_j22_cpu_rf_N313), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__31_ ( 
        .D(n29001), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[31]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_7_ ( .D(n71), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_uart_div0[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_3_ ( .D(
        j202_soc_core_wbqspiflash_00_N727), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_9_ ( 
        .D(j202_soc_core_wbqspiflash_00_N623), .DE(n29120), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_N614), .DE(n29120), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_8_ ( 
        .D(j202_soc_core_wbqspiflash_00_N622), .DE(n29120), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_N621), .DE(n29120), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_N620), .DE(n29120), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_N619), .DE(n29120), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_N618), .DE(n29120), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_N617), .DE(n29120), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_N616), .DE(n29120), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_N615), .DE(n29120), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_reset_counter[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_alt_ctrl_reg ( .D(
        j202_soc_core_wbqspiflash_00_N86), .DE(n29593), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_alt_ctrl) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_alt_cmd_reg ( .D(
        j202_soc_core_wbqspiflash_00_N85), .DE(n29593), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_alt_cmd) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_ctrl_reg ( .D(
        n28966), .DE(j202_soc_core_wbqspiflash_00_N743), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_ctrl) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_wr_reg ( .D(
        j202_soc_core_wbqspiflash_00_N734), .DE(
        j202_soc_core_wbqspiflash_00_N733), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_wr) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_0_ ( 
        .D(j202_soc_core_qspi_wb_addr[2]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_18_ ( 
        .D(j202_soc_core_qspi_wb_addr[20]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_16_ ( 
        .D(j202_soc_core_qspi_wb_addr[18]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_15_ ( 
        .D(j202_soc_core_qspi_wb_addr[17]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_14_ ( 
        .D(j202_soc_core_qspi_wb_addr[16]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_12_ ( 
        .D(j202_soc_core_qspi_wb_addr[14]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_11_ ( 
        .D(j202_soc_core_qspi_wb_addr[13]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_8_ ( 
        .D(j202_soc_core_qspi_wb_addr[10]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_7_ ( 
        .D(j202_soc_core_qspi_wb_addr[9]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_5_ ( 
        .D(j202_soc_core_qspi_wb_addr[7]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_4_ ( 
        .D(j202_soc_core_qspi_wb_addr[6]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_3_ ( 
        .D(j202_soc_core_qspi_wb_addr[5]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_2_ ( 
        .D(j202_soc_core_qspi_wb_addr[4]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_1_ ( 
        .D(j202_soc_core_qspi_wb_addr[3]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_4_ ( .D(
        j202_soc_core_wbqspiflash_00_N728), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_spd_reg ( .D(
        j202_soc_core_wbqspiflash_00_N592), .DE(
        j202_soc_core_wbqspiflash_00_N746), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_spd) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_spd_reg ( 
        .D(j202_soc_core_wbqspiflash_00_spi_spd), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N423), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_mod_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N356), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N354), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N358), .DE(n29237), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_interrupt_reg ( .D(
        j202_soc_core_wbqspiflash_00_N741), .DE(
        j202_soc_core_wbqspiflash_00_N740), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_int) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_20_ ( 
        .D(n29057), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[20])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N323), .DE(n29113), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N359), .DE(n29237), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N324), .DE(n29113), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N360), .DE(n29237), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N325), .DE(n29113), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N361), .DE(n29237), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N326), .DE(n29113), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_4_ ( 
        .D(n29216), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_4_ ( 
        .D(n29184), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_5_ ( 
        .D(n29205), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_5_ ( 
        .D(n29183), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_6_ ( 
        .D(n29215), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_6_ ( 
        .D(n29192), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_7_ ( 
        .D(n29199), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_7_ ( 
        .D(n29191), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_8_ ( 
        .D(n29198), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_8_ ( 
        .D(n29182), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_9_ ( 
        .D(n29202), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_9_ ( 
        .D(n29181), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_10_ ( 
        .D(n29197), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_10_ ( 
        .D(n29180), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_11_ ( 
        .D(n29201), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_11_ ( 
        .D(n29179), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_12_ ( 
        .D(n29218), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_12_ ( 
        .D(n29178), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_13_ ( 
        .D(n29219), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_13_ ( 
        .D(n29177), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_14_ ( 
        .D(n29214), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_14_ ( 
        .D(n29190), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_15_ ( 
        .D(n29200), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_15_ ( 
        .D(n29189), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_16_ ( 
        .D(n29196), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_16_ ( 
        .D(n29188), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_17_ ( 
        .D(n29213), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_17_ ( 
        .D(n29176), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_18_ ( 
        .D(n29195), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_18_ ( 
        .D(n29175), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_19_ ( 
        .D(n29212), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_19_ ( 
        .D(n29174), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_20_ ( 
        .D(n29211), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_20_ ( 
        .D(n29187), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_21_ ( 
        .D(n29194), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_21_ ( 
        .D(n29173), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_22_ ( 
        .D(n29210), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_22_ ( 
        .D(n29186), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_23_ ( 
        .D(n29217), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_23_ ( 
        .D(n29172), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_24_ ( 
        .D(n29193), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_24_ ( 
        .D(n29185), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_25_ ( 
        .D(n29209), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_25_ ( 
        .D(n29171), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_26_ ( 
        .D(n29208), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_26_ ( 
        .D(n29170), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_27_ ( 
        .D(n29207), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_27_ ( 
        .D(n29169), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_28_ ( 
        .D(n29206), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_28_ ( 
        .D(n29168), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_29_ ( 
        .D(n29204), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_29_ ( 
        .D(n29167), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_30_ ( 
        .D(n29203), .DE(n29237), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_out[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_30_ ( 
        .D(n29166), .DE(n29113), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_31_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N389), .DE(n29237), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_dir_reg ( .D(
        j202_soc_core_wbqspiflash_00_N594), .DE(
        j202_soc_core_wbqspiflash_00_N747), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_dir) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_dir_reg ( 
        .D(j202_soc_core_wbqspiflash_00_spi_dir), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N423), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_dir) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_mod_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N355), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N354), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_cmd_reg ( .D(
        j202_soc_core_wbqspiflash_00_N663), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_cmd) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_31_ ( 
        .D(j202_soc_core_qspi_wb_wdat[31]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_29_ ( 
        .D(j202_soc_core_qspi_wb_wdat[29]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_26_ ( 
        .D(j202_soc_core_qspi_wb_wdat[26]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_23_ ( 
        .D(j202_soc_core_qspi_wb_wdat[23]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_22_ ( 
        .D(j202_soc_core_qspi_wb_wdat[22]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_21_ ( 
        .D(j202_soc_core_qspi_wb_wdat[21]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_N718), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_20_ ( 
        .D(j202_soc_core_qspi_wb_wdat[20]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_N717), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_18_ ( 
        .D(j202_soc_core_qspi_wb_wdat[18]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_N715), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_15_ ( 
        .D(j202_soc_core_qspi_wb_wdat[15]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_N712), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_14_ ( 
        .D(j202_soc_core_qspi_wb_wdat[14]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_N711), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_13_ ( 
        .D(j202_soc_core_qspi_wb_wdat[13]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_12_ ( 
        .D(j202_soc_core_qspi_wb_wdat[12]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_10_ ( 
        .D(j202_soc_core_qspi_wb_wdat[10]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_8_ ( 
        .D(j202_soc_core_qspi_wb_wdat[8]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_7_ ( 
        .D(j202_soc_core_qspi_wb_wdat[7]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_6_ ( 
        .D(j202_soc_core_qspi_wb_wdat[6]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_6_ ( .D(
        n10531), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_5_ ( 
        .D(j202_soc_core_qspi_wb_wdat[5]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_4_ ( 
        .D(j202_soc_core_qspi_wb_wdat[4]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_4_ ( .D(
        n10533), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_3_ ( 
        .D(j202_soc_core_qspi_wb_wdat[3]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_2_ ( 
        .D(j202_soc_core_qspi_wb_wdat[2]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_2_ ( .D(
        n10535), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_0_ ( 
        .D(j202_soc_core_qspi_wb_wdat[0]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_0_ ( .D(
        j202_soc_core_wbqspiflash_00_N628), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_N611), .DE(
        j202_soc_core_wbqspiflash_00_N750), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_N612), .DE(
        j202_soc_core_wbqspiflash_00_N750), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_N605), .DE(n29358), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_last_status[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_N607), .DE(n29358), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_last_status[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_N608), .DE(n29358), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_last_status[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_N609), .DE(n29358), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_last_status[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_N613), .DE(n29358), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_last_status[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_N667), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_3_ ( .D(
        n10534), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_29_ ( 
        .D(j202_soc_core_wbqspiflash_00_N696), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_31_ ( 
        .D(j202_soc_core_wbqspiflash_00_N698), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_15_ ( 
        .D(n29031), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_13_ ( 
        .D(j202_soc_core_qspi_wb_addr[15]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_15_ ( .D(
        n29031), .DE(n29505), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3365), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3329), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3290), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2698), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2735), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[50]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2772), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[82]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2809), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[114]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2846), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[146]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2883), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[178]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2920), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[210]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2957), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[242]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2994), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[274]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3031), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[306]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3068), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[338]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3105), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[370]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3142), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[402]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3179), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[434]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3216), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[466]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3253), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[498]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2662), .DE(n29235), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_16_ ( .D(
        j202_soc_core_j22_cpu_ml_N319), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_16_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[16]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_16_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[16]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_16_ ( .D(
        j202_soc_core_j22_cpu_ml_N354), .DE(n29119), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ml_N412), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_16_ ( .D(
        j202_soc_core_j22_cpu_rf_N314), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__16_ ( 
        .D(n28984), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[16]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_16_ ( 
        .D(j202_soc_core_qspi_wb_wdat[16]), .CLK(wb_clk_i), .RESET_B(n29591), 
        .Q(j202_soc_core_bldc_core_00_wdata[16]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_0_ ( .D(n70), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_uart_div1[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_16_ ( 
        .D(j202_soc_core_qspi_wb_wdat[16]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_N713), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_8_ ( .D(
        j202_soc_core_j22_cpu_ml_N311), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_8_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[8]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_8_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[8]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__q_ ( .D(
        j202_soc_core_j22_cpu_rf_N2638), .DE(j202_soc_core_j22_cpu_rf_N2637), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__q_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_8_ ( .D(
        j202_soc_core_j22_cpu_ml_N420), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_8_ ( .D(
        j202_soc_core_j22_cpu_rf_N306), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__24_ ( 
        .D(n28993), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[24]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_0_ ( .D(n69), .CLK(
        wb_clk_i), .RESET_B(n12142), .Q(j202_soc_core_uart_div0[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_24_ ( 
        .D(j202_soc_core_qspi_wb_wdat[24]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_8_ ( .D(
        n29064), .DE(n11125), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_6_ ( 
        .D(j202_soc_core_qspi_wb_addr[8]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_8_ ( .D(
        n10529), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_8_ ( .D(
        n29064), .DE(n29505), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_CE__0_ ( .D(
        n29588), .DE(j202_soc_core_ahb2aqu_00_N95), .CLK(wb_clk_i), .Q(
        j202_soc_core_aquc_CE__0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_state_reg_1_ ( 
        .D(n29231), .CLK(wb_clk_i), .RESET_B(n12142), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_22_ ( 
        .D(n68), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_21_ ( 
        .D(n67), .CLK(wb_clk_i), .RESET_B(n29594), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_20_ ( 
        .D(n66), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_18_ ( 
        .D(n65), .CLK(wb_clk_i), .RESET_B(n29594), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_16_ ( 
        .D(n64), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_15_ ( 
        .D(n63), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_14_ ( 
        .D(n62), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_13_ ( 
        .D(n61), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_12_ ( 
        .D(n60), .CLK(wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_11_ ( 
        .D(n59), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_bldc_core_00_pwm_period[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_10_ ( 
        .D(n58), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_pwm_period[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_8_ ( 
        .D(n57), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_pwm_period[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_7_ ( 
        .D(n56), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_bldc_core_00_pwm_period[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_6_ ( 
        .D(n55), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_bldc_core_00_pwm_period[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_5_ ( 
        .D(n54), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_bldc_core_00_pwm_period[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_4_ ( 
        .D(n53), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_bldc_core_00_pwm_period[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_3_ ( 
        .D(n52), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_pwm_period[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_2_ ( 
        .D(n51), .CLK(wb_clk_i), .RESET_B(n29594), .Q(
        j202_soc_core_bldc_core_00_pwm_period[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_0_ ( 
        .D(n50), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_pwm_period[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_23_ ( 
        .D(n49), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bcr_00_reg_o_reg_0_ ( 
        .D(n48), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_pwm_en) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ccr_00_reg_o_reg_0_ ( 
        .D(n47), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_bldc_core_00_comm[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ccr_00_reg_o_reg_2_ ( 
        .D(n46), .CLK(wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_bldc_core_00_comm[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_00_reg_o_reg_0_ ( 
        .D(n45), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_wen_1_reg ( 
        .D(n29050), .CLK(wb_clk_i), .RESET_B(n12142), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_wen) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_00_reg_o_reg_0_ ( 
        .D(n44), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_reg_0_ ( 
        .D(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_nxt_latch_status_0_), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bldc_int_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_nxt_bldc_int), 
        .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_bldc_int) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_19_ ( 
        .D(n29051), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[19])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_14_ ( .D(
        j202_soc_core_j22_cpu_ml_N317), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_14_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[14]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_14_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[14]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_14_ ( .D(
        j202_soc_core_j22_cpu_ml_N426), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_14_ ( .D(
        j202_soc_core_j22_cpu_rf_N312), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__30_ ( 
        .D(n29000), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[30]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_6_ ( .D(n43), .CLK(
        wb_clk_i), .RESET_B(n29595), .Q(j202_soc_core_uart_div0[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_30_ ( 
        .D(j202_soc_core_qspi_wb_wdat[30]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3367), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3331), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3292), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2700), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2737), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[52]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2774), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[84]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2811), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[116]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2848), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[148]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2885), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[180]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2922), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[212]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2959), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[244]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2996), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[276]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3033), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[308]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3070), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[340]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3107), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[372]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3144), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[404]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3181), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[436]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3218), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[468]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3255), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[500]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_20_ ( .D(n13344), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_12_ ( .D(
        j202_soc_core_j22_cpu_ml_N315), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_12_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[12]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_12_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[12]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_12_ ( .D(
        j202_soc_core_j22_cpu_ml_N424), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_12_ ( .D(
        j202_soc_core_j22_cpu_rf_N310), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__28_ ( 
        .D(n28997), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[28]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_4_ ( .D(n42), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_uart_div0[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_28_ ( 
        .D(j202_soc_core_qspi_wb_wdat[28]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_02_state_reg_0_ ( .D(n11082), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2apb_02_state[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_02_state_reg_2_ ( .D(
        j202_soc_core_ahb2apb_02_N91), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_02_state[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_02_state_reg_1_ ( .D(
        j202_soc_core_ahb2apb_02_N90), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_02_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_2_ ( 
        .D(n12899), .DE(n10562), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_0_ ( .D(
        n29581), .DE(n12491), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_hsize_buf_reg_1_ ( .D(
        n29590), .DE(n12492), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_02_hsize_buf[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_hsize_buf_reg_0_ ( .D(
        n29578), .DE(n12491), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_02_hsize_buf[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_hwrite_buf_reg ( .D(
        n29489), .DE(n12492), .CLK(wb_clk_i), .Q(j202_soc_core_pwrite[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_7_ ( .D(
        n29579), .DE(n12491), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_6_ ( .D(
        n29584), .DE(n12492), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_5_ ( .D(
        n11081), .DE(n12491), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_4_ ( .D(
        n29582), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_3_ ( .D(
        n29583), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_2_ ( .D(
        n29580), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_1_ ( .D(
        n29575), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_31_ ( 
        .D(n29055), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_30_ ( 
        .D(n28929), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_29_ ( 
        .D(n28930), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_28_ ( 
        .D(n29054), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_26_ ( 
        .D(n28931), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_24_ ( 
        .D(n28932), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_23_ ( 
        .D(n28933), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_22_ ( 
        .D(n28934), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_21_ ( 
        .D(n28935), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_20_ ( 
        .D(n28936), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_18_ ( 
        .D(n28937), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_16_ ( 
        .D(n28938), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_15_ ( 
        .D(n28927), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_12_ ( 
        .D(n28939), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_10_ ( 
        .D(n28928), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_8_ ( 
        .D(n28940), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_7_ ( 
        .D(n28941), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_6_ ( 
        .D(n28942), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_5_ ( 
        .D(n28943), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_4_ ( 
        .D(n28944), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_2_ ( 
        .D(n28945), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_0_ ( 
        .D(n29086), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_31_ ( 
        .D(n29055), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_30_ ( 
        .D(n28929), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_29_ ( 
        .D(n28930), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_28_ ( 
        .D(n29054), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_26_ ( 
        .D(n28931), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_24_ ( 
        .D(n28932), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_23_ ( 
        .D(n28933), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_22_ ( 
        .D(n28934), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_21_ ( 
        .D(n28935), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_20_ ( 
        .D(n28936), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_18_ ( 
        .D(n28937), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_16_ ( 
        .D(n28938), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_15_ ( 
        .D(n28927), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_12_ ( 
        .D(n28939), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_10_ ( 
        .D(n28928), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_8_ ( 
        .D(n28940), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_7_ ( 
        .D(n28941), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_6_ ( 
        .D(n28942), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_5_ ( 
        .D(n28943), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_4_ ( 
        .D(n28944), .DE(n29315), .CLK(wb_clk_i), .Q(la_data_out[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_2_ ( 
        .D(n28945), .DE(n10676), .CLK(wb_clk_i), .Q(la_data_out[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_0_ ( 
        .D(n29086), .DE(n10676), .CLK(wb_clk_i), .Q(la_data_out[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_31_ ( 
        .D(n29055), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_30_ ( 
        .D(n28929), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_29_ ( 
        .D(n28930), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_28_ ( 
        .D(n29054), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_26_ ( 
        .D(n28931), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_24_ ( 
        .D(n28932), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_23_ ( 
        .D(n28933), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_22_ ( 
        .D(n28934), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_21_ ( 
        .D(n28935), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_20_ ( 
        .D(n28936), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_18_ ( 
        .D(n28937), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_16_ ( 
        .D(n28938), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_15_ ( 
        .D(n28927), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_12_ ( 
        .D(n28939), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_10_ ( 
        .D(n28928), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_8_ ( 
        .D(n28940), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_7_ ( 
        .D(n28941), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_6_ ( 
        .D(n28942), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_5_ ( 
        .D(n28943), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_4_ ( 
        .D(n28944), .DE(n29316), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_2_ ( 
        .D(n28945), .DE(n10674), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_0_ ( 
        .D(n29086), .DE(n10674), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_10_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N50), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_15_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N55), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_31_ ( 
        .D(n29055), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_31_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N71), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_31_ ( .D(
        j202_soc_core_ahb2apb_02_N159), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[63]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_30_ ( 
        .D(n28929), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_30_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N70), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_30_ ( .D(
        j202_soc_core_ahb2apb_02_N158), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[62]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_29_ ( 
        .D(n28930), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_29_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N69), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_29_ ( .D(
        j202_soc_core_ahb2apb_02_N157), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[61]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_28_ ( 
        .D(n29054), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_28_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N68), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_28_ ( .D(
        j202_soc_core_ahb2apb_02_N156), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[60]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_26_ ( 
        .D(n28931), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_26_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N66), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_26_ ( .D(
        j202_soc_core_ahb2apb_02_N154), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[58]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_24_ ( 
        .D(n28932), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_24_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N64), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_24_ ( .D(
        j202_soc_core_ahb2apb_02_N152), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[56]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_23_ ( 
        .D(n28933), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_23_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N63), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_23_ ( .D(
        j202_soc_core_ahb2apb_02_N151), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[55]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_22_ ( 
        .D(n28934), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_22_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N62), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_22_ ( .D(
        j202_soc_core_ahb2apb_02_N150), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[54]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_21_ ( 
        .D(n28935), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_21_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N61), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_21_ ( .D(
        j202_soc_core_ahb2apb_02_N149), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[53]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_20_ ( 
        .D(n28936), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_20_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N60), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_20_ ( .D(
        j202_soc_core_ahb2apb_02_N148), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[52]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_18_ ( 
        .D(n28937), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_18_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N58), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_18_ ( .D(
        j202_soc_core_ahb2apb_02_N146), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[50]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_16_ ( 
        .D(n28938), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_16_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N56), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_16_ ( .D(
        j202_soc_core_ahb2apb_02_N144), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[48]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_12_ ( 
        .D(n28939), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_12_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N52), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_12_ ( .D(
        j202_soc_core_ahb2apb_02_N140), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[44]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_8_ ( 
        .D(n28940), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_8_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N48), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_8_ ( .D(
        j202_soc_core_ahb2apb_02_N136), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[40]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_7_ ( 
        .D(n28941), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_7_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N47), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_7_ ( .D(
        j202_soc_core_ahb2apb_02_N135), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[39]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_6_ ( 
        .D(n28942), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_6_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N46), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_6_ ( .D(
        j202_soc_core_ahb2apb_02_N134), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[38]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_5_ ( 
        .D(n28943), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_5_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N45), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_5_ ( .D(
        j202_soc_core_ahb2apb_02_N133), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[37]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_4_ ( 
        .D(n28944), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_4_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N44), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_4_ ( .D(
        j202_soc_core_ahb2apb_02_N132), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[36]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_2_ ( 
        .D(n28945), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_2_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N42), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_2_ ( .D(
        j202_soc_core_ahb2apb_02_N130), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[34]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_0_ ( 
        .D(n29086), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N40), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_02_N128), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[32]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_1_ ( 
        .D(n29067), .DE(n10562), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_01_state_reg_0_ ( .D(n12274), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2apb_01_state[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_01_state_reg_2_ ( .D(
        j202_soc_core_ahb2apb_01_N91), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_01_state[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_01_state_reg_1_ ( .D(
        j202_soc_core_ahb2apb_01_N90), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_01_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_0_ ( .D(
        n12266), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_hsize_buf_reg_1_ ( .D(
        n12265), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_01_hsize_buf[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_hsize_buf_reg_0_ ( .D(
        n12228), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_01_hsize_buf[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_hwrite_buf_reg ( .D(
        n12236), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_pwrite[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_10_ ( .D(
        n12254), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_9_ ( .D(
        n12255), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_8_ ( .D(
        n12239), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_7_ ( .D(
        n12243), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_6_ ( .D(
        n12242), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_5_ ( .D(
        n12245), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_4_ ( .D(
        n12263), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_3_ ( .D(
        n12260), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_2_ ( .D(
        n12244), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_1_ ( .D(
        n12264), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_6_ ( .D(
        n29024), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_2_ ( .D(
        n29025), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_12_ ( 
        .D(n28948), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_10_ ( 
        .D(j202_soc_core_qspi_wb_addr[12]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_12_ ( .D(
        n28948), .DE(n29506), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_4_ ( .D(
        n29026), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_11_ ( .D(
        j202_soc_core_j22_cpu_ml_N314), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_11_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[11]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_11_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[11]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_11_ ( .D(
        j202_soc_core_j22_cpu_ml_N423), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_11_ ( .D(
        j202_soc_core_j22_cpu_rf_N309), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__27_ ( 
        .D(n28996), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[27]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_3_ ( .D(n41), .CLK(
        wb_clk_i), .RESET_B(n12142), .Q(j202_soc_core_uart_div0[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_clr_reg ( .D(
        j202_soc_core_uart_BRG_N21), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps_clr) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_0_ ( .D(
        j202_soc_core_uart_BRG_N12), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_1_ ( .D(
        j202_soc_core_uart_BRG_N13), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_2_ ( .D(
        j202_soc_core_uart_BRG_N14), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_3_ ( .D(
        j202_soc_core_uart_BRG_N15), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_4_ ( .D(
        j202_soc_core_uart_BRG_N16), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_5_ ( .D(
        j202_soc_core_uart_BRG_N17), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_6_ ( .D(
        j202_soc_core_uart_BRG_N18), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_7_ ( .D(
        j202_soc_core_uart_BRG_N19), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_27_ ( 
        .D(j202_soc_core_qspi_wb_wdat[27]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_27_ ( 
        .D(n28949), .DE(n10676), .CLK(wb_clk_i), .Q(la_data_out[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_27_ ( 
        .D(n28949), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_27_ ( 
        .D(n28949), .DE(n10674), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_27_ ( 
        .D(n28949), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_27_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N67), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_27_ ( .D(
        j202_soc_core_ahb2apb_02_N155), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[59]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_11_ ( .D(
        n13315), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_15__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_15__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_15_ ( 
        .D(n29046), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[15])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_14__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_14__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_14_ ( 
        .D(n29047), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[14])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_13__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_13__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_13_ ( 
        .D(n29049), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[13])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_12__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_12__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_12_ ( 
        .D(n29048), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[12])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_11__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_11__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_11_ ( 
        .D(n29060), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[11])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_10__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_10__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_10_ ( 
        .D(n29043), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[10])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_9__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_9__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_9_ ( 
        .D(n29044), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_8__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_8__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_8_ ( 
        .D(n29045), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_7__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_7__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_7_ ( 
        .D(n29042), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_6__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_6__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_6_ ( 
        .D(n29041), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_5__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_5__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_5_ ( 
        .D(n29039), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_4__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_4__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_4_ ( 
        .D(n29040), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_3__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_3__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_3_ ( 
        .D(n29037), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_2__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_2__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_2_ ( 
        .D(n29068), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_1__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_1__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_1_ ( 
        .D(n29052), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_0__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_0__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_0_ ( 
        .D(n29038), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[64]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[66]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[67]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[68]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[69]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[70]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[71]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[72]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[74]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[76]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[77]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[78]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[79]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[80]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[82]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[84]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[85]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[86]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[87]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[88]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[90]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[91]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[92]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[93]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[94]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[95]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[96]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[98]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[99]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[100]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[101]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[102]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[103]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[104]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[106]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[108]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[109]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[110]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[111]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[112]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[114]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[116]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[117]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[118]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[119]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[120]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[122]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[123]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[124]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[125]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[126]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[127]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[32]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[34]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[35]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[36]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[37]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[38]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[39]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[40]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[42]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[44]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[45]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[46]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[47]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[48]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[50]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[52]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[54]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[55]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[56]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[58]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[59]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[60]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[61]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[62]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[63]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[64]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[96]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[33]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[65]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[97]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[66]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[35]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[67]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[99]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[68]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[37]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[69]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[101]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[70]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[102]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[39]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[71]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[103]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[88]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[120]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[57]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[89]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[121]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[90]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[59]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[91]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[123]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[92]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[61]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[93]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[125]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[94]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[126]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[63]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[95]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[127]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[72]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[104]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[41]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[73]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[105]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[74]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[43]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[75]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[107]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[76]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[45]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[77]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[109]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[78]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[110]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[47]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[79]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[111]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[80]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[112]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[49]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[81]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[113]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[82]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[51]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[83]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[115]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[84]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[53]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[85]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[117]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[86]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[118]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[55]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[87]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[119]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_2_ ( .D(
        j202_soc_core_ahb2apb_01_N130), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[66]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_4_ ( .D(
        j202_soc_core_ahb2apb_01_N132), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[68]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_5_ ( .D(
        j202_soc_core_ahb2apb_01_N133), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[69]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_6_ ( .D(
        j202_soc_core_ahb2apb_01_N134), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[70]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_7_ ( .D(
        j202_soc_core_ahb2apb_01_N135), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[71]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_15_ ( .D(
        j202_soc_core_ahb2apb_01_N143), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[79]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_20_ ( .D(
        j202_soc_core_ahb2apb_01_N148), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[84]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_21_ ( .D(
        j202_soc_core_ahb2apb_01_N149), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[85]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_22_ ( .D(
        j202_soc_core_ahb2apb_01_N150), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[86]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_23_ ( .D(
        j202_soc_core_ahb2apb_01_N151), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[87]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_01_N128), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[64]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_10_ ( .D(
        j202_soc_core_ahb2apb_01_N138), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[74]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_24_ ( .D(
        j202_soc_core_ahb2apb_01_N152), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[88]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_26_ ( .D(
        j202_soc_core_ahb2apb_01_N154), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[90]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_27_ ( .D(
        j202_soc_core_ahb2apb_01_N155), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[91]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_28_ ( .D(
        j202_soc_core_ahb2apb_01_N156), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[92]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_29_ ( .D(
        j202_soc_core_ahb2apb_01_N157), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[93]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_30_ ( .D(
        j202_soc_core_ahb2apb_01_N158), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[94]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_31_ ( .D(
        j202_soc_core_ahb2apb_01_N159), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[95]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_15_ ( .D(
        n29074), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[15])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_13_ ( .D(
        n29019), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[13])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_11_ ( .D(
        n29020), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[11])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_9_ ( .D(
        n29078), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_7_ ( .D(
        n29023), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_5_ ( .D(
        n29016), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_3_ ( .D(
        n29073), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_11_ ( 
        .D(n29062), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_9_ ( 
        .D(j202_soc_core_qspi_wb_addr[11]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_11_ ( .D(
        n29062), .DE(n29505), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_12_ ( .D(
        n29017), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[12])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_10_ ( .D(
        n29022), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[10])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_8_ ( .D(
        n29021), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_17_ ( .D(
        j202_soc_core_j22_cpu_ml_N320), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_17_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[17]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_17_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[17]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_17_ ( .D(n12251), 
        .DE(n29119), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufb[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_17_ ( .D(
        j202_soc_core_j22_cpu_rf_N315), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ml_N413), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_1_ ( .D(
        j202_soc_core_j22_cpu_rf_N299), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3346), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__1_ ( .D(
        n28988), .DE(n29356), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_1_ ( 
        .D(j202_soc_core_qspi_wb_wdat[1]), .CLK(wb_clk_i), .RESET_B(n29591), 
        .Q(j202_soc_core_bldc_core_00_wdata[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ccr_00_reg_o_reg_1_ ( 
        .D(n40), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_bldc_core_00_comm[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bcr_00_reg_o_reg_1_ ( 
        .D(n39), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_bldc_core_00_adc_en) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_1_ ( 
        .D(n38), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_bldc_core_00_pwm_period[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_1_ ( .D(n37), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_uart_din_i[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__1_ ( .D(
        j202_soc_core_uart_din_i[1]), .DE(n29345), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__1_ ( .D(
        j202_soc_core_uart_din_i[1]), .DE(n29352), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__1_ ( .D(
        j202_soc_core_uart_din_i[1]), .DE(n29344), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__1_ ( .D(
        j202_soc_core_uart_din_i[1]), .DE(n29346), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_mem[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_1_ ( 
        .D(j202_soc_core_qspi_wb_wdat[1]), .CLK(wb_clk_i), .RESET_B(n29593), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_1_ ( 
        .D(n36), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_cmt_core_00_const1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_1_ ( 
        .D(n35), .CLK(wb_clk_i), .RESET_B(n29591), .Q(
        j202_soc_core_cmt_core_00_const0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_1_ ( 
        .D(n34), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_cks1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_1_ ( 
        .D(n33), .CLK(wb_clk_i), .RESET_B(n29593), .Q(
        j202_soc_core_cmt_core_00_cks0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[0]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[1]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[2]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[3]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[4]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[5]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[6]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[7]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[8]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[9]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmstr_reg_reg_o_reg_1_ ( 
        .D(n32), .CLK(wb_clk_i), .RESET_B(n29594), .Q(
        j202_soc_core_cmt_core_00_str1) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[9]), .CLK(wb_clk_i), .RESET_B(n29594), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[0]), .CLK(wb_clk_i), .RESET_B(n29594), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[2]), .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cnt1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[2]), .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[3]), .CLK(wb_clk_i), .RESET_B(n12142), .Q(j202_soc_core_cmt_core_00_cnt1[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[3]), .CLK(wb_clk_i), .RESET_B(n29591), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[4]), .CLK(wb_clk_i), .RESET_B(n12142), .Q(j202_soc_core_cmt_core_00_cnt1[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[4]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[5]), .CLK(wb_clk_i), .RESET_B(n12142), .Q(j202_soc_core_cmt_core_00_cnt1[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[5]), .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[6]), .CLK(wb_clk_i), .RESET_B(n12142), .Q(j202_soc_core_cmt_core_00_cnt1[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[6]), .CLK(wb_clk_i), .RESET_B(n29591), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[7]), .CLK(wb_clk_i), .RESET_B(n29591), .Q(j202_soc_core_cmt_core_00_cnt1[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[7]), .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[1]), .CLK(wb_clk_i), .RESET_B(n29594), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[2]), .CLK(wb_clk_i), .RESET_B(n29594), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[3]), .CLK(wb_clk_i), .RESET_B(n29594), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_4_ ( 
        .D(n29154), .CLK(wb_clk_i), .RESET_B(n29594), .Q(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[5]), .CLK(wb_clk_i), .RESET_B(n29594), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_6_ ( 
        .D(n29153), .CLK(wb_clk_i), .RESET_B(n29594), .Q(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[7]), .CLK(wb_clk_i), .RESET_B(n29594), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[8]), .CLK(wb_clk_i), .RESET_B(n29594), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[8]) );
  sky130_fd_sc_hd__dfstp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[0]), .CLK(wb_clk_i), .SET_B(n29593), .Q(j202_soc_core_cmt_core_00_cnt1[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[0]), .CLK(wb_clk_i), .RESET_B(n29591), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[8]), .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cnt1[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[8]), .CLK(wb_clk_i), .RESET_B(n29594), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[1]), .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cnt1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[1]), .CLK(wb_clk_i), .RESET_B(n29591), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_1_ ( 
        .D(j202_soc_core_qspi_wb_wdat[1]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_1_ ( .D(
        j202_soc_core_wbqspiflash_00_N629), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_quad_mode_enabled_reg ( 
        .D(j202_soc_core_wbqspiflash_00_N739), .DE(
        j202_soc_core_wbqspiflash_00_N738), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_27_ ( 
        .D(j202_soc_core_wbqspiflash_00_N694), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_N606), .DE(n29358), .CLK(wb_clk_i), 
        .Q(j202_soc_core_wbqspiflash_00_last_status[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[56]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[48]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[40]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[32]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[97]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[65]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[33]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_01_N129), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[65]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_1_ ( 
        .D(n28951), .DE(n10676), .CLK(wb_clk_i), .Q(la_data_out[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_1_ ( 
        .D(n28951), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_1_ ( 
        .D(n28951), .DE(n10674), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_1_ ( 
        .D(n28951), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_1_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N41), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_02_N129), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[33]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__17_ ( 
        .D(n28985), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[17]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_17_ ( 
        .D(j202_soc_core_qspi_wb_wdat[17]), .CLK(wb_clk_i), .RESET_B(n29592), 
        .Q(j202_soc_core_bldc_core_00_wdata[17]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_17_ ( 
        .D(n31), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_17_ ( 
        .D(j202_soc_core_qspi_wb_wdat[17]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_N714), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[60]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[52]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[44]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[36]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[113]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[81]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[49]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_17_ ( .D(
        j202_soc_core_ahb2apb_01_N145), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[81]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_17_ ( 
        .D(n28952), .DE(n10676), .CLK(wb_clk_i), .Q(la_data_out[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_17_ ( 
        .D(n28952), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_17_ ( 
        .D(n28952), .DE(n10674), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_17_ ( 
        .D(n28952), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_17_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N57), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_17_ ( .D(
        j202_soc_core_ahb2apb_02_N145), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[49]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_9_ ( .D(
        j202_soc_core_j22_cpu_rf_N307), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__25_ ( 
        .D(n28994), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_25_ ( 
        .D(j202_soc_core_qspi_wb_wdat[25]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[62]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[54]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[46]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[38]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[121]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[89]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[57]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_25_ ( .D(
        j202_soc_core_ahb2apb_01_N153), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[89]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_25_ ( 
        .D(n28953), .DE(n10676), .CLK(wb_clk_i), .Q(la_data_out[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_25_ ( 
        .D(n28953), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_25_ ( 
        .D(n28953), .DE(n10674), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_25_ ( 
        .D(n28953), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_25_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N65), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_25_ ( .D(
        j202_soc_core_ahb2apb_02_N153), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[57]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__9_ ( .D(
        n28974), .DE(n29356), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_9_ ( 
        .D(j202_soc_core_qspi_wb_wdat[9]), .CLK(wb_clk_i), .RESET_B(n29592), 
        .Q(j202_soc_core_bldc_core_00_wdata[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_9_ ( 
        .D(n30), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_pwm_period[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_9_ ( 
        .D(j202_soc_core_qspi_wb_wdat[9]), .CLK(wb_clk_i), .RESET_B(n29594), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_9_ ( 
        .D(n29), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_const1[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_9_ ( 
        .D(n28), .CLK(wb_clk_i), .RESET_B(n12142), .Q(
        j202_soc_core_cmt_core_00_const0[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[9]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cnt0[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[9]), .CLK(wb_clk_i), .RESET_B(n12142), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmf0_o_reg ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt0_to1), .CLK(
        wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmf0) );
  sky130_fd_sc_hd__dfstp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[0]), .CLK(wb_clk_i), .SET_B(n29593), .Q(j202_soc_core_cmt_core_00_cnt0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[0]), .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[0]), .CLK(wb_clk_i), 
        .RESET_B(n29592), .Q(j202_soc_core_prdata[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_00_N128), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[96]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[1]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cnt0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[1]), .CLK(wb_clk_i), .RESET_B(n29591), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[1]), .CLK(wb_clk_i), 
        .RESET_B(n29591), .Q(j202_soc_core_prdata[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_00_N129), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[97]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[2]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cnt0[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[2]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[2]), .CLK(wb_clk_i), 
        .RESET_B(n29594), .Q(j202_soc_core_prdata[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_2_ ( .D(
        j202_soc_core_ahb2apb_00_N130), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[98]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[3]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cnt0[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[3]), .CLK(wb_clk_i), .RESET_B(n29591), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[3]), .CLK(wb_clk_i), 
        .RESET_B(n29591), .Q(j202_soc_core_prdata[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_3_ ( .D(
        j202_soc_core_ahb2apb_00_N131), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[99]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[4]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cnt0[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[4]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[4]), .CLK(wb_clk_i), 
        .RESET_B(n29592), .Q(j202_soc_core_prdata[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_4_ ( .D(
        j202_soc_core_ahb2apb_00_N132), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[100])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[5]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cnt0[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[5]), .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[5]), .CLK(wb_clk_i), 
        .RESET_B(n29592), .Q(j202_soc_core_prdata[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_5_ ( .D(
        j202_soc_core_ahb2apb_00_N133), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[101])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[6]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cnt0[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[6]), .CLK(wb_clk_i), .RESET_B(n29591), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[6]), .CLK(wb_clk_i), 
        .RESET_B(n29591), .Q(j202_soc_core_prdata[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_6_ ( .D(
        j202_soc_core_ahb2apb_00_N134), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[102])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[7]), .CLK(wb_clk_i), .RESET_B(n29595), .Q(j202_soc_core_cmt_core_00_cnt0[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[7]), .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[8]), .CLK(wb_clk_i), .RESET_B(n12142), .Q(j202_soc_core_cmt_core_00_cnt0[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[8]), .CLK(wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[8]), .CLK(wb_clk_i), 
        .RESET_B(n29592), .Q(j202_soc_core_prdata[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_8_ ( .D(
        j202_soc_core_ahb2apb_00_N136), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[104])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[10]), .CLK(
        wb_clk_i), .RESET_B(n29595), .Q(j202_soc_core_cmt_core_00_cnt0[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[10]), .CLK(wb_clk_i), .RESET_B(
        n29593), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[11]), .CLK(
        wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cnt0[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[11]), .CLK(wb_clk_i), .RESET_B(
        n29592), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[11]), .CLK(wb_clk_i), .RESET_B(n29594), .Q(j202_soc_core_prdata[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_11_ ( .D(
        j202_soc_core_ahb2apb_00_N139), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[107])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[12]), .CLK(
        wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cnt0[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[12]), .CLK(wb_clk_i), .RESET_B(
        n29593), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[13]), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cnt0[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[13]), .CLK(wb_clk_i), .RESET_B(
        n29592), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[14]), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cnt0[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[14]), .CLK(wb_clk_i), .RESET_B(
        n29591), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[15]), .CLK(
        wb_clk_i), .RESET_B(n29591), .Q(j202_soc_core_cmt_core_00_cnt0[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[15]), .CLK(wb_clk_i), .RESET_B(
        n29591), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_9_ ( 
        .D(j202_soc_core_qspi_wb_wdat[9]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_9_ ( .D(
        n10528), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[58]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[50]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[42]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[34]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[105]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[73]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_9_ ( .D(
        j202_soc_core_ahb2apb_01_N137), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[73]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_9_ ( 
        .D(n28954), .DE(n10676), .CLK(wb_clk_i), .Q(la_data_out[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_9_ ( 
        .D(n28954), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_9_ ( 
        .D(n28954), .DE(n10674), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_9_ ( 
        .D(n28954), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_9_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N49), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_9_ ( .D(
        j202_soc_core_ahb2apb_02_N137), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[41]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3368), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3333), .DE(n29112), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3294), .DE(n23533), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gbr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2702), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2739), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[53]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2776), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[85]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2813), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[117]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2850), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[149]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2887), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[181]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2924), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[213]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2961), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[245]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2998), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[277]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3035), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[309]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3072), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[341]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3109), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[373]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3146), .DE(n29317), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[405]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3183), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[437]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3220), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[469]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3257), .DE(n13310), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_gpr[501]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_21_ ( .D(n12269), 
        .DE(n29235), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_3_ ( .D(
        j202_soc_core_ahb2apb_01_N131), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[67]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_3_ ( 
        .D(n28955), .DE(n10676), .CLK(wb_clk_i), .Q(la_data_out[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_3_ ( 
        .D(n28955), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_3_ ( 
        .D(n28955), .DE(n10674), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_3_ ( 
        .D(n28955), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_3_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N43), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_3_ ( .D(
        j202_soc_core_ahb2apb_02_N131), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[35]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__19_ ( 
        .D(n28987), .DE(n29356), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[19]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_19_ ( 
        .D(j202_soc_core_qspi_wb_wdat[19]), .CLK(wb_clk_i), .RESET_B(n12142), 
        .Q(j202_soc_core_bldc_core_00_wdata[19]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_19_ ( 
        .D(n27), .CLK(wb_clk_i), .RESET_B(n12142), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld_reg ( 
        .D(n26), .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_3_ ( .D(n25), .CLK(
        wb_clk_i), .RESET_B(n12142), .Q(j202_soc_core_uart_div1[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_19_ ( 
        .D(j202_soc_core_qspi_wb_wdat[19]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_N716), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[124]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[116]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[108]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[100]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[115]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[83]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[51]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_19_ ( .D(
        j202_soc_core_ahb2apb_01_N147), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[83]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_19_ ( 
        .D(n28956), .DE(n10676), .CLK(wb_clk_i), .Q(la_data_out[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_19_ ( 
        .D(n28956), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_19_ ( 
        .D(n28956), .DE(n10674), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_19_ ( 
        .D(n28956), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_19_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N59), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_19_ ( .D(
        j202_soc_core_ahb2apb_02_N147), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[51]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_29_ ( .D(
        j202_soc_core_j22_cpu_ml_N368), .DE(n29119), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_13_ ( .D(
        j202_soc_core_j22_cpu_ml_N425), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_25_ ( 
        .D(n29164), .DE(j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_24_ ( 
        .D(n29163), .DE(j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_23_ ( 
        .D(n29162), .DE(j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_22_ ( 
        .D(n29161), .DE(j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_21_ ( 
        .D(j202_soc_core_wbqspiflash_00_N688), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_20_ ( 
        .D(j202_soc_core_wbqspiflash_00_N687), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_19_ ( 
        .D(j202_soc_core_wbqspiflash_00_N686), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_18_ ( 
        .D(j202_soc_core_wbqspiflash_00_N685), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_17_ ( 
        .D(j202_soc_core_wbqspiflash_00_N684), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_16_ ( 
        .D(j202_soc_core_wbqspiflash_00_N683), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_15_ ( 
        .D(j202_soc_core_wbqspiflash_00_N682), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_14_ ( 
        .D(j202_soc_core_wbqspiflash_00_N681), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_13_ ( 
        .D(n29160), .DE(j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_12_ ( 
        .D(n29159), .DE(j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_11_ ( 
        .D(n29158), .DE(j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_10_ ( 
        .D(n29157), .DE(j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_9_ ( 
        .D(n29156), .DE(j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_8_ ( 
        .D(n29155), .DE(j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_N674), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_N673), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__6_ ( .D(
        n29324), .DE(n29357), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__6_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_N672), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_N671), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_N670), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_N669), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_N668), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_24_ ( .D(
        n10513), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_25_ ( .D(
        n10512), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_26_ ( .D(
        n10511), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_6_ ( .D(
        j202_soc_core_j22_cpu_ml_N418), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_22_ ( 
        .D(n28957), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_20_ ( 
        .D(j202_soc_core_qspi_wb_addr[22]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_8_ ( .D(
        j202_soc_core_ahb2apb_01_N136), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[72]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_31_ ( .D(
        j202_soc_core_j22_cpu_ml_N370), .DE(n29119), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_15_ ( .D(
        j202_soc_core_j22_cpu_ml_N427), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_32_ ( .D(
        j202_soc_core_j22_cpu_ml_N429), .DE(n29242), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[32]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_13_ ( .D(
        j202_soc_core_ahb2apb_01_N141), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[77]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_13_ ( 
        .D(n28958), .DE(n10676), .CLK(wb_clk_i), .Q(la_data_out[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_13_ ( 
        .D(n28958), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_13_ ( 
        .D(n28958), .DE(n10674), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_13_ ( 
        .D(n28958), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_13_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N53), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_13_ ( .D(
        j202_soc_core_ahb2apb_02_N141), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[45]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__4_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(n29350), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__3_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(n29350), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__2_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(n29350), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__1_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(n29350), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_mem[25]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_dpll_state_reg_1_ ( .D(n24), 
        .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_uart_TOP_dpll_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_cnt_reg_0_ ( .D(n29082), 
        .DE(j202_soc_core_uart_BRG_N55), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_cnt[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_cnt_reg_1_ ( .D(
        j202_soc_core_uart_BRG_N57), .DE(j202_soc_core_uart_BRG_N55), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_BRG_cnt[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_r_reg ( .D(n29090), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_BRG_sio_ce_r) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_reg ( .D(
        j202_soc_core_uart_BRG_N59), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_sio_ce) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_txf_empty_r_reg ( .D(
        j202_soc_core_uart_TOP_N16), .DE(n10679), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_txf_empty_r) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_load_reg ( .D(
        j202_soc_core_uart_TOP_N137), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_load) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_bit_cnt_reg_1_ ( .D(
        j202_soc_core_uart_TOP_N59), .DE(j202_soc_core_uart_TOP_N57), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_bit_cnt[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_bit_cnt_reg_3_ ( .D(
        j202_soc_core_uart_TOP_N61), .DE(j202_soc_core_uart_TOP_N57), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_bit_cnt[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_shift_en_reg ( .D(
        j202_soc_core_uart_TOP_N123), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_shift_en) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_shift_en_r_reg ( .D(n29080), 
        .DE(n10679), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_shift_en_r) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_bit_cnt_reg_0_ ( .D(
        j202_soc_core_uart_TOP_N58), .DE(j202_soc_core_uart_TOP_N57), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_bit_cnt[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_bit_cnt_reg_2_ ( .D(
        j202_soc_core_uart_TOP_N60), .DE(j202_soc_core_uart_TOP_N57), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_bit_cnt[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_tx_fifo_rp_reg_0_ ( .D(n23), 
        .CLK(wb_clk_i), .RESET_B(n29595), .Q(
        j202_soc_core_uart_TOP_tx_fifo_rp[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_tx_fifo_rp_reg_1_ ( .D(n22), 
        .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_uart_TOP_tx_fifo_rp[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_gb_reg ( .D(
        j202_soc_core_uart_TOP_tx_fifo_N42), .DE(
        j202_soc_core_uart_TOP_tx_fifo_N41), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_gb) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_8_ ( .D(
        j202_soc_core_uart_TOP_N33), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_7_ ( .D(
        j202_soc_core_uart_TOP_N32), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_6_ ( .D(
        j202_soc_core_uart_TOP_N31), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_5_ ( .D(
        j202_soc_core_uart_TOP_N30), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_4_ ( .D(
        j202_soc_core_uart_TOP_N29), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_3_ ( .D(
        j202_soc_core_uart_TOP_N28), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_2_ ( .D(
        j202_soc_core_uart_TOP_N27), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_1_ ( .D(
        j202_soc_core_uart_TOP_N26), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_0_ ( .D(
        j202_soc_core_uart_TOP_N25), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_txd_o_reg ( .D(
        j202_soc_core_uart_TOP_N43), .DE(n10679), .CLK(wb_clk_i), .Q(io_out[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_0_ ( .D(
        j202_soc_core_uart_BRG_N35), .DE(n10678), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_7_ ( .D(
        j202_soc_core_uart_BRG_N42), .DE(n10678), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_6_ ( .D(
        j202_soc_core_uart_BRG_N41), .DE(n10678), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_5_ ( .D(
        j202_soc_core_uart_BRG_N40), .DE(n10678), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_4_ ( .D(
        j202_soc_core_uart_BRG_N39), .DE(n10678), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_3_ ( .D(
        j202_soc_core_uart_BRG_N38), .DE(n10678), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_2_ ( .D(
        j202_soc_core_uart_BRG_N37), .DE(n10678), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_1_ ( .D(
        j202_soc_core_uart_BRG_N36), .DE(n10678), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_14_ ( .D(
        j202_soc_core_ahb2apb_01_N142), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[78]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_14_ ( 
        .D(n28959), .DE(n10676), .CLK(wb_clk_i), .Q(la_data_out[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_14_ ( 
        .D(n28959), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_14_ ( 
        .D(n28959), .DE(n10674), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_14_ ( 
        .D(n28959), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_14_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N54), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_14_ ( .D(
        j202_soc_core_ahb2apb_02_N142), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[46]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__i__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3392), .DE(j202_soc_core_j22_cpu_rf_N3391), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__i__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_7_ ( .D(
        j202_soc_core_j22_cpu_rf_N305), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_23_ ( 
        .D(n28960), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_21_ ( 
        .D(j202_soc_core_qspi_wb_addr[23]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[10]), .CLK(
        wb_clk_i), .RESET_B(n29593), .Q(j202_soc_core_cmt_core_00_cnt1[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[10]), .CLK(wb_clk_i), .RESET_B(
        n29592), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[10]), .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_prdata[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_10_ ( .D(
        j202_soc_core_ahb2apb_00_N138), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[106])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[12]), .CLK(
        wb_clk_i), .RESET_B(n29595), .Q(j202_soc_core_cmt_core_00_cnt1[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[12]), .CLK(wb_clk_i), .RESET_B(
        n29593), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[12]), .CLK(wb_clk_i), .RESET_B(n29595), .Q(j202_soc_core_prdata[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_12_ ( .D(
        j202_soc_core_ahb2apb_00_N140), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[108])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[13]), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cnt1[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[13]), .CLK(wb_clk_i), .RESET_B(
        n29592), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[13]), .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_prdata[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_13_ ( .D(
        j202_soc_core_ahb2apb_00_N141), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[109])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[14]), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cnt1[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[14]), .CLK(wb_clk_i), .RESET_B(
        n29591), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[14]), .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_prdata[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_14_ ( .D(
        j202_soc_core_ahb2apb_00_N142), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[110])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[15]), .CLK(
        wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_cmt_core_00_cnt1[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[15]), .CLK(wb_clk_i), .RESET_B(
        n29592), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[15]), .CLK(wb_clk_i), .RESET_B(n29592), .Q(j202_soc_core_prdata[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_15_ ( .D(
        j202_soc_core_ahb2apb_00_N143), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[111])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_11_ ( 
        .D(j202_soc_core_qspi_wb_wdat[11]), .DE(n29239), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[122]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[114]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[106]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[98]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[107]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[75]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[43]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_11_ ( .D(
        j202_soc_core_ahb2apb_01_N139), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[75]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_11_ ( 
        .D(n28961), .DE(n10676), .CLK(wb_clk_i), .Q(la_data_out[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_11_ ( 
        .D(n28961), .DE(n10675), .CLK(wb_clk_i), .Q(gpio_en_o[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_11_ ( 
        .D(n28961), .DE(n10674), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_11_ ( 
        .D(n28961), .DE(n29243), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_11_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N51), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_18_ ( 
        .D(n29058), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[18])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_18_ ( .D(
        j202_soc_core_ahb2apb_01_N146), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[82]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_11_ ( .D(
        j202_soc_core_ahb2apb_02_N139), .DE(n29234), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[43]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_18_ ( .D(
        j202_soc_core_j22_cpu_rf_N316), .DE(n29236), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_21_ ( 
        .D(n10939), .DE(n11125), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_19_ ( 
        .D(j202_soc_core_qspi_wb_addr[21]), .DE(n29240), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_29_ ( .D(
        n10508), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[29]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_nxt_latch_status_0_), 
        .CLK(wb_clk_i), .RESET_B(n29592), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[7]), .CLK(wb_clk_i), 
        .RESET_B(n29593), .Q(j202_soc_core_prdata[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_7_ ( .D(
        j202_soc_core_ahb2apb_00_N135), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[103])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N425), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N426), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N427), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N430), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N428), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N391), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N392), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N393), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N394), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N395), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_10_ ( .D(
        n10527), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_11_ ( .D(
        n10526), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_22_ ( .D(
        n10515), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_23_ ( .D(
        n10514), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_28_ ( .D(
        n10509), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_5_ ( .D(
        n10532), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N396), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N397), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_7_ ( .D(
        n10530), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N398), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_8_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N399), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_9_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N400), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_10_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N401), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_11_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N402), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_12_ ( .D(
        n10525), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_12_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N403), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_13_ ( .D(
        n10524), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_13_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N404), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_14_ ( .D(
        n10523), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_14_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N405), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_15_ ( .D(
        n10522), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_15_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N406), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_16_ ( .D(
        n10521), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_16_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N407), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_17_ ( .D(
        n10520), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_17_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N408), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_18_ ( .D(
        n10519), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_18_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N409), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_19_ ( .D(
        n10518), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_19_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N410), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_20_ ( .D(
        n10517), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_20_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N411), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_21_ ( .D(
        n10516), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_21_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N412), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_22_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N413), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_23_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N414), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_24_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N415), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_25_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N416), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_26_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N417), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_27_ ( .D(
        n10510), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_27_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N418), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_28_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N419), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_29_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N420), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_dat_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N317), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N315), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_30_ ( .D(
        n10507), .DE(n29361), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_30_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N421), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_31_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N422), .DE(n29244), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_dat_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N316), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N315), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_dat_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N319), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N315), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_dat_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N318), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N315), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_12_ ( .D(
        j202_soc_core_ahb2apb_01_N140), .DE(n29238), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[76]) );
  sky130_fd_sc_hd__fa_1 DP_OP_1508J1_126_2326_U6 ( .A(n29118), .B(
        DP_OP_1508J1_126_2326_n6), .CIN(DP_OP_1508J1_126_2326_n4), .COUT(
        DP_OP_1508J1_126_2326_n3), .SUM(U7_RSOP_1495_C3_DATA3_2) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_14_ ( .D(
        n29018), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[14])
         );
  sky130_fd_sc_hd__dfxtp_2 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__0_ ( .D(
        j202_soc_core_j22_cpu_ml_N152), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[10]) );
  sky130_fd_sc_hd__dfxtp_2 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[41]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[19]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_02_pstrb_o_reg_1_ ( .GATE(
        j202_soc_core_ahb2apb_02_N123), .D(n10905), .RESET_B(
        j202_soc_core_pwrite[2]), .Q(j202_soc_core_pstrb[1]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_02_pstrb_o_reg_3_ ( .GATE(
        j202_soc_core_ahb2apb_02_N123), .D(n10907), .RESET_B(
        j202_soc_core_pwrite[2]), .Q(j202_soc_core_pstrb[3]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_02_pstrb_o_reg_0_ ( .GATE(
        j202_soc_core_ahb2apb_02_N123), .D(n10904), .RESET_B(
        j202_soc_core_pwrite[2]), .Q(j202_soc_core_pstrb[0]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_02_pstrb_o_reg_2_ ( .GATE(
        j202_soc_core_ahb2apb_02_N123), .D(n10906), .RESET_B(
        j202_soc_core_pwrite[2]), .Q(j202_soc_core_pstrb[2]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_01_pstrb_o_reg_1_ ( .GATE(
        j202_soc_core_ahb2apb_01_N123), .D(n10746), .RESET_B(
        j202_soc_core_pwrite[1]), .Q(j202_soc_core_pstrb[5]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_01_pstrb_o_reg_3_ ( .GATE(
        j202_soc_core_ahb2apb_01_N123), .D(n10748), .RESET_B(
        j202_soc_core_pwrite[1]), .Q(j202_soc_core_pstrb[7]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_01_pstrb_o_reg_2_ ( .GATE(
        j202_soc_core_ahb2apb_01_N123), .D(n10747), .RESET_B(
        j202_soc_core_pwrite[1]), .Q(j202_soc_core_pstrb[6]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_01_pstrb_o_reg_0_ ( .GATE(
        j202_soc_core_ahb2apb_01_N123), .D(n10745), .RESET_B(
        j202_soc_core_pwrite[1]), .Q(j202_soc_core_pstrb[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_nega_o_reg ( 
        .D(n29089), .CLK(wb_clk_i), .RESET_B(n29591), .Q(io_out[17]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_posc_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posc), .CLK(wb_clk_i), .RESET_B(n29592), .Q(io_out[20]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_negb_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_negb), .CLK(wb_clk_i), .RESET_B(n29592), .Q(io_out[19]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_negc_o_reg ( 
        .D(n29088), .CLK(wb_clk_i), .RESET_B(n29591), .Q(io_out[21]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_posb_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posb), .CLK(wb_clk_i), .RESET_B(n29592), .Q(io_out[18]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_posa_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posa), .CLK(wb_clk_i), .RESET_B(n29591), .Q(io_out[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_wbqspiflash_00_spif_override_reg ( 
        .D(j202_soc_core_wbqspiflash_00_N742), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_override) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[53]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[2]) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_other__1_ ( 
        .D(n10489), .DE(n12514), .CLK(wb_clk_i), .Q(n12508), .Q_N(n12509) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_other__0_ ( 
        .D(n10490), .DE(n10584), .CLK(wb_clk_i), .Q(n12506), .Q_N(n12507) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_other__2_ ( 
        .D(n10488), .DE(n12513), .CLK(wb_clk_i), .Q(n12505), .Q_N() );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rm__0_ ( 
        .D(n29075), .DE(j202_soc_core_j22_cpu_id_idec_N857), .CLK(wb_clk_i), 
        .Q(n12431), .Q_N(n12432) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rm__1_ ( 
        .D(n29072), .DE(j202_soc_core_j22_cpu_id_idec_N857), .CLK(wb_clk_i), 
        .Q(n12429), .Q_N(n12430) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rm__3_ ( 
        .D(n12472), .DE(j202_soc_core_j22_cpu_id_idec_N857), .CLK(wb_clk_i), 
        .Q(n12427), .Q_N(n12428) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rm__2_ ( 
        .D(n12617), .DE(j202_soc_core_j22_cpu_id_idec_N857), .CLK(wb_clk_i), 
        .Q(n12425), .Q_N(n12426) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__1_ ( 
        .D(n10595), .DE(n29117), .CLK(wb_clk_i), .Q(n12381), .Q_N(n12382) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_We__0_ ( 
        .D(n10578), .DE(n10607), .CLK(wb_clk_i), .Q(n12365), .Q_N(n12366) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rb__0_ ( 
        .D(n10581), .DE(n29117), .CLK(wb_clk_i), .Q(n12350), .Q_N() );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[15]) );
  sky130_fd_sc_hd__dfxtp_2 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__3_ ( .D(
        j202_soc_core_j22_cpu_ml_N155), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_rst_reg ( .D(j202_soc_core_rst1), 
        .CLK(wb_clk_i), .Q(j202_soc_core_rst) );
  sky130_fd_sc_hd__dfxtp_2 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__4_ ( .D(
        j202_soc_core_j22_cpu_ml_N156), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[4]) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__11_ ( 
        .D(n10492), .DE(n12358), .CLK(wb_clk_i), .Q(n10989), .Q_N(n10990) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__10_ ( 
        .D(n10493), .DE(n12418), .CLK(wb_clk_i), .Q(n10987), .Q_N(n10988) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__9_ ( 
        .D(n10494), .DE(n12358), .CLK(wb_clk_i), .Q(n10985), .Q_N(n10986) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__8_ ( 
        .D(n10495), .DE(n29233), .CLK(wb_clk_i), .Q(n10984), .Q_N() );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__6_ ( 
        .D(n10497), .DE(n12497), .CLK(wb_clk_i), .Q(n10983), .Q_N() );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__4_ ( 
        .D(n10499), .DE(n29233), .CLK(wb_clk_i), .Q(n10981), .Q_N(n10982) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__0_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N917), .DE(n12497), .CLK(wb_clk_i), 
        .Q(n10979), .Q_N(n10980) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__5_ ( 
        .D(n10498), .DE(n12418), .CLK(wb_clk_i), .Q(n10977), .Q_N(n10978) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_ml_bufa_reg_4_ ( .D(
        j202_soc_core_j22_cpu_ml_N307), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(n10968), .Q_N(n10969) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_2_ ( .D(
        j202_soc_core_ahb2apb_00_N25), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(n10961), .Q_N() );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__1_ ( .D(
        n28976), .DE(j202_soc_core_ahb2aqu_00_N127), .CLK(wb_clk_i), .Q(n10960), .Q_N() );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_ahb2wbqspi_00_hwrite_temp_reg ( .D(
        n29066), .DE(n11125), .CLK(wb_clk_i), .Q(n10958), .Q_N(n10959) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__3_ ( 
        .D(n10500), .DE(n10585), .CLK(wb_clk_i), .Q(n10931), .Q_N() );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__2_ ( 
        .D(n10501), .DE(n10585), .CLK(wb_clk_i), .Q(n10929), .Q_N(n10930) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__1_ ( 
        .D(n10502), .DE(n12375), .CLK(wb_clk_i), .Q(n10922), .Q_N(n10923) );
  sky130_fd_sc_hd__edfxbp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__12_ ( 
        .D(n10491), .DE(n12375), .CLK(wb_clk_i), .Q(n10920), .Q_N(n10921) );
  sky130_fd_sc_hd__dfxtp_2 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__2_ ( .D(
        j202_soc_core_j22_cpu_ml_N154), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]) );
  sky130_fd_sc_hd__buf_4 U13283 ( .A(n23288), .X(n11125) );
  sky130_fd_sc_hd__nand2_1 U13285 ( .A(n11391), .B(n29594), .Y(n12491) );
  sky130_fd_sc_hd__nand2_1 U13286 ( .A(n11391), .B(n29594), .Y(
        j202_soc_core_ahb2apb_02_N22) );
  sky130_fd_sc_hd__clkbuf_1 U13287 ( .A(n24592), .X(n27234) );
  sky130_fd_sc_hd__inv_4 U13288 ( .A(n12168), .Y(n11122) );
  sky130_fd_sc_hd__buf_2 U13290 ( .A(n24638), .X(n24644) );
  sky130_fd_sc_hd__inv_2 U13291 ( .A(n11764), .Y(n27451) );
  sky130_fd_sc_hd__inv_2 U13292 ( .A(n11586), .Y(n12160) );
  sky130_fd_sc_hd__inv_4 U13293 ( .A(n12802), .Y(n26469) );
  sky130_fd_sc_hd__inv_4 U13294 ( .A(n11036), .Y(n11037) );
  sky130_fd_sc_hd__inv_1 U13295 ( .A(n11612), .Y(n24055) );
  sky130_fd_sc_hd__inv_4 U13296 ( .A(n24497), .Y(n26523) );
  sky130_fd_sc_hd__inv_2 U13297 ( .A(n23815), .Y(n12533) );
  sky130_fd_sc_hd__inv_4 U13298 ( .A(n11126), .Y(n11089) );
  sky130_fd_sc_hd__inv_2 U13299 ( .A(n23814), .Y(n11040) );
  sky130_fd_sc_hd__buf_2 U13300 ( .A(n25661), .X(n12473) );
  sky130_fd_sc_hd__inv_2 U13301 ( .A(n23552), .Y(n23553) );
  sky130_fd_sc_hd__buf_6 U13304 ( .A(n23814), .X(n11098) );
  sky130_fd_sc_hd__inv_2 U13306 ( .A(n11038), .Y(n11008) );
  sky130_fd_sc_hd__inv_2 U13307 ( .A(n11038), .Y(n11010) );
  sky130_fd_sc_hd__inv_6 U13308 ( .A(n12534), .Y(n11026) );
  sky130_fd_sc_hd__and3_1 U13310 ( .A(n27657), .B(n27656), .C(n27655), .X(
        n28874) );
  sky130_fd_sc_hd__nor2_1 U13311 ( .A(n27652), .B(n27653), .Y(n28876) );
  sky130_fd_sc_hd__nor2_1 U13312 ( .A(n27654), .B(n27653), .Y(n28875) );
  sky130_fd_sc_hd__buf_2 U13313 ( .A(n23167), .X(n29067) );
  sky130_fd_sc_hd__inv_2 U13314 ( .A(n11391), .Y(n12899) );
  sky130_fd_sc_hd__inv_2 U13315 ( .A(n25875), .Y(n26981) );
  sky130_fd_sc_hd__nor2_1 U13316 ( .A(n21030), .B(n25227), .Y(n29065) );
  sky130_fd_sc_hd__nand2_2 U13318 ( .A(n25156), .B(n25152), .Y(n12385) );
  sky130_fd_sc_hd__inv_2 U13319 ( .A(n23816), .Y(n23817) );
  sky130_fd_sc_hd__inv_2 U13320 ( .A(n12740), .Y(n11102) );
  sky130_fd_sc_hd__nand2b_1 U13322 ( .A_N(n24188), .B(n29011), .Y(n23814) );
  sky130_fd_sc_hd__buf_6 U13324 ( .A(n23552), .X(n10940) );
  sky130_fd_sc_hd__and2_2 U13329 ( .A(n23278), .B(n23277), .X(n13320) );
  sky130_fd_sc_hd__nor2_2 U13330 ( .A(n23114), .B(n23169), .Y(n27217) );
  sky130_fd_sc_hd__nor2_2 U13331 ( .A(n23131), .B(n23169), .Y(n27219) );
  sky130_fd_sc_hd__nor2_2 U13332 ( .A(n22998), .B(n23169), .Y(n27209) );
  sky130_fd_sc_hd__nand2b_1 U13335 ( .A_N(n12416), .B(n29032), .Y(n23812) );
  sky130_fd_sc_hd__nand2_1 U13336 ( .A(n25047), .B(n26722), .Y(n11697) );
  sky130_fd_sc_hd__inv_2 U13337 ( .A(n12411), .Y(n11036) );
  sky130_fd_sc_hd__or2_1 U13338 ( .A(n18916), .B(n25545), .X(n12123) );
  sky130_fd_sc_hd__inv_2 U13339 ( .A(n25116), .Y(n11551) );
  sky130_fd_sc_hd__nand2_1 U13340 ( .A(n12457), .B(n22669), .Y(n25227) );
  sky130_fd_sc_hd__o211a_2 U13341 ( .A1(n23014), .A2(n25159), .B1(n23035), 
        .C1(n23034), .X(n25152) );
  sky130_fd_sc_hd__nand3_1 U13343 ( .A(n22257), .B(n21901), .C(n21900), .Y(
        n28981) );
  sky130_fd_sc_hd__nor2_2 U13344 ( .A(n23123), .B(n23169), .Y(n27575) );
  sky130_fd_sc_hd__inv_2 U13347 ( .A(n24188), .Y(n11127) );
  sky130_fd_sc_hd__nor2_1 U13348 ( .A(n26516), .B(n26948), .Y(n24650) );
  sky130_fd_sc_hd__nand3_2 U13350 ( .A(n23229), .B(n23227), .C(n23228), .Y(
        n12487) );
  sky130_fd_sc_hd__clkbuf_1 U13352 ( .A(n27382), .X(n12645) );
  sky130_fd_sc_hd__nand2_1 U13354 ( .A(n11521), .B(n12666), .Y(n26557) );
  sky130_fd_sc_hd__a21oi_1 U13357 ( .A1(n26519), .A2(n26406), .B1(n24493), .Y(
        n11543) );
  sky130_fd_sc_hd__nand2_2 U13358 ( .A(n11521), .B(n23746), .Y(n27182) );
  sky130_fd_sc_hd__nand2_1 U13359 ( .A(n23268), .B(n23267), .Y(n27047) );
  sky130_fd_sc_hd__inv_2 U13363 ( .A(n12493), .Y(n26556) );
  sky130_fd_sc_hd__nand3_1 U13364 ( .A(n27261), .B(n11814), .C(n27957), .Y(
        n13233) );
  sky130_fd_sc_hd__nand2_1 U13367 ( .A(n26315), .B(n26542), .Y(n12374) );
  sky130_fd_sc_hd__nand2_1 U13368 ( .A(n19448), .B(n29535), .Y(n24590) );
  sky130_fd_sc_hd__nand2_1 U13369 ( .A(n13145), .B(n13143), .Y(n24636) );
  sky130_fd_sc_hd__nand2b_1 U13371 ( .A_N(n12714), .B(n29569), .Y(n23565) );
  sky130_fd_sc_hd__nand3_1 U13373 ( .A(n11983), .B(n11982), .C(n11981), .Y(
        n22242) );
  sky130_fd_sc_hd__a2bb2oi_1 U13374 ( .B1(n23777), .B2(n12175), .A1_N(n26312), 
        .A2_N(n29513), .Y(n26542) );
  sky130_fd_sc_hd__nor2_1 U13375 ( .A(n23162), .B(n11396), .Y(n27688) );
  sky130_fd_sc_hd__nand2_1 U13376 ( .A(n11128), .B(n26863), .Y(n21886) );
  sky130_fd_sc_hd__nor2_2 U13377 ( .A(n12065), .B(n24307), .Y(n12064) );
  sky130_fd_sc_hd__clkbuf_1 U13378 ( .A(n27566), .X(n12658) );
  sky130_fd_sc_hd__clkbuf_1 U13379 ( .A(n22278), .X(n29036) );
  sky130_fd_sc_hd__clkbuf_1 U13380 ( .A(n22274), .X(n12677) );
  sky130_fd_sc_hd__inv_2 U13381 ( .A(n23150), .Y(n11626) );
  sky130_fd_sc_hd__nor2_1 U13382 ( .A(n29077), .B(n12376), .Y(n23583) );
  sky130_fd_sc_hd__nand2_1 U13383 ( .A(n12154), .B(n12225), .Y(n11900) );
  sky130_fd_sc_hd__buf_4 U13384 ( .A(n13103), .X(n29075) );
  sky130_fd_sc_hd__and3_1 U13385 ( .A(n13234), .B(n20961), .C(n20963), .X(
        n12154) );
  sky130_fd_sc_hd__o21a_1 U13386 ( .A1(n17125), .A2(n26525), .B1(n17124), .X(
        n10957) );
  sky130_fd_sc_hd__nand3_1 U13387 ( .A(n15669), .B(n12198), .C(n15668), .Y(
        n28962) );
  sky130_fd_sc_hd__buf_2 U13389 ( .A(n28963), .X(n12735) );
  sky130_fd_sc_hd__nand2_1 U13391 ( .A(n16053), .B(n16052), .Y(n27720) );
  sky130_fd_sc_hd__nand2_1 U13394 ( .A(n14979), .B(n14978), .Y(n21916) );
  sky130_fd_sc_hd__nand2_1 U13396 ( .A(n11406), .B(n11397), .Y(n14979) );
  sky130_fd_sc_hd__nand2_1 U13398 ( .A(n18808), .B(n18809), .Y(n21499) );
  sky130_fd_sc_hd__nand2_1 U13399 ( .A(n12231), .B(n21318), .Y(n12734) );
  sky130_fd_sc_hd__inv_2 U13400 ( .A(n14849), .Y(n26812) );
  sky130_fd_sc_hd__nand2b_1 U13401 ( .A_N(n14847), .B(n23701), .Y(n21584) );
  sky130_fd_sc_hd__nand2_2 U13402 ( .A(n14852), .B(n11913), .Y(n14849) );
  sky130_fd_sc_hd__nor2_1 U13403 ( .A(n27187), .B(n18881), .Y(n22952) );
  sky130_fd_sc_hd__nand3_1 U13405 ( .A(n18879), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[0]), .C(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .Y(n25824) );
  sky130_fd_sc_hd__fa_2 U13409 ( .A(n18707), .B(n18706), .CIN(n18705), .COUT(
        n18765), .SUM(n18728) );
  sky130_fd_sc_hd__nand3_1 U13410 ( .A(n16457), .B(n16456), .C(n16455), .Y(
        n26971) );
  sky130_fd_sc_hd__fa_2 U13411 ( .A(n17949), .B(n17948), .CIN(n17947), .COUT(
        n17954), .SUM(n17958) );
  sky130_fd_sc_hd__fa_1 U13412 ( .A(n18323), .B(n18322), .CIN(n18321), .COUT(
        n18568), .SUM(n18573) );
  sky130_fd_sc_hd__fa_2 U13413 ( .A(n18017), .B(n18016), .CIN(n18015), .COUT(
        n18033), .SUM(n18026) );
  sky130_fd_sc_hd__a2bb2oi_1 U13415 ( .B1(n11162), .B2(n17369), .A1_N(n17378), 
        .A2_N(n11514), .Y(n17376) );
  sky130_fd_sc_hd__fa_2 U13416 ( .A(n17662), .B(n17660), .CIN(n17661), .COUT(
        n17686), .SUM(n17873) );
  sky130_fd_sc_hd__fa_1 U13418 ( .A(n17741), .B(n17740), .CIN(n17739), .COUT(
        n17875), .SUM(n17878) );
  sky130_fd_sc_hd__fa_1 U13419 ( .A(n17641), .B(n17640), .CIN(n17639), .COUT(
        n17645), .SUM(n17874) );
  sky130_fd_sc_hd__fa_2 U13420 ( .A(n18241), .B(n18240), .CIN(n18239), .COUT(
        n18565), .SUM(n18250) );
  sky130_fd_sc_hd__fa_1 U13421 ( .A(n17757), .B(n17756), .CIN(n17755), .COUT(
        n17760), .SUM(n17851) );
  sky130_fd_sc_hd__buf_2 U13422 ( .A(j202_soc_core_j22_cpu_ml_bufa[32]), .X(
        n22051) );
  sky130_fd_sc_hd__buf_4 U13423 ( .A(n13686), .X(n11115) );
  sky130_fd_sc_hd__or2_1 U13424 ( .A(n13638), .B(n23129), .X(n12163) );
  sky130_fd_sc_hd__or2_1 U13425 ( .A(n13638), .B(n23495), .X(n12185) );
  sky130_fd_sc_hd__nand2_1 U13426 ( .A(n13612), .B(n13750), .Y(n14466) );
  sky130_fd_sc_hd__fa_1 U13427 ( .A(n17594), .B(n17593), .CIN(n17592), .COUT(
        n17572), .SUM(n17903) );
  sky130_fd_sc_hd__a21oi_1 U13428 ( .A1(n18225), .A2(n18224), .B1(n18223), .Y(
        n12663) );
  sky130_fd_sc_hd__buf_4 U13429 ( .A(j202_soc_core_j22_cpu_ml_bufa[19]), .X(
        n22951) );
  sky130_fd_sc_hd__nor2_1 U13430 ( .A(n13688), .B(n13681), .Y(n13680) );
  sky130_fd_sc_hd__buf_2 U13431 ( .A(j202_soc_core_j22_cpu_ml_bufb[10]), .X(
        n18661) );
  sky130_fd_sc_hd__buf_2 U13432 ( .A(j202_soc_core_j22_cpu_ml_bufb[13]), .X(
        n18721) );
  sky130_fd_sc_hd__buf_2 U13433 ( .A(j202_soc_core_j22_cpu_ml_bufb[11]), .X(
        n18673) );
  sky130_fd_sc_hd__buf_2 U13434 ( .A(j202_soc_core_j22_cpu_ml_bufb[12]), .X(
        n18685) );
  sky130_fd_sc_hd__buf_4 U13435 ( .A(n17973), .X(n11159) );
  sky130_fd_sc_hd__xnor2_1 U13436 ( .A(j202_soc_core_j22_cpu_ml_bufa[5]), .B(
        n10969), .Y(n17427) );
  sky130_fd_sc_hd__buf_2 U13437 ( .A(j202_soc_core_j22_cpu_ml_bufb[7]), .X(
        n18649) );
  sky130_fd_sc_hd__buf_2 U13438 ( .A(j202_soc_core_j22_cpu_ml_bufb[4]), .X(
        n18479) );
  sky130_fd_sc_hd__buf_2 U13439 ( .A(j202_soc_core_j22_cpu_ml_bufb[32]), .X(
        n22052) );
  sky130_fd_sc_hd__buf_2 U13440 ( .A(j202_soc_core_j22_cpu_ml_bufb[9]), .X(
        n18708) );
  sky130_fd_sc_hd__buf_2 U13441 ( .A(j202_soc_core_j22_cpu_ml_bufb[3]), .X(
        n18466) );
  sky130_fd_sc_hd__buf_2 U13442 ( .A(j202_soc_core_j22_cpu_ml_bufb[2]), .X(
        n18426) );
  sky130_fd_sc_hd__buf_4 U13443 ( .A(j202_soc_core_j22_cpu_ml_bufa[5]), .X(
        n11440) );
  sky130_fd_sc_hd__buf_4 U13444 ( .A(j202_soc_core_j22_cpu_ml_bufa[9]), .X(
        n22919) );
  sky130_fd_sc_hd__nor2_1 U13445 ( .A(n20788), .B(n17274), .Y(n19125) );
  sky130_fd_sc_hd__buf_2 U13446 ( .A(j202_soc_core_j22_cpu_ml_bufb[0]), .X(
        n18353) );
  sky130_fd_sc_hd__clkbuf_1 U13447 ( .A(j202_soc_core_j22_cpu_ml_bufa[8]), .X(
        n25830) );
  sky130_fd_sc_hd__nor2_1 U13448 ( .A(n17277), .B(n11994), .Y(n16171) );
  sky130_fd_sc_hd__nand4bb_1 U13449 ( .A_N(n24385), .B_N(n24327), .C(n23187), 
        .D(n24402), .Y(n23188) );
  sky130_fd_sc_hd__nor2_1 U13450 ( .A(n23186), .B(n23185), .Y(n24327) );
  sky130_fd_sc_hd__nand3_1 U13453 ( .A(n11068), .B(n24135), .C(n29587), .Y(
        n21435) );
  sky130_fd_sc_hd__nand2_1 U13455 ( .A(n23233), .B(n26863), .Y(n24135) );
  sky130_fd_sc_hd__nand4_1 U13456 ( .A(n13050), .B(n13044), .C(n13043), .D(
        n23160), .Y(n10926) );
  sky130_fd_sc_hd__nand4_1 U13457 ( .A(n13050), .B(n13044), .C(n13043), .D(
        n23160), .Y(n24297) );
  sky130_fd_sc_hd__o21bai_1 U13460 ( .A1(n29075), .A2(n23184), .B1_N(n23183), 
        .Y(n23189) );
  sky130_fd_sc_hd__or2b_1 U13463 ( .A(n24328), .B_N(n23185), .X(n25811) );
  sky130_fd_sc_hd__clkinv_2 U13465 ( .A(n10940), .Y(n10932) );
  sky130_fd_sc_hd__a21oi_1 U13469 ( .A1(j202_soc_core_memory0_ram_dout0[321]), 
        .A2(n21593), .B1(n19926), .Y(n10933) );
  sky130_fd_sc_hd__nand3_1 U13473 ( .A(n22274), .B(n12733), .C(n13224), .Y(
        n12010) );
  sky130_fd_sc_hd__nor2_1 U13478 ( .A(n27523), .B(n11842), .Y(n27925) );
  sky130_fd_sc_hd__a21oi_2 U13480 ( .A1(n12068), .A2(n23493), .B1(n11535), .Y(
        n14852) );
  sky130_fd_sc_hd__inv_1 U13486 ( .A(n28960), .Y(n17150) );
  sky130_fd_sc_hd__or2_2 U13487 ( .A(n11956), .B(n11063), .X(n11043) );
  sky130_fd_sc_hd__nand2_2 U13488 ( .A(n15525), .B(n15524), .Y(n28919) );
  sky130_fd_sc_hd__nand3_1 U13489 ( .A(n17107), .B(n13314), .C(n21776), .Y(
        n13234) );
  sky130_fd_sc_hd__nand3_1 U13490 ( .A(n29519), .B(n24300), .C(n27550), .Y(
        n10938) );
  sky130_fd_sc_hd__nand3_1 U13491 ( .A(n12614), .B(n24300), .C(n27550), .Y(
        n27876) );
  sky130_fd_sc_hd__inv_1 U13492 ( .A(n28918), .Y(n21025) );
  sky130_fd_sc_hd__nor2_2 U13493 ( .A(n28918), .B(n28924), .Y(n17151) );
  sky130_fd_sc_hd__nand3_2 U13494 ( .A(n15669), .B(n12198), .C(n15668), .Y(
        n10939) );
  sky130_fd_sc_hd__nand3_2 U13496 ( .A(n17149), .B(n28920), .C(n28960), .Y(
        n11970) );
  sky130_fd_sc_hd__a21oi_2 U13497 ( .A1(n17262), .A2(n14120), .B1(n14119), .Y(
        n19415) );
  sky130_fd_sc_hd__nand2_1 U13498 ( .A(n21379), .B(n11065), .Y(n27428) );
  sky130_fd_sc_hd__nand2_2 U13499 ( .A(n13949), .B(n11978), .Y(n27409) );
  sky130_fd_sc_hd__a2bb2oi_1 U13500 ( .B1(n22715), .B2(n12175), .A1_N(n21915), 
        .A2_N(n29513), .Y(n21379) );
  sky130_fd_sc_hd__inv_2 U13501 ( .A(n26710), .Y(n25821) );
  sky130_fd_sc_hd__buf_8 U13508 ( .A(n23553), .X(n29245) );
  sky130_fd_sc_hd__buf_8 U13509 ( .A(n23553), .X(n12541) );
  sky130_fd_sc_hd__buf_8 U13511 ( .A(n29499), .X(n10943) );
  sky130_fd_sc_hd__buf_8 U13512 ( .A(n29499), .X(n10944) );
  sky130_fd_sc_hd__buf_8 U13514 ( .A(n23553), .X(n10945) );
  sky130_fd_sc_hd__buf_8 U13515 ( .A(n23553), .X(n10946) );
  sky130_fd_sc_hd__buf_8 U13516 ( .A(n23553), .X(n11091) );
  sky130_fd_sc_hd__buf_8 U13517 ( .A(n11040), .X(n10947) );
  sky130_fd_sc_hd__buf_8 U13518 ( .A(n11040), .X(n10948) );
  sky130_fd_sc_hd__buf_8 U13519 ( .A(n11040), .X(n10949) );
  sky130_fd_sc_hd__buf_8 U13520 ( .A(n11040), .X(n10950) );
  sky130_fd_sc_hd__inv_8 U13522 ( .A(n11098), .Y(n10952) );
  sky130_fd_sc_hd__inv_8 U13523 ( .A(n11098), .Y(n10953) );
  sky130_fd_sc_hd__inv_8 U13524 ( .A(n11098), .Y(n10954) );
  sky130_fd_sc_hd__inv_8 U13525 ( .A(n11098), .Y(n10955) );
  sky130_fd_sc_hd__nand3_2 U13527 ( .A(n11452), .B(n11451), .C(n11448), .Y(
        n23225) );
  sky130_fd_sc_hd__o21a_1 U13528 ( .A1(n17125), .A2(n26525), .B1(n17124), .X(
        n17148) );
  sky130_fd_sc_hd__nor2_2 U13529 ( .A(n12400), .B(n17148), .Y(n17130) );
  sky130_fd_sc_hd__xnor2_1 U13531 ( .A(n15305), .B(n10963), .Y(n25176) );
  sky130_fd_sc_hd__and2_1 U13532 ( .A(n15304), .B(n15953), .X(n10963) );
  sky130_fd_sc_hd__nand2_2 U13534 ( .A(n12587), .B(n20958), .Y(n12376) );
  sky130_fd_sc_hd__buf_2 U13537 ( .A(n13162), .X(n13159) );
  sky130_fd_sc_hd__nand3_1 U13538 ( .A(n12515), .B(n23583), .C(n23584), .Y(
        n13162) );
  sky130_fd_sc_hd__nor2b_1 U13539 ( .B_N(n29595), .A(n12122), .Y(n12457) );
  sky130_fd_sc_hd__inv_1 U13540 ( .A(n12629), .Y(n10967) );
  sky130_fd_sc_hd__nand2_2 U13542 ( .A(n12629), .B(n22581), .Y(n15669) );
  sky130_fd_sc_hd__nand2_2 U13543 ( .A(n11394), .B(n12588), .Y(n28957) );
  sky130_fd_sc_hd__nor3_1 U13544 ( .A(n17035), .B(n17075), .C(n14960), .Y(
        n15840) );
  sky130_fd_sc_hd__buf_8 U13545 ( .A(n10951), .X(n29246) );
  sky130_fd_sc_hd__nand2_1 U13546 ( .A(n23582), .B(n23565), .Y(n12842) );
  sky130_fd_sc_hd__nor2_1 U13547 ( .A(n10975), .B(n12501), .Y(n10970) );
  sky130_fd_sc_hd__nor2_1 U13548 ( .A(n10975), .B(n12501), .Y(n12642) );
  sky130_fd_sc_hd__nand2_1 U13549 ( .A(n17386), .B(n17385), .Y(n10971) );
  sky130_fd_sc_hd__nand2_1 U13550 ( .A(n17386), .B(n17385), .Y(n18068) );
  sky130_fd_sc_hd__xnor2_1 U13551 ( .A(n12194), .B(n10972), .Y(n23243) );
  sky130_fd_sc_hd__a21oi_1 U13552 ( .A1(n13330), .A2(n19249), .B1(n19248), .Y(
        n10972) );
  sky130_fd_sc_hd__nor2_1 U13554 ( .A(n10974), .B(n12501), .Y(n12394) );
  sky130_fd_sc_hd__nor2_2 U13555 ( .A(n29491), .B(n11869), .Y(n12093) );
  sky130_fd_sc_hd__nand3_1 U13556 ( .A(n12734), .B(n12716), .C(n21166), .Y(
        n10974) );
  sky130_fd_sc_hd__nand3_1 U13557 ( .A(n12734), .B(n12716), .C(n21166), .Y(
        n10975) );
  sky130_fd_sc_hd__nand2_2 U13559 ( .A(n22766), .B(n29535), .Y(n22767) );
  sky130_fd_sc_hd__a22oi_1 U13560 ( .A1(j202_soc_core_memory0_ram_dout0[137]), 
        .A2(n21592), .B1(n21734), .B2(j202_soc_core_memory0_ram_dout0[73]), 
        .Y(n20939) );
  sky130_fd_sc_hd__inv_1 U13561 ( .A(n22750), .Y(n21911) );
  sky130_fd_sc_hd__nand2_1 U13562 ( .A(n11964), .B(n23968), .Y(n10976) );
  sky130_fd_sc_hd__nand2_1 U13563 ( .A(n11964), .B(n23968), .Y(n12624) );
  sky130_fd_sc_hd__inv_6 U13564 ( .A(n12479), .Y(n10992) );
  sky130_fd_sc_hd__buf_8 U13566 ( .A(n29501), .X(n10991) );
  sky130_fd_sc_hd__buf_8 U13567 ( .A(n29501), .X(n11092) );
  sky130_fd_sc_hd__buf_8 U13568 ( .A(n29501), .X(n12403) );
  sky130_fd_sc_hd__buf_8 U13569 ( .A(n29501), .X(n12409) );
  sky130_fd_sc_hd__buf_8 U13570 ( .A(n29501), .X(n10997) );
  sky130_fd_sc_hd__inv_4 U13571 ( .A(n23813), .Y(n29250) );
  sky130_fd_sc_hd__inv_8 U13572 ( .A(n29250), .Y(n10993) );
  sky130_fd_sc_hd__inv_8 U13573 ( .A(n29250), .Y(n10994) );
  sky130_fd_sc_hd__inv_8 U13574 ( .A(n29250), .Y(n10995) );
  sky130_fd_sc_hd__inv_6 U13575 ( .A(n12479), .Y(n10996) );
  sky130_fd_sc_hd__buf_8 U13576 ( .A(n29501), .X(n10998) );
  sky130_fd_sc_hd__buf_8 U13577 ( .A(n29501), .X(n10999) );
  sky130_fd_sc_hd__buf_8 U13578 ( .A(n11122), .X(n11000) );
  sky130_fd_sc_hd__buf_8 U13579 ( .A(n11122), .X(n12405) );
  sky130_fd_sc_hd__buf_8 U13580 ( .A(n11122), .X(n12404) );
  sky130_fd_sc_hd__buf_8 U13581 ( .A(n11037), .X(n11001) );
  sky130_fd_sc_hd__buf_8 U13582 ( .A(n11037), .X(n11002) );
  sky130_fd_sc_hd__buf_8 U13583 ( .A(n11037), .X(n11123) );
  sky130_fd_sc_hd__buf_8 U13584 ( .A(n11122), .X(n12413) );
  sky130_fd_sc_hd__buf_8 U13585 ( .A(n11122), .X(n11018) );
  sky130_fd_sc_hd__buf_8 U13586 ( .A(n29494), .X(n11003) );
  sky130_fd_sc_hd__buf_8 U13587 ( .A(n29494), .X(n11004) );
  sky130_fd_sc_hd__buf_8 U13589 ( .A(n29488), .X(n11005) );
  sky130_fd_sc_hd__buf_8 U13591 ( .A(n29488), .X(n11006) );
  sky130_fd_sc_hd__buf_8 U13592 ( .A(n29488), .X(n11007) );
  sky130_fd_sc_hd__inv_6 U13593 ( .A(n11008), .Y(n11009) );
  sky130_fd_sc_hd__inv_6 U13594 ( .A(n11010), .Y(n11011) );
  sky130_fd_sc_hd__buf_8 U13598 ( .A(n29499), .X(n11014) );
  sky130_fd_sc_hd__buf_8 U13599 ( .A(n29499), .X(n11015) );
  sky130_fd_sc_hd__buf_8 U13600 ( .A(n29499), .X(n11101) );
  sky130_fd_sc_hd__buf_8 U13601 ( .A(n29499), .X(n11090) );
  sky130_fd_sc_hd__buf_8 U13602 ( .A(n29494), .X(n11016) );
  sky130_fd_sc_hd__buf_8 U13603 ( .A(n29494), .X(n11017) );
  sky130_fd_sc_hd__buf_8 U13604 ( .A(n29494), .X(n11121) );
  sky130_fd_sc_hd__buf_8 U13605 ( .A(n29494), .X(n11088) );
  sky130_fd_sc_hd__buf_8 U13606 ( .A(n29494), .X(n12539) );
  sky130_fd_sc_hd__buf_8 U13607 ( .A(n11122), .X(n11019) );
  sky130_fd_sc_hd__buf_8 U13608 ( .A(n11122), .X(n11097) );
  sky130_fd_sc_hd__buf_8 U13609 ( .A(n11037), .X(n11020) );
  sky130_fd_sc_hd__buf_8 U13610 ( .A(n11037), .X(n11021) );
  sky130_fd_sc_hd__inv_4 U13611 ( .A(n11089), .Y(n11022) );
  sky130_fd_sc_hd__inv_8 U13612 ( .A(n11089), .Y(n11023) );
  sky130_fd_sc_hd__inv_8 U13613 ( .A(n11089), .Y(n11024) );
  sky130_fd_sc_hd__inv_8 U13614 ( .A(n11089), .Y(n11025) );
  sky130_fd_sc_hd__inv_6 U13615 ( .A(n11026), .Y(n11027) );
  sky130_fd_sc_hd__inv_6 U13616 ( .A(n11026), .Y(n11028) );
  sky130_fd_sc_hd__inv_6 U13617 ( .A(n11026), .Y(n11029) );
  sky130_fd_sc_hd__inv_6 U13618 ( .A(n11026), .Y(n11030) );
  sky130_fd_sc_hd__buf_8 U13619 ( .A(n29488), .X(n11031) );
  sky130_fd_sc_hd__buf_8 U13620 ( .A(n29488), .X(n11087) );
  sky130_fd_sc_hd__buf_8 U13621 ( .A(n12533), .X(n11032) );
  sky130_fd_sc_hd__buf_8 U13622 ( .A(n12533), .X(n11033) );
  sky130_fd_sc_hd__buf_8 U13623 ( .A(n12533), .X(n11034) );
  sky130_fd_sc_hd__buf_8 U13624 ( .A(n12533), .X(n11035) );
  sky130_fd_sc_hd__clkinv_1 U13627 ( .A(n18672), .Y(n18229) );
  sky130_fd_sc_hd__clkinv_1 U13628 ( .A(n22685), .Y(n18142) );
  sky130_fd_sc_hd__inv_1 U13629 ( .A(n18599), .Y(n18337) );
  sky130_fd_sc_hd__clkinv_1 U13630 ( .A(n18681), .Y(n18531) );
  sky130_fd_sc_hd__clkinv_1 U13631 ( .A(n16578), .Y(n16881) );
  sky130_fd_sc_hd__clkinv_1 U13632 ( .A(n15423), .Y(n15424) );
  sky130_fd_sc_hd__inv_2 U13633 ( .A(n17063), .Y(n17064) );
  sky130_fd_sc_hd__clkinv_1 U13634 ( .A(n14862), .Y(n14895) );
  sky130_fd_sc_hd__clkinv_1 U13635 ( .A(n15845), .Y(n17044) );
  sky130_fd_sc_hd__clkinv_1 U13636 ( .A(n17082), .Y(n14903) );
  sky130_fd_sc_hd__nand2_2 U13637 ( .A(n17506), .B(n12139), .Y(n18515) );
  sky130_fd_sc_hd__buf_2 U13639 ( .A(j202_soc_core_j22_cpu_ml_bufb[8]), .X(
        n18654) );
  sky130_fd_sc_hd__clkinv_1 U13640 ( .A(n20442), .Y(n20527) );
  sky130_fd_sc_hd__clkinv_1 U13641 ( .A(n20526), .Y(n20515) );
  sky130_fd_sc_hd__clkinv_1 U13642 ( .A(n20668), .Y(n15469) );
  sky130_fd_sc_hd__clkinv_1 U13644 ( .A(n16564), .Y(n14860) );
  sky130_fd_sc_hd__clkinv_1 U13645 ( .A(n16911), .Y(n16947) );
  sky130_fd_sc_hd__clkinv_1 U13646 ( .A(n26427), .Y(n22734) );
  sky130_fd_sc_hd__buf_2 U13647 ( .A(j202_soc_core_j22_cpu_ml_bufb[15]), .X(
        n18651) );
  sky130_fd_sc_hd__buf_2 U13649 ( .A(j202_soc_core_j22_cpu_ml_bufb[14]), .X(
        n18687) );
  sky130_fd_sc_hd__clkinv_1 U13650 ( .A(n17382), .Y(n18628) );
  sky130_fd_sc_hd__inv_1 U13653 ( .A(n21102), .Y(n21103) );
  sky130_fd_sc_hd__clkinv_1 U13654 ( .A(n16688), .Y(n16764) );
  sky130_fd_sc_hd__clkinv_1 U13655 ( .A(n20648), .Y(n15695) );
  sky130_fd_sc_hd__clkinv_1 U13656 ( .A(n20479), .Y(n20678) );
  sky130_fd_sc_hd__clkinv_1 U13657 ( .A(n20499), .Y(n20583) );
  sky130_fd_sc_hd__clkinv_1 U13658 ( .A(n14859), .Y(n16095) );
  sky130_fd_sc_hd__clkinv_1 U13659 ( .A(n21606), .Y(n19298) );
  sky130_fd_sc_hd__clkinv_1 U13660 ( .A(n26326), .Y(n26415) );
  sky130_fd_sc_hd__clkinv_1 U13661 ( .A(n19125), .Y(n17283) );
  sky130_fd_sc_hd__nor2_1 U13662 ( .A(n19381), .B(n16845), .Y(n16180) );
  sky130_fd_sc_hd__clkinv_1 U13664 ( .A(n13388), .Y(n17037) );
  sky130_fd_sc_hd__inv_1 U13665 ( .A(n20054), .Y(n20302) );
  sky130_fd_sc_hd__clkinv_1 U13667 ( .A(n21270), .Y(n21041) );
  sky130_fd_sc_hd__clkinv_1 U13668 ( .A(n16159), .Y(n17161) );
  sky130_fd_sc_hd__clkinv_1 U13669 ( .A(n20377), .Y(n19985) );
  sky130_fd_sc_hd__nand2b_1 U13670 ( .A_N(n20747), .B(n20788), .Y(n21614) );
  sky130_fd_sc_hd__clkinv_1 U13671 ( .A(n20778), .Y(n21681) );
  sky130_fd_sc_hd__clkinv_1 U13672 ( .A(n19121), .Y(n17173) );
  sky130_fd_sc_hd__clkinv_1 U13673 ( .A(n17290), .Y(n17271) );
  sky130_fd_sc_hd__clkinv_1 U13674 ( .A(n25308), .Y(n26423) );
  sky130_fd_sc_hd__clkinv_1 U13676 ( .A(n26315), .Y(n11578) );
  sky130_fd_sc_hd__fa_1 U13677 ( .A(n17722), .B(n17721), .CIN(n17720), .COUT(
        n17745), .SUM(n17758) );
  sky130_fd_sc_hd__inv_1 U13679 ( .A(n12677), .Y(n13077) );
  sky130_fd_sc_hd__clkinv_1 U13681 ( .A(n25415), .Y(n26432) );
  sky130_fd_sc_hd__clkinv_1 U13682 ( .A(j202_soc_core_j22_cpu_regop_Ra__0_), 
        .Y(n13750) );
  sky130_fd_sc_hd__clkinv_1 U13684 ( .A(n16956), .Y(n20580) );
  sky130_fd_sc_hd__clkinv_1 U13686 ( .A(n21620), .Y(n21269) );
  sky130_fd_sc_hd__clkinv_1 U13688 ( .A(n20312), .Y(n20080) );
  sky130_fd_sc_hd__clkinv_1 U13690 ( .A(n20110), .Y(n19112) );
  sky130_fd_sc_hd__clkinv_1 U13691 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .Y(n12136) );
  sky130_fd_sc_hd__nand2b_1 U13692 ( .A_N(n17211), .B(n17173), .Y(n19971) );
  sky130_fd_sc_hd__clkinv_1 U13695 ( .A(n20247), .Y(n19901) );
  sky130_fd_sc_hd__clkinv_1 U13696 ( .A(n20118), .Y(n19847) );
  sky130_fd_sc_hd__clkinv_1 U13697 ( .A(n19969), .Y(n19830) );
  sky130_fd_sc_hd__clkinv_1 U13699 ( .A(j202_soc_core_j22_cpu_regop_Ra__1_), 
        .Y(n13751) );
  sky130_fd_sc_hd__clkinv_1 U13700 ( .A(n19483), .Y(n21881) );
  sky130_fd_sc_hd__inv_1 U13701 ( .A(n21449), .Y(n21450) );
  sky130_fd_sc_hd__nand2_1 U13702 ( .A(n27388), .B(n26323), .Y(n11570) );
  sky130_fd_sc_hd__inv_2 U13704 ( .A(n27690), .Y(n27692) );
  sky130_fd_sc_hd__inv_1 U13705 ( .A(n19736), .Y(n19719) );
  sky130_fd_sc_hd__clkinv_1 U13706 ( .A(n23109), .Y(n16471) );
  sky130_fd_sc_hd__nor2_1 U13707 ( .A(n22723), .B(n27428), .Y(n13142) );
  sky130_fd_sc_hd__clkinv_1 U13708 ( .A(n26971), .Y(n26702) );
  sky130_fd_sc_hd__nand2_1 U13709 ( .A(j202_soc_core_memory0_ram_dout0[144]), 
        .B(n21592), .Y(n11354) );
  sky130_fd_sc_hd__inv_1 U13710 ( .A(n24357), .Y(n24340) );
  sky130_fd_sc_hd__clkinv_1 U13711 ( .A(n21706), .Y(n19271) );
  sky130_fd_sc_hd__clkinv_1 U13712 ( .A(n20328), .Y(n20058) );
  sky130_fd_sc_hd__clkinv_1 U13714 ( .A(n20906), .Y(n20912) );
  sky130_fd_sc_hd__maj3_1 U13715 ( .A(j202_soc_core_intc_core_00_rg_ipr[71]), 
        .B(n27989), .C(n19507), .X(n19511) );
  sky130_fd_sc_hd__clkinv_1 U13716 ( .A(n13603), .Y(n11144) );
  sky130_fd_sc_hd__nand2_1 U13717 ( .A(j202_soc_core_memory0_ram_dout0[477]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12966) );
  sky130_fd_sc_hd__nand2_1 U13719 ( .A(n17154), .B(io_in[14]), .Y(n17137) );
  sky130_fd_sc_hd__clkinv_1 U13720 ( .A(n16090), .Y(n15384) );
  sky130_fd_sc_hd__o211ai_1 U13723 ( .A1(n26352), .A2(n27388), .B1(n26422), 
        .C1(n11570), .Y(n11569) );
  sky130_fd_sc_hd__inv_2 U13725 ( .A(n21524), .Y(n11986) );
  sky130_fd_sc_hd__clkinv_1 U13726 ( .A(n27364), .Y(n12111) );
  sky130_fd_sc_hd__inv_1 U13729 ( .A(n25538), .Y(n19821) );
  sky130_fd_sc_hd__maj3_1 U13730 ( .A(j202_soc_core_intc_core_00_rg_ipr[75]), 
        .B(n27509), .C(n19515), .X(n19519) );
  sky130_fd_sc_hd__clkinv_1 U13734 ( .A(n22187), .Y(n22520) );
  sky130_fd_sc_hd__clkinv_1 U13735 ( .A(j202_soc_core_j22_cpu_ml_bufa[28]), 
        .Y(n17370) );
  sky130_fd_sc_hd__clkinv_1 U13736 ( .A(n22951), .Y(n17417) );
  sky130_fd_sc_hd__clkinv_1 U13738 ( .A(n23850), .Y(n23851) );
  sky130_fd_sc_hd__o211a_2 U13739 ( .A1(n24088), .A2(n24087), .B1(n24086), 
        .C1(n24090), .X(n13196) );
  sky130_fd_sc_hd__nor2_2 U13740 ( .A(n13570), .B(n13571), .Y(n18865) );
  sky130_fd_sc_hd__inv_2 U13741 ( .A(n17827), .Y(n19425) );
  sky130_fd_sc_hd__nand2_1 U13743 ( .A(n11521), .B(n23789), .Y(n11486) );
  sky130_fd_sc_hd__clkinv_1 U13744 ( .A(n14725), .Y(n14288) );
  sky130_fd_sc_hd__nor2_1 U13747 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[1]), .B(
        n23000), .Y(n26539) );
  sky130_fd_sc_hd__o22ai_1 U13748 ( .A1(n29077), .A2(n27892), .B1(n27891), 
        .B2(n12581), .Y(n27897) );
  sky130_fd_sc_hd__inv_2 U13749 ( .A(n11758), .Y(n12670) );
  sky130_fd_sc_hd__a22oi_1 U13750 ( .A1(j202_soc_core_memory0_ram_dout0[393]), 
        .A2(n21597), .B1(n21735), .B2(j202_soc_core_memory0_ram_dout0[233]), 
        .Y(n20936) );
  sky130_fd_sc_hd__a22oi_1 U13751 ( .A1(j202_soc_core_memory0_ram_dout0[201]), 
        .A2(n21732), .B1(n21591), .B2(j202_soc_core_memory0_ram_dout0[105]), 
        .Y(n20938) );
  sky130_fd_sc_hd__nand2_1 U13754 ( .A(n21771), .B(n21677), .Y(n21738) );
  sky130_fd_sc_hd__inv_1 U13755 ( .A(n12895), .Y(n15752) );
  sky130_fd_sc_hd__inv_2 U13756 ( .A(n26847), .Y(n26849) );
  sky130_fd_sc_hd__inv_2 U13757 ( .A(n14852), .Y(n11907) );
  sky130_fd_sc_hd__nand3_1 U13758 ( .A(n13228), .B(n13227), .C(n22286), .Y(
        n13229) );
  sky130_fd_sc_hd__o31a_1 U13759 ( .A1(n25417), .A2(n26352), .A3(n12353), .B1(
        n25416), .X(n25418) );
  sky130_fd_sc_hd__clkinv_1 U13760 ( .A(n27856), .Y(n27097) );
  sky130_fd_sc_hd__clkinv_1 U13761 ( .A(n27864), .Y(n27764) );
  sky130_fd_sc_hd__clkinv_1 U13762 ( .A(n27850), .Y(n27760) );
  sky130_fd_sc_hd__clkinv_1 U13763 ( .A(n11584), .Y(n11583) );
  sky130_fd_sc_hd__o211ai_1 U13764 ( .A1(n26352), .A2(n27382), .B1(n26422), 
        .C1(n11765), .Y(n25047) );
  sky130_fd_sc_hd__clkinv_1 U13765 ( .A(n12079), .Y(n12078) );
  sky130_fd_sc_hd__nand2_1 U13766 ( .A(n11486), .B(n12352), .Y(n11463) );
  sky130_fd_sc_hd__inv_1 U13767 ( .A(n27415), .Y(n26893) );
  sky130_fd_sc_hd__inv_2 U13768 ( .A(n21887), .Y(n17585) );
  sky130_fd_sc_hd__nor2_1 U13769 ( .A(n23585), .B(n12480), .Y(n11839) );
  sky130_fd_sc_hd__inv_1 U13770 ( .A(n27774), .Y(n24421) );
  sky130_fd_sc_hd__clkinv_1 U13772 ( .A(n26840), .Y(n25770) );
  sky130_fd_sc_hd__nand3_1 U13773 ( .A(n11086), .B(n11543), .C(n11541), .Y(
        n11540) );
  sky130_fd_sc_hd__clkinv_1 U13774 ( .A(j202_soc_core_j22_cpu_regop_We__1_), 
        .Y(n23481) );
  sky130_fd_sc_hd__clkinv_1 U13775 ( .A(n25417), .Y(n23746) );
  sky130_fd_sc_hd__clkinv_1 U13777 ( .A(n27232), .Y(n11130) );
  sky130_fd_sc_hd__clkbuf_1 U13778 ( .A(n13152), .X(n11793) );
  sky130_fd_sc_hd__a22oi_1 U13780 ( .A1(j202_soc_core_memory0_ram_dout0[257]), 
        .A2(n21605), .B1(n21603), .B2(j202_soc_core_memory0_ram_dout0[289]), 
        .Y(n19927) );
  sky130_fd_sc_hd__a21oi_1 U13782 ( .A1(n19041), .A2(n16513), .B1(n14459), .Y(
        n26790) );
  sky130_fd_sc_hd__nand2_1 U13783 ( .A(n20712), .B(n12232), .Y(n12041) );
  sky130_fd_sc_hd__inv_2 U13784 ( .A(n26530), .Y(n12629) );
  sky130_fd_sc_hd__buf_4 U13785 ( .A(j202_soc_core_j22_cpu_ml_bufa[11]), .X(
        n18147) );
  sky130_fd_sc_hd__clkbuf_1 U13786 ( .A(j202_soc_core_j22_cpu_ml_bufa[26]), 
        .X(n25085) );
  sky130_fd_sc_hd__clkbuf_1 U13787 ( .A(n12052), .X(n12051) );
  sky130_fd_sc_hd__clkbuf_1 U13788 ( .A(n27388), .X(n12389) );
  sky130_fd_sc_hd__o22ai_1 U13789 ( .A1(n12618), .A2(n25218), .B1(n11713), 
        .B2(n25217), .Y(n25117) );
  sky130_fd_sc_hd__nor2_1 U13790 ( .A(n23557), .B(n23556), .Y(n26516) );
  sky130_fd_sc_hd__inv_2 U13791 ( .A(n11609), .Y(n11608) );
  sky130_fd_sc_hd__nor2_1 U13793 ( .A(n12380), .B(n23804), .Y(n24704) );
  sky130_fd_sc_hd__inv_1 U13794 ( .A(n20942), .Y(n20955) );
  sky130_fd_sc_hd__clkinv_1 U13795 ( .A(n24087), .Y(n11770) );
  sky130_fd_sc_hd__clkinv_1 U13796 ( .A(j202_soc_core_ahb2wbqspi_00_stb_o), 
        .Y(n26131) );
  sky130_fd_sc_hd__clkinv_1 U13797 ( .A(n26897), .Y(n11157) );
  sky130_fd_sc_hd__inv_2 U13801 ( .A(n12728), .Y(n12715) );
  sky130_fd_sc_hd__clkinv_1 U13802 ( .A(j202_soc_core_intc_core_00_rg_ipr[6]), 
        .Y(n27544) );
  sky130_fd_sc_hd__clkinv_1 U13803 ( .A(j202_soc_core_intc_core_00_rg_ipr[43]), 
        .Y(n25463) );
  sky130_fd_sc_hd__clkinv_1 U13804 ( .A(j202_soc_core_intc_core_00_rg_ipr[49]), 
        .Y(n25718) );
  sky130_fd_sc_hd__clkinv_1 U13805 ( .A(j202_soc_core_intc_core_00_rg_ipr[33]), 
        .Y(n25480) );
  sky130_fd_sc_hd__clkinv_1 U13806 ( .A(j202_soc_core_intc_core_00_rg_ipr[62]), 
        .Y(n25486) );
  sky130_fd_sc_hd__clkinv_1 U13807 ( .A(j202_soc_core_intc_core_00_rg_ipr[50]), 
        .Y(n25502) );
  sky130_fd_sc_hd__clkinv_1 U13808 ( .A(j202_soc_core_intc_core_00_rg_ipr[78]), 
        .Y(n27705) );
  sky130_fd_sc_hd__clkinv_1 U13809 ( .A(j202_soc_core_intc_core_00_rg_ipr[30]), 
        .Y(n27101) );
  sky130_fd_sc_hd__clkinv_1 U13811 ( .A(n27983), .Y(n27740) );
  sky130_fd_sc_hd__clkinv_1 U13812 ( .A(n28215), .Y(n28115) );
  sky130_fd_sc_hd__clkinv_1 U13813 ( .A(n28723), .Y(n28734) );
  sky130_fd_sc_hd__inv_1 U13814 ( .A(n27574), .Y(n11109) );
  sky130_fd_sc_hd__clkinv_1 U13815 ( .A(n27360), .Y(n27125) );
  sky130_fd_sc_hd__inv_2 U13817 ( .A(n24633), .Y(n24629) );
  sky130_fd_sc_hd__inv_2 U13818 ( .A(n11770), .Y(n27427) );
  sky130_fd_sc_hd__clkinv_1 U13819 ( .A(j202_soc_core_intr_req_), .Y(n25782)
         );
  sky130_fd_sc_hd__clkinv_1 U13820 ( .A(n29079), .Y(n11756) );
  sky130_fd_sc_hd__nand2_2 U13821 ( .A(n25293), .B(n23072), .Y(n12355) );
  sky130_fd_sc_hd__nand2b_1 U13822 ( .A_N(n23856), .B(n12365), .Y(n26946) );
  sky130_fd_sc_hd__clkinv_1 U13823 ( .A(n29237), .Y(n26240) );
  sky130_fd_sc_hd__clkinv_1 U13824 ( .A(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n28901) );
  sky130_fd_sc_hd__clkbuf_1 U13825 ( .A(n10674), .X(n29316) );
  sky130_fd_sc_hd__inv_1 U13828 ( .A(n12024), .Y(n28917) );
  sky130_fd_sc_hd__inv_1 U13832 ( .A(n29078), .Y(n10552) );
  sky130_fd_sc_hd__inv_2 U13836 ( .A(n23758), .Y(n11519) );
  sky130_fd_sc_hd__inv_2 U13837 ( .A(n23758), .Y(n11546) );
  sky130_fd_sc_hd__and2_1 U13838 ( .A(n14384), .B(n14382), .X(n11044) );
  sky130_fd_sc_hd__o21a_4 U13841 ( .A1(n26352), .A2(n24048), .B1(n11608), .X(
        n11047) );
  sky130_fd_sc_hd__and2_1 U13842 ( .A(n11839), .B(n11075), .X(n11048) );
  sky130_fd_sc_hd__nand2_1 U13843 ( .A(n26315), .B(n26553), .Y(n27395) );
  sky130_fd_sc_hd__inv_2 U13844 ( .A(n27566), .Y(n12475) );
  sky130_fd_sc_hd__and2_1 U13845 ( .A(n16034), .B(n16033), .X(n11049) );
  sky130_fd_sc_hd__or2_2 U13847 ( .A(n29535), .B(n27275), .X(n11051) );
  sky130_fd_sc_hd__o21a_1 U13850 ( .A1(n21892), .A2(n21889), .B1(n21890), .X(
        n11054) );
  sky130_fd_sc_hd__and2_1 U13851 ( .A(n22311), .B(n22310), .X(n11055) );
  sky130_fd_sc_hd__and2_1 U13852 ( .A(n20717), .B(n21750), .X(n11056) );
  sky130_fd_sc_hd__o211ai_1 U13853 ( .A1(n26703), .A2(n11143), .B1(n15411), 
        .C1(n15410), .Y(n11057) );
  sky130_fd_sc_hd__xor2_1 U13854 ( .A(j202_soc_core_j22_cpu_ml_bufa[19]), .B(
        j202_soc_core_j22_cpu_ml_bufa[18]), .X(n11058) );
  sky130_fd_sc_hd__and4_1 U13855 ( .A(n13170), .B(n13174), .C(n13166), .D(
        n20131), .X(n11059) );
  sky130_fd_sc_hd__and2_1 U13857 ( .A(n21814), .B(n21776), .X(n11061) );
  sky130_fd_sc_hd__and2_1 U13858 ( .A(n22505), .B(n12295), .X(n11062) );
  sky130_fd_sc_hd__a22o_1 U13859 ( .A1(n27347), .A2(n22515), .B1(n26887), .B2(
        n16824), .X(n11063) );
  sky130_fd_sc_hd__and2_1 U13860 ( .A(n14403), .B(n11044), .X(n11064) );
  sky130_fd_sc_hd__and2_1 U13862 ( .A(n21378), .B(n21377), .X(n11065) );
  sky130_fd_sc_hd__nand2_1 U13863 ( .A(n24335), .B(n24265), .Y(n24354) );
  sky130_fd_sc_hd__and2_1 U13864 ( .A(n12886), .B(n12885), .X(n11066) );
  sky130_fd_sc_hd__and2_1 U13866 ( .A(n24465), .B(n24464), .X(n12167) );
  sky130_fd_sc_hd__and3_2 U13868 ( .A(n19168), .B(n19166), .C(n19167), .X(
        n12451) );
  sky130_fd_sc_hd__and2_1 U13869 ( .A(n17131), .B(n17128), .X(n11067) );
  sky130_fd_sc_hd__and2_1 U13870 ( .A(n13145), .B(n13144), .X(n11068) );
  sky130_fd_sc_hd__nand3_2 U13871 ( .A(n21523), .B(n12690), .C(n21521), .Y(
        n12493) );
  sky130_fd_sc_hd__inv_1 U13872 ( .A(n26538), .Y(n23742) );
  sky130_fd_sc_hd__nor2_2 U13873 ( .A(n12559), .B(n23185), .Y(n12480) );
  sky130_fd_sc_hd__and2_1 U13874 ( .A(n10970), .B(n11675), .X(n11069) );
  sky130_fd_sc_hd__and3_1 U13875 ( .A(n27692), .B(n27691), .C(n29075), .X(
        n11070) );
  sky130_fd_sc_hd__and2_1 U13877 ( .A(n11533), .B(n24264), .X(n11071) );
  sky130_fd_sc_hd__and2_1 U13878 ( .A(n24656), .B(n24093), .X(n11072) );
  sky130_fd_sc_hd__and2_1 U13879 ( .A(n11839), .B(n11836), .X(n11073) );
  sky130_fd_sc_hd__and2_1 U13880 ( .A(n27781), .B(n27782), .X(n11074) );
  sky130_fd_sc_hd__and2_1 U13882 ( .A(n11833), .B(n13159), .X(n11075) );
  sky130_fd_sc_hd__inv_2 U13884 ( .A(n13189), .Y(n12395) );
  sky130_fd_sc_hd__and2_1 U13887 ( .A(n11937), .B(n11974), .X(n11079) );
  sky130_fd_sc_hd__buf_8 U13888 ( .A(n29501), .X(n12410) );
  sky130_fd_sc_hd__buf_8 U13889 ( .A(n29499), .X(n12402) );
  sky130_fd_sc_hd__buf_8 U13890 ( .A(n29499), .X(n12407) );
  sky130_fd_sc_hd__and3_1 U13896 ( .A(n11895), .B(n29035), .C(n12898), .X(
        n11081) );
  sky130_fd_sc_hd__and2_1 U13897 ( .A(n12899), .B(n12301), .X(n11082) );
  sky130_fd_sc_hd__inv_8 U13899 ( .A(n23817), .Y(n29248) );
  sky130_fd_sc_hd__buf_8 U13901 ( .A(n29488), .X(n29247) );
  sky130_fd_sc_hd__buf_8 U13902 ( .A(n29488), .X(n12401) );
  sky130_fd_sc_hd__buf_8 U13903 ( .A(n29488), .X(n12406) );
  sky130_fd_sc_hd__buf_8 U13904 ( .A(n11037), .X(n11099) );
  sky130_fd_sc_hd__buf_8 U13906 ( .A(n29494), .X(n12540) );
  sky130_fd_sc_hd__a21oi_2 U13911 ( .A1(n24001), .A2(n27045), .B1(n24000), .Y(
        n12124) );
  sky130_fd_sc_hd__a21o_1 U13912 ( .A1(n24480), .A2(n26407), .B1(n11544), .X(
        n11086) );
  sky130_fd_sc_hd__nand2_2 U13914 ( .A(n11546), .B(n12619), .Y(n26507) );
  sky130_fd_sc_hd__nor2_2 U13915 ( .A(n12516), .B(n25073), .Y(n12363) );
  sky130_fd_sc_hd__nor2_2 U13917 ( .A(n23147), .B(n23159), .Y(n13050) );
  sky130_fd_sc_hd__a21oi_2 U13918 ( .A1(n22398), .A2(n22103), .B1(n22102), .Y(
        n22892) );
  sky130_fd_sc_hd__nand2_2 U13919 ( .A(n21340), .B(n12233), .Y(n11811) );
  sky130_fd_sc_hd__o22ai_1 U13926 ( .A1(n27213), .A2(n11551), .B1(n27212), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N2817) );
  sky130_fd_sc_hd__nand3_1 U13929 ( .A(n27300), .B(n24102), .C(n11734), .Y(
        n10501) );
  sky130_fd_sc_hd__inv_2 U13931 ( .A(n12151), .Y(n11120) );
  sky130_fd_sc_hd__o22ai_1 U13932 ( .A1(n27333), .A2(n11551), .B1(n23178), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N3076) );
  sky130_fd_sc_hd__nor2_1 U13933 ( .A(n11050), .B(n25662), .Y(n25661) );
  sky130_fd_sc_hd__inv_4 U13934 ( .A(n24686), .Y(n27463) );
  sky130_fd_sc_hd__nor2_1 U13935 ( .A(n23188), .B(n23189), .Y(n24414) );
  sky130_fd_sc_hd__and2_1 U13936 ( .A(n26393), .B(n26450), .X(n12256) );
  sky130_fd_sc_hd__clkinv_1 U13938 ( .A(n24060), .Y(n21842) );
  sky130_fd_sc_hd__nand2_1 U13939 ( .A(n25326), .B(n29535), .Y(n11600) );
  sky130_fd_sc_hd__nand3_1 U13940 ( .A(n24464), .B(n22768), .C(n24465), .Y(
        n22551) );
  sky130_fd_sc_hd__nor2_1 U13942 ( .A(n25118), .B(n25117), .Y(n25193) );
  sky130_fd_sc_hd__a21oi_1 U13944 ( .A1(n24659), .A2(n25815), .B1(n24658), .Y(
        n25813) );
  sky130_fd_sc_hd__nor3_1 U13945 ( .A(n27883), .B(n27882), .C(n12679), .Y(
        n27884) );
  sky130_fd_sc_hd__clkinv_1 U13946 ( .A(n12423), .Y(n12424) );
  sky130_fd_sc_hd__nor3_1 U13947 ( .A(n22283), .B(n24409), .C(n24410), .Y(
        n22288) );
  sky130_fd_sc_hd__nand3_1 U13948 ( .A(n13065), .B(n24166), .C(n13064), .Y(
        n24465) );
  sky130_fd_sc_hd__inv_1 U13949 ( .A(n27882), .Y(n27229) );
  sky130_fd_sc_hd__clkinv_1 U13950 ( .A(n12581), .Y(n24387) );
  sky130_fd_sc_hd__nand2_1 U13951 ( .A(n23232), .B(n26863), .Y(n24700) );
  sky130_fd_sc_hd__nand2_1 U13952 ( .A(n23231), .B(n26863), .Y(n24166) );
  sky130_fd_sc_hd__a211oi_1 U13953 ( .A1(n12499), .A2(n22702), .B1(n12500), 
        .C1(n22610), .Y(n12498) );
  sky130_fd_sc_hd__inv_2 U13954 ( .A(n24639), .Y(n27297) );
  sky130_fd_sc_hd__inv_1 U13955 ( .A(n24367), .Y(n24369) );
  sky130_fd_sc_hd__xnor2_1 U13957 ( .A(n22529), .B(n22528), .Y(n23247) );
  sky130_fd_sc_hd__a21oi_1 U13958 ( .A1(n23829), .A2(n23828), .B1(n18916), .Y(
        n23852) );
  sky130_fd_sc_hd__or2_0 U13959 ( .A(n11141), .B(n27461), .X(n11647) );
  sky130_fd_sc_hd__clkinv_1 U13961 ( .A(n27823), .Y(n24119) );
  sky130_fd_sc_hd__inv_2 U13962 ( .A(n11589), .Y(n27401) );
  sky130_fd_sc_hd__inv_2 U13963 ( .A(n11611), .Y(n27461) );
  sky130_fd_sc_hd__o211ai_1 U13964 ( .A1(n23068), .A2(n18916), .B1(n23067), 
        .C1(n23066), .Y(n23069) );
  sky130_fd_sc_hd__o21ai_1 U13965 ( .A1(n21453), .A2(n22912), .B1(n21452), .Y(
        n21454) );
  sky130_fd_sc_hd__nand2_1 U13966 ( .A(n24437), .B(n23141), .Y(n24452) );
  sky130_fd_sc_hd__o211a_2 U13967 ( .A1(n26356), .A2(n18916), .B1(n26355), 
        .C1(n26354), .X(n26357) );
  sky130_fd_sc_hd__nand2_1 U13968 ( .A(n12351), .B(n23002), .Y(n23014) );
  sky130_fd_sc_hd__clkinv_1 U13969 ( .A(n23203), .Y(n23204) );
  sky130_fd_sc_hd__nand2_1 U13970 ( .A(n11519), .B(n26548), .Y(n12351) );
  sky130_fd_sc_hd__clkinv_1 U13971 ( .A(n13146), .Y(n13143) );
  sky130_fd_sc_hd__or2_0 U13973 ( .A(n21869), .B(n11457), .X(n11451) );
  sky130_fd_sc_hd__inv_2 U13974 ( .A(n23735), .Y(n12359) );
  sky130_fd_sc_hd__clkinv_1 U13975 ( .A(n19794), .Y(n19815) );
  sky130_fd_sc_hd__nand2_1 U13976 ( .A(n12587), .B(n20958), .Y(n29014) );
  sky130_fd_sc_hd__and2_1 U13977 ( .A(n11491), .B(n11489), .X(n19200) );
  sky130_fd_sc_hd__nor2_1 U13978 ( .A(n23201), .B(n24404), .Y(n23208) );
  sky130_fd_sc_hd__clkinv_1 U13979 ( .A(n19816), .Y(n19796) );
  sky130_fd_sc_hd__nand3_2 U13980 ( .A(n13234), .B(n13235), .C(n20963), .Y(
        n29009) );
  sky130_fd_sc_hd__nand3_1 U13982 ( .A(n11488), .B(n18889), .C(n21505), .Y(
        n11495) );
  sky130_fd_sc_hd__clkinv_1 U13983 ( .A(n22272), .Y(n12472) );
  sky130_fd_sc_hd__nor2_1 U13984 ( .A(n21498), .B(n18872), .Y(n22750) );
  sky130_fd_sc_hd__a21oi_1 U13985 ( .A1(n20955), .A2(n20956), .B1(n12191), .Y(
        n12496) );
  sky130_fd_sc_hd__nand3_2 U13986 ( .A(n20962), .B(n20960), .C(n20961), .Y(
        n29077) );
  sky130_fd_sc_hd__clkinv_1 U13987 ( .A(n27575), .Y(n11108) );
  sky130_fd_sc_hd__and2_0 U13988 ( .A(n11140), .B(n21792), .X(n12194) );
  sky130_fd_sc_hd__and2_0 U13989 ( .A(n21339), .B(n21750), .X(n12233) );
  sky130_fd_sc_hd__nand2b_1 U13990 ( .A_N(n27956), .B(n22026), .Y(n27947) );
  sky130_fd_sc_hd__a21oi_2 U13991 ( .A1(n18902), .A2(n18904), .B1(n18831), .Y(
        n22907) );
  sky130_fd_sc_hd__nor2_1 U13992 ( .A(n18819), .B(n12322), .Y(n21418) );
  sky130_fd_sc_hd__and2_1 U13993 ( .A(n20987), .B(n21776), .X(n11706) );
  sky130_fd_sc_hd__clkinv_1 U13995 ( .A(n21437), .Y(n21439) );
  sky130_fd_sc_hd__clkinv_1 U13996 ( .A(n21967), .Y(n22846) );
  sky130_fd_sc_hd__inv_1 U13998 ( .A(n20137), .Y(n20138) );
  sky130_fd_sc_hd__nand2_1 U13999 ( .A(n11498), .B(n11497), .Y(n13280) );
  sky130_fd_sc_hd__a21boi_0 U14000 ( .A1(n20802), .A2(n20801), .B1_N(n20800), 
        .Y(n20816) );
  sky130_fd_sc_hd__clkinv_1 U14001 ( .A(n18593), .Y(n11415) );
  sky130_fd_sc_hd__inv_1 U14002 ( .A(n21012), .Y(n15509) );
  sky130_fd_sc_hd__clkinv_1 U14003 ( .A(n18010), .Y(n12685) );
  sky130_fd_sc_hd__clkinv_1 U14004 ( .A(n17497), .Y(n17492) );
  sky130_fd_sc_hd__inv_2 U14005 ( .A(n23070), .Y(n26708) );
  sky130_fd_sc_hd__nand3_1 U14006 ( .A(n14154), .B(n12217), .C(n14153), .Y(
        n23070) );
  sky130_fd_sc_hd__clkinv_1 U14007 ( .A(n18587), .Y(n18561) );
  sky130_fd_sc_hd__inv_1 U14008 ( .A(n20329), .Y(n20104) );
  sky130_fd_sc_hd__clkinv_1 U14009 ( .A(n18588), .Y(n11416) );
  sky130_fd_sc_hd__a31o_1 U14010 ( .A1(n19381), .A2(n19380), .A3(n11994), .B1(
        n21043), .X(n19386) );
  sky130_fd_sc_hd__or2_0 U14011 ( .A(n20111), .B(n20110), .X(n20881) );
  sky130_fd_sc_hd__clkinv_1 U14012 ( .A(n16173), .Y(n16745) );
  sky130_fd_sc_hd__clkinv_1 U14013 ( .A(n20199), .Y(n20114) );
  sky130_fd_sc_hd__inv_2 U14014 ( .A(n12159), .Y(n18751) );
  sky130_fd_sc_hd__clkinv_1 U14015 ( .A(n15863), .Y(n16094) );
  sky130_fd_sc_hd__inv_2 U14016 ( .A(n14642), .Y(n11112) );
  sky130_fd_sc_hd__inv_2 U14017 ( .A(n14143), .Y(n11111) );
  sky130_fd_sc_hd__clkinv_1 U14018 ( .A(n20372), .Y(n19832) );
  sky130_fd_sc_hd__inv_2 U14019 ( .A(n15062), .Y(n11114) );
  sky130_fd_sc_hd__inv_2 U14020 ( .A(n15063), .Y(n11113) );
  sky130_fd_sc_hd__inv_2 U14021 ( .A(n14476), .Y(n11116) );
  sky130_fd_sc_hd__nor2_2 U14022 ( .A(n19413), .B(n24778), .Y(n26323) );
  sky130_fd_sc_hd__inv_1 U14023 ( .A(n13632), .Y(n13633) );
  sky130_fd_sc_hd__nand2_2 U14024 ( .A(n13577), .B(n17357), .Y(n27456) );
  sky130_fd_sc_hd__clkinv_1 U14025 ( .A(n17165), .Y(n17287) );
  sky130_fd_sc_hd__clkinv_1 U14026 ( .A(n20570), .Y(n20676) );
  sky130_fd_sc_hd__and2_0 U14027 ( .A(n18871), .B(n17357), .X(n12135) );
  sky130_fd_sc_hd__inv_4 U14028 ( .A(n12170), .Y(n11093) );
  sky130_fd_sc_hd__nand2_2 U14029 ( .A(n25219), .B(n17359), .Y(n26977) );
  sky130_fd_sc_hd__inv_2 U14030 ( .A(n14476), .Y(n11094) );
  sky130_fd_sc_hd__inv_2 U14032 ( .A(n13683), .Y(n23109) );
  sky130_fd_sc_hd__clkinv_1 U14033 ( .A(n18865), .Y(n13572) );
  sky130_fd_sc_hd__inv_2 U14035 ( .A(n14288), .Y(n11096) );
  sky130_fd_sc_hd__buf_2 U14036 ( .A(n13398), .X(n20687) );
  sky130_fd_sc_hd__and3_1 U14037 ( .A(n13751), .B(n13750), .C(
        j202_soc_core_intr_req_), .X(n13752) );
  sky130_fd_sc_hd__buf_4 U14038 ( .A(n17363), .X(n18719) );
  sky130_fd_sc_hd__nor2_1 U14039 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .B(n24282), .Y(n17356) );
  sky130_fd_sc_hd__inv_1 U14040 ( .A(j202_soc_core_j22_cpu_ml_bufa[20]), .Y(
        n22142) );
  sky130_fd_sc_hd__nor2_1 U14041 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[3]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[5]), .Y(n26682) );
  sky130_fd_sc_hd__buf_2 U14042 ( .A(j202_soc_core_j22_cpu_ml_bufa[30]), .X(
        n24505) );
  sky130_fd_sc_hd__a211oi_1 U14043 ( .A1(n27203), .A2(n26855), .B1(n29059), 
        .C1(n26854), .Y(n26856) );
  sky130_fd_sc_hd__inv_1 U14044 ( .A(n29069), .Y(n26902) );
  sky130_fd_sc_hd__nor2_1 U14045 ( .A(n11443), .B(n26976), .Y(n24065) );
  sky130_fd_sc_hd__and2_1 U14047 ( .A(n27273), .B(n12299), .X(n12157) );
  sky130_fd_sc_hd__and2_1 U14048 ( .A(n27273), .B(n12298), .X(n12156) );
  sky130_fd_sc_hd__buf_4 U14049 ( .A(n11083), .X(n29268) );
  sky130_fd_sc_hd__buf_4 U14050 ( .A(n11083), .X(n29267) );
  sky130_fd_sc_hd__and2_1 U14053 ( .A(n12355), .B(n26450), .X(n24561) );
  sky130_fd_sc_hd__nand3_1 U14055 ( .A(n22289), .B(n12377), .C(n22288), .Y(
        n28973) );
  sky130_fd_sc_hd__clkinv_1 U14057 ( .A(n24702), .Y(n24412) );
  sky130_fd_sc_hd__nand3_1 U14058 ( .A(n11465), .B(n11754), .C(n26103), .Y(
        n26105) );
  sky130_fd_sc_hd__inv_2 U14059 ( .A(n27441), .Y(n27448) );
  sky130_fd_sc_hd__and2_0 U14060 ( .A(n25075), .B(n25074), .X(n12516) );
  sky130_fd_sc_hd__clkinv_1 U14063 ( .A(n23010), .Y(n22687) );
  sky130_fd_sc_hd__clkbuf_1 U14064 ( .A(n26835), .X(n12125) );
  sky130_fd_sc_hd__or2_0 U14065 ( .A(n22221), .B(n25251), .X(n12262) );
  sky130_fd_sc_hd__nand2_1 U14066 ( .A(n23223), .B(n12177), .Y(n22228) );
  sky130_fd_sc_hd__clkinv_1 U14067 ( .A(n23015), .Y(n23009) );
  sky130_fd_sc_hd__clkinv_1 U14069 ( .A(n11848), .Y(n24424) );
  sky130_fd_sc_hd__inv_1 U14070 ( .A(n27550), .Y(n27555) );
  sky130_fd_sc_hd__a21oi_2 U14071 ( .A1(n23071), .A2(n23070), .B1(n23069), .Y(
        n25293) );
  sky130_fd_sc_hd__nand2_1 U14072 ( .A(n23230), .B(n26863), .Y(n24382) );
  sky130_fd_sc_hd__a21oi_1 U14073 ( .A1(n23241), .A2(n26863), .B1(n25027), .Y(
        n27275) );
  sky130_fd_sc_hd__clkbuf_1 U14074 ( .A(n23249), .X(n26321) );
  sky130_fd_sc_hd__inv_2 U14075 ( .A(n24328), .Y(n23182) );
  sky130_fd_sc_hd__nand2_1 U14076 ( .A(n23247), .B(n26863), .Y(n23978) );
  sky130_fd_sc_hd__and2_0 U14077 ( .A(n11465), .B(n11754), .X(n11464) );
  sky130_fd_sc_hd__nand3_1 U14078 ( .A(n11971), .B(n22671), .C(n22672), .Y(
        n23179) );
  sky130_fd_sc_hd__nand2_1 U14079 ( .A(n23242), .B(n26863), .Y(n18878) );
  sky130_fd_sc_hd__clkinv_1 U14080 ( .A(n25148), .Y(n22689) );
  sky130_fd_sc_hd__clkinv_1 U14081 ( .A(n24550), .Y(n26402) );
  sky130_fd_sc_hd__nand4_1 U14082 ( .A(n24091), .B(n27947), .C(n27256), .D(
        n27772), .Y(n23962) );
  sky130_fd_sc_hd__clkinv_1 U14083 ( .A(n22610), .Y(n11991) );
  sky130_fd_sc_hd__inv_2 U14084 ( .A(n12324), .Y(n22219) );
  sky130_fd_sc_hd__nand3_1 U14085 ( .A(n11653), .B(n12112), .C(n23046), .Y(
        n23071) );
  sky130_fd_sc_hd__xnor2_1 U14086 ( .A(n12481), .B(n18907), .Y(n23223) );
  sky130_fd_sc_hd__nand2_1 U14087 ( .A(n11661), .B(n26352), .Y(n11557) );
  sky130_fd_sc_hd__inv_1 U14089 ( .A(n24452), .Y(n24453) );
  sky130_fd_sc_hd__nor2_1 U14090 ( .A(n23570), .B(n12658), .Y(n23820) );
  sky130_fd_sc_hd__nor2_1 U14091 ( .A(n19198), .B(n25232), .Y(n22218) );
  sky130_fd_sc_hd__nand3_1 U14092 ( .A(n20980), .B(n20981), .C(n29593), .Y(
        n11914) );
  sky130_fd_sc_hd__inv_2 U14093 ( .A(n23014), .Y(n11104) );
  sky130_fd_sc_hd__inv_2 U14094 ( .A(n27957), .Y(n11105) );
  sky130_fd_sc_hd__o211a_2 U14095 ( .A1(n11564), .A2(n27395), .B1(n11562), 
        .C1(n11560), .X(n11559) );
  sky130_fd_sc_hd__inv_1 U14096 ( .A(n27421), .Y(n24592) );
  sky130_fd_sc_hd__inv_2 U14098 ( .A(n24350), .Y(n11106) );
  sky130_fd_sc_hd__inv_1 U14100 ( .A(n23583), .Y(n22284) );
  sky130_fd_sc_hd__and2_1 U14102 ( .A(n22669), .B(n29347), .X(n11973) );
  sky130_fd_sc_hd__clkinv_1 U14103 ( .A(n26831), .Y(n27207) );
  sky130_fd_sc_hd__nor2_1 U14104 ( .A(n24123), .B(n11942), .Y(n17133) );
  sky130_fd_sc_hd__nand4_1 U14105 ( .A(n13069), .B(n21917), .C(n13067), .D(
        n13066), .Y(n27453) );
  sky130_fd_sc_hd__nor2_1 U14106 ( .A(n21023), .B(n28919), .Y(n17129) );
  sky130_fd_sc_hd__inv_1 U14107 ( .A(n25771), .Y(n25772) );
  sky130_fd_sc_hd__clkbuf_1 U14108 ( .A(n19247), .X(n19160) );
  sky130_fd_sc_hd__nand3_1 U14109 ( .A(n29562), .B(n11494), .C(n11495), .Y(
        n11491) );
  sky130_fd_sc_hd__and2_1 U14110 ( .A(n11495), .B(n11494), .X(n21961) );
  sky130_fd_sc_hd__clkinv_1 U14112 ( .A(n22754), .Y(n21910) );
  sky130_fd_sc_hd__clkinv_1 U14113 ( .A(n23694), .Y(n29329) );
  sky130_fd_sc_hd__nor2_1 U14114 ( .A(n11153), .B(n22717), .Y(n12985) );
  sky130_fd_sc_hd__o22a_1 U14115 ( .A1(n26314), .A2(n26313), .B1(n26312), .B2(
        n26311), .X(n26555) );
  sky130_fd_sc_hd__and2_0 U14117 ( .A(n21814), .B(n22581), .X(n17004) );
  sky130_fd_sc_hd__nand2_1 U14118 ( .A(n28950), .B(n22712), .Y(n22717) );
  sky130_fd_sc_hd__clkinv_1 U14119 ( .A(n12877), .Y(n28971) );
  sky130_fd_sc_hd__clkinv_1 U14120 ( .A(n11747), .Y(n21793) );
  sky130_fd_sc_hd__inv_2 U14121 ( .A(n26536), .Y(n13068) );
  sky130_fd_sc_hd__nand2_1 U14122 ( .A(n11944), .B(n11943), .Y(n11942) );
  sky130_fd_sc_hd__clkinv_1 U14123 ( .A(n19444), .Y(n21804) );
  sky130_fd_sc_hd__clkinv_1 U14124 ( .A(n26535), .Y(n23763) );
  sky130_fd_sc_hd__clkinv_1 U14125 ( .A(n19481), .Y(n21874) );
  sky130_fd_sc_hd__clkinv_1 U14126 ( .A(n21788), .Y(n21789) );
  sky130_fd_sc_hd__clkinv_1 U14127 ( .A(n27213), .Y(n23106) );
  sky130_fd_sc_hd__nor2_1 U14128 ( .A(n18809), .B(n18808), .Y(n21498) );
  sky130_fd_sc_hd__clkinv_1 U14129 ( .A(n22243), .Y(n21518) );
  sky130_fd_sc_hd__clkinv_1 U14130 ( .A(n27221), .Y(n11136) );
  sky130_fd_sc_hd__or2_0 U14131 ( .A(n28590), .B(n24996), .X(n23442) );
  sky130_fd_sc_hd__o211a_2 U14132 ( .A1(n26581), .A2(n11143), .B1(n20996), 
        .C1(n20995), .X(n12213) );
  sky130_fd_sc_hd__nand2_1 U14136 ( .A(n29562), .B(n29574), .Y(n11489) );
  sky130_fd_sc_hd__clkinv_1 U14137 ( .A(n19482), .Y(n21873) );
  sky130_fd_sc_hd__clkinv_1 U14138 ( .A(n21909), .Y(n22753) );
  sky130_fd_sc_hd__inv_2 U14139 ( .A(n27124), .Y(n11141) );
  sky130_fd_sc_hd__nand3_2 U14140 ( .A(n23177), .B(n23038), .C(n23037), .Y(
        n23039) );
  sky130_fd_sc_hd__clkinv_1 U14141 ( .A(n22389), .Y(n22103) );
  sky130_fd_sc_hd__clkinv_1 U14143 ( .A(n21773), .Y(n19403) );
  sky130_fd_sc_hd__clkinv_1 U14145 ( .A(n21584), .Y(n16824) );
  sky130_fd_sc_hd__and2_0 U14146 ( .A(n24795), .B(n12694), .X(n11373) );
  sky130_fd_sc_hd__clkinv_1 U14147 ( .A(n22747), .Y(n22749) );
  sky130_fd_sc_hd__nor2_1 U14148 ( .A(n21805), .B(n21808), .Y(n11493) );
  sky130_fd_sc_hd__clkinv_1 U14149 ( .A(n15660), .Y(n15661) );
  sky130_fd_sc_hd__inv_2 U14150 ( .A(n22510), .Y(n11143) );
  sky130_fd_sc_hd__clkinv_1 U14151 ( .A(n20828), .Y(n20831) );
  sky130_fd_sc_hd__clkinv_1 U14152 ( .A(n19743), .Y(n19768) );
  sky130_fd_sc_hd__clkinv_1 U14153 ( .A(n22832), .Y(n22833) );
  sky130_fd_sc_hd__nor2_1 U14154 ( .A(n28590), .B(n14849), .Y(n12072) );
  sky130_fd_sc_hd__clkinv_1 U14155 ( .A(n17924), .Y(n12318) );
  sky130_fd_sc_hd__clkinv_1 U14156 ( .A(n17111), .Y(n16986) );
  sky130_fd_sc_hd__clkinv_1 U14157 ( .A(n20032), .Y(n20043) );
  sky130_fd_sc_hd__clkinv_1 U14158 ( .A(n22180), .Y(n22181) );
  sky130_fd_sc_hd__nor2_1 U14159 ( .A(n18273), .B(n18274), .Y(n21980) );
  sky130_fd_sc_hd__nand2_1 U14160 ( .A(n13280), .B(n12208), .Y(n17869) );
  sky130_fd_sc_hd__clkinv_1 U14161 ( .A(n19415), .Y(n21531) );
  sky130_fd_sc_hd__and3_1 U14162 ( .A(n13603), .B(
        j202_soc_core_j22_cpu_memop_Ma__0_), .C(n13649), .X(n22510) );
  sky130_fd_sc_hd__inv_1 U14163 ( .A(n15412), .Y(n15771) );
  sky130_fd_sc_hd__clkinv_1 U14164 ( .A(n21889), .Y(n21891) );
  sky130_fd_sc_hd__clkinv_1 U14165 ( .A(n20421), .Y(n20422) );
  sky130_fd_sc_hd__nor2_1 U14166 ( .A(n18833), .B(n18834), .Y(n22902) );
  sky130_fd_sc_hd__and2_0 U14167 ( .A(n15420), .B(n15419), .X(n15421) );
  sky130_fd_sc_hd__clkinv_1 U14168 ( .A(n16987), .Y(n16811) );
  sky130_fd_sc_hd__clkinv_1 U14169 ( .A(n18594), .Y(n11422) );
  sky130_fd_sc_hd__o2bb2ai_1 U14170 ( .B1(n11145), .B2(n26424), .A1_N(n26077), 
        .A2_N(n23070), .Y(n21831) );
  sky130_fd_sc_hd__clkinv_1 U14172 ( .A(n16651), .Y(n17115) );
  sky130_fd_sc_hd__clkinv_1 U14173 ( .A(n18455), .Y(n18458) );
  sky130_fd_sc_hd__clkinv_1 U14174 ( .A(n21446), .Y(n18842) );
  sky130_fd_sc_hd__and2_0 U14175 ( .A(n22305), .B(n22304), .X(n11625) );
  sky130_fd_sc_hd__or2_0 U14176 ( .A(n25835), .B(n25836), .X(n25837) );
  sky130_fd_sc_hd__or2_0 U14177 ( .A(n28590), .B(n24761), .X(n27312) );
  sky130_fd_sc_hd__or2_0 U14178 ( .A(n28590), .B(n24753), .X(n27676) );
  sky130_fd_sc_hd__inv_1 U14179 ( .A(n19173), .Y(n19179) );
  sky130_fd_sc_hd__or2_1 U14182 ( .A(n17864), .B(n17865), .X(n12208) );
  sky130_fd_sc_hd__clkinv_1 U14183 ( .A(n18852), .Y(n11503) );
  sky130_fd_sc_hd__nand2_1 U14184 ( .A(n22825), .B(n22824), .Y(n22826) );
  sky130_fd_sc_hd__or2_0 U14185 ( .A(n17860), .B(n17861), .X(n12364) );
  sky130_fd_sc_hd__clkinv_1 U14186 ( .A(n17496), .Y(n17493) );
  sky130_fd_sc_hd__clkinv_1 U14187 ( .A(n22397), .Y(n11478) );
  sky130_fd_sc_hd__nor2_1 U14188 ( .A(n11949), .B(n14388), .Y(n11948) );
  sky130_fd_sc_hd__or2_0 U14189 ( .A(n21969), .B(n21968), .X(n21970) );
  sky130_fd_sc_hd__inv_2 U14190 ( .A(n26724), .Y(n25128) );
  sky130_fd_sc_hd__clkinv_1 U14191 ( .A(n18600), .Y(n18338) );
  sky130_fd_sc_hd__a2bb2oi_1 U14192 ( .B1(n22731), .B2(n26724), .A1_N(n18916), 
        .A2_N(n22771), .Y(n22732) );
  sky130_fd_sc_hd__inv_1 U14193 ( .A(n21385), .Y(n21387) );
  sky130_fd_sc_hd__inv_2 U14194 ( .A(n26712), .Y(n27007) );
  sky130_fd_sc_hd__clkinv_1 U14195 ( .A(n19366), .Y(n19338) );
  sky130_fd_sc_hd__xnor3_1 U14196 ( .A(n12994), .B(n18072), .C(n18073), .X(
        n18032) );
  sky130_fd_sc_hd__nand3_1 U14197 ( .A(n16260), .B(n16259), .C(n16258), .Y(
        n26716) );
  sky130_fd_sc_hd__or2_0 U14198 ( .A(n22887), .B(n22893), .X(n22397) );
  sky130_fd_sc_hd__clkinv_1 U14199 ( .A(n22719), .Y(n17817) );
  sky130_fd_sc_hd__or2_0 U14200 ( .A(n20083), .B(n20082), .X(n20084) );
  sky130_fd_sc_hd__and2_0 U14201 ( .A(n13600), .B(n23487), .X(n11913) );
  sky130_fd_sc_hd__clkinv_1 U14202 ( .A(n20188), .Y(n19988) );
  sky130_fd_sc_hd__clkinv_1 U14203 ( .A(n24113), .Y(n24291) );
  sky130_fd_sc_hd__clkinv_1 U14204 ( .A(n19967), .Y(n17172) );
  sky130_fd_sc_hd__clkinv_1 U14205 ( .A(n21220), .Y(n21051) );
  sky130_fd_sc_hd__clkinv_1 U14206 ( .A(n20617), .Y(n20478) );
  sky130_fd_sc_hd__clkinv_1 U14207 ( .A(n16853), .Y(n16183) );
  sky130_fd_sc_hd__clkinv_1 U14208 ( .A(n21224), .Y(n21084) );
  sky130_fd_sc_hd__clkinv_1 U14209 ( .A(n16719), .Y(n16593) );
  sky130_fd_sc_hd__clkinv_1 U14210 ( .A(n15714), .Y(n15722) );
  sky130_fd_sc_hd__or2_0 U14211 ( .A(n20294), .B(n20349), .X(n20115) );
  sky130_fd_sc_hd__clkinv_1 U14212 ( .A(n21205), .Y(n21219) );
  sky130_fd_sc_hd__clkinv_1 U14213 ( .A(n16715), .Y(n16716) );
  sky130_fd_sc_hd__inv_2 U14214 ( .A(n17365), .Y(n22071) );
  sky130_fd_sc_hd__or2_0 U14215 ( .A(n20219), .B(n20918), .X(n20240) );
  sky130_fd_sc_hd__or2_0 U14216 ( .A(n22096), .B(n22097), .X(n22357) );
  sky130_fd_sc_hd__clkinv_1 U14217 ( .A(n20862), .Y(n20325) );
  sky130_fd_sc_hd__clkinv_1 U14218 ( .A(n16673), .Y(n16886) );
  sky130_fd_sc_hd__clkinv_1 U14219 ( .A(n21632), .Y(n21715) );
  sky130_fd_sc_hd__or2_0 U14220 ( .A(n22422), .B(n22423), .X(n22679) );
  sky130_fd_sc_hd__or2_0 U14221 ( .A(n22420), .B(n22418), .X(n22474) );
  sky130_fd_sc_hd__or2_0 U14222 ( .A(n22390), .B(n22391), .X(n22553) );
  sky130_fd_sc_hd__or2_0 U14223 ( .A(n20096), .B(n20058), .X(n20113) );
  sky130_fd_sc_hd__clkinv_1 U14224 ( .A(n20099), .Y(n17223) );
  sky130_fd_sc_hd__or2_0 U14225 ( .A(n16787), .B(n16620), .X(n16715) );
  sky130_fd_sc_hd__or2_0 U14226 ( .A(n20348), .B(n20114), .X(n20900) );
  sky130_fd_sc_hd__clkinv_1 U14227 ( .A(n20380), .Y(n17220) );
  sky130_fd_sc_hd__a22o_1 U14228 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[13]), .B1(n18183), .B2(
        j202_soc_core_j22_cpu_ml_macl[29]), .X(n18322) );
  sky130_fd_sc_hd__clkinv_1 U14229 ( .A(n21287), .Y(n17288) );
  sky130_fd_sc_hd__clkinv_1 U14230 ( .A(n15853), .Y(n14870) );
  sky130_fd_sc_hd__clkinv_1 U14231 ( .A(n16905), .Y(n16783) );
  sky130_fd_sc_hd__clkinv_1 U14232 ( .A(n20007), .Y(n19898) );
  sky130_fd_sc_hd__clkinv_1 U14233 ( .A(n16858), .Y(n16873) );
  sky130_fd_sc_hd__nor2_1 U14234 ( .A(n18295), .B(n23253), .Y(n17365) );
  sky130_fd_sc_hd__clkinv_1 U14235 ( .A(n20219), .Y(n19878) );
  sky130_fd_sc_hd__or2_0 U14236 ( .A(n22466), .B(n13278), .X(n22468) );
  sky130_fd_sc_hd__clkinv_1 U14237 ( .A(n17735), .Y(n11623) );
  sky130_fd_sc_hd__clkinv_1 U14238 ( .A(n20117), .Y(n20301) );
  sky130_fd_sc_hd__or2_0 U14239 ( .A(n16094), .B(n15864), .X(n15879) );
  sky130_fd_sc_hd__clkinv_1 U14240 ( .A(n20664), .Y(n20448) );
  sky130_fd_sc_hd__clkinv_1 U14241 ( .A(n21184), .Y(n21268) );
  sky130_fd_sc_hd__clkinv_1 U14242 ( .A(n17049), .Y(n15874) );
  sky130_fd_sc_hd__nand2b_1 U14243 ( .A_N(n21206), .B(n20623), .Y(n20884) );
  sky130_fd_sc_hd__or2_0 U14244 ( .A(n12159), .B(n22465), .X(n13278) );
  sky130_fd_sc_hd__clkinv_1 U14245 ( .A(n16840), .Y(n16562) );
  sky130_fd_sc_hd__and2_0 U14246 ( .A(n23322), .B(n24293), .X(n12147) );
  sky130_fd_sc_hd__inv_2 U14247 ( .A(n15062), .Y(n11150) );
  sky130_fd_sc_hd__inv_2 U14248 ( .A(n14143), .Y(n11151) );
  sky130_fd_sc_hd__clkinv_1 U14249 ( .A(n20376), .Y(n20917) );
  sky130_fd_sc_hd__inv_2 U14250 ( .A(n14642), .Y(n11152) );
  sky130_fd_sc_hd__o2bb2ai_1 U14251 ( .B1(n11156), .B2(n23172), .A1_N(n23080), 
        .A2_N(n23174), .Y(n23081) );
  sky130_fd_sc_hd__clkinv_1 U14252 ( .A(n17167), .Y(n17164) );
  sky130_fd_sc_hd__o22ai_1 U14253 ( .A1(n17972), .A2(n17405), .B1(n17441), 
        .B2(n11159), .Y(n17411) );
  sky130_fd_sc_hd__clkinv_1 U14254 ( .A(n18861), .Y(n17360) );
  sky130_fd_sc_hd__o2bb2ai_1 U14255 ( .B1(n11164), .B2(n23172), .A1_N(n23104), 
        .A2_N(n23174), .Y(n23105) );
  sky130_fd_sc_hd__or2_0 U14256 ( .A(n23011), .B(n24778), .X(n26407) );
  sky130_fd_sc_hd__o2bb2ai_1 U14257 ( .B1(n11165), .B2(n23172), .A1_N(n23036), 
        .A2_N(n23174), .Y(n22998) );
  sky130_fd_sc_hd__clkinv_1 U14258 ( .A(n17376), .Y(n11481) );
  sky130_fd_sc_hd__buf_6 U14259 ( .A(n23130), .X(n11110) );
  sky130_fd_sc_hd__clkinv_1 U14260 ( .A(n16078), .Y(n14922) );
  sky130_fd_sc_hd__inv_1 U14261 ( .A(n14950), .Y(n16172) );
  sky130_fd_sc_hd__clkinv_1 U14262 ( .A(n15789), .Y(n14921) );
  sky130_fd_sc_hd__o22ai_1 U14263 ( .A1(n17719), .A2(n17972), .B1(n17718), 
        .B2(n11159), .Y(n11499) );
  sky130_fd_sc_hd__and2_0 U14264 ( .A(n20632), .B(n11994), .X(n15437) );
  sky130_fd_sc_hd__clkinv_1 U14265 ( .A(n15818), .Y(n15846) );
  sky130_fd_sc_hd__clkinv_1 U14266 ( .A(n14902), .Y(n14880) );
  sky130_fd_sc_hd__clkinv_1 U14267 ( .A(n20665), .Y(n15688) );
  sky130_fd_sc_hd__inv_4 U14268 ( .A(n23076), .Y(n11156) );
  sky130_fd_sc_hd__inv_1 U14269 ( .A(n14877), .Y(n14885) );
  sky130_fd_sc_hd__o22ai_1 U14270 ( .A1(n17972), .A2(n17695), .B1(n17708), 
        .B2(n11159), .Y(n17724) );
  sky130_fd_sc_hd__clkinv_1 U14271 ( .A(n14951), .Y(n14856) );
  sky130_fd_sc_hd__and2_0 U14272 ( .A(n22034), .B(n14752), .X(n11915) );
  sky130_fd_sc_hd__inv_2 U14273 ( .A(n14288), .Y(n11160) );
  sky130_fd_sc_hd__or2_0 U14274 ( .A(n25231), .B(n25338), .X(n12298) );
  sky130_fd_sc_hd__or2_0 U14275 ( .A(n25339), .B(n25338), .X(n12299) );
  sky130_fd_sc_hd__clkinv_1 U14276 ( .A(n16516), .Y(n16005) );
  sky130_fd_sc_hd__clkinv_1 U14278 ( .A(n15557), .Y(n15630) );
  sky130_fd_sc_hd__nand3_2 U14279 ( .A(n23922), .B(n18916), .C(n23927), .Y(
        n24778) );
  sky130_fd_sc_hd__inv_2 U14280 ( .A(n12186), .Y(n16363) );
  sky130_fd_sc_hd__clkinv_1 U14281 ( .A(n16170), .Y(n15458) );
  sky130_fd_sc_hd__clkinv_1 U14282 ( .A(n20626), .Y(n13429) );
  sky130_fd_sc_hd__clkinv_1 U14283 ( .A(n11514), .Y(n11513) );
  sky130_fd_sc_hd__clkinv_1 U14284 ( .A(n14898), .Y(n14879) );
  sky130_fd_sc_hd__o22ai_1 U14285 ( .A1(n18750), .A2(n18230), .B1(n18229), 
        .B2(n18747), .Y(n18330) );
  sky130_fd_sc_hd__buf_4 U14286 ( .A(n18515), .X(n18424) );
  sky130_fd_sc_hd__or2b_4 U14287 ( .A(n26682), .B_N(n26691), .X(n18916) );
  sky130_fd_sc_hd__nor2b_1 U14290 ( .B_N(n18353), .A(n12367), .Y(n17454) );
  sky130_fd_sc_hd__clkinv_1 U14291 ( .A(n19013), .Y(n13725) );
  sky130_fd_sc_hd__a22oi_1 U14292 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__15_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__15_), .Y(n20977) );
  sky130_fd_sc_hd__inv_4 U14293 ( .A(n12171), .Y(n11165) );
  sky130_fd_sc_hd__inv_4 U14294 ( .A(n12172), .Y(n11164) );
  sky130_fd_sc_hd__clkinv_1 U14295 ( .A(n16126), .Y(n14881) );
  sky130_fd_sc_hd__or2_0 U14296 ( .A(j202_soc_core_qspi_wb_addr[14]), .B(
        n23385), .X(n23387) );
  sky130_fd_sc_hd__or2_0 U14297 ( .A(j202_soc_core_qspi_wb_addr[13]), .B(
        n23383), .X(n23384) );
  sky130_fd_sc_hd__or2_0 U14298 ( .A(j202_soc_core_qspi_wb_addr[18]), .B(
        n23418), .X(n23420) );
  sky130_fd_sc_hd__or2_0 U14299 ( .A(j202_soc_core_qspi_wb_addr[12]), .B(
        n23396), .X(n23397) );
  sky130_fd_sc_hd__buf_2 U14300 ( .A(n17393), .X(n17805) );
  sky130_fd_sc_hd__or2_0 U14301 ( .A(j202_soc_core_qspi_wb_addr[11]), .B(
        n23398), .X(n23400) );
  sky130_fd_sc_hd__or2_0 U14302 ( .A(j202_soc_core_qspi_wb_addr[4]), .B(n23374), .X(n23373) );
  sky130_fd_sc_hd__or2_0 U14303 ( .A(j202_soc_core_qspi_wb_addr[16]), .B(
        n23411), .X(n23413) );
  sky130_fd_sc_hd__clkinv_1 U14304 ( .A(n22487), .Y(n18302) );
  sky130_fd_sc_hd__clkinv_1 U14305 ( .A(n13702), .Y(n13699) );
  sky130_fd_sc_hd__or2_0 U14306 ( .A(j202_soc_core_qspi_wb_addr[3]), .B(n23470), .X(n23376) );
  sky130_fd_sc_hd__or2_0 U14307 ( .A(j202_soc_core_qspi_wb_addr[22]), .B(
        n23432), .X(n23434) );
  sky130_fd_sc_hd__or2_0 U14308 ( .A(j202_soc_core_qspi_wb_addr[10]), .B(
        n23390), .X(n23391) );
  sky130_fd_sc_hd__clkinv_1 U14309 ( .A(n18863), .Y(n23252) );
  sky130_fd_sc_hd__clkbuf_1 U14310 ( .A(j202_soc_core_j22_cpu_ml_bufa[16]), 
        .X(n12577) );
  sky130_fd_sc_hd__or2_0 U14311 ( .A(j202_soc_core_qspi_wb_addr[20]), .B(
        n23425), .X(n23427) );
  sky130_fd_sc_hd__or2_0 U14312 ( .A(j202_soc_core_qspi_wb_addr[9]), .B(n23392), .X(n23393) );
  sky130_fd_sc_hd__or2_0 U14313 ( .A(j202_soc_core_qspi_wb_addr[6]), .B(n23361), .X(n23360) );
  sky130_fd_sc_hd__clkinv_1 U14316 ( .A(n19508), .Y(n19510) );
  sky130_fd_sc_hd__or2_0 U14317 ( .A(j202_soc_core_qspi_wb_addr[8]), .B(n23352), .X(n23354) );
  sky130_fd_sc_hd__or2_0 U14318 ( .A(j202_soc_core_qspi_wb_addr[7]), .B(n23358), .X(n23355) );
  sky130_fd_sc_hd__clkinv_1 U14319 ( .A(j202_soc_core_j22_cpu_regop_Rn__1_), 
        .Y(n13614) );
  sky130_fd_sc_hd__clkinv_1 U14320 ( .A(n13698), .Y(n13563) );
  sky130_fd_sc_hd__clkinv_1 U14321 ( .A(n24019), .Y(n11166) );
  sky130_fd_sc_hd__or2_0 U14322 ( .A(j202_soc_core_qspi_wb_addr[19]), .B(
        n23344), .X(n23345) );
  sky130_fd_sc_hd__or2_1 U14323 ( .A(n13665), .B(n13684), .X(n12172) );
  sky130_fd_sc_hd__or2_0 U14324 ( .A(j202_soc_core_qspi_wb_addr[21]), .B(
        n23341), .X(n23343) );
  sky130_fd_sc_hd__inv_1 U14325 ( .A(j202_soc_core_j22_cpu_ml_bufa[6]), .Y(
        n25339) );
  sky130_fd_sc_hd__or2_0 U14326 ( .A(j202_soc_core_qspi_wb_addr[15]), .B(
        n23349), .X(n23351) );
  sky130_fd_sc_hd__or2_0 U14327 ( .A(j202_soc_core_qspi_wb_addr[5]), .B(n23371), .X(n23363) );
  sky130_fd_sc_hd__or2_0 U14328 ( .A(j202_soc_core_qspi_wb_addr[17]), .B(
        n23346), .X(n23348) );
  sky130_fd_sc_hd__nor2_1 U14329 ( .A(j202_soc_core_j22_cpu_macop_MAC_[3]), 
        .B(j202_soc_core_j22_cpu_macop_MAC_[2]), .Y(n24019) );
  sky130_fd_sc_hd__clkinv_1 U14330 ( .A(j202_soc_core_ahb2apb_01_state[1]), 
        .Y(n24320) );
  sky130_fd_sc_hd__or2_0 U14331 ( .A(start_n_reg[1]), .B(wb_rst_i), .X(n470)
         );
  sky130_fd_sc_hd__inv_2 U14333 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .Y(n15454) );
  sky130_fd_sc_hd__buf_6 U14334 ( .A(j202_soc_core_rst), .X(n28590) );
  sky130_fd_sc_hd__buf_6 U14335 ( .A(n24181), .X(n29259) );
  sky130_fd_sc_hd__buf_6 U14336 ( .A(n24181), .X(n29260) );
  sky130_fd_sc_hd__nand2_1 U14337 ( .A(n28981), .B(n24225), .Y(n24180) );
  sky130_fd_sc_hd__inv_2 U14338 ( .A(n13014), .Y(n27203) );
  sky130_fd_sc_hd__clkinv_1 U14339 ( .A(n11459), .Y(n11458) );
  sky130_fd_sc_hd__a21oi_1 U14340 ( .A1(n13000), .A2(
        j202_soc_core_j22_cpu_ml_macl[13]), .B1(n25286), .Y(n25288) );
  sky130_fd_sc_hd__a21oi_1 U14341 ( .A1(n13000), .A2(
        j202_soc_core_j22_cpu_ml_macl[7]), .B1(n24741), .Y(n24744) );
  sky130_fd_sc_hd__nand3_1 U14342 ( .A(n11756), .B(n27981), .C(n11755), .Y(
        n10593) );
  sky130_fd_sc_hd__and2_1 U14345 ( .A(n12802), .B(n26450), .X(n12271) );
  sky130_fd_sc_hd__inv_1 U14346 ( .A(n29016), .Y(n10548) );
  sky130_fd_sc_hd__inv_1 U14347 ( .A(n29028), .Y(n10544) );
  sky130_fd_sc_hd__inv_2 U14348 ( .A(n29020), .Y(n10554) );
  sky130_fd_sc_hd__inv_1 U14349 ( .A(n29017), .Y(n10555) );
  sky130_fd_sc_hd__nand2_1 U14350 ( .A(n13021), .B(n13023), .Y(n13015) );
  sky130_fd_sc_hd__inv_1 U14351 ( .A(n29025), .Y(n10545) );
  sky130_fd_sc_hd__inv_2 U14352 ( .A(n29073), .Y(n10546) );
  sky130_fd_sc_hd__inv_1 U14353 ( .A(n29019), .Y(n10556) );
  sky130_fd_sc_hd__inv_1 U14354 ( .A(n29026), .Y(n10547) );
  sky130_fd_sc_hd__inv_2 U14356 ( .A(n29018), .Y(n10557) );
  sky130_fd_sc_hd__inv_2 U14357 ( .A(n29074), .Y(n10558) );
  sky130_fd_sc_hd__inv_1 U14358 ( .A(n29021), .Y(n10551) );
  sky130_fd_sc_hd__inv_4 U14359 ( .A(n11778), .Y(n12161) );
  sky130_fd_sc_hd__and2_1 U14360 ( .A(n26881), .B(n26450), .X(n12272) );
  sky130_fd_sc_hd__inv_2 U14361 ( .A(n29023), .Y(n10550) );
  sky130_fd_sc_hd__inv_1 U14363 ( .A(n12355), .Y(n27462) );
  sky130_fd_sc_hd__nand3_1 U14364 ( .A(n22246), .B(n22371), .C(n11714), .Y(
        n29005) );
  sky130_fd_sc_hd__clkinv_1 U14365 ( .A(n24371), .Y(n24373) );
  sky130_fd_sc_hd__nand3_1 U14367 ( .A(n22309), .B(n22551), .C(n22308), .Y(
        n28977) );
  sky130_fd_sc_hd__nand3_1 U14368 ( .A(n22319), .B(n22220), .C(n12262), .Y(
        n28986) );
  sky130_fd_sc_hd__nand3_1 U14369 ( .A(n11991), .B(n21581), .C(n11990), .Y(
        n28982) );
  sky130_fd_sc_hd__and2_1 U14370 ( .A(n26105), .B(n26450), .X(n13322) );
  sky130_fd_sc_hd__nand3_1 U14372 ( .A(n11073), .B(n24341), .C(n11834), .Y(
        n24342) );
  sky130_fd_sc_hd__nand2_1 U14373 ( .A(n23072), .B(n25293), .Y(n27459) );
  sky130_fd_sc_hd__nand2_1 U14376 ( .A(n24050), .B(n24051), .Y(n24371) );
  sky130_fd_sc_hd__clkinv_1 U14377 ( .A(n24997), .Y(n25002) );
  sky130_fd_sc_hd__inv_1 U14378 ( .A(n13320), .Y(n23280) );
  sky130_fd_sc_hd__nand3_1 U14379 ( .A(n22245), .B(n22768), .C(n22244), .Y(
        n22371) );
  sky130_fd_sc_hd__and2_0 U14380 ( .A(n25111), .B(n13287), .X(n13335) );
  sky130_fd_sc_hd__and2_1 U14382 ( .A(n24686), .B(n26450), .X(n12267) );
  sky130_fd_sc_hd__and2_1 U14383 ( .A(n26514), .B(n24495), .X(n12738) );
  sky130_fd_sc_hd__nand3_1 U14384 ( .A(n11791), .B(n29495), .C(n11509), .Y(
        n11504) );
  sky130_fd_sc_hd__clkinv_1 U14385 ( .A(n11791), .Y(n12153) );
  sky130_fd_sc_hd__clkinv_1 U14387 ( .A(n27571), .Y(n11681) );
  sky130_fd_sc_hd__nand2_2 U14388 ( .A(n25711), .B(n24632), .Y(n25705) );
  sky130_fd_sc_hd__or2_0 U14389 ( .A(n23306), .B(n23305), .X(n13287) );
  sky130_fd_sc_hd__nand3_1 U14390 ( .A(n11470), .B(n11045), .C(n11469), .Y(
        n24997) );
  sky130_fd_sc_hd__nor2_1 U14391 ( .A(n11803), .B(n27595), .Y(n27596) );
  sky130_fd_sc_hd__nor2_1 U14392 ( .A(n27783), .B(n27784), .Y(n11640) );
  sky130_fd_sc_hd__and2_0 U14393 ( .A(n23854), .B(n23853), .X(n23855) );
  sky130_fd_sc_hd__clkbuf_1 U14394 ( .A(n22270), .X(n12387) );
  sky130_fd_sc_hd__nand3_1 U14395 ( .A(n11711), .B(n22239), .C(n22240), .Y(
        n22241) );
  sky130_fd_sc_hd__nor2_1 U14396 ( .A(n29535), .B(n25270), .Y(n11584) );
  sky130_fd_sc_hd__inv_2 U14397 ( .A(n28973), .Y(n11124) );
  sky130_fd_sc_hd__clkinv_1 U14398 ( .A(n23270), .Y(n23271) );
  sky130_fd_sc_hd__clkinv_1 U14399 ( .A(n25744), .Y(n25745) );
  sky130_fd_sc_hd__nand3_1 U14400 ( .A(n11808), .B(n11807), .C(n11806), .Y(
        n11805) );
  sky130_fd_sc_hd__a22o_1 U14401 ( .A1(n12617), .A2(n12035), .B1(n25811), .B2(
        n29072), .X(n24111) );
  sky130_fd_sc_hd__clkinv_1 U14402 ( .A(n24106), .Y(n12114) );
  sky130_fd_sc_hd__and2_1 U14404 ( .A(n25810), .B(n26450), .X(n12268) );
  sky130_fd_sc_hd__or2_0 U14406 ( .A(n27441), .B(n27381), .X(n12252) );
  sky130_fd_sc_hd__or2_0 U14407 ( .A(n27441), .B(n27376), .X(n13277) );
  sky130_fd_sc_hd__or2_0 U14408 ( .A(n27441), .B(n27387), .X(n12253) );
  sky130_fd_sc_hd__a22oi_1 U14409 ( .A1(n25538), .A2(n19820), .B1(n25524), 
        .B2(n19819), .Y(n19826) );
  sky130_fd_sc_hd__or2_0 U14410 ( .A(n27441), .B(n27440), .X(n12251) );
  sky130_fd_sc_hd__and2_0 U14412 ( .A(n27693), .B(n13081), .X(n12278) );
  sky130_fd_sc_hd__nand2_1 U14413 ( .A(n18878), .B(n18877), .Y(n24138) );
  sky130_fd_sc_hd__o21a_1 U14414 ( .A1(n22221), .A2(n25250), .B1(n22217), .X(
        n22220) );
  sky130_fd_sc_hd__nand3_1 U14415 ( .A(n25710), .B(n25709), .C(n25708), .Y(
        n24634) );
  sky130_fd_sc_hd__inv_2 U14416 ( .A(n23225), .Y(n11128) );
  sky130_fd_sc_hd__inv_2 U14417 ( .A(n27883), .Y(n23818) );
  sky130_fd_sc_hd__clkinv_1 U14419 ( .A(n11472), .Y(n11471) );
  sky130_fd_sc_hd__buf_6 U14420 ( .A(n11936), .X(n11129) );
  sky130_fd_sc_hd__o21ai_1 U14421 ( .A1(n26322), .A2(n26321), .B1(n26320), .Y(
        n26359) );
  sky130_fd_sc_hd__nand3_1 U14422 ( .A(n25663), .B(n25665), .C(n25664), .Y(
        n25703) );
  sky130_fd_sc_hd__nor2_1 U14423 ( .A(n23820), .B(n11809), .Y(n11808) );
  sky130_fd_sc_hd__clkinv_1 U14424 ( .A(n24166), .Y(n24167) );
  sky130_fd_sc_hd__clkinv_1 U14426 ( .A(n24382), .Y(n22460) );
  sky130_fd_sc_hd__nand3_1 U14427 ( .A(n26108), .B(n26107), .C(n26106), .Y(
        n26510) );
  sky130_fd_sc_hd__nand2_1 U14428 ( .A(n13197), .B(n13196), .Y(n25662) );
  sky130_fd_sc_hd__clkinv_1 U14429 ( .A(n23975), .Y(n23976) );
  sky130_fd_sc_hd__clkinv_1 U14430 ( .A(n24368), .Y(n12673) );
  sky130_fd_sc_hd__clkinv_1 U14431 ( .A(n24798), .Y(n24771) );
  sky130_fd_sc_hd__nand3_1 U14432 ( .A(n11558), .B(n26718), .C(n11557), .Y(
        n11556) );
  sky130_fd_sc_hd__nand3_1 U14433 ( .A(n25322), .B(n25321), .C(n25320), .Y(
        n25332) );
  sky130_fd_sc_hd__clkinv_1 U14435 ( .A(n23569), .Y(n27788) );
  sky130_fd_sc_hd__a2bb2oi_1 U14436 ( .B1(n25077), .B2(n26948), .A1_N(n25714), 
        .A2_N(n11102), .Y(n25078) );
  sky130_fd_sc_hd__and2_0 U14438 ( .A(n24031), .B(n26329), .X(n12240) );
  sky130_fd_sc_hd__o22ai_1 U14442 ( .A1(n27386), .A2(n27438), .B1(n27450), 
        .B2(n11551), .Y(n27387) );
  sky130_fd_sc_hd__and2_0 U14443 ( .A(n12035), .B(n25815), .X(n12037) );
  sky130_fd_sc_hd__inv_1 U14444 ( .A(n13159), .Y(n13161) );
  sky130_fd_sc_hd__nand2_1 U14445 ( .A(n11815), .B(n27553), .Y(n27776) );
  sky130_fd_sc_hd__nor2_1 U14446 ( .A(n12938), .B(n12935), .Y(n25273) );
  sky130_fd_sc_hd__and2_0 U14447 ( .A(n27952), .B(n27902), .X(n12284) );
  sky130_fd_sc_hd__nand3_1 U14448 ( .A(n12438), .B(n24455), .C(n23185), .Y(
        n11819) );
  sky130_fd_sc_hd__nand3_1 U14449 ( .A(n11520), .B(n25138), .C(n25139), .Y(
        n25191) );
  sky130_fd_sc_hd__and2_0 U14450 ( .A(n18918), .B(n18917), .X(n12177) );
  sky130_fd_sc_hd__and2_1 U14451 ( .A(n26099), .B(n12707), .X(n11754) );
  sky130_fd_sc_hd__inv_2 U14452 ( .A(n22458), .Y(n21843) );
  sky130_fd_sc_hd__o21ba_2 U14453 ( .A1(n22980), .A2(n24066), .B1_N(n22979), 
        .X(n22981) );
  sky130_fd_sc_hd__clkinv_1 U14454 ( .A(n11454), .Y(n11453) );
  sky130_fd_sc_hd__nor2_1 U14456 ( .A(n11554), .B(n11409), .Y(n11553) );
  sky130_fd_sc_hd__xnor2_1 U14457 ( .A(n21455), .B(n21454), .Y(n23248) );
  sky130_fd_sc_hd__nand3_1 U14458 ( .A(n19443), .B(n19441), .C(n19442), .Y(
        n11703) );
  sky130_fd_sc_hd__nand3_1 U14459 ( .A(n11456), .B(n21869), .C(n22619), .Y(
        n11454) );
  sky130_fd_sc_hd__clkinv_1 U14460 ( .A(n12325), .Y(n25241) );
  sky130_fd_sc_hd__o211ai_1 U14462 ( .A1(n27340), .A2(n26859), .B1(n24481), 
        .C1(n23917), .Y(n11483) );
  sky130_fd_sc_hd__nand2_1 U14463 ( .A(n11463), .B(n11548), .Y(n25138) );
  sky130_fd_sc_hd__clkinv_1 U14464 ( .A(n24108), .Y(n23801) );
  sky130_fd_sc_hd__clkinv_1 U14465 ( .A(n23274), .Y(n22614) );
  sky130_fd_sc_hd__nand3_1 U14466 ( .A(n12372), .B(n24661), .C(n12373), .Y(
        n24682) );
  sky130_fd_sc_hd__and2_0 U14467 ( .A(n27899), .B(n27969), .X(n27952) );
  sky130_fd_sc_hd__and2_0 U14468 ( .A(n25225), .B(n17158), .X(n12237) );
  sky130_fd_sc_hd__clkinv_1 U14469 ( .A(n24125), .Y(n17159) );
  sky130_fd_sc_hd__a21oi_1 U14470 ( .A1(n22410), .A2(n26872), .B1(n22409), .Y(
        n23262) );
  sky130_fd_sc_hd__nand3_1 U14471 ( .A(n11053), .B(n11508), .C(n11507), .Y(
        n11506) );
  sky130_fd_sc_hd__nand3_1 U14473 ( .A(n11937), .B(n29515), .C(n17128), .Y(
        n17142) );
  sky130_fd_sc_hd__nor2_1 U14474 ( .A(n21028), .B(n21029), .Y(n22671) );
  sky130_fd_sc_hd__clkinv_1 U14475 ( .A(n20978), .Y(n25225) );
  sky130_fd_sc_hd__nand3_1 U14476 ( .A(n11577), .B(n11576), .C(n11575), .Y(
        n25298) );
  sky130_fd_sc_hd__inv_2 U14477 ( .A(n12744), .Y(n11132) );
  sky130_fd_sc_hd__nor2_1 U14478 ( .A(n23589), .B(n27958), .Y(n11659) );
  sky130_fd_sc_hd__xor2_1 U14479 ( .A(n26508), .B(n26507), .X(n26100) );
  sky130_fd_sc_hd__clkinv_1 U14481 ( .A(n27565), .Y(n24261) );
  sky130_fd_sc_hd__clkinv_1 U14482 ( .A(n12742), .Y(n23800) );
  sky130_fd_sc_hd__xnor2_1 U14483 ( .A(n19225), .B(n19224), .Y(n22410) );
  sky130_fd_sc_hd__nand2_1 U14485 ( .A(n27421), .B(n19440), .Y(n19441) );
  sky130_fd_sc_hd__o211ai_1 U14486 ( .A1(n24680), .A2(n18916), .B1(n24679), 
        .C1(n24678), .Y(n24681) );
  sky130_fd_sc_hd__clkinv_1 U14487 ( .A(n27128), .Y(n27129) );
  sky130_fd_sc_hd__o211a_2 U14488 ( .A1(n26875), .A2(n26398), .B1(n22490), 
        .C1(n22489), .X(n22491) );
  sky130_fd_sc_hd__clkinv_1 U14489 ( .A(n22710), .Y(n22673) );
  sky130_fd_sc_hd__nand2_2 U14490 ( .A(n11521), .B(n12593), .Y(n26064) );
  sky130_fd_sc_hd__nand3_1 U14491 ( .A(n17132), .B(n13292), .C(n17133), .Y(
        n11930) );
  sky130_fd_sc_hd__nand2_1 U14492 ( .A(n21408), .B(n21409), .Y(n13146) );
  sky130_fd_sc_hd__nor2_1 U14493 ( .A(n26773), .B(n26772), .Y(n11727) );
  sky130_fd_sc_hd__clkinv_1 U14494 ( .A(n29030), .Y(n22668) );
  sky130_fd_sc_hd__inv_1 U14495 ( .A(n26901), .Y(n26903) );
  sky130_fd_sc_hd__clkinv_1 U14496 ( .A(n19820), .Y(n25537) );
  sky130_fd_sc_hd__clkinv_1 U14498 ( .A(n19819), .Y(n25523) );
  sky130_fd_sc_hd__and2_0 U14499 ( .A(n13271), .B(n27980), .X(n12227) );
  sky130_fd_sc_hd__clkinv_1 U14500 ( .A(n12421), .Y(n21024) );
  sky130_fd_sc_hd__clkinv_1 U14501 ( .A(n27204), .Y(n25775) );
  sky130_fd_sc_hd__nor2_1 U14503 ( .A(n11043), .B(n11920), .Y(n17138) );
  sky130_fd_sc_hd__a21oi_1 U14504 ( .A1(n22661), .A2(n19230), .B1(n19229), .Y(
        n19231) );
  sky130_fd_sc_hd__nand3_1 U14506 ( .A(n21338), .B(n12196), .C(n21337), .Y(
        n29030) );
  sky130_fd_sc_hd__nand2_1 U14507 ( .A(n12493), .B(n21550), .Y(n11981) );
  sky130_fd_sc_hd__inv_2 U14508 ( .A(n11792), .Y(n12060) );
  sky130_fd_sc_hd__a21o_1 U14509 ( .A1(n21797), .A2(n21788), .B1(n11747), .X(
        n19248) );
  sky130_fd_sc_hd__a2bb2oi_1 U14510 ( .B1(n19800), .B2(n19785), .A1_N(n19794), 
        .A2_N(n19816), .Y(n19792) );
  sky130_fd_sc_hd__inv_2 U14511 ( .A(n27523), .Y(n11133) );
  sky130_fd_sc_hd__clkinv_1 U14512 ( .A(n26689), .Y(n26692) );
  sky130_fd_sc_hd__inv_4 U14513 ( .A(n21511), .Y(n22944) );
  sky130_fd_sc_hd__clkinv_1 U14514 ( .A(n28922), .Y(n21027) );
  sky130_fd_sc_hd__and2_0 U14515 ( .A(n21790), .B(n21788), .X(n13330) );
  sky130_fd_sc_hd__o22ai_1 U14516 ( .A1(n26314), .A2(n23697), .B1(n26312), 
        .B2(n26538), .Y(n12079) );
  sky130_fd_sc_hd__clkinv_1 U14517 ( .A(n12083), .Y(n12082) );
  sky130_fd_sc_hd__nand3_1 U14518 ( .A(n11491), .B(n11489), .C(n11367), .Y(
        n11366) );
  sky130_fd_sc_hd__nand3_1 U14519 ( .A(n12690), .B(n21523), .C(n21521), .Y(
        n27408) );
  sky130_fd_sc_hd__and2_0 U14520 ( .A(n21796), .B(n21790), .X(n21799) );
  sky130_fd_sc_hd__or2_0 U14521 ( .A(n29072), .B(n29071), .X(n12277) );
  sky130_fd_sc_hd__clkinv_1 U14522 ( .A(n26883), .Y(n26884) );
  sky130_fd_sc_hd__o21ba_2 U14523 ( .A1(n21511), .A2(n12780), .B1_N(n22909), 
        .X(n22911) );
  sky130_fd_sc_hd__inv_2 U14524 ( .A(n27258), .Y(n11134) );
  sky130_fd_sc_hd__clkinv_1 U14525 ( .A(n23697), .Y(n29327) );
  sky130_fd_sc_hd__inv_2 U14526 ( .A(n19160), .Y(n21797) );
  sky130_fd_sc_hd__nand2_1 U14528 ( .A(n25071), .B(n25072), .Y(n11554) );
  sky130_fd_sc_hd__nand2_1 U14529 ( .A(n23742), .B(n26539), .Y(n11545) );
  sky130_fd_sc_hd__nand2_1 U14530 ( .A(n23731), .B(n26539), .Y(n11768) );
  sky130_fd_sc_hd__clkinv_1 U14531 ( .A(n23695), .Y(n29325) );
  sky130_fd_sc_hd__nand2_1 U14533 ( .A(n12024), .B(
        j202_soc_core_j22_cpu_ma_M_address[1]), .Y(n13105) );
  sky130_fd_sc_hd__nand2_1 U14534 ( .A(n12510), .B(n21814), .Y(n26537) );
  sky130_fd_sc_hd__nand2b_1 U14535 ( .A_N(n23695), .B(n22712), .Y(n21816) );
  sky130_fd_sc_hd__a21oi_1 U14536 ( .A1(n26096), .A2(n12158), .B1(n11057), .Y(
        n12588) );
  sky130_fd_sc_hd__clkinv_1 U14537 ( .A(n26387), .Y(n26388) );
  sky130_fd_sc_hd__clkinv_1 U14538 ( .A(n24404), .Y(n24405) );
  sky130_fd_sc_hd__clkinv_1 U14539 ( .A(n27720), .Y(
        j202_soc_core_j22_cpu_ifetch) );
  sky130_fd_sc_hd__clkinv_1 U14540 ( .A(n19804), .Y(n19806) );
  sky130_fd_sc_hd__clkinv_1 U14541 ( .A(n19785), .Y(n19801) );
  sky130_fd_sc_hd__clkinv_1 U14542 ( .A(n11700), .Y(n26843) );
  sky130_fd_sc_hd__a21oi_1 U14543 ( .A1(n26710), .A2(n26085), .B1(n11565), .Y(
        n11562) );
  sky130_fd_sc_hd__clkinv_1 U14544 ( .A(n22797), .Y(n22800) );
  sky130_fd_sc_hd__clkinv_1 U14545 ( .A(n22358), .Y(n22133) );
  sky130_fd_sc_hd__clkinv_1 U14546 ( .A(n22798), .Y(n22799) );
  sky130_fd_sc_hd__nand2b_1 U14547 ( .A_N(n26538), .B(n22714), .Y(n21521) );
  sky130_fd_sc_hd__nand2_1 U14549 ( .A(n18816), .B(n22750), .Y(n19246) );
  sky130_fd_sc_hd__clkinv_1 U14550 ( .A(n22940), .Y(n22943) );
  sky130_fd_sc_hd__nand2b_1 U14551 ( .A_N(n23696), .B(n22712), .Y(n19166) );
  sky130_fd_sc_hd__clkinv_1 U14552 ( .A(n22941), .Y(n22942) );
  sky130_fd_sc_hd__clkinv_1 U14553 ( .A(n11959), .Y(n11955) );
  sky130_fd_sc_hd__clkinv_1 U14554 ( .A(n27264), .Y(n27572) );
  sky130_fd_sc_hd__clkbuf_1 U14555 ( .A(n12496), .X(n12771) );
  sky130_fd_sc_hd__nand2_1 U14557 ( .A(n12969), .B(n12130), .Y(n12510) );
  sky130_fd_sc_hd__nor2_1 U14558 ( .A(n20430), .B(n20560), .Y(n28926) );
  sky130_fd_sc_hd__clkbuf_1 U14559 ( .A(n11488), .X(n18886) );
  sky130_fd_sc_hd__clkinv_1 U14560 ( .A(n29034), .Y(n27634) );
  sky130_fd_sc_hd__and2_1 U14561 ( .A(n12616), .B(n26539), .X(n11424) );
  sky130_fd_sc_hd__clkinv_1 U14562 ( .A(n22890), .Y(n22105) );
  sky130_fd_sc_hd__a21o_1 U14563 ( .A1(n25838), .A2(n25837), .B1(n13342), .X(
        n26745) );
  sky130_fd_sc_hd__inv_2 U14564 ( .A(n21448), .Y(n21451) );
  sky130_fd_sc_hd__clkinv_1 U14565 ( .A(n23696), .Y(n29326) );
  sky130_fd_sc_hd__clkinv_1 U14566 ( .A(n12741), .Y(n19480) );
  sky130_fd_sc_hd__clkinv_1 U14567 ( .A(n25147), .Y(n25150) );
  sky130_fd_sc_hd__or2_1 U14568 ( .A(n26548), .B(n26531), .X(n12152) );
  sky130_fd_sc_hd__and3_1 U14569 ( .A(n27942), .B(n27954), .C(n27941), .X(
        n12471) );
  sky130_fd_sc_hd__and2_0 U14570 ( .A(n22471), .B(n22480), .X(n22482) );
  sky130_fd_sc_hd__clkinv_1 U14571 ( .A(n27949), .Y(n23966) );
  sky130_fd_sc_hd__clkinv_1 U14572 ( .A(n21498), .Y(n21500) );
  sky130_fd_sc_hd__o21ai_2 U14573 ( .A1(n24113), .A2(n23560), .B1(n24650), .Y(
        j202_soc_core_j22_cpu_rf_N3371) );
  sky130_fd_sc_hd__a21oi_1 U14574 ( .A1(n22398), .A2(n22165), .B1(n22164), .Y(
        n22941) );
  sky130_fd_sc_hd__clkinv_1 U14575 ( .A(n24703), .Y(n24270) );
  sky130_fd_sc_hd__clkinv_1 U14576 ( .A(n22910), .Y(n12780) );
  sky130_fd_sc_hd__clkbuf_1 U14577 ( .A(n11941), .X(n12616) );
  sky130_fd_sc_hd__clkinv_1 U14578 ( .A(n27977), .Y(n27970) );
  sky130_fd_sc_hd__nand2_1 U14579 ( .A(n22471), .B(n22470), .Y(n22680) );
  sky130_fd_sc_hd__clkinv_1 U14580 ( .A(n22612), .Y(n21578) );
  sky130_fd_sc_hd__inv_1 U14581 ( .A(n11944), .Y(n11889) );
  sky130_fd_sc_hd__clkinv_1 U14582 ( .A(n11963), .Y(n11962) );
  sky130_fd_sc_hd__clkinv_1 U14583 ( .A(n27967), .Y(n24254) );
  sky130_fd_sc_hd__o21ai_1 U14584 ( .A1(n21329), .A2(n21373), .B1(n21328), .Y(
        n21347) );
  sky130_fd_sc_hd__o21ba_2 U14585 ( .A1(n21357), .A2(n21373), .B1_N(n21358), 
        .X(n21363) );
  sky130_fd_sc_hd__clkinv_1 U14586 ( .A(n23693), .Y(n29324) );
  sky130_fd_sc_hd__a21oi_1 U14587 ( .A1(n11493), .A2(n19444), .B1(n11492), .Y(
        n11364) );
  sky130_fd_sc_hd__nand2_2 U14588 ( .A(n19663), .B(n19662), .Y(n27202) );
  sky130_fd_sc_hd__or2_0 U14589 ( .A(n27980), .B(n27796), .X(n12129) );
  sky130_fd_sc_hd__nand2_1 U14591 ( .A(n23703), .B(n23699), .Y(n23705) );
  sky130_fd_sc_hd__clkinv_1 U14592 ( .A(n25526), .Y(n25527) );
  sky130_fd_sc_hd__inv_2 U14593 ( .A(n23757), .Y(n11135) );
  sky130_fd_sc_hd__clkinv_1 U14594 ( .A(n12578), .Y(n21877) );
  sky130_fd_sc_hd__clkinv_1 U14595 ( .A(n27217), .Y(n23115) );
  sky130_fd_sc_hd__clkinv_1 U14596 ( .A(n21873), .Y(n19484) );
  sky130_fd_sc_hd__inv_1 U14597 ( .A(n23753), .Y(n26528) );
  sky130_fd_sc_hd__and2_0 U14599 ( .A(n21751), .B(n21776), .X(n12084) );
  sky130_fd_sc_hd__clkinv_1 U14600 ( .A(n27466), .Y(n23091) );
  sky130_fd_sc_hd__o21ai_2 U14601 ( .A1(n23532), .A2(n23531), .B1(n23530), .Y(
        n23533) );
  sky130_fd_sc_hd__clkinv_1 U14602 ( .A(n27209), .Y(n23073) );
  sky130_fd_sc_hd__clkinv_1 U14603 ( .A(n26948), .Y(n26070) );
  sky130_fd_sc_hd__o21ai_2 U14604 ( .A1(n23540), .A2(n23538), .B1(n23039), .Y(
        j202_soc_core_j22_cpu_rf_N2746) );
  sky130_fd_sc_hd__nor2_1 U14605 ( .A(n11980), .B(n11979), .Y(n21373) );
  sky130_fd_sc_hd__clkinv_1 U14606 ( .A(n11958), .Y(n11957) );
  sky130_fd_sc_hd__and2_1 U14607 ( .A(n20145), .B(n21750), .X(n12230) );
  sky130_fd_sc_hd__inv_1 U14608 ( .A(n27980), .Y(n12065) );
  sky130_fd_sc_hd__clkinv_1 U14609 ( .A(n27969), .Y(n27972) );
  sky130_fd_sc_hd__clkinv_1 U14610 ( .A(n12579), .Y(n21981) );
  sky130_fd_sc_hd__clkinv_1 U14611 ( .A(n27979), .Y(n27599) );
  sky130_fd_sc_hd__clkinv_1 U14612 ( .A(n27942), .Y(n24100) );
  sky130_fd_sc_hd__clkinv_1 U14613 ( .A(n27778), .Y(n27796) );
  sky130_fd_sc_hd__clkinv_1 U14614 ( .A(n27947), .Y(n24408) );
  sky130_fd_sc_hd__and2_0 U14615 ( .A(n11473), .B(n22396), .X(n22478) );
  sky130_fd_sc_hd__clkinv_1 U14616 ( .A(n25873), .Y(n25877) );
  sky130_fd_sc_hd__nor2_1 U14617 ( .A(n12107), .B(n12106), .Y(n12105) );
  sky130_fd_sc_hd__inv_2 U14618 ( .A(n26313), .Y(n29328) );
  sky130_fd_sc_hd__and2_1 U14619 ( .A(n28965), .B(
        j202_soc_core_ahbcs_6__HREADY_), .X(n29116) );
  sky130_fd_sc_hd__inv_2 U14621 ( .A(n22905), .Y(n21975) );
  sky130_fd_sc_hd__clkinv_1 U14622 ( .A(n27219), .Y(n23132) );
  sky130_fd_sc_hd__clkinv_1 U14623 ( .A(n12071), .Y(n28515) );
  sky130_fd_sc_hd__and2_0 U14624 ( .A(n20145), .B(n22715), .X(n12220) );
  sky130_fd_sc_hd__clkinv_1 U14625 ( .A(n22831), .Y(n21982) );
  sky130_fd_sc_hd__clkinv_1 U14627 ( .A(n25335), .Y(n26067) );
  sky130_fd_sc_hd__nor2_1 U14628 ( .A(n21785), .B(n21794), .Y(n18824) );
  sky130_fd_sc_hd__clkinv_1 U14629 ( .A(n26889), .Y(n26890) );
  sky130_fd_sc_hd__o21ai_1 U14630 ( .A1(n21420), .A2(n21418), .B1(n21419), .Y(
        n21791) );
  sky130_fd_sc_hd__nand2b_1 U14631 ( .A_N(n19199), .B(n21431), .Y(n12317) );
  sky130_fd_sc_hd__clkinv_1 U14632 ( .A(n27220), .Y(n26374) );
  sky130_fd_sc_hd__clkinv_1 U14633 ( .A(n21870), .Y(n21872) );
  sky130_fd_sc_hd__clkinv_1 U14634 ( .A(n27216), .Y(n25819) );
  sky130_fd_sc_hd__o21ai_2 U14635 ( .A1(n23541), .A2(n23538), .B1(n27212), .Y(
        j202_soc_core_j22_cpu_rf_N2820) );
  sky130_fd_sc_hd__and2_0 U14636 ( .A(n18902), .B(n18901), .X(n12481) );
  sky130_fd_sc_hd__o21ai_2 U14637 ( .A1(n23539), .A2(n23538), .B1(n27465), .Y(
        j202_soc_core_j22_cpu_rf_N2783) );
  sky130_fd_sc_hd__inv_1 U14638 ( .A(n18872), .Y(n18874) );
  sky130_fd_sc_hd__clkinv_1 U14639 ( .A(j202_soc_core_j22_cpu_rf_N2627), .Y(
        n26814) );
  sky130_fd_sc_hd__nor2_1 U14641 ( .A(n17125), .B(n12914), .Y(n11940) );
  sky130_fd_sc_hd__inv_1 U14642 ( .A(n27956), .Y(n27932) );
  sky130_fd_sc_hd__clkinv_1 U14643 ( .A(n27927), .Y(n27950) );
  sky130_fd_sc_hd__clkinv_1 U14644 ( .A(n28518), .Y(n28510) );
  sky130_fd_sc_hd__nand3_1 U14645 ( .A(n11312), .B(n11313), .C(n11311), .Y(
        n20718) );
  sky130_fd_sc_hd__clkinv_1 U14646 ( .A(n22751), .Y(n22752) );
  sky130_fd_sc_hd__clkinv_1 U14647 ( .A(n25539), .Y(n26908) );
  sky130_fd_sc_hd__clkinv_1 U14648 ( .A(n25756), .Y(n26911) );
  sky130_fd_sc_hd__clkinv_1 U14649 ( .A(n24594), .Y(n24595) );
  sky130_fd_sc_hd__clkinv_1 U14650 ( .A(n23484), .Y(n24471) );
  sky130_fd_sc_hd__clkinv_1 U14651 ( .A(n27218), .Y(n26369) );
  sky130_fd_sc_hd__nor2_1 U14652 ( .A(n11339), .B(n11338), .Y(n11337) );
  sky130_fd_sc_hd__nor2_1 U14653 ( .A(n21418), .B(n19159), .Y(n21788) );
  sky130_fd_sc_hd__clkinv_1 U14655 ( .A(n15659), .Y(n15662) );
  sky130_fd_sc_hd__clkinv_1 U14656 ( .A(n10565), .Y(n23692) );
  sky130_fd_sc_hd__o21ai_1 U14657 ( .A1(n21575), .A2(n18908), .B1(n18909), .Y(
        n22835) );
  sky130_fd_sc_hd__and2_0 U14659 ( .A(n20832), .B(n21776), .X(n13288) );
  sky130_fd_sc_hd__clkinv_1 U14660 ( .A(n18908), .Y(n18910) );
  sky130_fd_sc_hd__clkinv_1 U14661 ( .A(n27928), .Y(n11138) );
  sky130_fd_sc_hd__clkinv_1 U14662 ( .A(n21574), .Y(n21576) );
  sky130_fd_sc_hd__clkinv_1 U14663 ( .A(n25840), .Y(n25847) );
  sky130_fd_sc_hd__clkinv_1 U14664 ( .A(n11943), .Y(n11890) );
  sky130_fd_sc_hd__clkinv_1 U14665 ( .A(n19228), .Y(n19469) );
  sky130_fd_sc_hd__and2_0 U14666 ( .A(n16533), .B(n16553), .X(n16556) );
  sky130_fd_sc_hd__o21ai_2 U14667 ( .A1(n23540), .A2(n23537), .B1(n27227), .Y(
        j202_soc_core_j22_cpu_rf_N3190) );
  sky130_fd_sc_hd__clkinv_1 U14668 ( .A(n27334), .Y(n26803) );
  sky130_fd_sc_hd__o21ai_2 U14669 ( .A1(n23539), .A2(n23537), .B1(n27210), .Y(
        j202_soc_core_j22_cpu_rf_N3227) );
  sky130_fd_sc_hd__clkinv_1 U14670 ( .A(n21420), .Y(n21421) );
  sky130_fd_sc_hd__clkinv_1 U14671 ( .A(n25451), .Y(n26907) );
  sky130_fd_sc_hd__clkinv_1 U14672 ( .A(n19221), .Y(n21441) );
  sky130_fd_sc_hd__clkinv_1 U14673 ( .A(n19227), .Y(n19467) );
  sky130_fd_sc_hd__clkinv_1 U14674 ( .A(n26813), .Y(n26798) );
  sky130_fd_sc_hd__o21a_1 U14675 ( .A1(n15663), .A2(n15660), .B1(n15664), .X(
        n15416) );
  sky130_fd_sc_hd__clkinv_1 U14676 ( .A(n25235), .Y(n25236) );
  sky130_fd_sc_hd__nor2_1 U14677 ( .A(n11408), .B(n11407), .Y(n11406) );
  sky130_fd_sc_hd__a2bb2oi_1 U14678 ( .B1(n19786), .B2(n19788), .A1_N(n19757), 
        .A2_N(n19768), .Y(n19758) );
  sky130_fd_sc_hd__nor2_1 U14679 ( .A(n22397), .B(n22389), .Y(n22470) );
  sky130_fd_sc_hd__nand2_1 U14680 ( .A(n11413), .B(n11415), .Y(n11412) );
  sky130_fd_sc_hd__clkinv_1 U14681 ( .A(n26000), .Y(n26124) );
  sky130_fd_sc_hd__and2_0 U14682 ( .A(n14978), .B(n21776), .X(n12283) );
  sky130_fd_sc_hd__clkinv_1 U14683 ( .A(n23490), .Y(n24468) );
  sky130_fd_sc_hd__nand2_1 U14684 ( .A(n23508), .B(n23555), .Y(n23558) );
  sky130_fd_sc_hd__clkinv_1 U14685 ( .A(n19159), .Y(n21422) );
  sky130_fd_sc_hd__a21oi_1 U14686 ( .A1(n18846), .A2(n19228), .B1(n18845), .Y(
        n18847) );
  sky130_fd_sc_hd__nor2_1 U14688 ( .A(n12045), .B(n18812), .Y(n21909) );
  sky130_fd_sc_hd__nand3_2 U14689 ( .A(n23177), .B(n23111), .C(n23110), .Y(
        n27216) );
  sky130_fd_sc_hd__inv_2 U14690 ( .A(n23177), .Y(n23169) );
  sky130_fd_sc_hd__and2_1 U14691 ( .A(n18981), .B(n22581), .X(n11726) );
  sky130_fd_sc_hd__clkinv_1 U14692 ( .A(n19222), .Y(n21440) );
  sky130_fd_sc_hd__nand3_2 U14693 ( .A(n23177), .B(n23096), .C(n23095), .Y(
        n27220) );
  sky130_fd_sc_hd__and2_0 U14695 ( .A(n12072), .B(j202_soc_core_j22_cpu_intack), .X(n12071) );
  sky130_fd_sc_hd__nand2_2 U14696 ( .A(n21584), .B(n13603), .Y(n22596) );
  sky130_fd_sc_hd__o21ai_2 U14697 ( .A1(n23528), .A2(n24113), .B1(n27124), .Y(
        j202_soc_core_j22_cpu_rf_N2709) );
  sky130_fd_sc_hd__nand2_2 U14698 ( .A(n22592), .B(n22590), .Y(n22515) );
  sky130_fd_sc_hd__and2_0 U14699 ( .A(n20954), .B(n20953), .X(n12191) );
  sky130_fd_sc_hd__nor2_1 U14700 ( .A(n18908), .B(n21574), .Y(n22831) );
  sky130_fd_sc_hd__nand3_2 U14701 ( .A(n23177), .B(n23128), .C(n23127), .Y(
        n27218) );
  sky130_fd_sc_hd__clkinv_1 U14702 ( .A(n24645), .Y(n24646) );
  sky130_fd_sc_hd__clkinv_1 U14703 ( .A(n21805), .Y(n19445) );
  sky130_fd_sc_hd__inv_2 U14704 ( .A(n21794), .Y(n11140) );
  sky130_fd_sc_hd__o21ai_2 U14705 ( .A1(n23543), .A2(n23540), .B1(n27222), .Y(
        j202_soc_core_j22_cpu_rf_N3042) );
  sky130_fd_sc_hd__inv_2 U14706 ( .A(n17125), .Y(n22581) );
  sky130_fd_sc_hd__clkinv_1 U14707 ( .A(n26754), .Y(n26761) );
  sky130_fd_sc_hd__clkinv_1 U14708 ( .A(n26763), .Y(n26766) );
  sky130_fd_sc_hd__nor2_1 U14709 ( .A(n22902), .B(n22908), .Y(n19227) );
  sky130_fd_sc_hd__clkinv_1 U14710 ( .A(n26753), .Y(n26762) );
  sky130_fd_sc_hd__clkinv_1 U14711 ( .A(n22908), .Y(n21973) );
  sky130_fd_sc_hd__clkinv_1 U14712 ( .A(n27921), .Y(n27930) );
  sky130_fd_sc_hd__and2_0 U14713 ( .A(n20042), .B(n20043), .X(n12287) );
  sky130_fd_sc_hd__o21ai_1 U14714 ( .A1(n14132), .A2(n19415), .B1(n14131), .Y(
        n18998) );
  sky130_fd_sc_hd__inv_2 U14715 ( .A(n17109), .Y(n16989) );
  sky130_fd_sc_hd__nand2_1 U14716 ( .A(n18270), .B(n18269), .Y(n21575) );
  sky130_fd_sc_hd__clkinv_1 U14718 ( .A(n22590), .Y(n17120) );
  sky130_fd_sc_hd__nor2_1 U14719 ( .A(n18818), .B(n18817), .Y(n19159) );
  sky130_fd_sc_hd__inv_1 U14720 ( .A(n21480), .Y(n21481) );
  sky130_fd_sc_hd__clkinv_1 U14721 ( .A(n21980), .Y(n22834) );
  sky130_fd_sc_hd__clkinv_1 U14722 ( .A(n21479), .Y(n21482) );
  sky130_fd_sc_hd__nand4_1 U14723 ( .A(n13042), .B(n13041), .C(n13040), .D(
        n13153), .Y(n11301) );
  sky130_fd_sc_hd__clkinv_1 U14724 ( .A(n19802), .Y(n19803) );
  sky130_fd_sc_hd__clkinv_1 U14725 ( .A(n19809), .Y(n19810) );
  sky130_fd_sc_hd__clkinv_1 U14726 ( .A(n19817), .Y(n19818) );
  sky130_fd_sc_hd__clkinv_1 U14727 ( .A(n19789), .Y(n19791) );
  sky130_fd_sc_hd__clkinv_1 U14728 ( .A(n19555), .Y(n19566) );
  sky130_fd_sc_hd__a21oi_1 U14729 ( .A1(n13280), .A2(n21460), .B1(n11496), .Y(
        n17868) );
  sky130_fd_sc_hd__o21a_1 U14730 ( .A1(n19769), .A2(n13028), .B1(n19770), .X(
        n13027) );
  sky130_fd_sc_hd__clkinv_1 U14731 ( .A(n22902), .Y(n22904) );
  sky130_fd_sc_hd__clkinv_1 U14732 ( .A(n22182), .Y(n22186) );
  sky130_fd_sc_hd__clkinv_1 U14733 ( .A(n19651), .Y(n19665) );
  sky130_fd_sc_hd__and2_0 U14734 ( .A(n20709), .B(n21776), .X(n12289) );
  sky130_fd_sc_hd__clkinv_1 U14735 ( .A(n11420), .Y(n11417) );
  sky130_fd_sc_hd__clkinv_1 U14736 ( .A(n26764), .Y(n26765) );
  sky130_fd_sc_hd__nand3_1 U14737 ( .A(n13603), .B(
        j202_soc_core_j22_cpu_memop_Ma__0_), .C(
        j202_soc_core_j22_cpu_memop_Ma__1_), .Y(n17125) );
  sky130_fd_sc_hd__clkinv_1 U14738 ( .A(n26610), .Y(n11961) );
  sky130_fd_sc_hd__clkinv_1 U14739 ( .A(n16538), .Y(n16148) );
  sky130_fd_sc_hd__clkinv_1 U14740 ( .A(n16532), .Y(n16149) );
  sky130_fd_sc_hd__clkinv_1 U14741 ( .A(n17242), .Y(n17257) );
  sky130_fd_sc_hd__nor2_1 U14742 ( .A(n19470), .B(n18844), .Y(n18846) );
  sky130_fd_sc_hd__clkinv_1 U14743 ( .A(n22325), .Y(n22326) );
  sky130_fd_sc_hd__clkinv_1 U14744 ( .A(n21869), .Y(n11449) );
  sky130_fd_sc_hd__o21ai_1 U14745 ( .A1(n22093), .A2(n22182), .B1(n22092), .Y(
        n22130) );
  sky130_fd_sc_hd__clkinv_1 U14746 ( .A(n21808), .Y(n21810) );
  sky130_fd_sc_hd__nor2_1 U14747 ( .A(n22093), .B(n22180), .Y(n22131) );
  sky130_fd_sc_hd__and3_1 U14748 ( .A(n19143), .B(n19156), .C(n19154), .X(
        n19144) );
  sky130_fd_sc_hd__clkinv_1 U14749 ( .A(n21478), .Y(n22327) );
  sky130_fd_sc_hd__and3_1 U14750 ( .A(n20137), .B(n20130), .C(n20141), .X(
        n20131) );
  sky130_fd_sc_hd__clkinv_1 U14751 ( .A(n19769), .Y(n19771) );
  sky130_fd_sc_hd__clkinv_1 U14752 ( .A(n20410), .Y(n20420) );
  sky130_fd_sc_hd__clkinv_1 U14753 ( .A(n19775), .Y(n19777) );
  sky130_fd_sc_hd__clkinv_1 U14754 ( .A(n21324), .Y(n21329) );
  sky130_fd_sc_hd__clkinv_1 U14755 ( .A(n21327), .Y(n21328) );
  sky130_fd_sc_hd__clkinv_1 U14756 ( .A(n16138), .Y(n16139) );
  sky130_fd_sc_hd__clkinv_1 U14757 ( .A(n17262), .Y(n20279) );
  sky130_fd_sc_hd__clkinv_1 U14758 ( .A(n22161), .Y(n22162) );
  sky130_fd_sc_hd__nand2_1 U14759 ( .A(n18086), .B(n18085), .Y(n18093) );
  sky130_fd_sc_hd__clkinv_1 U14760 ( .A(n21894), .Y(n19464) );
  sky130_fd_sc_hd__inv_1 U14761 ( .A(n21526), .Y(n21528) );
  sky130_fd_sc_hd__clkinv_1 U14762 ( .A(n22160), .Y(n22163) );
  sky130_fd_sc_hd__clkinv_1 U14763 ( .A(n19322), .Y(n19323) );
  sky130_fd_sc_hd__clkinv_1 U14764 ( .A(n15899), .Y(n15304) );
  sky130_fd_sc_hd__clkinv_1 U14765 ( .A(n21013), .Y(n15508) );
  sky130_fd_sc_hd__clkinv_1 U14766 ( .A(n21504), .Y(n18887) );
  sky130_fd_sc_hd__and3_1 U14767 ( .A(n17350), .B(n17337), .C(n17349), .X(
        n17338) );
  sky130_fd_sc_hd__and2_0 U14768 ( .A(n17096), .B(n17097), .X(n11676) );
  sky130_fd_sc_hd__clkinv_1 U14769 ( .A(n22329), .Y(n22331) );
  sky130_fd_sc_hd__o21ai_1 U14770 ( .A1(n14063), .A2(n21919), .B1(n21920), .Y(
        n17262) );
  sky130_fd_sc_hd__clkinv_1 U14771 ( .A(n19319), .Y(n19320) );
  sky130_fd_sc_hd__clkinv_1 U14773 ( .A(n21330), .Y(n21346) );
  sky130_fd_sc_hd__clkinv_1 U14774 ( .A(n16531), .Y(n16152) );
  sky130_fd_sc_hd__clkinv_1 U14775 ( .A(n21345), .Y(n21331) );
  sky130_fd_sc_hd__clkinv_1 U14776 ( .A(n16536), .Y(n15956) );
  sky130_fd_sc_hd__inv_1 U14777 ( .A(n16535), .Y(n16024) );
  sky130_fd_sc_hd__clkinv_1 U14778 ( .A(n21332), .Y(n21334) );
  sky130_fd_sc_hd__clkinv_1 U14779 ( .A(n22587), .Y(n18999) );
  sky130_fd_sc_hd__inv_1 U14780 ( .A(n19418), .Y(n19420) );
  sky130_fd_sc_hd__inv_1 U14781 ( .A(n20286), .Y(n19417) );
  sky130_fd_sc_hd__clkinv_1 U14782 ( .A(n21357), .Y(n21371) );
  sky130_fd_sc_hd__clkinv_1 U14783 ( .A(n22763), .Y(n21962) );
  sky130_fd_sc_hd__clkinv_1 U14784 ( .A(n20275), .Y(n20277) );
  sky130_fd_sc_hd__inv_1 U14785 ( .A(n19416), .Y(n20287) );
  sky130_fd_sc_hd__clkinv_1 U14787 ( .A(n21359), .Y(n21361) );
  sky130_fd_sc_hd__clkinv_1 U14788 ( .A(n19466), .Y(n18841) );
  sky130_fd_sc_hd__clkinv_1 U14789 ( .A(n21370), .Y(n21358) );
  sky130_fd_sc_hd__clkinv_1 U14790 ( .A(n16818), .Y(n16820) );
  sky130_fd_sc_hd__o2bb2ai_1 U14791 ( .B1(n26713), .B2(n26424), .A1_N(n26077), 
        .A2_N(n26722), .Y(n19185) );
  sky130_fd_sc_hd__mux2_2 U14792 ( .A0(n19642), .A1(n19643), .S(n26840), .X(
        n19769) );
  sky130_fd_sc_hd__clkinv_1 U14793 ( .A(n15512), .Y(n15514) );
  sky130_fd_sc_hd__inv_1 U14794 ( .A(n22511), .Y(n20998) );
  sky130_fd_sc_hd__inv_1 U14795 ( .A(n20999), .Y(n21001) );
  sky130_fd_sc_hd__clkinv_1 U14796 ( .A(n20997), .Y(n22512) );
  sky130_fd_sc_hd__inv_1 U14798 ( .A(n26418), .Y(n25131) );
  sky130_fd_sc_hd__inv_1 U14799 ( .A(n16994), .Y(n16996) );
  sky130_fd_sc_hd__clkinv_1 U14800 ( .A(n15194), .Y(n14843) );
  sky130_fd_sc_hd__and2_0 U14801 ( .A(n26872), .B(n24805), .X(n11462) );
  sky130_fd_sc_hd__a2bb2oi_1 U14802 ( .B1(n26718), .B2(n26077), .A1_N(n25403), 
        .A2_N(n26424), .Y(n24787) );
  sky130_fd_sc_hd__clkinv_1 U14803 ( .A(n19470), .Y(n19226) );
  sky130_fd_sc_hd__clkinv_1 U14804 ( .A(n15663), .Y(n15665) );
  sky130_fd_sc_hd__nand3_1 U14805 ( .A(n19696), .B(n19695), .C(n19694), .Y(
        n26825) );
  sky130_fd_sc_hd__clkinv_1 U14806 ( .A(n26588), .Y(n26667) );
  sky130_fd_sc_hd__clkinv_1 U14807 ( .A(n21867), .Y(n18854) );
  sky130_fd_sc_hd__inv_1 U14808 ( .A(n15952), .Y(n15210) );
  sky130_fd_sc_hd__clkinv_1 U14809 ( .A(n15772), .Y(n15774) );
  sky130_fd_sc_hd__a2bb2oi_1 U14810 ( .B1(n26061), .B2(n26077), .A1_N(n26581), 
        .A2_N(n26424), .Y(n24141) );
  sky130_fd_sc_hd__inv_1 U14811 ( .A(n21919), .Y(n21921) );
  sky130_fd_sc_hd__nor2_1 U14812 ( .A(n21359), .B(n21357), .Y(n21324) );
  sky130_fd_sc_hd__clkinv_1 U14813 ( .A(n26349), .Y(n24665) );
  sky130_fd_sc_hd__inv_2 U14814 ( .A(n17867), .Y(n11498) );
  sky130_fd_sc_hd__clkinv_1 U14815 ( .A(n16657), .Y(n16659) );
  sky130_fd_sc_hd__clkinv_1 U14816 ( .A(n17114), .Y(n16652) );
  sky130_fd_sc_hd__clkinv_1 U14817 ( .A(n16982), .Y(n16983) );
  sky130_fd_sc_hd__clkinv_1 U14818 ( .A(n15418), .Y(n15420) );
  sky130_fd_sc_hd__clkinv_1 U14819 ( .A(n16979), .Y(n16980) );
  sky130_fd_sc_hd__clkinv_1 U14820 ( .A(n16643), .Y(n16644) );
  sky130_fd_sc_hd__nor2_1 U14821 ( .A(n14830), .B(n14831), .Y(n21014) );
  sky130_fd_sc_hd__nand2_1 U14822 ( .A(n19598), .B(n19597), .Y(n26840) );
  sky130_fd_sc_hd__clkinv_1 U14823 ( .A(n22238), .Y(n22239) );
  sky130_fd_sc_hd__clkinv_1 U14824 ( .A(n22222), .Y(n22223) );
  sky130_fd_sc_hd__nor2_1 U14825 ( .A(n14560), .B(n14561), .Y(n21359) );
  sky130_fd_sc_hd__nor2_1 U14826 ( .A(n14558), .B(n14559), .Y(n21357) );
  sky130_fd_sc_hd__clkinv_1 U14827 ( .A(n22774), .Y(n22775) );
  sky130_fd_sc_hd__xor2_1 U14828 ( .A(n18399), .B(n11742), .X(n18606) );
  sky130_fd_sc_hd__clkinv_1 U14829 ( .A(n25769), .Y(n26836) );
  sky130_fd_sc_hd__clkinv_1 U14830 ( .A(n22303), .Y(n22304) );
  sky130_fd_sc_hd__clkinv_1 U14831 ( .A(n19786), .Y(n19787) );
  sky130_fd_sc_hd__o21ai_1 U14832 ( .A1(n19756), .A2(n19693), .B1(n19754), .Y(
        n19696) );
  sky130_fd_sc_hd__clkinv_1 U14833 ( .A(n18840), .Y(n11430) );
  sky130_fd_sc_hd__nor2_1 U14834 ( .A(n18838), .B(n18837), .Y(n19473) );
  sky130_fd_sc_hd__clkinv_1 U14835 ( .A(n18839), .Y(n11431) );
  sky130_fd_sc_hd__clkinv_1 U14836 ( .A(n22010), .Y(n21396) );
  sky130_fd_sc_hd__clkinv_1 U14837 ( .A(n21489), .Y(n18853) );
  sky130_fd_sc_hd__clkinv_1 U14838 ( .A(n22263), .Y(n22264) );
  sky130_fd_sc_hd__clkinv_1 U14839 ( .A(n19772), .Y(n19773) );
  sky130_fd_sc_hd__nand2b_1 U14840 ( .A_N(n18851), .B(n11503), .Y(n21490) );
  sky130_fd_sc_hd__nor2_1 U14841 ( .A(n14828), .B(n14829), .Y(n20999) );
  sky130_fd_sc_hd__clkinv_1 U14842 ( .A(n19778), .Y(n19779) );
  sky130_fd_sc_hd__clkinv_1 U14843 ( .A(n21923), .Y(n14063) );
  sky130_fd_sc_hd__clkinv_1 U14844 ( .A(n27306), .Y(n27307) );
  sky130_fd_sc_hd__clkinv_1 U14845 ( .A(n28594), .Y(n28595) );
  sky130_fd_sc_hd__clkinv_1 U14846 ( .A(n23016), .Y(n19028) );
  sky130_fd_sc_hd__clkinv_1 U14847 ( .A(n26615), .Y(n24033) );
  sky130_fd_sc_hd__clkinv_1 U14848 ( .A(n25584), .Y(n25589) );
  sky130_fd_sc_hd__clkinv_1 U14849 ( .A(n23919), .Y(n19023) );
  sky130_fd_sc_hd__clkinv_1 U14850 ( .A(n18084), .Y(n11581) );
  sky130_fd_sc_hd__clkinv_1 U14851 ( .A(n21515), .Y(n17841) );
  sky130_fd_sc_hd__clkinv_1 U14852 ( .A(n27399), .Y(n25165) );
  sky130_fd_sc_hd__clkinv_1 U14853 ( .A(n26700), .Y(n26743) );
  sky130_fd_sc_hd__clkinv_1 U14854 ( .A(n22183), .Y(n22184) );
  sky130_fd_sc_hd__inv_1 U14855 ( .A(n18256), .Y(n12440) );
  sky130_fd_sc_hd__clkinv_1 U14856 ( .A(n22069), .Y(n22185) );
  sky130_fd_sc_hd__clkinv_1 U14857 ( .A(n19026), .Y(n19027) );
  sky130_fd_sc_hd__inv_2 U14858 ( .A(n18602), .Y(n12762) );
  sky130_fd_sc_hd__and2_0 U14859 ( .A(n22477), .B(n11478), .X(n11476) );
  sky130_fd_sc_hd__a21oi_1 U14860 ( .A1(n11475), .A2(n22477), .B1(n22476), .Y(
        n11474) );
  sky130_fd_sc_hd__clkinv_1 U14861 ( .A(n16923), .Y(n16790) );
  sky130_fd_sc_hd__nand2_1 U14862 ( .A(n19638), .B(n19637), .Y(n25769) );
  sky130_fd_sc_hd__clkinv_1 U14863 ( .A(n19393), .Y(n17325) );
  sky130_fd_sc_hd__clkinv_1 U14865 ( .A(n21821), .Y(n21823) );
  sky130_fd_sc_hd__clkinv_1 U14866 ( .A(n22519), .Y(n22082) );
  sky130_fd_sc_hd__clkinv_1 U14867 ( .A(n26887), .Y(n24998) );
  sky130_fd_sc_hd__clkinv_1 U14868 ( .A(n26634), .Y(n19018) );
  sky130_fd_sc_hd__inv_1 U14870 ( .A(n26827), .Y(n26828) );
  sky130_fd_sc_hd__and2_0 U14871 ( .A(n27308), .B(n29594), .X(n27857) );
  sky130_fd_sc_hd__clkinv_1 U14872 ( .A(n27405), .Y(n26082) );
  sky130_fd_sc_hd__clkinv_1 U14873 ( .A(n27443), .Y(n24612) );
  sky130_fd_sc_hd__inv_1 U14874 ( .A(n18255), .Y(n12441) );
  sky130_fd_sc_hd__clkinv_1 U14875 ( .A(n22469), .Y(n22429) );
  sky130_fd_sc_hd__clkinv_1 U14876 ( .A(n22475), .Y(n22428) );
  sky130_fd_sc_hd__clkinv_1 U14877 ( .A(n27365), .Y(n26582) );
  sky130_fd_sc_hd__clkinv_1 U14878 ( .A(n27412), .Y(n26569) );
  sky130_fd_sc_hd__clkinv_1 U14879 ( .A(n27383), .Y(n25057) );
  sky130_fd_sc_hd__xnor2_1 U14880 ( .A(n11743), .B(n18400), .Y(n11742) );
  sky130_fd_sc_hd__clkinv_1 U14881 ( .A(n27347), .Y(n26885) );
  sky130_fd_sc_hd__clkinv_1 U14882 ( .A(n27357), .Y(n26579) );
  sky130_fd_sc_hd__clkinv_1 U14883 ( .A(n27389), .Y(n25121) );
  sky130_fd_sc_hd__clkinv_1 U14884 ( .A(n27419), .Y(n24518) );
  sky130_fd_sc_hd__clkinv_1 U14885 ( .A(n27447), .Y(n26580) );
  sky130_fd_sc_hd__clkinv_1 U14886 ( .A(n27425), .Y(n24072) );
  sky130_fd_sc_hd__clkinv_1 U14887 ( .A(n25024), .Y(n25025) );
  sky130_fd_sc_hd__clkinv_1 U14888 ( .A(n24613), .Y(n27439) );
  sky130_fd_sc_hd__clkinv_1 U14889 ( .A(n24671), .Y(n27375) );
  sky130_fd_sc_hd__clkinv_1 U14890 ( .A(n22794), .Y(n22796) );
  sky130_fd_sc_hd__clkinv_1 U14891 ( .A(n24052), .Y(n24038) );
  sky130_fd_sc_hd__nor2_1 U14893 ( .A(n22075), .B(n22076), .Y(n22187) );
  sky130_fd_sc_hd__nor2_1 U14895 ( .A(n17860), .B(n17861), .Y(n22843) );
  sky130_fd_sc_hd__clkinv_1 U14896 ( .A(n27392), .Y(n23834) );
  sky130_fd_sc_hd__clkinv_1 U14897 ( .A(n25122), .Y(n27386) );
  sky130_fd_sc_hd__clkinv_1 U14898 ( .A(n26720), .Y(n26336) );
  sky130_fd_sc_hd__clkinv_1 U14899 ( .A(n27354), .Y(n26566) );
  sky130_fd_sc_hd__clkinv_1 U14900 ( .A(n23547), .Y(n23548) );
  sky130_fd_sc_hd__clkinv_1 U14901 ( .A(n27361), .Y(n26564) );
  sky130_fd_sc_hd__nand2_1 U14902 ( .A(n19734), .B(n19733), .Y(n26827) );
  sky130_fd_sc_hd__clkinv_1 U14903 ( .A(n21259), .Y(n21106) );
  sky130_fd_sc_hd__clkinv_1 U14904 ( .A(n26916), .Y(n26917) );
  sky130_fd_sc_hd__clkinv_1 U14906 ( .A(n26919), .Y(n25575) );
  sky130_fd_sc_hd__clkinv_1 U14907 ( .A(n11715), .Y(n11714) );
  sky130_fd_sc_hd__clkinv_1 U14908 ( .A(n27455), .Y(n23982) );
  sky130_fd_sc_hd__nand2_1 U14909 ( .A(n22268), .B(n22824), .Y(n12296) );
  sky130_fd_sc_hd__clkinv_1 U14911 ( .A(n27474), .Y(n27481) );
  sky130_fd_sc_hd__clkinv_1 U14912 ( .A(n27377), .Y(n24667) );
  sky130_fd_sc_hd__clkinv_1 U14913 ( .A(n27372), .Y(n26413) );
  sky130_fd_sc_hd__clkinv_1 U14914 ( .A(n25586), .Y(n25587) );
  sky130_fd_sc_hd__clkinv_1 U14915 ( .A(n19311), .Y(n19312) );
  sky130_fd_sc_hd__clkinv_1 U14916 ( .A(n27396), .Y(n23832) );
  sky130_fd_sc_hd__clkinv_1 U14917 ( .A(n25560), .Y(n25561) );
  sky130_fd_sc_hd__a21oi_1 U14919 ( .A1(n22357), .A2(n22099), .B1(n22098), .Y(
        n22100) );
  sky130_fd_sc_hd__clkinv_1 U14920 ( .A(n22396), .Y(n11475) );
  sky130_fd_sc_hd__clkinv_1 U14921 ( .A(n27432), .Y(n26572) );
  sky130_fd_sc_hd__clkinv_1 U14922 ( .A(n22157), .Y(n22159) );
  sky130_fd_sc_hd__clkinv_1 U14924 ( .A(n25094), .Y(n25095) );
  sky130_fd_sc_hd__clkinv_1 U14925 ( .A(n27380), .Y(n25061) );
  sky130_fd_sc_hd__clkinv_1 U14926 ( .A(n25230), .Y(n19198) );
  sky130_fd_sc_hd__clkinv_1 U14927 ( .A(n20083), .Y(n20055) );
  sky130_fd_sc_hd__clkinv_1 U14928 ( .A(n20195), .Y(n19106) );
  sky130_fd_sc_hd__clkinv_1 U14929 ( .A(n27469), .Y(n26290) );
  sky130_fd_sc_hd__nand3_1 U14930 ( .A(n11916), .B(n16014), .C(n11915), .Y(
        n13551) );
  sky130_fd_sc_hd__a31o_1 U14931 ( .A1(n20006), .A2(n12165), .A3(n20374), .B1(
        n20927), .X(n17199) );
  sky130_fd_sc_hd__clkinv_1 U14932 ( .A(n27269), .Y(n24115) );
  sky130_fd_sc_hd__clkinv_1 U14933 ( .A(n22361), .Y(n22129) );
  sky130_fd_sc_hd__clkinv_1 U14934 ( .A(n22359), .Y(n22099) );
  sky130_fd_sc_hd__inv_2 U14935 ( .A(n17902), .Y(n12752) );
  sky130_fd_sc_hd__clkinv_1 U14936 ( .A(n19883), .Y(n19884) );
  sky130_fd_sc_hd__clkinv_1 U14937 ( .A(n23531), .Y(n23444) );
  sky130_fd_sc_hd__nand3_2 U14938 ( .A(n13786), .B(n13785), .C(n13784), .Y(
        n23920) );
  sky130_fd_sc_hd__a21o_1 U14939 ( .A1(n20639), .A2(n20529), .B1(n20651), .X(
        n20530) );
  sky130_fd_sc_hd__nand3_1 U14940 ( .A(n12211), .B(n13296), .C(n14769), .Y(
        n26724) );
  sky130_fd_sc_hd__clkinv_1 U14941 ( .A(n21278), .Y(n21619) );
  sky130_fd_sc_hd__nand3_2 U14942 ( .A(n14592), .B(n12188), .C(n14591), .Y(
        n26719) );
  sky130_fd_sc_hd__nand3_2 U14943 ( .A(n13648), .B(n12190), .C(n13647), .Y(
        n26717) );
  sky130_fd_sc_hd__clkinv_1 U14944 ( .A(n20243), .Y(n20244) );
  sky130_fd_sc_hd__clkinv_1 U14945 ( .A(n26205), .Y(n23914) );
  sky130_fd_sc_hd__clkinv_1 U14946 ( .A(n19843), .Y(n19992) );
  sky130_fd_sc_hd__clkinv_1 U14947 ( .A(n26791), .Y(n27422) );
  sky130_fd_sc_hd__nand3_2 U14948 ( .A(n13975), .B(n12189), .C(n13974), .Y(
        n27415) );
  sky130_fd_sc_hd__nand3_1 U14949 ( .A(n13845), .B(n12201), .C(n13844), .Y(
        n26712) );
  sky130_fd_sc_hd__clkinv_1 U14950 ( .A(n29347), .Y(n27722) );
  sky130_fd_sc_hd__clkinv_1 U14951 ( .A(n25290), .Y(n23041) );
  sky130_fd_sc_hd__inv_2 U14952 ( .A(n26600), .Y(n11145) );
  sky130_fd_sc_hd__clkinv_1 U14953 ( .A(n21217), .Y(n21067) );
  sky130_fd_sc_hd__nand3_1 U14954 ( .A(n14485), .B(n14484), .C(n14483), .Y(
        n26721) );
  sky130_fd_sc_hd__nor2_1 U14955 ( .A(n11674), .B(n11672), .Y(n11671) );
  sky130_fd_sc_hd__clkinv_1 U14956 ( .A(n27488), .Y(n26304) );
  sky130_fd_sc_hd__nand3_1 U14957 ( .A(n11679), .B(n17013), .C(n14915), .Y(
        n14871) );
  sky130_fd_sc_hd__clkinv_1 U14958 ( .A(n18166), .Y(n18168) );
  sky130_fd_sc_hd__clkinv_1 U14959 ( .A(n16738), .Y(n16736) );
  sky130_fd_sc_hd__clkinv_1 U14960 ( .A(n10562), .Y(n27601) );
  sky130_fd_sc_hd__clkinv_1 U14961 ( .A(n24133), .Y(n21427) );
  sky130_fd_sc_hd__clkinv_1 U14962 ( .A(n27640), .Y(n27641) );
  sky130_fd_sc_hd__clkinv_1 U14963 ( .A(n20852), .Y(n20061) );
  sky130_fd_sc_hd__clkinv_1 U14964 ( .A(n21713), .Y(n20755) );
  sky130_fd_sc_hd__clkinv_1 U14965 ( .A(n20239), .Y(n20223) );
  sky130_fd_sc_hd__clkinv_1 U14966 ( .A(n19278), .Y(n19280) );
  sky130_fd_sc_hd__clkinv_1 U14967 ( .A(n22094), .Y(n22089) );
  sky130_fd_sc_hd__clkinv_1 U14968 ( .A(n20865), .Y(n20891) );
  sky130_fd_sc_hd__clkinv_1 U14969 ( .A(n21133), .Y(n21138) );
  sky130_fd_sc_hd__clkinv_1 U14970 ( .A(n21626), .Y(n11995) );
  sky130_fd_sc_hd__clkinv_1 U14971 ( .A(n15374), .Y(n15619) );
  sky130_fd_sc_hd__clkinv_1 U14972 ( .A(n16681), .Y(n16683) );
  sky130_fd_sc_hd__clkinv_1 U14973 ( .A(n18484), .Y(n12776) );
  sky130_fd_sc_hd__clkinv_1 U14974 ( .A(n16189), .Y(n16190) );
  sky130_fd_sc_hd__clkinv_1 U14975 ( .A(n20366), .Y(n20330) );
  sky130_fd_sc_hd__clkinv_1 U14976 ( .A(n23857), .Y(n23614) );
  sky130_fd_sc_hd__and2_0 U14977 ( .A(n21927), .B(n21926), .X(n24602) );
  sky130_fd_sc_hd__clkinv_1 U14978 ( .A(n26288), .Y(n26281) );
  sky130_fd_sc_hd__clkinv_1 U14979 ( .A(n26183), .Y(n23320) );
  sky130_fd_sc_hd__clkinv_1 U14980 ( .A(n20229), .Y(n20014) );
  sky130_fd_sc_hd__clkinv_1 U14981 ( .A(n15856), .Y(n11679) );
  sky130_fd_sc_hd__clkinv_1 U14982 ( .A(n20550), .Y(n20555) );
  sky130_fd_sc_hd__clkinv_1 U14983 ( .A(n26446), .Y(n16649) );
  sky130_fd_sc_hd__clkinv_1 U14984 ( .A(n27985), .Y(n24252) );
  sky130_fd_sc_hd__clkinv_1 U14985 ( .A(n20365), .Y(n19105) );
  sky130_fd_sc_hd__clkinv_1 U14986 ( .A(n19307), .Y(n19317) );
  sky130_fd_sc_hd__clkinv_1 U14987 ( .A(n21654), .Y(n19360) );
  sky130_fd_sc_hd__clkinv_1 U14988 ( .A(n26069), .Y(n26071) );
  sky130_fd_sc_hd__clkinv_1 U14989 ( .A(n25578), .Y(n25579) );
  sky130_fd_sc_hd__a21o_1 U14990 ( .A1(n13591), .A2(n13592), .B1(n11538), .X(
        n11536) );
  sky130_fd_sc_hd__clkinv_1 U14991 ( .A(n16908), .Y(n16909) );
  sky130_fd_sc_hd__clkinv_1 U14992 ( .A(n16560), .Y(n16561) );
  sky130_fd_sc_hd__clkinv_1 U14993 ( .A(n20650), .Y(n20654) );
  sky130_fd_sc_hd__clkinv_1 U14994 ( .A(n19900), .Y(n20018) );
  sky130_fd_sc_hd__clkinv_1 U14995 ( .A(n21187), .Y(n19301) );
  sky130_fd_sc_hd__clkinv_1 U14996 ( .A(n16750), .Y(n16757) );
  sky130_fd_sc_hd__clkinv_1 U14997 ( .A(n26283), .Y(n25583) );
  sky130_fd_sc_hd__or2_0 U14998 ( .A(n19175), .B(n19174), .X(n19177) );
  sky130_fd_sc_hd__clkinv_1 U14999 ( .A(n24173), .Y(n23454) );
  sky130_fd_sc_hd__clkinv_1 U15000 ( .A(n15732), .Y(n15734) );
  sky130_fd_sc_hd__clkinv_1 U15001 ( .A(n20500), .Y(n20642) );
  sky130_fd_sc_hd__clkinv_1 U15002 ( .A(n20810), .Y(n21679) );
  sky130_fd_sc_hd__clkinv_1 U15003 ( .A(n19600), .Y(n19591) );
  sky130_fd_sc_hd__clkinv_1 U15004 ( .A(n15568), .Y(n15314) );
  sky130_fd_sc_hd__clkinv_1 U15005 ( .A(n20675), .Y(n20608) );
  sky130_fd_sc_hd__clkinv_1 U15006 ( .A(n13437), .Y(n13416) );
  sky130_fd_sc_hd__clkinv_1 U15007 ( .A(n20461), .Y(n20464) );
  sky130_fd_sc_hd__clkinv_1 U15008 ( .A(n13412), .Y(n13414) );
  sky130_fd_sc_hd__nor4b_1 U15009 ( .D_N(n14961), .A(n16095), .B(n17076), .C(
        n15865), .Y(n16105) );
  sky130_fd_sc_hd__clkinv_1 U15010 ( .A(n18880), .Y(n18881) );
  sky130_fd_sc_hd__clkinv_1 U15011 ( .A(n19652), .Y(n19654) );
  sky130_fd_sc_hd__or2_0 U15012 ( .A(n21925), .B(n21924), .X(n21927) );
  sky130_fd_sc_hd__o22ai_1 U15013 ( .A1(n18882), .A2(n22841), .B1(n22926), 
        .B2(n18307), .Y(n17749) );
  sky130_fd_sc_hd__clkinv_1 U15014 ( .A(n21279), .Y(n19335) );
  sky130_fd_sc_hd__clkinv_1 U15015 ( .A(n16856), .Y(n16699) );
  sky130_fd_sc_hd__clkinv_1 U15016 ( .A(n21641), .Y(n20758) );
  sky130_fd_sc_hd__o22ai_1 U15017 ( .A1(n18882), .A2(n18295), .B1(n17589), 
        .B2(n18307), .Y(n17617) );
  sky130_fd_sc_hd__clkinv_1 U15018 ( .A(n19113), .Y(n19970) );
  sky130_fd_sc_hd__clkinv_1 U15019 ( .A(n28637), .Y(n20985) );
  sky130_fd_sc_hd__clkinv_1 U15020 ( .A(n21711), .Y(n19347) );
  sky130_fd_sc_hd__clkinv_1 U15022 ( .A(n20300), .Y(n19995) );
  sky130_fd_sc_hd__clkinv_1 U15023 ( .A(n20016), .Y(n20177) );
  sky130_fd_sc_hd__clkinv_1 U15024 ( .A(n21115), .Y(n21173) );
  sky130_fd_sc_hd__clkinv_1 U15025 ( .A(n16198), .Y(n16165) );
  sky130_fd_sc_hd__clkinv_1 U15026 ( .A(n21045), .Y(n19359) );
  sky130_fd_sc_hd__clkinv_1 U15027 ( .A(n21657), .Y(n20739) );
  sky130_fd_sc_hd__clkinv_1 U15028 ( .A(n21615), .Y(n21233) );
  sky130_fd_sc_hd__clkinv_1 U15029 ( .A(n21070), .Y(n19274) );
  sky130_fd_sc_hd__inv_1 U15030 ( .A(n21245), .Y(n21719) );
  sky130_fd_sc_hd__clkinv_1 U15031 ( .A(n21097), .Y(n19283) );
  sky130_fd_sc_hd__clkinv_1 U15032 ( .A(n21617), .Y(n21683) );
  sky130_fd_sc_hd__clkinv_1 U15033 ( .A(n21684), .Y(n21686) );
  sky130_fd_sc_hd__clkinv_1 U15034 ( .A(n24249), .Y(n24248) );
  sky130_fd_sc_hd__clkinv_1 U15035 ( .A(n19639), .Y(n19622) );
  sky130_fd_sc_hd__clkinv_1 U15036 ( .A(n16843), .Y(n16850) );
  sky130_fd_sc_hd__clkinv_1 U15037 ( .A(n16889), .Y(n16893) );
  sky130_fd_sc_hd__clkinv_1 U15038 ( .A(n19625), .Y(n19649) );
  sky130_fd_sc_hd__clkinv_1 U15039 ( .A(n23785), .Y(n25151) );
  sky130_fd_sc_hd__clkinv_1 U15040 ( .A(n18564), .Y(n12949) );
  sky130_fd_sc_hd__clkinv_1 U15041 ( .A(n21108), .Y(n21111) );
  sky130_fd_sc_hd__clkinv_1 U15042 ( .A(n15383), .Y(n15342) );
  sky130_fd_sc_hd__clkinv_1 U15043 ( .A(n15226), .Y(n15313) );
  sky130_fd_sc_hd__clkinv_1 U15044 ( .A(n21618), .Y(n21075) );
  sky130_fd_sc_hd__clkinv_1 U15045 ( .A(n15833), .Y(n15834) );
  sky130_fd_sc_hd__clkinv_1 U15046 ( .A(n21213), .Y(n21061) );
  sky130_fd_sc_hd__clkinv_1 U15047 ( .A(n22177), .Y(n22179) );
  sky130_fd_sc_hd__clkinv_1 U15048 ( .A(n16875), .Y(n16678) );
  sky130_fd_sc_hd__clkinv_1 U15049 ( .A(n28107), .Y(n10533) );
  sky130_fd_sc_hd__clkinv_1 U15050 ( .A(n22472), .Y(n22473) );
  sky130_fd_sc_hd__clkinv_1 U15051 ( .A(n22887), .Y(n22889) );
  sky130_fd_sc_hd__clkinv_1 U15052 ( .A(n16697), .Y(n16894) );
  sky130_fd_sc_hd__clkinv_1 U15053 ( .A(n22678), .Y(n22424) );
  sky130_fd_sc_hd__clkinv_1 U15054 ( .A(n21651), .Y(n20811) );
  sky130_fd_sc_hd__clkinv_1 U15055 ( .A(n20481), .Y(n15692) );
  sky130_fd_sc_hd__clkinv_1 U15056 ( .A(n12200), .Y(n11538) );
  sky130_fd_sc_hd__clkinv_1 U15057 ( .A(n22681), .Y(n22425) );
  sky130_fd_sc_hd__clkinv_1 U15058 ( .A(n28118), .Y(n10531) );
  sky130_fd_sc_hd__clkinv_1 U15059 ( .A(n16720), .Y(n16725) );
  sky130_fd_sc_hd__clkinv_1 U15060 ( .A(n16721), .Y(n16724) );
  sky130_fd_sc_hd__clkinv_1 U15061 ( .A(n16617), .Y(n16709) );
  sky130_fd_sc_hd__clkinv_1 U15062 ( .A(n19540), .Y(n19541) );
  sky130_fd_sc_hd__clkinv_1 U15063 ( .A(n22655), .Y(n22657) );
  sky130_fd_sc_hd__clkinv_1 U15064 ( .A(n21718), .Y(n20785) );
  sky130_fd_sc_hd__clkinv_1 U15065 ( .A(n19549), .Y(n19550) );
  sky130_fd_sc_hd__clkinv_1 U15066 ( .A(n16918), .Y(n16585) );
  sky130_fd_sc_hd__clkinv_1 U15067 ( .A(n22554), .Y(n22393) );
  sky130_fd_sc_hd__clkinv_1 U15068 ( .A(n22552), .Y(n22392) );
  sky130_fd_sc_hd__clkinv_1 U15069 ( .A(n20294), .Y(n20295) );
  sky130_fd_sc_hd__clkinv_1 U15070 ( .A(n22937), .Y(n22939) );
  sky130_fd_sc_hd__clkinv_1 U15071 ( .A(n26204), .Y(n26206) );
  sky130_fd_sc_hd__clkinv_1 U15072 ( .A(n19356), .Y(n17275) );
  sky130_fd_sc_hd__clkinv_1 U15073 ( .A(n22555), .Y(n22388) );
  sky130_fd_sc_hd__clkinv_1 U15074 ( .A(n24542), .Y(n24543) );
  sky130_fd_sc_hd__clkinv_1 U15075 ( .A(n19376), .Y(n17331) );
  sky130_fd_sc_hd__clkinv_1 U15076 ( .A(n22356), .Y(n22098) );
  sky130_fd_sc_hd__clkinv_1 U15077 ( .A(n20679), .Y(n15455) );
  sky130_fd_sc_hd__clkinv_1 U15078 ( .A(j202_soc_core_wbqspiflash_00_N710), 
        .Y(n27123) );
  sky130_fd_sc_hd__clkinv_1 U15079 ( .A(n19747), .Y(n19748) );
  sky130_fd_sc_hd__clkinv_1 U15080 ( .A(n15696), .Y(n20647) );
  sky130_fd_sc_hd__clkinv_1 U15081 ( .A(n20252), .Y(n20844) );
  sky130_fd_sc_hd__clkinv_1 U15082 ( .A(n29358), .Y(n25983) );
  sky130_fd_sc_hd__clkinv_1 U15083 ( .A(n28743), .Y(n26209) );
  sky130_fd_sc_hd__clkinv_1 U15084 ( .A(n20111), .Y(n20841) );
  sky130_fd_sc_hd__clkinv_1 U15085 ( .A(n20653), .Y(n15735) );
  sky130_fd_sc_hd__inv_6 U15086 ( .A(n18183), .Y(n18307) );
  sky130_fd_sc_hd__clkinv_1 U15087 ( .A(n15713), .Y(n20641) );
  sky130_fd_sc_hd__and2_0 U15088 ( .A(n15560), .B(n15534), .X(n13464) );
  sky130_fd_sc_hd__clkinv_1 U15089 ( .A(n19744), .Y(n19745) );
  sky130_fd_sc_hd__clkinv_1 U15090 ( .A(n15332), .Y(n15228) );
  sky130_fd_sc_hd__clkinv_1 U15091 ( .A(n26287), .Y(n26285) );
  sky130_fd_sc_hd__clkinv_1 U15092 ( .A(n16175), .Y(n16785) );
  sky130_fd_sc_hd__clkinv_1 U15094 ( .A(n21068), .Y(n21069) );
  sky130_fd_sc_hd__clkinv_1 U15095 ( .A(n25329), .Y(n25330) );
  sky130_fd_sc_hd__clkinv_1 U15096 ( .A(n20773), .Y(n21132) );
  sky130_fd_sc_hd__clkinv_1 U15097 ( .A(n21078), .Y(n21716) );
  sky130_fd_sc_hd__clkinv_1 U15098 ( .A(n21704), .Y(n21707) );
  sky130_fd_sc_hd__and2_0 U15099 ( .A(n13948), .B(n13947), .X(n11978) );
  sky130_fd_sc_hd__clkinv_1 U15100 ( .A(n19544), .Y(n19547) );
  sky130_fd_sc_hd__clkinv_1 U15101 ( .A(n11614), .Y(n26878) );
  sky130_fd_sc_hd__clkinv_1 U15102 ( .A(n23858), .Y(n23191) );
  sky130_fd_sc_hd__clkinv_1 U15103 ( .A(n19752), .Y(n19718) );
  sky130_fd_sc_hd__nand3_1 U15104 ( .A(n13305), .B(n15844), .C(n14870), .Y(
        n16118) );
  sky130_fd_sc_hd__clkinv_1 U15105 ( .A(n16620), .Y(n16195) );
  sky130_fd_sc_hd__clkinv_1 U15106 ( .A(n24244), .Y(n24245) );
  sky130_fd_sc_hd__clkinv_1 U15107 ( .A(n19628), .Y(n19640) );
  sky130_fd_sc_hd__clkinv_1 U15108 ( .A(n19722), .Y(n19740) );
  sky130_fd_sc_hd__clkinv_1 U15109 ( .A(n19539), .Y(n19543) );
  sky130_fd_sc_hd__clkinv_1 U15110 ( .A(n19656), .Y(n19621) );
  sky130_fd_sc_hd__clkinv_1 U15111 ( .A(n19724), .Y(n19735) );
  sky130_fd_sc_hd__clkinv_1 U15112 ( .A(n27915), .Y(n27916) );
  sky130_fd_sc_hd__clkinv_1 U15113 ( .A(n16914), .Y(n16916) );
  sky130_fd_sc_hd__clkinv_1 U15114 ( .A(n20611), .Y(n20458) );
  sky130_fd_sc_hd__clkinv_1 U15115 ( .A(n16059), .Y(n16062) );
  sky130_fd_sc_hd__nor2_1 U15116 ( .A(n11403), .B(n11398), .Y(n11397) );
  sky130_fd_sc_hd__clkinv_1 U15117 ( .A(n20121), .Y(n20170) );
  sky130_fd_sc_hd__nor2_1 U15118 ( .A(n12100), .B(n12095), .Y(n12094) );
  sky130_fd_sc_hd__clkinv_1 U15119 ( .A(n18958), .Y(n21198) );
  sky130_fd_sc_hd__clkinv_1 U15120 ( .A(n15691), .Y(n15471) );
  sky130_fd_sc_hd__clkinv_1 U15121 ( .A(n19690), .Y(n19698) );
  sky130_fd_sc_hd__clkinv_1 U15122 ( .A(n16112), .Y(n16115) );
  sky130_fd_sc_hd__clkinv_1 U15123 ( .A(n19114), .Y(n19897) );
  sky130_fd_sc_hd__clkinv_1 U15124 ( .A(n26233), .Y(n23912) );
  sky130_fd_sc_hd__clkinv_1 U15125 ( .A(n20323), .Y(n20008) );
  sky130_fd_sc_hd__fa_1 U15126 ( .A(n18731), .B(n18729), .CIN(n18730), .COUT(
        n18726), .SUM(n18806) );
  sky130_fd_sc_hd__clkinv_1 U15127 ( .A(n16114), .Y(n14872) );
  sky130_fd_sc_hd__clkinv_1 U15128 ( .A(n16776), .Y(n16687) );
  sky130_fd_sc_hd__clkinv_1 U15129 ( .A(n20646), .Y(n20531) );
  sky130_fd_sc_hd__clkinv_1 U15130 ( .A(n15560), .Y(n15563) );
  sky130_fd_sc_hd__clkinv_1 U15131 ( .A(n15556), .Y(n15559) );
  sky130_fd_sc_hd__clkinv_1 U15132 ( .A(n18966), .Y(n21645) );
  sky130_fd_sc_hd__clkinv_1 U15133 ( .A(n15544), .Y(n15549) );
  sky130_fd_sc_hd__clkinv_1 U15134 ( .A(n20336), .Y(n19951) );
  sky130_fd_sc_hd__clkinv_1 U15135 ( .A(n21215), .Y(n19353) );
  sky130_fd_sc_hd__clkinv_1 U15136 ( .A(n15331), .Y(n15333) );
  sky130_fd_sc_hd__inv_2 U15137 ( .A(n17599), .Y(n17555) );
  sky130_fd_sc_hd__clkinv_1 U15138 ( .A(n21613), .Y(n19387) );
  sky130_fd_sc_hd__clkinv_1 U15139 ( .A(n24799), .Y(n15519) );
  sky130_fd_sc_hd__clkinv_1 U15140 ( .A(n15457), .Y(n15693) );
  sky130_fd_sc_hd__clkinv_1 U15141 ( .A(n17219), .Y(n20358) );
  sky130_fd_sc_hd__clkinv_1 U15142 ( .A(n16917), .Y(n16599) );
  sky130_fd_sc_hd__clkinv_1 U15143 ( .A(n17042), .Y(n17043) );
  sky130_fd_sc_hd__nor2_1 U15144 ( .A(n12794), .B(n12799), .Y(n17355) );
  sky130_fd_sc_hd__clkinv_1 U15145 ( .A(n20349), .Y(n20063) );
  sky130_fd_sc_hd__clkinv_1 U15146 ( .A(n16935), .Y(n16867) );
  sky130_fd_sc_hd__clkinv_1 U15147 ( .A(n21714), .Y(n21174) );
  sky130_fd_sc_hd__clkinv_1 U15148 ( .A(n15310), .Y(n13413) );
  sky130_fd_sc_hd__clkinv_1 U15149 ( .A(n15220), .Y(n15363) );
  sky130_fd_sc_hd__clkinv_1 U15150 ( .A(n20096), .Y(n19879) );
  sky130_fd_sc_hd__clkinv_1 U15151 ( .A(n20462), .Y(n20569) );
  sky130_fd_sc_hd__clkinv_1 U15152 ( .A(n15361), .Y(n15368) );
  sky130_fd_sc_hd__and2_0 U15153 ( .A(n20736), .B(n19284), .X(n21185) );
  sky130_fd_sc_hd__clkinv_1 U15154 ( .A(n16890), .Y(n16565) );
  sky130_fd_sc_hd__clkinv_1 U15155 ( .A(n11597), .Y(n11595) );
  sky130_fd_sc_hd__clkinv_1 U15156 ( .A(n21265), .Y(n21266) );
  sky130_fd_sc_hd__clkinv_1 U15157 ( .A(n13415), .Y(n15381) );
  sky130_fd_sc_hd__nor2_1 U15158 ( .A(n11333), .B(n11328), .Y(n11327) );
  sky130_fd_sc_hd__clkinv_1 U15159 ( .A(n18937), .Y(n19286) );
  sky130_fd_sc_hd__clkinv_1 U15160 ( .A(n20897), .Y(n20196) );
  sky130_fd_sc_hd__clkinv_1 U15161 ( .A(n15254), .Y(n15255) );
  sky130_fd_sc_hd__clkinv_1 U15162 ( .A(n24585), .Y(n29354) );
  sky130_fd_sc_hd__clkinv_1 U15163 ( .A(n21656), .Y(n21257) );
  sky130_fd_sc_hd__clkinv_1 U15164 ( .A(n20514), .Y(n15470) );
  sky130_fd_sc_hd__clkinv_1 U15165 ( .A(n19997), .Y(n20241) );
  sky130_fd_sc_hd__clkinv_1 U15166 ( .A(n18083), .Y(n11580) );
  sky130_fd_sc_hd__clkinv_1 U15167 ( .A(n16835), .Y(n16766) );
  sky130_fd_sc_hd__clkinv_1 U15168 ( .A(n16558), .Y(n16836) );
  sky130_fd_sc_hd__clkinv_1 U15169 ( .A(n19754), .Y(n19755) );
  sky130_fd_sc_hd__clkinv_1 U15170 ( .A(n21190), .Y(n17292) );
  sky130_fd_sc_hd__clkinv_1 U15171 ( .A(n20883), .Y(n17221) );
  sky130_fd_sc_hd__clkinv_1 U15172 ( .A(n21093), .Y(n21100) );
  sky130_fd_sc_hd__clkinv_1 U15173 ( .A(n29059), .Y(n27018) );
  sky130_fd_sc_hd__clkinv_1 U15174 ( .A(n27166), .Y(n24394) );
  sky130_fd_sc_hd__clkinv_1 U15175 ( .A(n22479), .Y(n22418) );
  sky130_fd_sc_hd__clkinv_1 U15176 ( .A(n22229), .Y(n22230) );
  sky130_fd_sc_hd__clkinv_1 U15177 ( .A(n14944), .Y(n14866) );
  sky130_fd_sc_hd__clkinv_1 U15178 ( .A(n23523), .Y(n23528) );
  sky130_fd_sc_hd__clkinv_1 U15179 ( .A(n15319), .Y(n15550) );
  sky130_fd_sc_hd__clkinv_1 U15180 ( .A(n15596), .Y(n15364) );
  sky130_fd_sc_hd__clkinv_1 U15181 ( .A(n15258), .Y(n15530) );
  sky130_fd_sc_hd__clkinv_1 U15182 ( .A(n20634), .Y(n20662) );
  sky130_fd_sc_hd__clkinv_1 U15183 ( .A(n22235), .Y(n22237) );
  sky130_fd_sc_hd__clkinv_1 U15184 ( .A(n16844), .Y(n16962) );
  sky130_fd_sc_hd__clkinv_1 U15185 ( .A(n11442), .Y(n22247) );
  sky130_fd_sc_hd__clkinv_1 U15186 ( .A(n20502), .Y(n20506) );
  sky130_fd_sc_hd__clkinv_1 U15187 ( .A(n16868), .Y(n16741) );
  sky130_fd_sc_hd__clkinv_1 U15188 ( .A(n25781), .Y(n25783) );
  sky130_fd_sc_hd__nand2_1 U15189 ( .A(n19676), .B(n19675), .Y(n19686) );
  sky130_fd_sc_hd__clkinv_1 U15190 ( .A(n18773), .Y(n11437) );
  sky130_fd_sc_hd__clkinv_1 U15191 ( .A(n22615), .Y(n11147) );
  sky130_fd_sc_hd__clkinv_1 U15192 ( .A(n26351), .Y(n24067) );
  sky130_fd_sc_hd__clkinv_1 U15193 ( .A(n14904), .Y(n14865) );
  sky130_fd_sc_hd__clkinv_1 U15194 ( .A(n28238), .Y(n28073) );
  sky130_fd_sc_hd__clkinv_1 U15195 ( .A(n28078), .Y(n28093) );
  sky130_fd_sc_hd__clkinv_1 U15196 ( .A(n28187), .Y(n28172) );
  sky130_fd_sc_hd__o2bb2ai_1 U15197 ( .B1(n11110), .B2(n23172), .A1_N(n23129), 
        .A2_N(n23174), .Y(n23131) );
  sky130_fd_sc_hd__clkinv_1 U15198 ( .A(n22007), .Y(n22009) );
  sky130_fd_sc_hd__clkinv_1 U15199 ( .A(n18758), .Y(n11784) );
  sky130_fd_sc_hd__clkinv_1 U15200 ( .A(n22394), .Y(n22391) );
  sky130_fd_sc_hd__clkinv_1 U15201 ( .A(n15359), .Y(n15266) );
  sky130_fd_sc_hd__clkinv_1 U15202 ( .A(n16685), .Y(n16610) );
  sky130_fd_sc_hd__clkinv_1 U15203 ( .A(n26846), .Y(n26848) );
  sky130_fd_sc_hd__clkinv_1 U15205 ( .A(n22387), .Y(n22395) );
  sky130_fd_sc_hd__clkinv_1 U15206 ( .A(n25188), .Y(n25189) );
  sky130_fd_sc_hd__clkinv_1 U15207 ( .A(n19737), .Y(n19738) );
  sky130_fd_sc_hd__clkinv_1 U15208 ( .A(n27829), .Y(n24845) );
  sky130_fd_sc_hd__inv_1 U15209 ( .A(n20582), .Y(n20521) );
  sky130_fd_sc_hd__and2_0 U15210 ( .A(n20384), .B(n20884), .X(n20331) );
  sky130_fd_sc_hd__clkinv_1 U15211 ( .A(n28628), .Y(n28030) );
  sky130_fd_sc_hd__clkinv_1 U15212 ( .A(n15880), .Y(n14900) );
  sky130_fd_sc_hd__clkinv_1 U15213 ( .A(n22422), .Y(n22385) );
  sky130_fd_sc_hd__clkinv_1 U15214 ( .A(n15545), .Y(n15570) );
  sky130_fd_sc_hd__clkinv_1 U15215 ( .A(n22096), .Y(n22095) );
  sky130_fd_sc_hd__clkinv_1 U15216 ( .A(n14942), .Y(n15817) );
  sky130_fd_sc_hd__clkinv_1 U15217 ( .A(n20440), .Y(n20612) );
  sky130_fd_sc_hd__clkinv_1 U15218 ( .A(n19729), .Y(n19753) );
  sky130_fd_sc_hd__clkinv_1 U15219 ( .A(n20354), .Y(n20075) );
  sky130_fd_sc_hd__clkinv_1 U15220 ( .A(n25300), .Y(n25302) );
  sky130_fd_sc_hd__and2_0 U15221 ( .A(n21243), .B(n21286), .X(n21258) );
  sky130_fd_sc_hd__clkinv_1 U15222 ( .A(n15609), .Y(n13467) );
  sky130_fd_sc_hd__clkinv_1 U15223 ( .A(n15498), .Y(n15499) );
  sky130_fd_sc_hd__clkinv_1 U15224 ( .A(n22074), .Y(n22097) );
  sky130_fd_sc_hd__clkinv_1 U15226 ( .A(n21985), .Y(n25791) );
  sky130_fd_sc_hd__clkinv_1 U15227 ( .A(n19489), .Y(n26327) );
  sky130_fd_sc_hd__clkinv_1 U15228 ( .A(n20884), .Y(n20888) );
  sky130_fd_sc_hd__clkinv_1 U15229 ( .A(n22950), .Y(n22221) );
  sky130_fd_sc_hd__clkinv_1 U15230 ( .A(n20477), .Y(n15672) );
  sky130_fd_sc_hd__clkinv_1 U15231 ( .A(n22086), .Y(n22079) );
  sky130_fd_sc_hd__clkinv_1 U15232 ( .A(n19741), .Y(n19721) );
  sky130_fd_sc_hd__clkinv_1 U15233 ( .A(n22420), .Y(n22427) );
  sky130_fd_sc_hd__clkinv_1 U15234 ( .A(n22390), .Y(n22050) );
  sky130_fd_sc_hd__clkinv_1 U15235 ( .A(n19184), .Y(n22731) );
  sky130_fd_sc_hd__clkinv_1 U15236 ( .A(n22426), .Y(n22423) );
  sky130_fd_sc_hd__clkinv_1 U15237 ( .A(n22088), .Y(n22087) );
  sky130_fd_sc_hd__clkinv_1 U15238 ( .A(n17085), .Y(n17086) );
  sky130_fd_sc_hd__clkinv_1 U15239 ( .A(n19647), .Y(n11699) );
  sky130_fd_sc_hd__clkinv_1 U15240 ( .A(n28737), .Y(n28649) );
  sky130_fd_sc_hd__clkinv_1 U15241 ( .A(n17243), .Y(n17246) );
  sky130_fd_sc_hd__clkinv_1 U15242 ( .A(n21098), .Y(n21230) );
  sky130_fd_sc_hd__clkinv_1 U15243 ( .A(n28739), .Y(n28731) );
  sky130_fd_sc_hd__clkinv_1 U15244 ( .A(n19588), .Y(n19599) );
  sky130_fd_sc_hd__clkinv_1 U15245 ( .A(n19991), .Y(n19943) );
  sky130_fd_sc_hd__clkinv_1 U15246 ( .A(n15757), .Y(n15758) );
  sky130_fd_sc_hd__clkinv_1 U15247 ( .A(n17244), .Y(n17245) );
  sky130_fd_sc_hd__and2_0 U15248 ( .A(n15609), .B(n15340), .X(n15531) );
  sky130_fd_sc_hd__clkinv_1 U15249 ( .A(n19633), .Y(n19657) );
  sky130_fd_sc_hd__inv_2 U15250 ( .A(n20842), .Y(n20924) );
  sky130_fd_sc_hd__and2_0 U15251 ( .A(n20305), .B(n20047), .X(n13302) );
  sky130_fd_sc_hd__clkinv_1 U15252 ( .A(n21286), .Y(n17319) );
  sky130_fd_sc_hd__clkinv_1 U15254 ( .A(n20082), .Y(n17206) );
  sky130_fd_sc_hd__clkinv_1 U15255 ( .A(n15689), .Y(n15680) );
  sky130_fd_sc_hd__clkinv_1 U15256 ( .A(n16576), .Y(n16205) );
  sky130_fd_sc_hd__clkinv_1 U15257 ( .A(n21688), .Y(n19350) );
  sky130_fd_sc_hd__clkinv_1 U15258 ( .A(n28647), .Y(n25011) );
  sky130_fd_sc_hd__clkinv_1 U15259 ( .A(n20574), .Y(n15706) );
  sky130_fd_sc_hd__clkinv_1 U15260 ( .A(n19641), .Y(n19642) );
  sky130_fd_sc_hd__clkinv_1 U15261 ( .A(n11635), .Y(n11633) );
  sky130_fd_sc_hd__clkinv_1 U15262 ( .A(n19644), .Y(n19646) );
  sky130_fd_sc_hd__clkinv_1 U15263 ( .A(n19650), .Y(n19624) );
  sky130_fd_sc_hd__clkinv_1 U15264 ( .A(n14006), .Y(n14007) );
  sky130_fd_sc_hd__and2_0 U15265 ( .A(n15533), .B(n15564), .X(n15601) );
  sky130_fd_sc_hd__clkinv_1 U15266 ( .A(n15366), .Y(n15367) );
  sky130_fd_sc_hd__clkinv_1 U15267 ( .A(n16201), .Y(n16619) );
  sky130_fd_sc_hd__clkinv_1 U15268 ( .A(n25938), .Y(n23463) );
  sky130_fd_sc_hd__clkinv_1 U15269 ( .A(n16769), .Y(n16778) );
  sky130_fd_sc_hd__clkinv_1 U15270 ( .A(n16770), .Y(n16196) );
  sky130_fd_sc_hd__clkinv_1 U15271 ( .A(n19272), .Y(n20801) );
  sky130_fd_sc_hd__clkinv_1 U15272 ( .A(n20004), .Y(n19891) );
  sky130_fd_sc_hd__clkinv_1 U15273 ( .A(n17027), .Y(n15787) );
  sky130_fd_sc_hd__and2_0 U15274 ( .A(n19969), .B(n20080), .X(n20228) );
  sky130_fd_sc_hd__and2_0 U15275 ( .A(n19971), .B(n20375), .X(n20896) );
  sky130_fd_sc_hd__clkinv_1 U15276 ( .A(n28581), .Y(n24233) );
  sky130_fd_sc_hd__clkinv_1 U15277 ( .A(n15347), .Y(n15348) );
  sky130_fd_sc_hd__clkinv_1 U15278 ( .A(n17016), .Y(n15798) );
  sky130_fd_sc_hd__clkinv_1 U15279 ( .A(n17903), .Y(n17595) );
  sky130_fd_sc_hd__clkinv_1 U15280 ( .A(n26260), .Y(n26262) );
  sky130_fd_sc_hd__nand2b_1 U15281 ( .A_N(n14009), .B(n13790), .Y(n16322) );
  sky130_fd_sc_hd__clkinv_1 U15282 ( .A(n20305), .Y(n20010) );
  sky130_fd_sc_hd__clkinv_1 U15283 ( .A(n21243), .Y(n21249) );
  sky130_fd_sc_hd__clkinv_1 U15284 ( .A(n15350), .Y(n15253) );
  sky130_fd_sc_hd__clkinv_1 U15285 ( .A(n15866), .Y(n16104) );
  sky130_fd_sc_hd__inv_1 U15286 ( .A(n20306), .Y(n20011) );
  sky130_fd_sc_hd__clkinv_1 U15287 ( .A(n16882), .Y(n16904) );
  sky130_fd_sc_hd__clkinv_1 U15288 ( .A(n15407), .Y(n15656) );
  sky130_fd_sc_hd__and2_0 U15289 ( .A(n20221), .B(n20350), .X(n20052) );
  sky130_fd_sc_hd__clkinv_1 U15290 ( .A(n24687), .Y(n23780) );
  sky130_fd_sc_hd__nor2_1 U15291 ( .A(n17290), .B(n17278), .Y(n20778) );
  sky130_fd_sc_hd__clkinv_1 U15292 ( .A(n21203), .Y(n20751) );
  sky130_fd_sc_hd__clkinv_1 U15293 ( .A(n21206), .Y(n21208) );
  sky130_fd_sc_hd__clkinv_1 U15294 ( .A(n15801), .Y(n14875) );
  sky130_fd_sc_hd__clkinv_1 U15295 ( .A(n17024), .Y(n16101) );
  sky130_fd_sc_hd__and2_0 U15296 ( .A(n15613), .B(n15340), .X(n15222) );
  sky130_fd_sc_hd__clkinv_1 U15297 ( .A(n28615), .Y(n28945) );
  sky130_fd_sc_hd__clkinv_1 U15299 ( .A(n20772), .Y(n18936) );
  sky130_fd_sc_hd__clkinv_1 U15300 ( .A(n13430), .Y(n13432) );
  sky130_fd_sc_hd__clkinv_1 U15301 ( .A(n28606), .Y(n28938) );
  sky130_fd_sc_hd__clkinv_1 U15302 ( .A(n19382), .Y(n21040) );
  sky130_fd_sc_hd__clkinv_1 U15303 ( .A(n25529), .Y(n21585) );
  sky130_fd_sc_hd__clkinv_1 U15304 ( .A(n20045), .Y(n21646) );
  sky130_fd_sc_hd__clkinv_1 U15305 ( .A(n16677), .Y(n16592) );
  sky130_fd_sc_hd__clkinv_1 U15306 ( .A(n15321), .Y(n15592) );
  sky130_fd_sc_hd__clkinv_1 U15307 ( .A(n20411), .Y(n20413) );
  sky130_fd_sc_hd__and2_0 U15308 ( .A(n17010), .B(n16078), .X(n13305) );
  sky130_fd_sc_hd__clkinv_1 U15309 ( .A(n16714), .Y(n16961) );
  sky130_fd_sc_hd__clkinv_1 U15310 ( .A(n17048), .Y(n14878) );
  sky130_fd_sc_hd__clkinv_1 U15311 ( .A(n28245), .Y(n28247) );
  sky130_fd_sc_hd__and2_0 U15312 ( .A(n20885), .B(n21206), .X(n19088) );
  sky130_fd_sc_hd__clkinv_1 U15313 ( .A(n21319), .Y(n21341) );
  sky130_fd_sc_hd__clkinv_1 U15314 ( .A(n21631), .Y(n21109) );
  sky130_fd_sc_hd__and2_0 U15316 ( .A(n17007), .B(n15796), .X(n14915) );
  sky130_fd_sc_hd__clkinv_1 U15317 ( .A(n20601), .Y(n20630) );
  sky130_fd_sc_hd__clkinv_1 U15318 ( .A(n17007), .Y(n15852) );
  sky130_fd_sc_hd__inv_2 U15319 ( .A(n15723), .Y(n20680) );
  sky130_fd_sc_hd__clkinv_1 U15320 ( .A(n14926), .Y(n16117) );
  sky130_fd_sc_hd__clkinv_1 U15321 ( .A(n15340), .Y(n13438) );
  sky130_fd_sc_hd__clkinv_1 U15322 ( .A(n15671), .Y(n15724) );
  sky130_fd_sc_hd__clkinv_1 U15323 ( .A(n24738), .Y(n23776) );
  sky130_fd_sc_hd__clkinv_1 U15324 ( .A(n28629), .Y(n28630) );
  sky130_fd_sc_hd__clkinv_1 U15325 ( .A(n23940), .Y(n24494) );
  sky130_fd_sc_hd__clkinv_1 U15326 ( .A(n15369), .Y(n13479) );
  sky130_fd_sc_hd__clkinv_1 U15327 ( .A(n22004), .Y(n22932) );
  sky130_fd_sc_hd__inv_1 U15328 ( .A(n18755), .Y(n18702) );
  sky130_fd_sc_hd__clkinv_1 U15329 ( .A(n28551), .Y(n28549) );
  sky130_fd_sc_hd__clkinv_1 U15330 ( .A(n15537), .Y(n13390) );
  sky130_fd_sc_hd__clkinv_1 U15331 ( .A(n19841), .Y(n19842) );
  sky130_fd_sc_hd__clkinv_1 U15332 ( .A(n20606), .Y(n15738) );
  sky130_fd_sc_hd__clkinv_1 U15333 ( .A(n20637), .Y(n20661) );
  sky130_fd_sc_hd__clkinv_1 U15334 ( .A(n21228), .Y(n19334) );
  sky130_fd_sc_hd__clkinv_1 U15335 ( .A(n15612), .Y(n15622) );
  sky130_fd_sc_hd__clkinv_1 U15336 ( .A(n18952), .Y(n17333) );
  sky130_fd_sc_hd__clkinv_1 U15337 ( .A(n20602), .Y(n15733) );
  sky130_fd_sc_hd__clkinv_1 U15338 ( .A(n17070), .Y(n16100) );
  sky130_fd_sc_hd__and2_0 U15339 ( .A(n26977), .B(n11713), .X(n22956) );
  sky130_fd_sc_hd__clkinv_1 U15340 ( .A(n17030), .Y(n14864) );
  sky130_fd_sc_hd__clkinv_1 U15341 ( .A(n14946), .Y(n14947) );
  sky130_fd_sc_hd__clkinv_1 U15342 ( .A(n14954), .Y(n15882) );
  sky130_fd_sc_hd__clkinv_1 U15343 ( .A(n17014), .Y(n16102) );
  sky130_fd_sc_hd__clkinv_1 U15344 ( .A(n25858), .Y(n28932) );
  sky130_fd_sc_hd__or2_0 U15345 ( .A(n18237), .B(n18236), .X(n18321) );
  sky130_fd_sc_hd__inv_2 U15346 ( .A(n18700), .Y(n18676) );
  sky130_fd_sc_hd__clkinv_1 U15347 ( .A(n20843), .Y(n20168) );
  sky130_fd_sc_hd__clkinv_1 U15348 ( .A(n15741), .Y(n15707) );
  sky130_fd_sc_hd__clkinv_1 U15349 ( .A(n16953), .Y(n20513) );
  sky130_fd_sc_hd__clkinv_1 U15351 ( .A(n22456), .Y(n22459) );
  sky130_fd_sc_hd__clkinv_1 U15352 ( .A(n14897), .Y(n17035) );
  sky130_fd_sc_hd__clkinv_1 U15353 ( .A(n28028), .Y(n28031) );
  sky130_fd_sc_hd__clkinv_1 U15354 ( .A(n21267), .Y(n21627) );
  sky130_fd_sc_hd__clkinv_1 U15355 ( .A(n15814), .Y(n14901) );
  sky130_fd_sc_hd__clkinv_1 U15356 ( .A(n15589), .Y(n15623) );
  sky130_fd_sc_hd__clkinv_1 U15357 ( .A(n15482), .Y(n15484) );
  sky130_fd_sc_hd__and2_0 U15358 ( .A(n18866), .B(n18892), .X(n11684) );
  sky130_fd_sc_hd__clkinv_1 U15359 ( .A(n24142), .Y(n18884) );
  sky130_fd_sc_hd__nand2_2 U15360 ( .A(n17361), .B(n17360), .Y(n23253) );
  sky130_fd_sc_hd__clkinv_1 U15361 ( .A(n17010), .Y(n17011) );
  sky130_fd_sc_hd__inv_1 U15362 ( .A(n17073), .Y(n14861) );
  sky130_fd_sc_hd__clkinv_1 U15363 ( .A(n20532), .Y(n15676) );
  sky130_fd_sc_hd__clkinv_1 U15364 ( .A(n26277), .Y(n26278) );
  sky130_fd_sc_hd__clkinv_1 U15365 ( .A(n23049), .Y(n21888) );
  sky130_fd_sc_hd__clkinv_1 U15366 ( .A(n25905), .Y(n28213) );
  sky130_fd_sc_hd__clkinv_1 U15367 ( .A(n24507), .Y(n24509) );
  sky130_fd_sc_hd__clkinv_1 U15368 ( .A(n27817), .Y(n27901) );
  sky130_fd_sc_hd__clkinv_1 U15369 ( .A(n26298), .Y(n26297) );
  sky130_fd_sc_hd__clkinv_1 U15370 ( .A(n25779), .Y(n25780) );
  sky130_fd_sc_hd__clkinv_1 U15371 ( .A(n26102), .Y(n25181) );
  sky130_fd_sc_hd__clkinv_1 U15372 ( .A(n27951), .Y(n24432) );
  sky130_fd_sc_hd__clkinv_1 U15373 ( .A(n28261), .Y(n28069) );
  sky130_fd_sc_hd__clkinv_1 U15374 ( .A(n28061), .Y(n28062) );
  sky130_fd_sc_hd__clkinv_1 U15375 ( .A(n16177), .Y(n16164) );
  sky130_fd_sc_hd__clkinv_1 U15376 ( .A(n16182), .Y(n16692) );
  sky130_fd_sc_hd__clkinv_1 U15377 ( .A(n24905), .Y(n24906) );
  sky130_fd_sc_hd__nor2_1 U15378 ( .A(n19873), .B(n17168), .Y(n20110) );
  sky130_fd_sc_hd__clkinv_1 U15379 ( .A(n20214), .Y(n17228) );
  sky130_fd_sc_hd__clkinv_1 U15380 ( .A(n19822), .Y(n19823) );
  sky130_fd_sc_hd__clkinv_1 U15381 ( .A(n28550), .Y(n28171) );
  sky130_fd_sc_hd__clkinv_1 U15382 ( .A(n26475), .Y(n26162) );
  sky130_fd_sc_hd__clkinv_1 U15383 ( .A(n23701), .Y(n23702) );
  sky130_fd_sc_hd__clkinv_1 U15384 ( .A(n23698), .Y(n23700) );
  sky130_fd_sc_hd__clkinv_1 U15385 ( .A(n20375), .Y(n17227) );
  sky130_fd_sc_hd__clkinv_1 U15386 ( .A(n16879), .Y(n16207) );
  sky130_fd_sc_hd__inv_2 U15387 ( .A(n12169), .Y(n16248) );
  sky130_fd_sc_hd__clkinv_1 U15388 ( .A(n28096), .Y(n26192) );
  sky130_fd_sc_hd__inv_2 U15389 ( .A(n15063), .Y(n16325) );
  sky130_fd_sc_hd__clkinv_1 U15390 ( .A(n16857), .Y(n16675) );
  sky130_fd_sc_hd__clkinv_1 U15391 ( .A(n23957), .Y(n23198) );
  sky130_fd_sc_hd__o2bb2ai_1 U15392 ( .B1(n23089), .B2(n23172), .A1_N(n23088), 
        .A2_N(n23174), .Y(n23090) );
  sky130_fd_sc_hd__o2bb2ai_1 U15393 ( .B1(n23113), .B2(n23172), .A1_N(n23112), 
        .A2_N(n23174), .Y(n23114) );
  sky130_fd_sc_hd__clkinv_1 U15394 ( .A(n23462), .Y(n23464) );
  sky130_fd_sc_hd__clkinv_1 U15395 ( .A(n16598), .Y(n16842) );
  sky130_fd_sc_hd__a21oi_2 U15396 ( .A1(n19511), .A2(n19510), .B1(n19509), .Y(
        n26846) );
  sky130_fd_sc_hd__clkinv_1 U15397 ( .A(n25763), .Y(n29359) );
  sky130_fd_sc_hd__clkinv_1 U15398 ( .A(n26200), .Y(n26201) );
  sky130_fd_sc_hd__clkinv_1 U15399 ( .A(n28640), .Y(n25009) );
  sky130_fd_sc_hd__clkinv_1 U15400 ( .A(n16849), .Y(n16216) );
  sky130_fd_sc_hd__clkinv_1 U15401 ( .A(n28083), .Y(n28248) );
  sky130_fd_sc_hd__a2bb2oi_1 U15402 ( .B1(n22965), .B2(n24505), .A1_N(n26398), 
        .A2_N(n24507), .Y(n22630) );
  sky130_fd_sc_hd__clkinv_1 U15403 ( .A(n23575), .Y(n23576) );
  sky130_fd_sc_hd__nor2_1 U15404 ( .A(n11912), .B(n23706), .Y(n11911) );
  sky130_fd_sc_hd__clkinv_1 U15405 ( .A(n25885), .Y(n23479) );
  sky130_fd_sc_hd__clkinv_1 U15406 ( .A(n16767), .Y(n16837) );
  sky130_fd_sc_hd__clkinv_1 U15407 ( .A(n26014), .Y(n26015) );
  sky130_fd_sc_hd__clkinv_1 U15408 ( .A(n26247), .Y(n25989) );
  sky130_fd_sc_hd__clkinv_1 U15409 ( .A(n16903), .Y(n16735) );
  sky130_fd_sc_hd__clkinv_1 U15410 ( .A(n24481), .Y(n19411) );
  sky130_fd_sc_hd__clkinv_1 U15411 ( .A(n14059), .Y(n11887) );
  sky130_fd_sc_hd__clkinv_1 U15412 ( .A(n14939), .Y(n17076) );
  sky130_fd_sc_hd__clkinv_1 U15413 ( .A(n14934), .Y(n14935) );
  sky130_fd_sc_hd__clkinv_1 U15414 ( .A(n28250), .Y(n28103) );
  sky130_fd_sc_hd__clkinv_1 U15415 ( .A(n24874), .Y(n24873) );
  sky130_fd_sc_hd__clkinv_1 U15416 ( .A(n24951), .Y(n24957) );
  sky130_fd_sc_hd__clkinv_1 U15417 ( .A(n24831), .Y(n24827) );
  sky130_fd_sc_hd__clkinv_1 U15418 ( .A(n24393), .Y(n24395) );
  sky130_fd_sc_hd__clkinv_1 U15419 ( .A(n28211), .Y(n28254) );
  sky130_fd_sc_hd__clkinv_1 U15420 ( .A(n25247), .Y(n25248) );
  sky130_fd_sc_hd__clkinv_1 U15421 ( .A(n16872), .Y(n16713) );
  sky130_fd_sc_hd__clkinv_1 U15422 ( .A(n26013), .Y(n26016) );
  sky130_fd_sc_hd__clkinv_1 U15423 ( .A(n23500), .Y(n23501) );
  sky130_fd_sc_hd__clkinv_1 U15424 ( .A(n22601), .Y(n25676) );
  sky130_fd_sc_hd__clkinv_1 U15425 ( .A(n26194), .Y(n26195) );
  sky130_fd_sc_hd__and2_0 U15426 ( .A(n25344), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n12300) );
  sky130_fd_sc_hd__and2_0 U15427 ( .A(n20632), .B(n16616), .X(n20592) );
  sky130_fd_sc_hd__clkinv_1 U15428 ( .A(n25897), .Y(n25898) );
  sky130_fd_sc_hd__a21oi_2 U15429 ( .A1(n19585), .A2(n19584), .B1(n19583), .Y(
        n26842) );
  sky130_fd_sc_hd__clkinv_1 U15430 ( .A(n23525), .Y(n23526) );
  sky130_fd_sc_hd__clkinv_1 U15431 ( .A(n23524), .Y(n23527) );
  sky130_fd_sc_hd__clkinv_1 U15432 ( .A(n15431), .Y(n15429) );
  sky130_fd_sc_hd__clkinv_1 U15433 ( .A(n23564), .Y(n23859) );
  sky130_fd_sc_hd__clkinv_1 U15434 ( .A(n23255), .Y(n23267) );
  sky130_fd_sc_hd__clkinv_1 U15435 ( .A(n16073), .Y(n16074) );
  sky130_fd_sc_hd__clkinv_1 U15437 ( .A(n20683), .Y(n20533) );
  sky130_fd_sc_hd__clkinv_1 U15438 ( .A(n28620), .Y(n28621) );
  sky130_fd_sc_hd__clkinv_1 U15439 ( .A(n19858), .Y(n17201) );
  sky130_fd_sc_hd__clkinv_1 U15440 ( .A(n17203), .Y(n20164) );
  sky130_fd_sc_hd__clkinv_1 U15441 ( .A(n23699), .Y(n23483) );
  sky130_fd_sc_hd__clkinv_1 U15442 ( .A(n25900), .Y(n28090) );
  sky130_fd_sc_hd__clkinv_1 U15443 ( .A(n26050), .Y(n28119) );
  sky130_fd_sc_hd__clkinv_1 U15444 ( .A(n23518), .Y(n23519) );
  sky130_fd_sc_hd__and2_0 U15445 ( .A(n25344), .B(n11440), .X(n11443) );
  sky130_fd_sc_hd__clkinv_1 U15446 ( .A(n20632), .Y(n15737) );
  sky130_fd_sc_hd__clkinv_1 U15447 ( .A(n25993), .Y(n26155) );
  sky130_fd_sc_hd__inv_2 U15448 ( .A(n12185), .Y(n16273) );
  sky130_fd_sc_hd__and2_0 U15449 ( .A(n28751), .B(n29594), .X(n29220) );
  sky130_fd_sc_hd__clkinv_1 U15450 ( .A(n20633), .Y(n16942) );
  sky130_fd_sc_hd__clkinv_1 U15451 ( .A(n26251), .Y(n24579) );
  sky130_fd_sc_hd__clkinv_1 U15452 ( .A(n26115), .Y(n25026) );
  sky130_fd_sc_hd__clkinv_1 U15453 ( .A(n15703), .Y(n15726) );
  sky130_fd_sc_hd__clkinv_1 U15454 ( .A(n15586), .Y(n15588) );
  sky130_fd_sc_hd__clkinv_1 U15455 ( .A(n17276), .Y(n17285) );
  sky130_fd_sc_hd__clkinv_1 U15456 ( .A(n22965), .Y(n22850) );
  sky130_fd_sc_hd__clkinv_1 U15457 ( .A(n16951), .Y(n16952) );
  sky130_fd_sc_hd__inv_2 U15458 ( .A(n18635), .Y(n18762) );
  sky130_fd_sc_hd__clkinv_1 U15459 ( .A(n23860), .Y(n27955) );
  sky130_fd_sc_hd__clkinv_1 U15460 ( .A(n16035), .Y(n16036) );
  sky130_fd_sc_hd__clkinv_1 U15461 ( .A(n15493), .Y(n20693) );
  sky130_fd_sc_hd__clkinv_1 U15462 ( .A(n26167), .Y(n25948) );
  sky130_fd_sc_hd__clkinv_1 U15463 ( .A(n28086), .Y(n28249) );
  sky130_fd_sc_hd__clkinv_1 U15464 ( .A(n26225), .Y(n26214) );
  sky130_fd_sc_hd__clkinv_1 U15465 ( .A(n13577), .Y(n13578) );
  sky130_fd_sc_hd__clkinv_1 U15466 ( .A(n14943), .Y(n14945) );
  sky130_fd_sc_hd__clkinv_1 U15467 ( .A(n28633), .Y(n12) );
  sky130_fd_sc_hd__inv_1 U15468 ( .A(n23513), .Y(n23514) );
  sky130_fd_sc_hd__o2bb2ai_1 U15469 ( .B1(n23098), .B2(n23172), .A1_N(n23097), 
        .A2_N(n23174), .Y(n23099) );
  sky130_fd_sc_hd__clkinv_1 U15470 ( .A(n27164), .Y(n24475) );
  sky130_fd_sc_hd__and2_0 U15471 ( .A(n15870), .B(n15818), .X(n16119) );
  sky130_fd_sc_hd__clkinv_1 U15472 ( .A(n17047), .Y(n15790) );
  sky130_fd_sc_hd__clkinv_1 U15473 ( .A(n16202), .Y(n16161) );
  sky130_fd_sc_hd__clkinv_1 U15474 ( .A(n28199), .Y(n28157) );
  sky130_fd_sc_hd__clkinv_1 U15475 ( .A(n28751), .Y(n26184) );
  sky130_fd_sc_hd__clkinv_1 U15476 ( .A(n24695), .Y(n24693) );
  sky130_fd_sc_hd__clkinv_1 U15477 ( .A(n26173), .Y(n28234) );
  sky130_fd_sc_hd__clkinv_1 U15478 ( .A(n25982), .Y(n27039) );
  sky130_fd_sc_hd__clkinv_1 U15479 ( .A(n23022), .Y(n24783) );
  sky130_fd_sc_hd__clkinv_1 U15480 ( .A(n25614), .Y(n25609) );
  sky130_fd_sc_hd__inv_2 U15481 ( .A(n26323), .Y(n11153) );
  sky130_fd_sc_hd__clkinv_1 U15482 ( .A(n14941), .Y(n16055) );
  sky130_fd_sc_hd__clkinv_1 U15483 ( .A(n25582), .Y(n25572) );
  sky130_fd_sc_hd__clkinv_1 U15484 ( .A(n14929), .Y(n15857) );
  sky130_fd_sc_hd__clkinv_1 U15485 ( .A(n14894), .Y(n15786) );
  sky130_fd_sc_hd__inv_2 U15486 ( .A(n12185), .Y(n14744) );
  sky130_fd_sc_hd__o22ai_1 U15487 ( .A1(n18713), .A2(n18664), .B1(n18688), 
        .B2(n18716), .Y(n11789) );
  sky130_fd_sc_hd__clkinv_1 U15488 ( .A(n16964), .Y(n16924) );
  sky130_fd_sc_hd__clkinv_1 U15489 ( .A(n26242), .Y(n26246) );
  sky130_fd_sc_hd__clkinv_1 U15490 ( .A(n22877), .Y(n22957) );
  sky130_fd_sc_hd__clkinv_1 U15491 ( .A(n17045), .Y(n17051) );
  sky130_fd_sc_hd__clkinv_1 U15492 ( .A(n28026), .Y(n28023) );
  sky130_fd_sc_hd__clkinv_1 U15493 ( .A(n22875), .Y(n22958) );
  sky130_fd_sc_hd__clkinv_1 U15494 ( .A(n27660), .Y(n27655) );
  sky130_fd_sc_hd__clkinv_1 U15495 ( .A(n28063), .Y(n23321) );
  sky130_fd_sc_hd__clkinv_1 U15496 ( .A(n28066), .Y(n26114) );
  sky130_fd_sc_hd__clkinv_1 U15497 ( .A(n22712), .Y(n19404) );
  sky130_fd_sc_hd__clkinv_1 U15499 ( .A(n28221), .Y(n28126) );
  sky130_fd_sc_hd__clkinv_1 U15500 ( .A(n16029), .Y(n21009) );
  sky130_fd_sc_hd__clkinv_1 U15501 ( .A(n15869), .Y(n15850) );
  sky130_fd_sc_hd__clkinv_1 U15502 ( .A(n28097), .Y(n28099) );
  sky130_fd_sc_hd__clkinv_1 U15503 ( .A(n14918), .Y(n15837) );
  sky130_fd_sc_hd__clkinv_1 U15504 ( .A(n28601), .Y(n28954) );
  sky130_fd_sc_hd__o22ai_1 U15505 ( .A1(n18660), .A2(n18485), .B1(n18473), 
        .B2(n12991), .Y(n18501) );
  sky130_fd_sc_hd__inv_2 U15506 ( .A(n12163), .Y(n11154) );
  sky130_fd_sc_hd__inv_1 U15507 ( .A(n23495), .Y(n23496) );
  sky130_fd_sc_hd__clkinv_1 U15508 ( .A(n18867), .Y(n18869) );
  sky130_fd_sc_hd__clkinv_1 U15509 ( .A(n26243), .Y(n26128) );
  sky130_fd_sc_hd__clkinv_1 U15510 ( .A(n26456), .Y(n29054) );
  sky130_fd_sc_hd__inv_2 U15511 ( .A(n13986), .Y(n14414) );
  sky130_fd_sc_hd__clkinv_1 U15512 ( .A(n15855), .Y(n14858) );
  sky130_fd_sc_hd__clkinv_1 U15513 ( .A(n28228), .Y(n26040) );
  sky130_fd_sc_hd__or2_1 U15514 ( .A(n13638), .B(n23121), .X(n12174) );
  sky130_fd_sc_hd__clkinv_1 U15515 ( .A(n16180), .Y(n16181) );
  sky130_fd_sc_hd__nand3_1 U15516 ( .A(n18867), .B(n22055), .C(n17356), .Y(
        n18871) );
  sky130_fd_sc_hd__inv_2 U15518 ( .A(n14668), .Y(n11155) );
  sky130_fd_sc_hd__clkinv_1 U15519 ( .A(n17273), .Y(n17078) );
  sky130_fd_sc_hd__clkinv_1 U15520 ( .A(n25725), .Y(n29360) );
  sky130_fd_sc_hd__o211ai_1 U15521 ( .A1(j202_soc_core_intc_core_00_rg_ipr[46]), .A2(n25449), .B1(n19668), .C1(n19667), .Y(n19670) );
  sky130_fd_sc_hd__clkinv_1 U15522 ( .A(n29058), .Y(n26818) );
  sky130_fd_sc_hd__clkinv_1 U15523 ( .A(n15830), .Y(n17094) );
  sky130_fd_sc_hd__ha_1 U15524 ( .A(n17814), .B(n17813), .COUT(n17809), .SUM(
        n17816) );
  sky130_fd_sc_hd__clkinv_1 U15525 ( .A(n25985), .Y(n26165) );
  sky130_fd_sc_hd__clkinv_1 U15526 ( .A(n26141), .Y(n23466) );
  sky130_fd_sc_hd__clkinv_1 U15527 ( .A(n15870), .Y(n14873) );
  sky130_fd_sc_hd__clkinv_1 U15528 ( .A(n26127), .Y(n23441) );
  sky130_fd_sc_hd__clkinv_1 U15530 ( .A(n23509), .Y(n23510) );
  sky130_fd_sc_hd__clkinv_1 U15531 ( .A(n23554), .Y(n23560) );
  sky130_fd_sc_hd__clkinv_1 U15532 ( .A(n28614), .Y(n28955) );
  sky130_fd_sc_hd__clkinv_1 U15533 ( .A(n16611), .Y(n16919) );
  sky130_fd_sc_hd__clkinv_1 U15534 ( .A(n28232), .Y(n26185) );
  sky130_fd_sc_hd__o22ai_1 U15535 ( .A1(n17805), .A2(n17785), .B1(n24137), 
        .B2(n17802), .Y(n17807) );
  sky130_fd_sc_hd__clkinv_1 U15537 ( .A(n23596), .Y(n23192) );
  sky130_fd_sc_hd__clkinv_1 U15539 ( .A(n26202), .Y(n23546) );
  sky130_fd_sc_hd__inv_2 U15540 ( .A(n12186), .Y(n16448) );
  sky130_fd_sc_hd__clkinv_1 U15541 ( .A(n28597), .Y(n28959) );
  sky130_fd_sc_hd__o22ai_1 U15542 ( .A1(n18067), .A2(n17465), .B1(n17533), 
        .B2(n18068), .Y(n17535) );
  sky130_fd_sc_hd__clkinv_1 U15543 ( .A(n28230), .Y(n26252) );
  sky130_fd_sc_hd__clkinv_1 U15545 ( .A(n28602), .Y(n28952) );
  sky130_fd_sc_hd__or2_1 U15546 ( .A(n13638), .B(n23097), .X(n12187) );
  sky130_fd_sc_hd__clkinv_1 U15547 ( .A(n28607), .Y(n28927) );
  sky130_fd_sc_hd__clkinv_1 U15548 ( .A(n25891), .Y(n23468) );
  sky130_fd_sc_hd__clkinv_1 U15549 ( .A(n25890), .Y(n25906) );
  sky130_fd_sc_hd__clkinv_1 U15550 ( .A(n17067), .Y(n14857) );
  sky130_fd_sc_hd__clkinv_1 U15551 ( .A(n28496), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N33) );
  sky130_fd_sc_hd__o21a_1 U15552 ( .A1(n13572), .A2(n18868), .B1(n24285), .X(
        n13577) );
  sky130_fd_sc_hd__clkinv_1 U15553 ( .A(n13556), .Y(n13557) );
  sky130_fd_sc_hd__clkinv_1 U15554 ( .A(n25573), .Y(n25574) );
  sky130_fd_sc_hd__clkinv_1 U15555 ( .A(n28504), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N34) );
  sky130_fd_sc_hd__clkinv_1 U15556 ( .A(n19086), .Y(n17162) );
  sky130_fd_sc_hd__o22ai_1 U15557 ( .A1(n11514), .A2(n18341), .B1(n18719), 
        .B2(n18342), .Y(n18391) );
  sky130_fd_sc_hd__clkinv_1 U15558 ( .A(n24955), .Y(n24953) );
  sky130_fd_sc_hd__clkinv_1 U15559 ( .A(n28603), .Y(n28951) );
  sky130_fd_sc_hd__clkinv_1 U15560 ( .A(n20663), .Y(n20465) );
  sky130_fd_sc_hd__clkinv_1 U15561 ( .A(n28609), .Y(n28928) );
  sky130_fd_sc_hd__clkinv_1 U15562 ( .A(n28462), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N29) );
  sky130_fd_sc_hd__clkinv_1 U15563 ( .A(n28470), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N30) );
  sky130_fd_sc_hd__clkinv_1 U15564 ( .A(n27108), .Y(n27042) );
  sky130_fd_sc_hd__clkinv_1 U15565 ( .A(n13394), .Y(n13395) );
  sky130_fd_sc_hd__clkinv_1 U15566 ( .A(n28454), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N28) );
  sky130_fd_sc_hd__clkinv_1 U15567 ( .A(n28596), .Y(n28961) );
  sky130_fd_sc_hd__clkinv_1 U15568 ( .A(n29052), .Y(n25748) );
  sky130_fd_sc_hd__clkinv_1 U15569 ( .A(n28488), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N32) );
  sky130_fd_sc_hd__nand2b_1 U15570 ( .A_N(n25219), .B(n23252), .Y(n23255) );
  sky130_fd_sc_hd__clkinv_1 U15571 ( .A(n29057), .Y(n26481) );
  sky130_fd_sc_hd__clkinv_1 U15572 ( .A(n17281), .Y(n17329) );
  sky130_fd_sc_hd__clkinv_1 U15573 ( .A(n24469), .Y(n22026) );
  sky130_fd_sc_hd__clkinv_1 U15574 ( .A(n23323), .Y(n23324) );
  sky130_fd_sc_hd__clkinv_1 U15575 ( .A(n29037), .Y(n25279) );
  sky130_fd_sc_hd__clkinv_1 U15576 ( .A(n19163), .Y(n18922) );
  sky130_fd_sc_hd__clkinv_1 U15577 ( .A(n28231), .Y(n28089) );
  sky130_fd_sc_hd__clkinv_1 U15578 ( .A(n19661), .Y(n19662) );
  sky130_fd_sc_hd__clkinv_1 U15579 ( .A(n29038), .Y(n25353) );
  sky130_fd_sc_hd__clkinv_1 U15580 ( .A(n29068), .Y(n27197) );
  sky130_fd_sc_hd__clkinv_1 U15581 ( .A(n27351), .Y(n24022) );
  sky130_fd_sc_hd__clkinv_1 U15582 ( .A(n19380), .Y(n21170) );
  sky130_fd_sc_hd__clkinv_1 U15583 ( .A(n21915), .Y(n22714) );
  sky130_fd_sc_hd__clkinv_1 U15584 ( .A(n28969), .Y(n23691) );
  sky130_fd_sc_hd__clkinv_1 U15585 ( .A(n22033), .Y(n22867) );
  sky130_fd_sc_hd__clkinv_1 U15586 ( .A(n29042), .Y(n25440) );
  sky130_fd_sc_hd__clkinv_1 U15587 ( .A(n29041), .Y(n25433) );
  sky130_fd_sc_hd__clkinv_1 U15588 ( .A(n28598), .Y(n28958) );
  sky130_fd_sc_hd__or2_0 U15589 ( .A(n25231), .B(n25824), .X(n11460) );
  sky130_fd_sc_hd__clkinv_1 U15590 ( .A(n24241), .Y(n24235) );
  sky130_fd_sc_hd__clkinv_1 U15591 ( .A(n29039), .Y(n25361) );
  sky130_fd_sc_hd__clkinv_1 U15592 ( .A(n29040), .Y(n25367) );
  sky130_fd_sc_hd__o22ai_1 U15593 ( .A1(n18660), .A2(n18019), .B1(n17970), 
        .B2(n12991), .Y(n11668) );
  sky130_fd_sc_hd__clkinv_1 U15594 ( .A(n19124), .Y(n17300) );
  sky130_fd_sc_hd__clkinv_1 U15595 ( .A(n26494), .Y(n28934) );
  sky130_fd_sc_hd__clkinv_1 U15596 ( .A(n25427), .Y(n28935) );
  sky130_fd_sc_hd__clkinv_1 U15597 ( .A(n28604), .Y(n28936) );
  sky130_fd_sc_hd__clkinv_1 U15598 ( .A(n13436), .Y(n13431) );
  sky130_fd_sc_hd__clkinv_1 U15599 ( .A(n26254), .Y(n26119) );
  sky130_fd_sc_hd__clkinv_1 U15600 ( .A(n28605), .Y(n28937) );
  sky130_fd_sc_hd__clkinv_1 U15601 ( .A(n14863), .Y(n13389) );
  sky130_fd_sc_hd__clkinv_1 U15602 ( .A(n28600), .Y(n28956) );
  sky130_fd_sc_hd__clkinv_1 U15603 ( .A(n19765), .Y(n19766) );
  sky130_fd_sc_hd__clkinv_1 U15604 ( .A(n28608), .Y(n28939) );
  sky130_fd_sc_hd__clkinv_1 U15605 ( .A(n19762), .Y(n19763) );
  sky130_fd_sc_hd__clkinv_1 U15606 ( .A(n29051), .Y(n25685) );
  sky130_fd_sc_hd__clkinv_1 U15607 ( .A(n22858), .Y(n21847) );
  sky130_fd_sc_hd__clkinv_1 U15608 ( .A(n15704), .Y(n15439) );
  sky130_fd_sc_hd__clkinv_1 U15609 ( .A(n28599), .Y(n28940) );
  sky130_fd_sc_hd__clkinv_1 U15610 ( .A(n16176), .Y(n16160) );
  sky130_fd_sc_hd__clkinv_1 U15611 ( .A(n13553), .Y(n13536) );
  sky130_fd_sc_hd__clkinv_1 U15612 ( .A(n28610), .Y(n28941) );
  sky130_fd_sc_hd__clkinv_1 U15613 ( .A(n28611), .Y(n28942) );
  sky130_fd_sc_hd__clkinv_1 U15614 ( .A(n28612), .Y(n28943) );
  sky130_fd_sc_hd__clkinv_1 U15615 ( .A(n23326), .Y(n23328) );
  sky130_fd_sc_hd__clkinv_1 U15616 ( .A(n22824), .Y(n23292) );
  sky130_fd_sc_hd__clkinv_1 U15617 ( .A(n23322), .Y(n23332) );
  sky130_fd_sc_hd__clkinv_1 U15618 ( .A(n22318), .Y(n11158) );
  sky130_fd_sc_hd__clkinv_1 U15619 ( .A(n26783), .Y(n26605) );
  sky130_fd_sc_hd__clkinv_1 U15620 ( .A(n28613), .Y(n28944) );
  sky130_fd_sc_hd__clkinv_1 U15621 ( .A(n27037), .Y(n26130) );
  sky130_fd_sc_hd__clkinv_1 U15622 ( .A(n25203), .Y(n28953) );
  sky130_fd_sc_hd__clkinv_1 U15623 ( .A(n27081), .Y(n29055) );
  sky130_fd_sc_hd__clkinv_1 U15624 ( .A(n26314), .Y(n23777) );
  sky130_fd_sc_hd__clkinv_1 U15625 ( .A(n25649), .Y(n28949) );
  sky130_fd_sc_hd__clkinv_1 U15626 ( .A(n28432), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N25) );
  sky130_fd_sc_hd__clkinv_1 U15627 ( .A(n28034), .Y(n28626) );
  sky130_fd_sc_hd__clkinv_1 U15628 ( .A(n28424), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N24) );
  sky130_fd_sc_hd__clkinv_1 U15629 ( .A(n28414), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N23) );
  sky130_fd_sc_hd__clkinv_1 U15630 ( .A(n22039), .Y(n23302) );
  sky130_fd_sc_hd__clkinv_1 U15631 ( .A(n28407), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N22) );
  sky130_fd_sc_hd__clkinv_1 U15632 ( .A(n25972), .Y(n26154) );
  sky130_fd_sc_hd__clkinv_1 U15633 ( .A(n27095), .Y(n28929) );
  sky130_fd_sc_hd__clkinv_1 U15634 ( .A(n26959), .Y(n28930) );
  sky130_fd_sc_hd__clkinv_1 U15635 ( .A(n15428), .Y(n15426) );
  sky130_fd_sc_hd__clkinv_1 U15636 ( .A(n28021), .Y(n28024) );
  sky130_fd_sc_hd__clkinv_1 U15637 ( .A(n28399), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N21) );
  sky130_fd_sc_hd__clkinv_1 U15638 ( .A(n27028), .Y(n28933) );
  sky130_fd_sc_hd__clkinv_1 U15639 ( .A(n25097), .Y(n28931) );
  sky130_fd_sc_hd__clkinv_1 U15640 ( .A(n16162), .Y(n16163) );
  sky130_fd_sc_hd__clkinv_1 U15641 ( .A(n15584), .Y(n15616) );
  sky130_fd_sc_hd__clkinv_1 U15642 ( .A(n13417), .Y(n13401) );
  sky130_fd_sc_hd__clkinv_1 U15643 ( .A(n16616), .Y(n13468) );
  sky130_fd_sc_hd__clkinv_1 U15644 ( .A(n26312), .Y(n23762) );
  sky130_fd_sc_hd__clkinv_1 U15645 ( .A(n13794), .Y(n23094) );
  sky130_fd_sc_hd__and2_0 U15646 ( .A(n12142), .B(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .X(n20983) );
  sky130_fd_sc_hd__clkinv_1 U15647 ( .A(n25994), .Y(n25995) );
  sky130_fd_sc_hd__nor2_1 U15648 ( .A(j202_soc_core_j22_cpu_regop_Rn__3_), .B(
        n13635), .Y(n13627) );
  sky130_fd_sc_hd__clkinv_1 U15649 ( .A(n28056), .Y(n23318) );
  sky130_fd_sc_hd__clkinv_1 U15650 ( .A(n12577), .Y(n22531) );
  sky130_fd_sc_hd__and2_4 U15651 ( .A(n13706), .B(n19045), .X(n16012) );
  sky130_fd_sc_hd__clkinv_1 U15652 ( .A(n23281), .Y(n23282) );
  sky130_fd_sc_hd__clkinv_1 U15653 ( .A(n15838), .Y(n14937) );
  sky130_fd_sc_hd__and2_0 U15654 ( .A(n23545), .B(n12142), .X(n25010) );
  sky130_fd_sc_hd__clkinv_1 U15655 ( .A(n15673), .Y(n15422) );
  sky130_fd_sc_hd__clkinv_1 U15657 ( .A(n27651), .Y(n23316) );
  sky130_fd_sc_hd__clkinv_1 U15658 ( .A(n24969), .Y(n24011) );
  sky130_fd_sc_hd__clkinv_1 U15659 ( .A(n25085), .Y(n22408) );
  sky130_fd_sc_hd__clkinv_1 U15660 ( .A(n23668), .Y(n23648) );
  sky130_fd_sc_hd__clkinv_1 U15661 ( .A(n26198), .Y(n25012) );
  sky130_fd_sc_hd__clkinv_1 U15662 ( .A(n24818), .Y(n24811) );
  sky130_fd_sc_hd__clkinv_1 U15663 ( .A(n17021), .Y(n15831) );
  sky130_fd_sc_hd__buf_2 U15664 ( .A(n17358), .X(n18867) );
  sky130_fd_sc_hd__clkinv_1 U15665 ( .A(n27648), .Y(n27650) );
  sky130_fd_sc_hd__clkinv_1 U15666 ( .A(n17356), .Y(n13584) );
  sky130_fd_sc_hd__clkinv_1 U15667 ( .A(n23597), .Y(n22276) );
  sky130_fd_sc_hd__clkinv_1 U15668 ( .A(n26017), .Y(n28251) );
  sky130_fd_sc_hd__clkinv_1 U15669 ( .A(n18147), .Y(n21459) );
  sky130_fd_sc_hd__clkinv_1 U15670 ( .A(n29029), .Y(n24377) );
  sky130_fd_sc_hd__or2_1 U15671 ( .A(n13638), .B(n23171), .X(n12186) );
  sky130_fd_sc_hd__nor2b_1 U15672 ( .B_N(n18353), .A(n18370), .Y(n17536) );
  sky130_fd_sc_hd__clkinv_1 U15673 ( .A(n24376), .Y(n24379) );
  sky130_fd_sc_hd__clkinv_1 U15674 ( .A(n26781), .Y(n25834) );
  sky130_fd_sc_hd__clkinv_1 U15675 ( .A(n25961), .Y(n28100) );
  sky130_fd_sc_hd__clkinv_1 U15676 ( .A(n11912), .Y(n11909) );
  sky130_fd_sc_hd__clkinv_1 U15677 ( .A(n26049), .Y(n26052) );
  sky130_fd_sc_hd__inv_2 U15678 ( .A(n24132), .Y(n24137) );
  sky130_fd_sc_hd__or2_0 U15679 ( .A(j202_soc_core_j22_cpu_memop_MEM__0_), .B(
        n16054), .X(n13601) );
  sky130_fd_sc_hd__clkinv_1 U15680 ( .A(n15725), .Y(n15447) );
  sky130_fd_sc_hd__clkinv_1 U15681 ( .A(n24021), .Y(n24017) );
  sky130_fd_sc_hd__and4_1 U15682 ( .A(n13541), .B(n13540), .C(n13539), .D(
        n13538), .X(n13542) );
  sky130_fd_sc_hd__and2_0 U15683 ( .A(io_in[29]), .B(n12142), .X(n29143) );
  sky130_fd_sc_hd__and2_0 U15684 ( .A(io_in[30]), .B(n12142), .X(n29142) );
  sky130_fd_sc_hd__and2_0 U15685 ( .A(io_in[31]), .B(n12142), .X(n29141) );
  sky130_fd_sc_hd__and2_0 U15686 ( .A(io_in[32]), .B(n12142), .X(n29140) );
  sky130_fd_sc_hd__and2_0 U15687 ( .A(io_in[33]), .B(n12142), .X(n29139) );
  sky130_fd_sc_hd__and2_0 U15688 ( .A(io_in[34]), .B(n12142), .X(n29138) );
  sky130_fd_sc_hd__clkinv_1 U15689 ( .A(n23196), .Y(n14850) );
  sky130_fd_sc_hd__and2_0 U15690 ( .A(io_in[35]), .B(n12142), .X(n29137) );
  sky130_fd_sc_hd__o211ai_1 U15691 ( .A1(j202_soc_core_intc_core_00_rg_ipr[2]), 
        .A2(n27544), .B1(n19579), .C1(n19578), .Y(n19581) );
  sky130_fd_sc_hd__and2_0 U15692 ( .A(io_in[36]), .B(n12142), .X(n29136) );
  sky130_fd_sc_hd__clkinv_1 U15693 ( .A(n28243), .Y(n28079) );
  sky130_fd_sc_hd__clkinv_1 U15694 ( .A(n25980), .Y(n28229) );
  sky130_fd_sc_hd__clkinv_1 U15695 ( .A(n13385), .Y(n13451) );
  sky130_fd_sc_hd__and2_0 U15696 ( .A(n16706), .B(n17277), .X(n15309) );
  sky130_fd_sc_hd__clkinv_1 U15697 ( .A(n23194), .Y(n27905) );
  sky130_fd_sc_hd__clkinv_1 U15698 ( .A(n27908), .Y(n27911) );
  sky130_fd_sc_hd__clkinv_1 U15699 ( .A(n20149), .Y(n28915) );
  sky130_fd_sc_hd__clkinv_1 U15700 ( .A(n25954), .Y(n25920) );
  sky130_fd_sc_hd__clkinv_1 U15701 ( .A(n26188), .Y(n26039) );
  sky130_fd_sc_hd__and2_0 U15702 ( .A(n15838), .B(n17277), .X(n13294) );
  sky130_fd_sc_hd__clkinv_1 U15703 ( .A(n20548), .Y(n20273) );
  sky130_fd_sc_hd__clkinv_1 U15704 ( .A(n28019), .Y(n28016) );
  sky130_fd_sc_hd__clkinv_1 U15705 ( .A(n16054), .Y(n23299) );
  sky130_fd_sc_hd__clkinv_1 U15706 ( .A(n28775), .Y(n28003) );
  sky130_fd_sc_hd__mux2i_1 U15707 ( .A0(j202_soc_core_aquc_ADR__3_), .A1(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[3]), .S(n20149), 
        .Y(n25677) );
  sky130_fd_sc_hd__clkinv_1 U15708 ( .A(n18898), .Y(n18899) );
  sky130_fd_sc_hd__clkinv_1 U15709 ( .A(n26148), .Y(n25949) );
  sky130_fd_sc_hd__clkinv_1 U15710 ( .A(n24260), .Y(n23863) );
  sky130_fd_sc_hd__clkinv_1 U15711 ( .A(n14965), .Y(n17098) );
  sky130_fd_sc_hd__clkinv_1 U15712 ( .A(n13789), .Y(n13790) );
  sky130_fd_sc_hd__clkinv_1 U15713 ( .A(n26149), .Y(n28225) );
  sky130_fd_sc_hd__clkinv_1 U15714 ( .A(n19076), .Y(n21762) );
  sky130_fd_sc_hd__clkinv_1 U15715 ( .A(n25971), .Y(n25988) );
  sky130_fd_sc_hd__clkinv_1 U15716 ( .A(n24956), .Y(n24958) );
  sky130_fd_sc_hd__clkinv_1 U15717 ( .A(n15297), .Y(n15298) );
  sky130_fd_sc_hd__clkinv_1 U15718 ( .A(n19410), .Y(n19004) );
  sky130_fd_sc_hd__clkinv_1 U15719 ( .A(n28208), .Y(n25996) );
  sky130_fd_sc_hd__clkinv_1 U15720 ( .A(n19631), .Y(n19632) );
  sky130_fd_sc_hd__clkinv_1 U15721 ( .A(n13350), .Y(n13351) );
  sky130_fd_sc_hd__inv_2 U15722 ( .A(n12137), .Y(n17175) );
  sky130_fd_sc_hd__and2_0 U15723 ( .A(io_in[0]), .B(n12142), .X(n29152) );
  sky130_fd_sc_hd__and2_0 U15724 ( .A(io_in[1]), .B(n12142), .X(n29151) );
  sky130_fd_sc_hd__and2_0 U15725 ( .A(io_in[2]), .B(n12142), .X(n29150) );
  sky130_fd_sc_hd__clkinv_1 U15726 ( .A(n19534), .Y(n19504) );
  sky130_fd_sc_hd__and2_0 U15727 ( .A(io_in[3]), .B(n12142), .X(n29149) );
  sky130_fd_sc_hd__clkinv_1 U15728 ( .A(n13494), .Y(n13495) );
  sky130_fd_sc_hd__and2_0 U15729 ( .A(io_in[4]), .B(n12142), .X(n29148) );
  sky130_fd_sc_hd__and2_0 U15730 ( .A(io_in[7]), .B(n12142), .X(n29147) );
  sky130_fd_sc_hd__and2_0 U15731 ( .A(io_in[26]), .B(n12142), .X(n29146) );
  sky130_fd_sc_hd__clkinv_1 U15732 ( .A(n28560), .Y(n29087) );
  sky130_fd_sc_hd__and2_0 U15733 ( .A(io_in[27]), .B(n12142), .X(n29145) );
  sky130_fd_sc_hd__and2_0 U15734 ( .A(io_in[28]), .B(n12142), .X(n29144) );
  sky130_fd_sc_hd__and3_1 U15735 ( .A(n24774), .B(n26750), .C(n27910), .X(
        n13724) );
  sky130_fd_sc_hd__clkinv_1 U15736 ( .A(n29081), .Y(n28008) );
  sky130_fd_sc_hd__clkinv_1 U15737 ( .A(n27196), .Y(n27013) );
  sky130_fd_sc_hd__and2_0 U15738 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15]), .X(n29226) );
  sky130_fd_sc_hd__and2_0 U15739 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14]), .X(n29227) );
  sky130_fd_sc_hd__clkinv_1 U15740 ( .A(n13791), .Y(n13732) );
  sky130_fd_sc_hd__clkinv_1 U15741 ( .A(n17066), .Y(n14886) );
  sky130_fd_sc_hd__clkinv_1 U15742 ( .A(n26008), .Y(n28080) );
  sky130_fd_sc_hd__inv_2 U15743 ( .A(n12176), .Y(n15983) );
  sky130_fd_sc_hd__clkinv_1 U15744 ( .A(n25921), .Y(n26116) );
  sky130_fd_sc_hd__and2_0 U15745 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[12]), .X(n29084) );
  sky130_fd_sc_hd__and2_0 U15746 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[11]), .X(n29222) );
  sky130_fd_sc_hd__clkinv_1 U15747 ( .A(n19727), .Y(n19728) );
  sky130_fd_sc_hd__and2_0 U15748 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[10]), .X(n29228) );
  sky130_fd_sc_hd__and2_0 U15749 ( .A(n19354), .B(n17277), .X(n12181) );
  sky130_fd_sc_hd__clkinv_1 U15750 ( .A(n16706), .Y(n15432) );
  sky130_fd_sc_hd__and2_0 U15751 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[9]), .X(n29229) );
  sky130_fd_sc_hd__nand2_1 U15752 ( .A(n16706), .B(n20787), .Y(n16162) );
  sky130_fd_sc_hd__clkinv_1 U15753 ( .A(n23290), .Y(n23289) );
  sky130_fd_sc_hd__and2_0 U15755 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[2]), .X(n29225) );
  sky130_fd_sc_hd__and2_0 U15756 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]), .X(n29223) );
  sky130_fd_sc_hd__inv_2 U15757 ( .A(n12176), .Y(n15164) );
  sky130_fd_sc_hd__and2_0 U15758 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]), .X(n29230) );
  sky130_fd_sc_hd__and2_0 U15759 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]), .X(n29224) );
  sky130_fd_sc_hd__clkinv_1 U15760 ( .A(n20806), .Y(n17313) );
  sky130_fd_sc_hd__clkinv_1 U15761 ( .A(n25830), .Y(n25823) );
  sky130_fd_sc_hd__clkinv_1 U15762 ( .A(n25746), .Y(n25514) );
  sky130_fd_sc_hd__clkinv_1 U15763 ( .A(n23329), .Y(n23331) );
  sky130_fd_sc_hd__and2_0 U15764 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[23]), .X(n29085) );
  sky130_fd_sc_hd__clkinv_1 U15765 ( .A(n20547), .Y(n20549) );
  sky130_fd_sc_hd__clkinv_1 U15766 ( .A(j202_soc_core_uart_TOP_N24), .Y(n28781) );
  sky130_fd_sc_hd__clkinv_1 U15767 ( .A(n26147), .Y(n26152) );
  sky130_fd_sc_hd__clkinv_1 U15768 ( .A(n18659), .Y(n13201) );
  sky130_fd_sc_hd__clkinv_1 U15769 ( .A(n20991), .Y(n20992) );
  sky130_fd_sc_hd__clkinv_1 U15770 ( .A(n22715), .Y(n11161) );
  sky130_fd_sc_hd__clkinv_1 U15771 ( .A(n18915), .Y(n23297) );
  sky130_fd_sc_hd__clkinv_1 U15772 ( .A(n19072), .Y(n18914) );
  sky130_fd_sc_hd__buf_4 U15773 ( .A(n17403), .X(n18151) );
  sky130_fd_sc_hd__clkinv_1 U15774 ( .A(n26232), .Y(n26227) );
  sky130_fd_sc_hd__buf_4 U15775 ( .A(n17371), .X(n18750) );
  sky130_fd_sc_hd__clkinv_1 U15776 ( .A(n19025), .Y(n26747) );
  sky130_fd_sc_hd__clkinv_1 U15777 ( .A(n19575), .Y(n19576) );
  sky130_fd_sc_hd__clkinv_1 U15778 ( .A(n25916), .Y(n23473) );
  sky130_fd_sc_hd__clkinv_1 U15779 ( .A(n23336), .Y(n22508) );
  sky130_fd_sc_hd__clkinv_1 U15780 ( .A(n28236), .Y(n25003) );
  sky130_fd_sc_hd__clkinv_1 U15781 ( .A(n23927), .Y(n19007) );
  sky130_fd_sc_hd__buf_4 U15782 ( .A(n17939), .X(n18660) );
  sky130_fd_sc_hd__clkinv_1 U15784 ( .A(n27909), .Y(n14011) );
  sky130_fd_sc_hd__clkinv_1 U15785 ( .A(n27066), .Y(n28880) );
  sky130_fd_sc_hd__clkinv_1 U15786 ( .A(n20284), .Y(n21904) );
  sky130_fd_sc_hd__clkinv_1 U15787 ( .A(n28207), .Y(n28209) );
  sky130_fd_sc_hd__and2_0 U15788 ( .A(j202_soc_core_memory0_ram_dout0[507]), 
        .B(n21771), .X(n17106) );
  sky130_fd_sc_hd__clkinv_1 U15791 ( .A(n13503), .Y(n13504) );
  sky130_fd_sc_hd__clkinv_1 U15792 ( .A(n26782), .Y(n26776) );
  sky130_fd_sc_hd__clkinv_1 U15793 ( .A(n19003), .Y(n26738) );
  sky130_fd_sc_hd__inv_2 U15794 ( .A(n12136), .Y(n12137) );
  sky130_fd_sc_hd__clkinv_1 U15795 ( .A(n25951), .Y(n23471) );
  sky130_fd_sc_hd__xnor2_1 U15796 ( .A(j202_soc_core_j22_cpu_ml_bufa[32]), .B(
        n22487), .Y(n12303) );
  sky130_fd_sc_hd__and2_0 U15797 ( .A(n24317), .B(n24316), .X(n12301) );
  sky130_fd_sc_hd__inv_1 U15798 ( .A(n11716), .Y(n25231) );
  sky130_fd_sc_hd__clkinv_1 U15799 ( .A(n14752), .Y(n14156) );
  sky130_fd_sc_hd__clkinv_1 U15800 ( .A(n24960), .Y(n23649) );
  sky130_fd_sc_hd__clkinv_1 U15801 ( .A(n26046), .Y(n25926) );
  sky130_fd_sc_hd__clkinv_1 U15802 ( .A(n23283), .Y(n13545) );
  sky130_fd_sc_hd__clkinv_1 U15803 ( .A(n24429), .Y(n13560) );
  sky130_fd_sc_hd__clkinv_1 U15804 ( .A(n19714), .Y(n19716) );
  sky130_fd_sc_hd__clkinv_1 U15805 ( .A(n19054), .Y(n19051) );
  sky130_fd_sc_hd__inv_2 U15807 ( .A(n13638), .Y(n11163) );
  sky130_fd_sc_hd__clkinv_1 U15808 ( .A(n13687), .Y(n11884) );
  sky130_fd_sc_hd__clkinv_1 U15809 ( .A(n13688), .Y(n11883) );
  sky130_fd_sc_hd__clkinv_1 U15810 ( .A(n23536), .Y(n23544) );
  sky130_fd_sc_hd__clkinv_1 U15811 ( .A(n26749), .Y(n27912) );
  sky130_fd_sc_hd__clkinv_1 U15812 ( .A(n26682), .Y(n13651) );
  sky130_fd_sc_hd__inv_2 U15813 ( .A(n13666), .Y(n13681) );
  sky130_fd_sc_hd__and2_0 U15814 ( .A(n17289), .B(
        j202_soc_core_bootrom_00_address_w[11]), .X(n13293) );
  sky130_fd_sc_hd__clkinv_1 U15815 ( .A(n24572), .Y(n25112) );
  sky130_fd_sc_hd__inv_1 U15816 ( .A(n13624), .Y(n13636) );
  sky130_fd_sc_hd__clkinv_1 U15817 ( .A(n13677), .Y(n13678) );
  sky130_fd_sc_hd__clkinv_1 U15819 ( .A(n13547), .Y(n13546) );
  sky130_fd_sc_hd__clkinv_1 U15820 ( .A(n19516), .Y(n19518) );
  sky130_fd_sc_hd__clkinv_1 U15821 ( .A(n26398), .Y(n11713) );
  sky130_fd_sc_hd__clkinv_1 U15822 ( .A(n21771), .Y(n20830) );
  sky130_fd_sc_hd__nor2_1 U15823 ( .A(j202_soc_core_j22_cpu_regop_Rn__1_), .B(
        n13624), .Y(n13626) );
  sky130_fd_sc_hd__clkinv_1 U15824 ( .A(n24428), .Y(n23532) );
  sky130_fd_sc_hd__clkinv_1 U15825 ( .A(n25991), .Y(n25992) );
  sky130_fd_sc_hd__clkinv_1 U15826 ( .A(n23020), .Y(n23918) );
  sky130_fd_sc_hd__clkinv_1 U15827 ( .A(n23327), .Y(n13579) );
  sky130_fd_sc_hd__clkinv_1 U15828 ( .A(n21352), .Y(n21353) );
  sky130_fd_sc_hd__inv_1 U15829 ( .A(n12725), .Y(n22338) );
  sky130_fd_sc_hd__clkinv_1 U15830 ( .A(n24774), .Y(n24775) );
  sky130_fd_sc_hd__clkinv_1 U15831 ( .A(n28749), .Y(n25019) );
  sky130_fd_sc_hd__clkinv_1 U15832 ( .A(n25590), .Y(n25581) );
  sky130_fd_sc_hd__clkinv_1 U15833 ( .A(n19674), .Y(n19675) );
  sky130_fd_sc_hd__xor2_1 U15834 ( .A(n22052), .B(n22487), .X(n17369) );
  sky130_fd_sc_hd__clkinv_1 U15835 ( .A(j202_soc_core_intc_core_00_rg_ipr[53]), 
        .Y(n25375) );
  sky130_fd_sc_hd__clkinv_1 U15836 ( .A(j202_soc_core_intc_core_00_rg_itgt[86]), .Y(n25099) );
  sky130_fd_sc_hd__clkinv_1 U15837 ( .A(j202_soc_core_cmt_core_00_cnt1[1]), 
        .Y(n24938) );
  sky130_fd_sc_hd__clkinv_1 U15838 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]), .Y(n23341) );
  sky130_fd_sc_hd__clkinv_1 U15839 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[1]), 
        .Y(n23685) );
  sky130_fd_sc_hd__clkinv_1 U15840 ( .A(j202_soc_core_j22_cpu_rf_gpr[15]), .Y(
        n14647) );
  sky130_fd_sc_hd__clkinv_1 U15841 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[6]), .Y(n27549) );
  sky130_fd_sc_hd__clkinv_1 U15842 ( .A(j202_soc_core_intc_core_00_rg_itgt[87]), .Y(n27098) );
  sky130_fd_sc_hd__clkinv_1 U15843 ( .A(j202_soc_core_uart_sio_ce_x4), .Y(
        n28559) );
  sky130_fd_sc_hd__clkinv_1 U15844 ( .A(j202_soc_core_j22_cpu_rf_tmp[15]), .Y(
        n19066) );
  sky130_fd_sc_hd__clkinv_1 U15845 ( .A(j202_soc_core_uart_BRG_ps[6]), .Y(
        n28029) );
  sky130_fd_sc_hd__clkinv_1 U15846 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .Y(n17061) );
  sky130_fd_sc_hd__clkinv_1 U15847 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[5]), .Y(n26945) );
  sky130_fd_sc_hd__clkinv_1 U15848 ( .A(j202_soc_core_j22_cpu_opst[4]), .Y(
        n22275) );
  sky130_fd_sc_hd__clkinv_1 U15849 ( .A(j202_soc_core_j22_cpu_rf_vbr[30]), .Y(
        n22602) );
  sky130_fd_sc_hd__clkinv_1 U15850 ( .A(j202_soc_core_uart_BRG_ps[4]), .Y(
        n28022) );
  sky130_fd_sc_hd__inv_2 U15851 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), 
        .Y(n22055) );
  sky130_fd_sc_hd__clkinv_1 U15852 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[12]), .Y(n23396) );
  sky130_fd_sc_hd__clkinv_1 U15853 ( .A(j202_soc_core_intc_core_00_rg_ipr[55]), 
        .Y(n27020) );
  sky130_fd_sc_hd__clkinv_1 U15854 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[0]), 
        .Y(n23000) );
  sky130_fd_sc_hd__clkinv_1 U15855 ( .A(j202_soc_core_intc_core_00_rg_ipr[3]), 
        .Y(n24746) );
  sky130_fd_sc_hd__clkinv_1 U15856 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__2_), 
        .Y(n23534) );
  sky130_fd_sc_hd__clkinv_1 U15857 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[2]), .Y(n23656) );
  sky130_fd_sc_hd__clkinv_1 U15858 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[10]), .Y(n28345) );
  sky130_fd_sc_hd__clkinv_1 U15859 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[0]), .Y(n13518) );
  sky130_fd_sc_hd__clkinv_1 U15860 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[23]), .Y(n23618) );
  sky130_fd_sc_hd__clkinv_1 U15861 ( .A(j202_soc_core_cmt_core_00_cnt1[4]), 
        .Y(n25599) );
  sky130_fd_sc_hd__clkinv_1 U15862 ( .A(j202_soc_core_uart_BRG_br_clr), .Y(
        n28035) );
  sky130_fd_sc_hd__clkinv_1 U15863 ( .A(j202_soc_core_j22_cpu_opst[1]), .Y(
        n23195) );
  sky130_fd_sc_hd__clkinv_1 U15864 ( .A(j202_soc_core_qspi_wb_wdat[10]), .Y(
        n28339) );
  sky130_fd_sc_hd__clkinv_1 U15865 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[16]), .Y(n28700) );
  sky130_fd_sc_hd__clkinv_1 U15866 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[11]), .Y(n27237) );
  sky130_fd_sc_hd__clkinv_1 U15867 ( .A(j202_soc_core_cmt_core_00_cnt1[2]), 
        .Y(n24944) );
  sky130_fd_sc_hd__clkinv_1 U15868 ( .A(j202_soc_core_cmt_core_00_cnt1[8]), 
        .Y(n25613) );
  sky130_fd_sc_hd__clkinv_1 U15869 ( .A(j202_soc_core_cmt_core_00_cnt1[6]), 
        .Y(n25603) );
  sky130_fd_sc_hd__clkinv_1 U15870 ( .A(j202_soc_core_intc_core_00_rg_itgt[55]), .Y(n26961) );
  sky130_fd_sc_hd__clkinv_1 U15871 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .Y(n23432) );
  sky130_fd_sc_hd__clkinv_1 U15872 ( .A(j202_soc_core_intc_core_00_rg_ipr[7]), 
        .Y(n24745) );
  sky130_fd_sc_hd__clkinv_1 U15873 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[2]), .Y(n13576) );
  sky130_fd_sc_hd__clkinv_1 U15874 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .Y(n23470) );
  sky130_fd_sc_hd__clkinv_1 U15875 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[0]), .Y(n28127) );
  sky130_fd_sc_hd__clkinv_1 U15876 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[3]), .Y(n27834) );
  sky130_fd_sc_hd__clkinv_1 U15877 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[14]), .Y(n28694) );
  sky130_fd_sc_hd__clkinv_1 U15878 ( .A(j202_soc_core_memory0_ram_dout0[484]), 
        .Y(n21770) );
  sky130_fd_sc_hd__clkinv_1 U15879 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[5]), .Y(n28310) );
  sky130_fd_sc_hd__clkinv_1 U15880 ( .A(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[0]), .Y(n20155) );
  sky130_fd_sc_hd__clkinv_1 U15881 ( .A(j202_soc_core_j22_cpu_rf_pr[12]), .Y(
        n19495) );
  sky130_fd_sc_hd__clkinv_1 U15882 ( .A(j202_soc_core_bldc_core_00_pwm_en), 
        .Y(n28582) );
  sky130_fd_sc_hd__clkinv_1 U15883 ( .A(j202_soc_core_intc_core_00_rg_ipr[2]), 
        .Y(n24987) );
  sky130_fd_sc_hd__clkinv_1 U15884 ( .A(j202_soc_core_cmt_core_00_reg_addr[3]), 
        .Y(n24895) );
  sky130_fd_sc_hd__clkinv_1 U15885 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[9]), .Y(n23392) );
  sky130_fd_sc_hd__clkinv_1 U15886 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__1_), 
        .Y(n23494) );
  sky130_fd_sc_hd__clkinv_1 U15887 ( .A(j202_soc_core_j22_cpu_rf_gpr[510]), 
        .Y(n22603) );
  sky130_fd_sc_hd__clkinv_1 U15888 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[18]), .Y(n28400) );
  sky130_fd_sc_hd__clkinv_1 U15889 ( .A(j202_soc_core_j22_cpu_rf_tmp[12]), .Y(
        n19498) );
  sky130_fd_sc_hd__clkinv_1 U15890 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[17]), .Y(n28388) );
  sky130_fd_sc_hd__clkinv_1 U15891 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[22]), .Y(n23627) );
  sky130_fd_sc_hd__clkinv_1 U15892 ( .A(j202_soc_core_intc_core_00_rg_itgt[20]), .Y(n26486) );
  sky130_fd_sc_hd__clkinv_1 U15893 ( .A(j202_soc_core_ahb2apb_02_state[1]), 
        .Y(n24315) );
  sky130_fd_sc_hd__clkinv_1 U15894 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[122]), .Y(n27244) );
  sky130_fd_sc_hd__clkinv_1 U15895 ( .A(j202_soc_core_wbqspiflash_00_spi_wr), 
        .Y(n25880) );
  sky130_fd_sc_hd__clkinv_1 U15896 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[118]), .Y(n25651) );
  sky130_fd_sc_hd__clkinv_1 U15897 ( .A(j202_soc_core_cmt_core_00_cnt1[15]), 
        .Y(n27501) );
  sky130_fd_sc_hd__clkinv_1 U15898 ( .A(j202_soc_core_intc_core_00_rg_ipr[0]), 
        .Y(n24606) );
  sky130_fd_sc_hd__clkinv_1 U15899 ( .A(j202_soc_core_j22_cpu_regop_imm__7_), 
        .Y(n14363) );
  sky130_fd_sc_hd__clkinv_1 U15900 ( .A(j202_soc_core_bldc_core_00_comm[0]), 
        .Y(n28586) );
  sky130_fd_sc_hd__clkinv_1 U15901 ( .A(j202_soc_core_j22_cpu_regop_Wm__0_), 
        .Y(n24444) );
  sky130_fd_sc_hd__clkinv_1 U15902 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .Y(n23344) );
  sky130_fd_sc_hd__clkinv_1 U15903 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[7]), .Y(n23358) );
  sky130_fd_sc_hd__clkinv_1 U15904 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[1]), .Y(n24824) );
  sky130_fd_sc_hd__clkinv_1 U15905 ( .A(j202_soc_core_wbqspiflash_00_spif_req), 
        .Y(n26125) );
  sky130_fd_sc_hd__clkinv_1 U15906 ( .A(j202_soc_core_intc_core_00_rg_itgt[22]), .Y(n25860) );
  sky130_fd_sc_hd__clkinv_1 U15907 ( .A(j202_soc_core_qspi_wb_wdat[30]), .Y(
        n27109) );
  sky130_fd_sc_hd__clkinv_1 U15908 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16]), .Y(n28381) );
  sky130_fd_sc_hd__clkinv_1 U15909 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[3]), .Y(n24829) );
  sky130_fd_sc_hd__clkinv_1 U15910 ( .A(j202_soc_core_j22_cpu_ml_mach[31]), 
        .Y(n22464) );
  sky130_fd_sc_hd__clkinv_1 U15911 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[6]), .Y(n24833) );
  sky130_fd_sc_hd__clkinv_1 U15912 ( .A(
        j202_soc_core_intc_core_00_in_intreq[7]), .Y(n27309) );
  sky130_fd_sc_hd__clkinv_1 U15913 ( .A(j202_soc_core_j22_cpu_ml_macl[30]), 
        .Y(n22628) );
  sky130_fd_sc_hd__clkinv_1 U15914 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[10]), .Y(n28682) );
  sky130_fd_sc_hd__clkinv_1 U15916 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[9]), .Y(n23651) );
  sky130_fd_sc_hd__clkinv_1 U15917 ( .A(j202_soc_core_intc_core_00_rg_ipr[13]), 
        .Y(n25296) );
  sky130_fd_sc_hd__clkinv_1 U15918 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[8]), .Y(n24839) );
  sky130_fd_sc_hd__clkinv_1 U15919 ( .A(j202_soc_core_intc_core_00_rg_ipr[8]), 
        .Y(n25359) );
  sky130_fd_sc_hd__clkinv_1 U15920 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .Y(n26679) );
  sky130_fd_sc_hd__clkinv_1 U15921 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[24]), .Y(n28443) );
  sky130_fd_sc_hd__clkinv_1 U15922 ( .A(j202_soc_core_wbqspiflash_00_spi_in[9]), .Y(n28679) );
  sky130_fd_sc_hd__clkinv_1 U15923 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[6]), .Y(n23361) );
  sky130_fd_sc_hd__clkinv_1 U15924 ( .A(j202_soc_core_intr_vec__0_), .Y(n25452) );
  sky130_fd_sc_hd__clkinv_1 U15925 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[7]), .Y(n23650) );
  sky130_fd_sc_hd__clkinv_1 U15926 ( .A(j202_soc_core_j22_cpu_ml_macl[14]), 
        .Y(n23949) );
  sky130_fd_sc_hd__clkinv_1 U15927 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[4]), .Y(n28178) );
  sky130_fd_sc_hd__clkinv_1 U15928 ( .A(j202_soc_core_j22_cpu_rf_gbr[4]), .Y(
        n19452) );
  sky130_fd_sc_hd__clkinv_1 U15929 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[17]), .Y(n23626) );
  sky130_fd_sc_hd__clkinv_1 U15930 ( .A(j202_soc_core_uart_TOP_rx_fifo_wp[0]), 
        .Y(n27135) );
  sky130_fd_sc_hd__clkinv_1 U15931 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13]), .Y(n28359) );
  sky130_fd_sc_hd__clkinv_1 U15932 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[19]), .Y(n23630) );
  sky130_fd_sc_hd__clkinv_1 U15933 ( .A(j202_soc_core_j22_cpu_ml_macl[12]), 
        .Y(n23947) );
  sky130_fd_sc_hd__clkinv_1 U15934 ( .A(j202_soc_core_uart_TOP_rx_fifo_gb), 
        .Y(n23309) );
  sky130_fd_sc_hd__clkinv_1 U15935 ( .A(j202_soc_core_j22_cpu_macop_MAC_[4]), 
        .Y(n24293) );
  sky130_fd_sc_hd__clkinv_1 U15936 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[5]), .Y(n23371) );
  sky130_fd_sc_hd__clkinv_1 U15937 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[16]), .Y(n28383) );
  sky130_fd_sc_hd__clkinv_1 U15938 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[0]), 
        .Y(n28623) );
  sky130_fd_sc_hd__clkinv_1 U15939 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[3]), .Y(n28552) );
  sky130_fd_sc_hd__clkinv_1 U15940 ( .A(j202_soc_core_j22_cpu_rf_gpr[511]), 
        .Y(n22493) );
  sky130_fd_sc_hd__clkinv_1 U15941 ( .A(j202_soc_core_intr_vec__1_), .Y(n28511) );
  sky130_fd_sc_hd__clkinv_1 U15942 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[1]), .Y(n28512) );
  sky130_fd_sc_hd__clkinv_1 U15943 ( .A(j202_soc_core_intc_core_00_rg_ipr[54]), 
        .Y(n25503) );
  sky130_fd_sc_hd__clkinv_1 U15944 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[9]), .Y(n25619) );
  sky130_fd_sc_hd__clkinv_1 U15945 ( .A(j202_soc_core_intc_core_00_rg_ipr[23]), 
        .Y(n25432) );
  sky130_fd_sc_hd__clkinv_1 U15946 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[21]), .Y(n23622) );
  sky130_fd_sc_hd__clkinv_1 U15947 ( .A(j202_soc_core_intr_vec__2_), .Y(n28513) );
  sky130_fd_sc_hd__clkinv_1 U15948 ( .A(j202_soc_core_j22_cpu_rf_pr[14]), .Y(
        n21566) );
  sky130_fd_sc_hd__clkinv_1 U15949 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[7]), .Y(n28324) );
  sky130_fd_sc_hd__clkinv_1 U15950 ( .A(j202_soc_core_intc_core_00_rg_ie[11]), 
        .Y(n27015) );
  sky130_fd_sc_hd__clkinv_1 U15951 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[28]), .Y(n28475) );
  sky130_fd_sc_hd__clkinv_1 U15952 ( .A(j202_soc_core_intc_core_00_rg_ipr[9]), 
        .Y(n24030) );
  sky130_fd_sc_hd__clkinv_1 U15953 ( .A(j202_soc_core_wbqspiflash_00_spi_in[4]), .Y(n28664) );
  sky130_fd_sc_hd__clkinv_1 U15954 ( .A(j202_soc_core_qspi_wb_wdat[28]), .Y(
        n26466) );
  sky130_fd_sc_hd__clkinv_1 U15955 ( .A(j202_soc_core_uart_TOP_rx_fifo_wp[1]), 
        .Y(n27134) );
  sky130_fd_sc_hd__clkinv_1 U15956 ( .A(j202_soc_core_cmt_core_00_cnt1[14]), 
        .Y(n27495) );
  sky130_fd_sc_hd__clkinv_1 U15957 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[7]), .Y(n28200) );
  sky130_fd_sc_hd__clkinv_1 U15958 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[4]), .Y(n24832) );
  sky130_fd_sc_hd__clkinv_1 U15959 ( .A(j202_soc_core_j22_cpu_rf_vbr[31]), .Y(
        n22494) );
  sky130_fd_sc_hd__clkinv_1 U15960 ( .A(j202_soc_core_qspi_wb_addr[5]), .Y(
        n28113) );
  sky130_fd_sc_hd__clkinv_1 U15961 ( .A(j202_soc_core_wbqspiflash_00_spi_in[8]), .Y(n28676) );
  sky130_fd_sc_hd__clkinv_1 U15962 ( .A(j202_soc_core_intc_core_00_rg_ipr[14]), 
        .Y(n25533) );
  sky130_fd_sc_hd__clkinv_1 U15963 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[27]), .Y(n28471) );
  sky130_fd_sc_hd__clkinv_1 U15964 ( .A(j202_soc_core_intr_vec__3_), .Y(n28516) );
  sky130_fd_sc_hd__clkinv_1 U15965 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[1]), .Y(n28158) );
  sky130_fd_sc_hd__clkinv_1 U15966 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[119]), .Y(n27083) );
  sky130_fd_sc_hd__clkinv_1 U15967 ( .A(j202_soc_core_uart_TOP_dpll_state[1]), 
        .Y(n21784) );
  sky130_fd_sc_hd__clkinv_1 U15968 ( .A(j202_soc_core_cmt_core_00_cnt0[3]), 
        .Y(n25567) );
  sky130_fd_sc_hd__clkinv_1 U15969 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]), .Y(n28325) );
  sky130_fd_sc_hd__clkinv_1 U15970 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]), .Y(n23340) );
  sky130_fd_sc_hd__clkinv_1 U15971 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[2]), .Y(n28163) );
  sky130_fd_sc_hd__clkinv_1 U15972 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[6]), .Y(n28317) );
  sky130_fd_sc_hd__clkinv_1 U15973 ( .A(
        j202_soc_core_bldc_core_00_pwm_duty[10]), .Y(n26488) );
  sky130_fd_sc_hd__clkinv_1 U15974 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[11]), .Y(n28685) );
  sky130_fd_sc_hd__clkinv_1 U15975 ( .A(j202_soc_core_j22_cpu_rf_gpr[17]), .Y(
        n14751) );
  sky130_fd_sc_hd__clkinv_1 U15976 ( .A(j202_soc_core_j22_cpu_rf_tmp[17]), .Y(
        n14750) );
  sky130_fd_sc_hd__clkinv_1 U15977 ( .A(j202_soc_core_qspi_wb_wdat[24]), .Y(
        n25870) );
  sky130_fd_sc_hd__clkinv_1 U15978 ( .A(gpio_en_o[28]), .Y(n28480) );
  sky130_fd_sc_hd__clkinv_1 U15979 ( .A(j202_soc_core_intc_core_00_rg_itgt[81]), .Y(n27536) );
  sky130_fd_sc_hd__clkinv_1 U15980 ( .A(j202_soc_core_bldc_core_00_wdata[1]), 
        .Y(n27618) );
  sky130_fd_sc_hd__clkinv_1 U15981 ( .A(j202_soc_core_intc_core_00_rg_ipr[59]), 
        .Y(n25642) );
  sky130_fd_sc_hd__clkinv_1 U15982 ( .A(j202_soc_core_qspi_wb_wdat[20]), .Y(
        n27594) );
  sky130_fd_sc_hd__clkinv_1 U15983 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[10]), .Y(n27984) );
  sky130_fd_sc_hd__clkinv_1 U15984 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[10]), .Y(n27279) );
  sky130_fd_sc_hd__clkinv_1 U15985 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]), .Y(n23385) );
  sky130_fd_sc_hd__clkinv_1 U15986 ( .A(j202_soc_core_j22_cpu_rf_pr[3]), .Y(
        n21411) );
  sky130_fd_sc_hd__clkinv_1 U15987 ( .A(j202_soc_core_intc_core_00_rg_ipr[79]), 
        .Y(n27509) );
  sky130_fd_sc_hd__clkinv_1 U15988 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[106]), .Y(n27246) );
  sky130_fd_sc_hd__clkinv_1 U15989 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[22]), .Y(n28433) );
  sky130_fd_sc_hd__clkinv_1 U15990 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[11]), .Y(n27242) );
  sky130_fd_sc_hd__clkinv_1 U15991 ( .A(j202_soc_core_intc_core_00_rg_ipr[47]), 
        .Y(n25462) );
  sky130_fd_sc_hd__clkinv_1 U15992 ( .A(j202_soc_core_qspi_wb_addr[7]), .Y(
        n28122) );
  sky130_fd_sc_hd__clkinv_1 U15993 ( .A(j202_soc_core_wbqspiflash_00_spi_in[7]), .Y(n28673) );
  sky130_fd_sc_hd__clkinv_1 U15994 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[12]), .Y(n28688) );
  sky130_fd_sc_hd__clkinv_1 U15995 ( .A(j202_soc_core_j22_cpu_memop_Ma__1_), 
        .Y(n13649) );
  sky130_fd_sc_hd__clkinv_1 U15996 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[2]), .Y(n28289) );
  sky130_fd_sc_hd__clkinv_1 U15997 ( .A(j202_soc_core_intc_core_00_rg_ipr[107]), .Y(n28528) );
  sky130_fd_sc_hd__clkinv_1 U15998 ( .A(j202_soc_core_wbqspiflash_00_spi_busy), 
        .Y(n25944) );
  sky130_fd_sc_hd__clkinv_1 U15999 ( .A(j202_soc_core_intc_core_00_rg_ipr[65]), 
        .Y(n27665) );
  sky130_fd_sc_hd__clkinv_1 U16000 ( .A(j202_soc_core_intc_core_00_rg_ipr[74]), 
        .Y(n27283) );
  sky130_fd_sc_hd__clkinv_1 U16001 ( .A(j202_soc_core_qspi_wb_wdat[18]), .Y(
        n25256) );
  sky130_fd_sc_hd__clkinv_1 U16002 ( .A(j202_soc_core_bldc_core_00_pwm_duty[0]), .Y(n26275) );
  sky130_fd_sc_hd__clkinv_1 U16003 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .Y(n24230) );
  sky130_fd_sc_hd__clkinv_1 U16004 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[15]), .Y(n27503) );
  sky130_fd_sc_hd__clkinv_1 U16005 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[10]), .Y(n23390) );
  sky130_fd_sc_hd__inv_2 U16006 ( .A(j202_soc_core_j22_cpu_regop_Rn__2_), .Y(
        n13625) );
  sky130_fd_sc_hd__clkinv_1 U16007 ( .A(j202_soc_core_intc_core_00_rg_itgt[49]), .Y(n26933) );
  sky130_fd_sc_hd__clkinv_1 U16008 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[112]), .Y(n28522) );
  sky130_fd_sc_hd__clkinv_1 U16009 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[7]), .Y(n27326) );
  sky130_fd_sc_hd__clkinv_1 U16010 ( .A(j202_soc_core_j22_cpu_rf_tmp[2]), .Y(
        n19204) );
  sky130_fd_sc_hd__clkinv_1 U16011 ( .A(j202_soc_core_intc_core_00_rg_itgt[80]), .Y(n24978) );
  sky130_fd_sc_hd__clkinv_1 U16012 ( .A(j202_soc_core_cmt_core_00_cmf1), .Y(
        n27323) );
  sky130_fd_sc_hd__clkinv_1 U16013 ( .A(j202_soc_core_qspi_wb_wdat[11]), .Y(
        n28346) );
  sky130_fd_sc_hd__clkinv_1 U16014 ( .A(j202_soc_core_j22_cpu_regop_Rs__0_), 
        .Y(n13530) );
  sky130_fd_sc_hd__clkinv_1 U16015 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[4]), .Y(n24237) );
  sky130_fd_sc_hd__clkinv_1 U16016 ( .A(j202_soc_core_j22_cpu_rf_tmp[8]), .Y(
        n21997) );
  sky130_fd_sc_hd__clkinv_1 U16017 ( .A(j202_soc_core_bldc_core_00_pwm_duty[1]), .Y(n27804) );
  sky130_fd_sc_hd__clkinv_1 U16018 ( .A(j202_soc_core_j22_cpu_memop_MEM__1_), 
        .Y(n27268) );
  sky130_fd_sc_hd__clkinv_1 U16019 ( .A(j202_soc_core_bldc_core_00_pwm_duty[2]), .Y(n27704) );
  sky130_fd_sc_hd__clkinv_1 U16020 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .Y(n13574) );
  sky130_fd_sc_hd__clkinv_1 U16021 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[21]), .Y(n25392) );
  sky130_fd_sc_hd__clkinv_1 U16022 ( .A(
        j202_soc_core_intc_core_00_in_intreq[0]), .Y(n27765) );
  sky130_fd_sc_hd__clkinv_1 U16023 ( .A(j202_soc_core_intc_core_00_rg_ipr[35]), 
        .Y(n25484) );
  sky130_fd_sc_hd__clkinv_1 U16024 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[26]), .Y(n28463) );
  sky130_fd_sc_hd__clkinv_1 U16025 ( .A(j202_soc_core_intc_core_00_rg_ipr[70]), 
        .Y(n25521) );
  sky130_fd_sc_hd__clkinv_1 U16026 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[3]), .Y(n27846) );
  sky130_fd_sc_hd__clkinv_1 U16027 ( .A(j202_soc_core_bldc_core_00_pwm_duty[3]), .Y(n27508) );
  sky130_fd_sc_hd__clkinv_1 U16028 ( .A(j202_soc_core_intc_core_00_rg_itgt[98]), .Y(n27243) );
  sky130_fd_sc_hd__clkinv_1 U16029 ( .A(j202_soc_core_cmt_core_00_cnt0[2]), 
        .Y(n25562) );
  sky130_fd_sc_hd__clkinv_1 U16030 ( .A(j202_soc_core_intc_core_00_rg_ipr[34]), 
        .Y(n24967) );
  sky130_fd_sc_hd__clkinv_1 U16031 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]), .Y(n13575) );
  sky130_fd_sc_hd__clkinv_1 U16032 ( .A(j202_soc_core_j22_cpu_rf_gbr[1]), .Y(
        n22781) );
  sky130_fd_sc_hd__clkinv_1 U16033 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[20]), .Y(n27110) );
  sky130_fd_sc_hd__clkinv_1 U16034 ( .A(j202_soc_core_bldc_core_00_pwm_duty[4]), .Y(n27051) );
  sky130_fd_sc_hd__clkinv_1 U16035 ( .A(j202_soc_core_j22_cpu_rfuo_sr__s_), 
        .Y(n24273) );
  sky130_fd_sc_hd__clkinv_1 U16036 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[14]), .Y(n28373) );
  sky130_fd_sc_hd__clkinv_1 U16037 ( .A(j202_soc_core_intc_core_00_rg_ipr[67]), 
        .Y(n27989) );
  sky130_fd_sc_hd__clkinv_1 U16038 ( .A(j202_soc_core_bldc_core_00_pwm_duty[6]), .Y(n25258) );
  sky130_fd_sc_hd__clkinv_1 U16039 ( .A(j202_soc_core_qspi_wb_wdat[14]), .Y(
        n28367) );
  sky130_fd_sc_hd__clkinv_1 U16040 ( .A(j202_soc_core_j22_cpu_rf_tmp[11]), .Y(
        n21471) );
  sky130_fd_sc_hd__clkinv_1 U16041 ( .A(j202_soc_core_j22_cpu_rf_gpr[1]), .Y(
        n14000) );
  sky130_fd_sc_hd__clkinv_1 U16042 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[9]), .Y(n25624) );
  sky130_fd_sc_hd__clkinv_1 U16043 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[1]), .Y(n24886) );
  sky130_fd_sc_hd__clkinv_1 U16044 ( .A(j202_soc_core_bldc_core_00_pwm_duty[8]), .Y(n27578) );
  sky130_fd_sc_hd__clkinv_1 U16045 ( .A(j202_soc_core_rst), .Y(n28562) );
  sky130_fd_sc_hd__clkinv_1 U16046 ( .A(j202_soc_core_j22_cpu_rf_pr[11]), .Y(
        n21468) );
  sky130_fd_sc_hd__clkinv_1 U16047 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[14]), .Y(n28150) );
  sky130_fd_sc_hd__clkinv_1 U16048 ( .A(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[0]), .Y(n22600) );
  sky130_fd_sc_hd__clkinv_1 U16049 ( .A(j202_soc_core_intc_core_00_rg_ipr[71]), 
        .Y(n27313) );
  sky130_fd_sc_hd__clkinv_1 U16050 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[2]), .Y(n24966) );
  sky130_fd_sc_hd__clkinv_1 U16051 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[3]), .Y(n24116) );
  sky130_fd_sc_hd__clkinv_1 U16052 ( .A(j202_soc_core_j22_cpu_pc[1]), .Y(
        n22782) );
  sky130_fd_sc_hd__clkinv_1 U16053 ( .A(j202_soc_core_wbqspiflash_00_spi_in[6]), .Y(n28670) );
  sky130_fd_sc_hd__clkinv_1 U16054 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[6]), .Y(n11919) );
  sky130_fd_sc_hd__clkinv_1 U16055 ( .A(j202_soc_core_bldc_core_00_pwm_duty[9]), .Y(n25374) );
  sky130_fd_sc_hd__clkinv_1 U16056 ( .A(j202_soc_core_intc_core_00_rg_itgt[23]), .Y(n26458) );
  sky130_fd_sc_hd__clkinv_1 U16057 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[18]), .Y(n28180) );
  sky130_fd_sc_hd__clkinv_1 U16058 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[8]), .Y(n27145) );
  sky130_fd_sc_hd__clkinv_1 U16059 ( .A(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[2]), .Y(n24808) );
  sky130_fd_sc_hd__clkinv_1 U16060 ( .A(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .Y(n18864) );
  sky130_fd_sc_hd__clkinv_1 U16061 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[11]), .Y(n23398) );
  sky130_fd_sc_hd__clkinv_1 U16062 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[15]), .Y(n27111) );
  sky130_fd_sc_hd__clkinv_1 U16063 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[8]), .Y(n27150) );
  sky130_fd_sc_hd__clkinv_1 U16064 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[4]), .Y(n28298) );
  sky130_fd_sc_hd__clkinv_1 U16065 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]), .Y(n23346) );
  sky130_fd_sc_hd__clkinv_1 U16066 ( .A(j202_soc_core_intc_core_00_rg_ipr[51]), 
        .Y(n25672) );
  sky130_fd_sc_hd__clkinv_1 U16067 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]), .Y(n23425) );
  sky130_fd_sc_hd__clkinv_1 U16068 ( .A(j202_soc_core_j22_cpu_opst[3]), .Y(
        n23862) );
  sky130_fd_sc_hd__clkinv_1 U16069 ( .A(j202_soc_core_qspi_wb_wdat[15]), .Y(
        n28374) );
  sky130_fd_sc_hd__clkinv_1 U16070 ( .A(j202_soc_core_j22_cpu_opst[2]), .Y(
        n22024) );
  sky130_fd_sc_hd__clkinv_1 U16071 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]), .Y(n28290) );
  sky130_fd_sc_hd__clkinv_1 U16072 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[15]), .Y(n28380) );
  sky130_fd_sc_hd__clkinv_1 U16073 ( .A(j202_soc_core_j22_cpu_regop_Wm__3_), 
        .Y(n24442) );
  sky130_fd_sc_hd__clkinv_1 U16074 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[117]), .Y(n27030) );
  sky130_fd_sc_hd__clkinv_1 U16075 ( .A(j202_soc_core_qspi_wb_wdat[16]), .Y(
        n27062) );
  sky130_fd_sc_hd__clkinv_1 U16076 ( .A(j202_soc_core_wbqspiflash_00_spi_in[5]), .Y(n28667) );
  sky130_fd_sc_hd__clkinv_1 U16077 ( .A(j202_soc_core_intc_core_00_rg_itgt[85]), .Y(n26496) );
  sky130_fd_sc_hd__clkinv_1 U16078 ( .A(j202_soc_core_j22_cpu_regop_Wm__2_), 
        .Y(n24433) );
  sky130_fd_sc_hd__clkinv_1 U16079 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[15]), .Y(n23349) );
  sky130_fd_sc_hd__clkbuf_1 U16080 ( .A(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[4]), .X(n13571) );
  sky130_fd_sc_hd__clkinv_1 U16081 ( .A(gpio_en_o[20]), .Y(n28417) );
  sky130_fd_sc_hd__clkinv_1 U16082 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[4]), .Y(n23374) );
  sky130_fd_sc_hd__clkinv_1 U16083 ( .A(j202_soc_core_intc_core_00_rg_itgt[53]), .Y(n25383) );
  sky130_fd_sc_hd__clkinv_1 U16084 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[24]), .Y(n23617) );
  sky130_fd_sc_hd__clkinv_1 U16085 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[20]), .Y(n28415) );
  sky130_fd_sc_hd__clkinv_1 U16086 ( .A(
        j202_soc_core_bldc_core_00_pwm_duty[11]), .Y(n24571) );
  sky130_fd_sc_hd__clkinv_1 U16087 ( .A(j202_soc_core_uart_BRG_ps[2]), .Y(
        n28015) );
  sky130_fd_sc_hd__clkinv_1 U16088 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]), .Y(n28282) );
  sky130_fd_sc_hd__clkinv_1 U16089 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__0_), 
        .Y(n23499) );
  sky130_fd_sc_hd__clkinv_1 U16090 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[31]), .Y(n28505) );
  sky130_fd_sc_hd__clkinv_1 U16091 ( .A(j202_soc_core_bldc_core_00_wdata[0]), 
        .Y(n27741) );
  sky130_fd_sc_hd__clkinv_1 U16092 ( .A(j202_soc_core_j22_cpu_regop_Wm__1_), 
        .Y(n24441) );
  sky130_fd_sc_hd__clkinv_1 U16093 ( .A(j202_soc_core_uart_BRG_ps_clr), .Y(
        n28012) );
  sky130_fd_sc_hd__clkinv_1 U16094 ( .A(j202_soc_core_intc_core_00_rg_itgt[84]), .Y(n28537) );
  sky130_fd_sc_hd__clkinv_1 U16095 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[15]), .Y(n28697) );
  sky130_fd_sc_hd__clkinv_1 U16096 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[16]), .Y(n28165) );
  sky130_fd_sc_hd__clkinv_1 U16097 ( .A(j202_soc_core_qspi_wb_wdat[17]), .Y(
        n28389) );
  sky130_fd_sc_hd__buf_4 U16098 ( .A(j202_soc_core_j22_cpu_ml_bufb[1]), .X(
        n18367) );
  sky130_fd_sc_hd__clkinv_1 U16099 ( .A(
        j202_soc_core_bldc_core_00_hall_value[0]), .Y(n27726) );
  sky130_fd_sc_hd__clkinv_1 U16100 ( .A(j202_soc_core_cmt_core_00_cnt1[12]), 
        .Y(n26305) );
  sky130_fd_sc_hd__clkinv_1 U16101 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[13]), .Y(n23383) );
  sky130_fd_sc_hd__clkinv_1 U16102 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[4]), .Y(n26992) );
  sky130_fd_sc_hd__clkinv_1 U16103 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[31]), .Y(n28503) );
  sky130_fd_sc_hd__clkinv_1 U16104 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[8]), .Y(n23352) );
  sky130_fd_sc_hd__clkinv_1 U16105 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__0_), 
        .Y(n23505) );
  sky130_fd_sc_hd__clkinv_1 U16106 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[14]), .Y(n27699) );
  sky130_fd_sc_hd__clkinv_1 U16107 ( .A(j202_soc_core_j22_cpu_rf_tmp[5]), .Y(
        n21860) );
  sky130_fd_sc_hd__clkinv_1 U16108 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[115]), .Y(n27512) );
  sky130_fd_sc_hd__clkinv_1 U16109 ( .A(j202_soc_core_intc_core_00_rg_ipr[57]), 
        .Y(n25195) );
  sky130_fd_sc_hd__or2_0 U16110 ( .A(start_n_reg[0]), .B(wb_rst_i), .X(n4) );
  sky130_fd_sc_hd__clkinv_1 U16111 ( .A(j202_soc_core_qspi_wb_wdat[1]), .Y(
        n28273) );
  sky130_fd_sc_hd__clkinv_1 U16112 ( .A(j202_soc_core_j22_cpu_rf_pr[15]), .Y(
        n19064) );
  sky130_fd_sc_hd__clkinv_1 U16113 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[21]), .Y(n28423) );
  sky130_fd_sc_hd__clkinv_1 U16114 ( .A(j202_soc_core_uart_TOP_dpll_state[0]), 
        .Y(n28556) );
  sky130_fd_sc_hd__clkinv_1 U16115 ( .A(j202_soc_core_j22_cpu_rf_gbr[0]), .Y(
        n21951) );
  sky130_fd_sc_hd__clkinv_1 U16116 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[30]), .Y(n28497) );
  sky130_fd_sc_hd__clkinv_1 U16117 ( .A(j202_soc_core_intr_level__4_), .Y(
        n23284) );
  sky130_fd_sc_hd__clkinv_1 U16118 ( .A(j202_soc_core_intc_core_00_rg_itgt[83]), .Y(n27708) );
  sky130_fd_sc_hd__clkinv_1 U16119 ( .A(j202_soc_core_qspi_wb_wdat[23]), .Y(
        n24574) );
  sky130_fd_sc_hd__clkinv_1 U16120 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[5]), .Y(n26930) );
  sky130_fd_sc_hd__clkinv_1 U16121 ( .A(j202_soc_core_j22_cpu_memop_MEM__3_), 
        .Y(n24280) );
  sky130_fd_sc_hd__clkinv_1 U16122 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .Y(n23418) );
  sky130_fd_sc_hd__clkinv_1 U16123 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[0]), .Y(n27742) );
  sky130_fd_sc_hd__clkinv_1 U16124 ( .A(j202_soc_core_cmt_core_00_cnt1[0]), 
        .Y(n24939) );
  sky130_fd_sc_hd__clkinv_1 U16125 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[13]), .Y(n27799) );
  sky130_fd_sc_hd__inv_2 U16126 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]), 
        .Y(n13570) );
  sky130_fd_sc_hd__clkinv_1 U16127 ( .A(j202_soc_core_intc_core_00_rg_itgt[82]), .Y(n27286) );
  sky130_fd_sc_hd__clkinv_1 U16128 ( .A(j202_soc_core_j22_cpu_rf_tmp[10]), .Y(
        n19216) );
  sky130_fd_sc_hd__clkinv_1 U16129 ( .A(j202_soc_core_intc_core_00_rg_ipr[56]), 
        .Y(n25854) );
  sky130_fd_sc_hd__clkinv_1 U16130 ( .A(j202_soc_core_j22_cpu_rf_gbr[7]), .Y(
        n19047) );
  sky130_fd_sc_hd__clkinv_1 U16131 ( .A(j202_soc_core_j22_cpu_rf_gbr[9]), .Y(
        n22859) );
  sky130_fd_sc_hd__clkinv_1 U16132 ( .A(j202_soc_core_j22_cpu_rf_pr[10]), .Y(
        n19214) );
  sky130_fd_sc_hd__clkinv_1 U16133 ( .A(j202_soc_core_qspi_wb_wdat[21]), .Y(
        n25391) );
  sky130_fd_sc_hd__clkinv_1 U16134 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[21]), .Y(n28425) );
  sky130_fd_sc_hd__clkinv_1 U16135 ( .A(j202_soc_core_intc_core_00_rg_ipr[64]), 
        .Y(n19521) );
  sky130_fd_sc_hd__clkinv_1 U16136 ( .A(j202_soc_core_j22_cpu_rfuo_sr__m_), 
        .Y(n22857) );
  sky130_fd_sc_hd__clkinv_1 U16137 ( .A(j202_soc_core_j22_cpu_rf_gpr[0]), .Y(
        n21955) );
  sky130_fd_sc_hd__clkinv_1 U16138 ( .A(
        j202_soc_core_bldc_core_00_hall_value[1]), .Y(n27607) );
  sky130_fd_sc_hd__clkinv_1 U16139 ( .A(j202_soc_core_intc_core_00_rg_ipr[58]), 
        .Y(n25087) );
  sky130_fd_sc_hd__clkinv_1 U16140 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[29]), .Y(n28489) );
  sky130_fd_sc_hd__clkinv_1 U16141 ( .A(j202_soc_core_j22_cpu_memop_Ma__0_), 
        .Y(n13656) );
  sky130_fd_sc_hd__clkinv_1 U16142 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[13]), .Y(n28691) );
  sky130_fd_sc_hd__clkinv_1 U16143 ( .A(j202_soc_core_j22_cpu_rf_pr[0]), .Y(
        n21950) );
  sky130_fd_sc_hd__clkinv_1 U16144 ( .A(j202_soc_core_j22_cpu_rf_gpr[9]), .Y(
        n14541) );
  sky130_fd_sc_hd__clkinv_1 U16145 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[6]), .Y(n27533) );
  sky130_fd_sc_hd__clkinv_1 U16146 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[11]), .Y(n28352) );
  sky130_fd_sc_hd__clkinv_1 U16147 ( .A(j202_soc_core_uart_BRG_br_cnt[2]), .Y(
        n28040) );
  sky130_fd_sc_hd__clkinv_1 U16148 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__3_), 
        .Y(n23507) );
  sky130_fd_sc_hd__clkinv_1 U16149 ( .A(j202_soc_core_intc_core_00_rg_ipr[75]), 
        .Y(n25535) );
  sky130_fd_sc_hd__clkinv_1 U16150 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__2_), 
        .Y(n13559) );
  sky130_fd_sc_hd__clkinv_1 U16151 ( .A(j202_soc_core_uart_BRG_br_cnt[4]), .Y(
        n28043) );
  sky130_fd_sc_hd__clkinv_1 U16152 ( .A(j202_soc_core_j22_cpu_rf_tmp[0]), .Y(
        n21954) );
  sky130_fd_sc_hd__clkinv_1 U16153 ( .A(j202_soc_core_wbqspiflash_00_state[1]), 
        .Y(n25984) );
  sky130_fd_sc_hd__clkinv_1 U16154 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[113]), .Y(n27304) );
  sky130_fd_sc_hd__clkinv_1 U16155 ( .A(j202_soc_core_uart_BRG_br_cnt[6]), .Y(
        n28036) );
  sky130_fd_sc_hd__clkinv_1 U16156 ( .A(j202_soc_core_intc_core_00_rg_ipr[63]), 
        .Y(n25501) );
  sky130_fd_sc_hd__clkinv_1 U16157 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[7]), .Y(n27332) );
  sky130_fd_sc_hd__clkinv_1 U16158 ( .A(j202_soc_core_qspi_wb_wdat[27]), .Y(
        n25659) );
  sky130_fd_sc_hd__clkinv_1 U16159 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]), .Y(n24240) );
  sky130_fd_sc_hd__clkinv_1 U16160 ( .A(j202_soc_core_j22_cpu_pc[0]), .Y(
        n23720) );
  sky130_fd_sc_hd__clkinv_1 U16161 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]), .Y(n23411) );
  sky130_fd_sc_hd__clkinv_1 U16162 ( .A(wbs_dat_o[0]), .Y(n10487) );
  sky130_fd_sc_hd__clkinv_1 U16163 ( .A(j202_soc_core_j22_cpu_pc[20]), .Y(
        n13720) );
  sky130_fd_sc_hd__clkinv_1 U16164 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .Y(n23469) );
  sky130_fd_sc_hd__clkinv_1 U16165 ( .A(j202_soc_core_pwrite[2]), .Y(n27649)
         );
  sky130_fd_sc_hd__clkinv_1 U16166 ( .A(j202_soc_core_j22_cpu_ml_mach[2]), .Y(
        n17429) );
  sky130_fd_sc_hd__clkinv_1 U16167 ( .A(j202_soc_core_intc_core_00_bs_addr[7]), 
        .Y(n24751) );
  sky130_fd_sc_hd__clkinv_1 U16168 ( .A(j202_soc_core_intc_core_00_rg_ie[19]), 
        .Y(n25689) );
  sky130_fd_sc_hd__clkinv_1 U16169 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[9]), .Y(n28338) );
  sky130_fd_sc_hd__clkinv_1 U16170 ( .A(j202_soc_core_aquc_ADR__0_), .Y(n13453) );
  sky130_fd_sc_hd__buf_4 U16171 ( .A(j202_soc_core_j22_cpu_ml_bufa[27]), .X(
        n22685) );
  sky130_fd_sc_hd__clkinv_1 U16172 ( .A(j202_soc_core_intc_core_00_rg_ipr[66]), 
        .Y(n24968) );
  sky130_fd_sc_hd__clkinv_1 U16173 ( .A(j202_soc_core_intc_core_00_bs_addr[5]), 
        .Y(n28892) );
  sky130_fd_sc_hd__clkinv_1 U16174 ( .A(j202_soc_core_intc_core_00_rg_ipr[68]), 
        .Y(n24599) );
  sky130_fd_sc_hd__clkinv_1 U16175 ( .A(j202_soc_core_intc_core_00_rg_ipr[72]), 
        .Y(n27151) );
  sky130_fd_sc_hd__clkinv_1 U16176 ( .A(j202_soc_core_gpio_core_00_reg_addr[4]), .Y(n23453) );
  sky130_fd_sc_hd__clkinv_1 U16177 ( .A(j202_soc_core_intc_core_00_rg_itgt[72]), .Y(n24981) );
  sky130_fd_sc_hd__clkinv_1 U16178 ( .A(j202_soc_core_wbqspiflash_00_spi_in[2]), .Y(n28658) );
  sky130_fd_sc_hd__clkinv_1 U16179 ( .A(j202_soc_core_intc_core_00_rg_itgt[15]), .Y(n25492) );
  sky130_fd_sc_hd__clkinv_1 U16180 ( .A(j202_soc_core_memory0_ram_dout0_sel[1]), .Y(n13375) );
  sky130_fd_sc_hd__clkinv_1 U16181 ( .A(j202_soc_core_intc_core_00_rg_itgt[14]), .Y(n25493) );
  sky130_fd_sc_hd__clkinv_1 U16182 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[0]), .Y(n23619) );
  sky130_fd_sc_hd__clkinv_1 U16183 ( .A(j202_soc_core_gpio_core_00_reg_addr[2]), .Y(n23452) );
  sky130_fd_sc_hd__clkinv_1 U16184 ( .A(j202_soc_core_intc_core_00_rg_ie[25]), 
        .Y(n25202) );
  sky130_fd_sc_hd__clkinv_1 U16185 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .Y(n23455) );
  sky130_fd_sc_hd__clkinv_1 U16186 ( .A(j202_soc_core_bldc_core_00_comm[2]), 
        .Y(n22996) );
  sky130_fd_sc_hd__clkinv_1 U16187 ( .A(j202_soc_core_aquc_ADR__2_), .Y(n20157) );
  sky130_fd_sc_hd__clkinv_1 U16188 ( .A(j202_soc_core_intc_core_00_rg_ipr[80]), 
        .Y(n24600) );
  sky130_fd_sc_hd__clkinv_1 U16189 ( .A(j202_soc_core_intc_core_00_rg_itgt[12]), .Y(n25510) );
  sky130_fd_sc_hd__clkinv_1 U16190 ( .A(j202_soc_core_intc_core_00_rg_ipr[37]), 
        .Y(n25479) );
  sky130_fd_sc_hd__clkinv_1 U16191 ( .A(j202_soc_core_intc_core_00_rg_ipr[82]), 
        .Y(n25522) );
  sky130_fd_sc_hd__clkinv_1 U16192 ( .A(j202_soc_core_intc_core_00_bs_addr[8]), 
        .Y(n24756) );
  sky130_fd_sc_hd__clkinv_1 U16193 ( .A(j202_soc_core_intc_core_00_rg_itgt[10]), .Y(n25458) );
  sky130_fd_sc_hd__clkinv_1 U16194 ( .A(j202_soc_core_j22_cpu_rf_gpr[4]), .Y(
        n19457) );
  sky130_fd_sc_hd__clkinv_1 U16195 ( .A(j202_soc_core_intc_core_00_rg_ie[16]), 
        .Y(n25767) );
  sky130_fd_sc_hd__clkinv_1 U16196 ( .A(j202_soc_core_intc_core_00_rg_ipr[127]), .Y(n27078) );
  sky130_fd_sc_hd__clkinv_1 U16197 ( .A(j202_soc_core_intc_core_00_rg_ipr[84]), 
        .Y(n27579) );
  sky130_fd_sc_hd__clkinv_1 U16198 ( .A(j202_soc_core_intc_core_00_rg_itgt[8]), 
        .Y(n25472) );
  sky130_fd_sc_hd__and2_0 U16199 ( .A(j202_soc_core_j22_cpu_ml_bufb[31]), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .X(n27350) );
  sky130_fd_sc_hd__clkinv_1 U16200 ( .A(j202_soc_core_intc_core_00_rg_ipr[85]), 
        .Y(n25376) );
  sky130_fd_sc_hd__clkinv_1 U16201 ( .A(j202_soc_core_j22_cpu_rf_tmp[4]), .Y(
        n19456) );
  sky130_fd_sc_hd__clkinv_1 U16202 ( .A(j202_soc_core_intc_core_00_rg_itgt[13]), .Y(n25511) );
  sky130_fd_sc_hd__clkinv_1 U16203 ( .A(j202_soc_core_j22_cpu_macop_MAC_[2]), 
        .Y(n27338) );
  sky130_fd_sc_hd__clkinv_1 U16204 ( .A(j202_soc_core_gpio_core_00_reg_addr[3]), .Y(n27659) );
  sky130_fd_sc_hd__clkinv_1 U16205 ( .A(j202_soc_core_intc_core_00_rg_ipr[86]), 
        .Y(n26498) );
  sky130_fd_sc_hd__clkinv_1 U16206 ( .A(j202_soc_core_intc_core_00_rg_itgt[11]), .Y(n27009) );
  sky130_fd_sc_hd__clkinv_1 U16207 ( .A(j202_soc_core_j22_cpu_macop_MAC_[3]), 
        .Y(n24278) );
  sky130_fd_sc_hd__clkinv_1 U16208 ( .A(j202_soc_core_intc_core_00_rg_itgt[9]), 
        .Y(n25465) );
  sky130_fd_sc_hd__clkinv_1 U16209 ( .A(j202_soc_core_intc_core_00_rg_ipr[89]), 
        .Y(n25197) );
  sky130_fd_sc_hd__clkinv_1 U16210 ( .A(j202_soc_core_intc_core_00_rg_ipr[87]), 
        .Y(n27022) );
  sky130_fd_sc_hd__clkinv_1 U16211 ( .A(j202_soc_core_j22_cpu_ml_mach[26]), 
        .Y(n22384) );
  sky130_fd_sc_hd__clkinv_1 U16212 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[17]), .Y(n25740) );
  sky130_fd_sc_hd__clkinv_1 U16213 ( .A(
        j202_soc_core_wbqspiflash_00_w_qspi_sck), .Y(n28635) );
  sky130_fd_sc_hd__clkinv_1 U16214 ( .A(j202_soc_core_intc_core_00_rg_ie[13]), 
        .Y(n25516) );
  sky130_fd_sc_hd__clkinv_1 U16215 ( .A(j202_soc_core_uart_TOP_load), .Y(
        n28001) );
  sky130_fd_sc_hd__clkinv_1 U16216 ( .A(j202_soc_core_memory0_ram_dout0_sel[5]), .Y(n13372) );
  sky130_fd_sc_hd__clkinv_1 U16217 ( .A(j202_soc_core_intc_core_00_rg_ipr[121]), .Y(n25200) );
  sky130_fd_sc_hd__clkinv_1 U16218 ( .A(j202_soc_core_intc_core_00_rg_ipr[126]), .Y(n27092) );
  sky130_fd_sc_hd__clkinv_1 U16219 ( .A(j202_soc_core_intc_core_00_rg_ipr[83]), 
        .Y(n25536) );
  sky130_fd_sc_hd__clkinv_1 U16220 ( .A(j202_soc_core_j22_cpu_ml_macl[7]), .Y(
        n19008) );
  sky130_fd_sc_hd__clkinv_1 U16221 ( .A(j202_soc_core_j22_cpu_ml_mach[3]), .Y(
        n17455) );
  sky130_fd_sc_hd__clkinv_1 U16222 ( .A(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[0]), .Y(n23643) );
  sky130_fd_sc_hd__clkinv_1 U16223 ( .A(j202_soc_core_intc_core_00_rg_ipr[115]), .Y(n25675) );
  sky130_fd_sc_hd__clkinv_1 U16224 ( .A(j202_soc_core_intc_core_00_rg_ipr[125]), .Y(n26956) );
  sky130_fd_sc_hd__clkinv_1 U16225 ( .A(j202_soc_core_j22_cpu_ml_mach[23]), 
        .Y(n22049) );
  sky130_fd_sc_hd__clkinv_1 U16226 ( .A(j202_soc_core_j22_cpu_rf_pr[4]), .Y(
        n19450) );
  sky130_fd_sc_hd__clkinv_1 U16227 ( .A(j202_soc_core_intc_core_00_rg_ipr[124]), .Y(n26454) );
  sky130_fd_sc_hd__clkinv_1 U16228 ( .A(j202_soc_core_intc_core_00_rg_itgt[38]), .Y(n25198) );
  sky130_fd_sc_hd__clkinv_1 U16229 ( .A(j202_soc_core_cmt_core_00_reg_addr[6]), 
        .Y(n23646) );
  sky130_fd_sc_hd__clkinv_1 U16230 ( .A(j202_soc_core_intc_core_00_rg_ipr[123]), .Y(n25646) );
  sky130_fd_sc_hd__clkinv_1 U16231 ( .A(j202_soc_core_j22_cpu_ml_macl[23]), 
        .Y(n22030) );
  sky130_fd_sc_hd__clkinv_1 U16232 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[100]), .Y(n25673) );
  sky130_fd_sc_hd__clkinv_1 U16233 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[127]), .Y(n27077) );
  sky130_fd_sc_hd__clkinv_1 U16234 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__0_), 
        .Y(n19451) );
  sky130_fd_sc_hd__clkinv_1 U16235 ( .A(j202_soc_core_intc_core_00_rg_ipr[122]), .Y(n25092) );
  sky130_fd_sc_hd__clkinv_1 U16236 ( .A(j202_soc_core_cmt_core_00_reg_addr[7]), 
        .Y(n23645) );
  sky130_fd_sc_hd__clkinv_1 U16237 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[108]), .Y(n28543) );
  sky130_fd_sc_hd__clkinv_1 U16238 ( .A(j202_soc_core_cmt_core_00_reg_addr[1]), 
        .Y(n23644) );
  sky130_fd_sc_hd__clkinv_1 U16239 ( .A(j202_soc_core_qspi_wb_cyc), .Y(n23459)
         );
  sky130_fd_sc_hd__clkinv_1 U16240 ( .A(j202_soc_core_gpio_core_00_reg_addr[0]), .Y(n27633) );
  sky130_fd_sc_hd__clkinv_1 U16241 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[116]), .Y(n25674) );
  sky130_fd_sc_hd__clkinv_1 U16242 ( .A(j202_soc_core_intc_core_00_rg_itgt[95]), .Y(n27091) );
  sky130_fd_sc_hd__clkinv_1 U16243 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .Y(n25495) );
  sky130_fd_sc_hd__clkinv_1 U16244 ( .A(j202_soc_core_qspi_wb_wdat[0]), .Y(
        n28271) );
  sky130_fd_sc_hd__clkinv_1 U16245 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]), .Y(n28514) );
  sky130_fd_sc_hd__clkinv_1 U16246 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[3]), .Y(n28517) );
  sky130_fd_sc_hd__clkinv_1 U16247 ( .A(j202_soc_core_j22_cpu_ml_macl[6]), .Y(
        n21537) );
  sky130_fd_sc_hd__clkinv_1 U16248 ( .A(j202_soc_core_intc_core_00_rg_itgt[45]), .Y(n25380) );
  sky130_fd_sc_hd__clkinv_1 U16249 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[4]), .Y(n23628) );
  sky130_fd_sc_hd__clkinv_1 U16250 ( .A(j202_soc_core_j22_cpu_ml_mach[28]), 
        .Y(n22416) );
  sky130_fd_sc_hd__clkinv_1 U16251 ( .A(j202_soc_core_intc_core_00_rg_ie[21]), 
        .Y(n25381) );
  sky130_fd_sc_hd__clkinv_1 U16252 ( .A(j202_soc_core_intc_core_00_rg_itgt[76]), .Y(n28532) );
  sky130_fd_sc_hd__clkinv_1 U16253 ( .A(
        j202_soc_core_wbqspiflash_00_write_protect), .Y(n26467) );
  sky130_fd_sc_hd__clkinv_1 U16254 ( .A(j202_soc_core_intc_core_00_rg_itgt[7]), 
        .Y(n25445) );
  sky130_fd_sc_hd__clkinv_1 U16255 ( .A(j202_soc_core_intc_core_00_rg_itgt[6]), 
        .Y(n25438) );
  sky130_fd_sc_hd__clkinv_1 U16256 ( .A(j202_soc_core_intc_core_00_rg_itgt[4]), 
        .Y(n25372) );
  sky130_fd_sc_hd__clkinv_1 U16257 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[1]), .Y(n27647) );
  sky130_fd_sc_hd__clkinv_1 U16258 ( .A(j202_soc_core_intc_core_00_rg_ie[22]), 
        .Y(n26493) );
  sky130_fd_sc_hd__clkinv_1 U16259 ( .A(j202_soc_core_intc_core_00_rg_itgt[2]), 
        .Y(n27153) );
  sky130_fd_sc_hd__clkinv_1 U16260 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[6]), .Y(n23633) );
  sky130_fd_sc_hd__clkinv_1 U16261 ( .A(j202_soc_core_intc_core_00_rg_ie[23]), 
        .Y(n27027) );
  sky130_fd_sc_hd__clkinv_1 U16262 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[29]), .Y(n28730) );
  sky130_fd_sc_hd__clkinv_1 U16263 ( .A(j202_soc_core_j22_cpu_rf_pr[7]), .Y(
        n19042) );
  sky130_fd_sc_hd__clkinv_1 U16264 ( .A(j202_soc_core_j22_cpu_rf_gpr[7]), .Y(
        n14454) );
  sky130_fd_sc_hd__clkinv_1 U16265 ( .A(j202_soc_core_intc_core_00_rg_ie[24]), 
        .Y(n25857) );
  sky130_fd_sc_hd__clkinv_1 U16266 ( .A(j202_soc_core_intc_core_00_rg_itgt[0]), 
        .Y(n27761) );
  sky130_fd_sc_hd__clkinv_1 U16267 ( .A(j202_soc_core_j22_cpu_rf_tmp[7]), .Y(
        n14453) );
  sky130_fd_sc_hd__clkinv_1 U16268 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[19]), .Y(n28709) );
  sky130_fd_sc_hd__clkinv_1 U16269 ( .A(j202_soc_core_intc_core_00_rg_ie[26]), 
        .Y(n25096) );
  sky130_fd_sc_hd__clkinv_1 U16270 ( .A(j202_soc_core_intc_core_00_rg_ie[27]), 
        .Y(n25648) );
  sky130_fd_sc_hd__clkinv_1 U16271 ( .A(j202_soc_core_intc_core_00_rg_itgt[5]), 
        .Y(n25366) );
  sky130_fd_sc_hd__clkinv_1 U16272 ( .A(j202_soc_core_cmt_core_00_cmf0), .Y(
        n27321) );
  sky130_fd_sc_hd__clkinv_1 U16273 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[5]), .Y(n23631) );
  sky130_fd_sc_hd__clkinv_1 U16274 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__1_), 
        .Y(n21856) );
  sky130_fd_sc_hd__clkinv_1 U16275 ( .A(j202_soc_core_intc_core_00_rg_ie[28]), 
        .Y(n26455) );
  sky130_fd_sc_hd__clkinv_1 U16276 ( .A(j202_soc_core_j22_cpu_ml_mach[22]), 
        .Y(n22048) );
  sky130_fd_sc_hd__clkinv_1 U16277 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__3_), 
        .Y(n19043) );
  sky130_fd_sc_hd__clkinv_1 U16278 ( .A(j202_soc_core_j22_cpu_ml_macl[10]), 
        .Y(n19239) );
  sky130_fd_sc_hd__clkinv_1 U16279 ( .A(j202_soc_core_intc_core_00_rg_itgt[3]), 
        .Y(n25284) );
  sky130_fd_sc_hd__clkinv_1 U16280 ( .A(j202_soc_core_intc_core_00_rg_itgt[1]), 
        .Y(n26997) );
  sky130_fd_sc_hd__clkinv_1 U16281 ( .A(j202_soc_core_intc_core_00_rg_ie[29]), 
        .Y(n26958) );
  sky130_fd_sc_hd__clkinv_1 U16282 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[19]), .Y(n28408) );
  sky130_fd_sc_hd__clkinv_1 U16283 ( .A(j202_soc_core_intc_core_00_rg_ie[30]), 
        .Y(n27094) );
  sky130_fd_sc_hd__clkinv_1 U16284 ( .A(j202_soc_core_j22_cpu_ml_macl[26]), 
        .Y(n22407) );
  sky130_fd_sc_hd__clkinv_1 U16285 ( .A(j202_soc_core_intc_core_00_rg_ie[31]), 
        .Y(n27080) );
  sky130_fd_sc_hd__clkinv_1 U16286 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[107]), .Y(n27514) );
  sky130_fd_sc_hd__clkinv_1 U16287 ( .A(j202_soc_core_intc_core_00_rg_ipr[60]), 
        .Y(n26451) );
  sky130_fd_sc_hd__clkinv_1 U16288 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[5]), .Y(n13386) );
  sky130_fd_sc_hd__clkinv_1 U16289 ( .A(j202_soc_core_intc_core_00_rg_ipr[4]), 
        .Y(n24601) );
  sky130_fd_sc_hd__clkinv_1 U16290 ( .A(j202_soc_core_intc_core_00_rg_ipr[52]), 
        .Y(n25520) );
  sky130_fd_sc_hd__clkinv_1 U16291 ( .A(j202_soc_core_intc_core_00_rg_itgt[75]), .Y(n27710) );
  sky130_fd_sc_hd__clkinv_1 U16292 ( .A(j202_soc_core_j22_cpu_rf_gpr[5]), .Y(
        n21861) );
  sky130_fd_sc_hd__clkinv_1 U16293 ( .A(j202_soc_core_j22_cpu_pc[22]), .Y(
        n15408) );
  sky130_fd_sc_hd__clkinv_1 U16294 ( .A(j202_soc_core_j22_cpu_ml_mach[1]), .Y(
        n17467) );
  sky130_fd_sc_hd__clkinv_1 U16295 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[17]), .Y(n28395) );
  sky130_fd_sc_hd__clkinv_1 U16296 ( .A(j202_soc_core_j22_cpu_ml_mach[27]), 
        .Y(n22419) );
  sky130_fd_sc_hd__clkinv_1 U16297 ( .A(j202_soc_core_j22_cpu_rf_pr[5]), .Y(
        n21855) );
  sky130_fd_sc_hd__clkinv_1 U16298 ( .A(j202_soc_core_intc_core_00_rg_ipr[12]), 
        .Y(n25358) );
  sky130_fd_sc_hd__clkinv_1 U16299 ( .A(j202_soc_core_intc_core_00_rg_ipr[40]), 
        .Y(n25459) );
  sky130_fd_sc_hd__clkinv_1 U16300 ( .A(j202_soc_core_intc_core_00_rg_itgt[43]), .Y(n27809) );
  sky130_fd_sc_hd__clkinv_1 U16301 ( .A(j202_soc_core_j22_cpu_pc[19]), .Y(
        n15767) );
  sky130_fd_sc_hd__clkinv_1 U16302 ( .A(j202_soc_core_j22_cpu_ma_M_area[0]), 
        .Y(n13381) );
  sky130_fd_sc_hd__clkinv_1 U16303 ( .A(j202_soc_core_intc_core_00_rg_itgt[74]), .Y(n27288) );
  sky130_fd_sc_hd__clkinv_1 U16304 ( .A(j202_soc_core_memory0_ram_dout0_sel[3]), .Y(n13373) );
  sky130_fd_sc_hd__clkinv_1 U16305 ( .A(j202_soc_core_aquc_WE_), .Y(n22296) );
  sky130_fd_sc_hd__clkinv_1 U16306 ( .A(j202_soc_core_uart_TOP_tx_bit_cnt[2]), 
        .Y(n28625) );
  sky130_fd_sc_hd__clkinv_1 U16307 ( .A(j202_soc_core_intc_core_00_bs_addr[2]), 
        .Y(n24026) );
  sky130_fd_sc_hd__clkinv_1 U16308 ( .A(j202_soc_core_j22_cpu_ml_bufa[18]), 
        .Y(n22202) );
  sky130_fd_sc_hd__clkinv_1 U16309 ( .A(j202_soc_core_j22_cpu_ml_macl[9]), .Y(
        n22926) );
  sky130_fd_sc_hd__clkinv_1 U16310 ( .A(j202_soc_core_bldc_core_00_pwm_duty[5]), .Y(n25742) );
  sky130_fd_sc_hd__clkinv_1 U16311 ( .A(j202_soc_core_j22_cpu_ml_macl[25]), 
        .Y(n22841) );
  sky130_fd_sc_hd__clkinv_1 U16312 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[105]), .Y(n28527) );
  sky130_fd_sc_hd__clkinv_1 U16313 ( .A(j202_soc_core_intc_core_00_rg_itgt[73]), .Y(n27538) );
  sky130_fd_sc_hd__clkinv_1 U16314 ( .A(
        j202_soc_core_intc_core_00_in_intreq[19]), .Y(n25692) );
  sky130_fd_sc_hd__clkinv_1 U16315 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[1]), .Y(n23625) );
  sky130_fd_sc_hd__clkinv_1 U16316 ( .A(j202_soc_core_intc_core_00_bs_addr[4]), 
        .Y(n28890) );
  sky130_fd_sc_hd__clkinv_1 U16317 ( .A(j202_soc_core_intc_core_00_rg_ipr[18]), 
        .Y(n25360) );
  sky130_fd_sc_hd__clkinv_1 U16318 ( .A(j202_soc_core_qspi_wb_wdat[9]), .Y(
        n28332) );
  sky130_fd_sc_hd__clkinv_1 U16319 ( .A(j202_soc_core_intc_core_00_rg_ipr[20]), 
        .Y(n25430) );
  sky130_fd_sc_hd__clkinv_1 U16320 ( .A(j202_soc_core_intc_core_00_rg_ie[8]), 
        .Y(n25476) );
  sky130_fd_sc_hd__clkinv_1 U16321 ( .A(j202_soc_core_intc_core_00_rg_itgt[41]), .Y(n26935) );
  sky130_fd_sc_hd__clkinv_1 U16322 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[104]), .Y(n27849) );
  sky130_fd_sc_hd__xnor2_1 U16323 ( .A(j202_soc_core_j22_cpu_ml_bufa[28]), .B(
        j202_soc_core_j22_cpu_ml_bufa[27]), .Y(n17371) );
  sky130_fd_sc_hd__clkinv_1 U16324 ( .A(j202_soc_core_j22_cpu_rf_pr[6]), .Y(
        n21552) );
  sky130_fd_sc_hd__clkinv_1 U16325 ( .A(j202_soc_core_j22_cpu_ifetchl), .Y(
        n24474) );
  sky130_fd_sc_hd__clkinv_1 U16326 ( .A(j202_soc_core_j22_cpu_pc[16]), .Y(
        n20994) );
  sky130_fd_sc_hd__clkinv_1 U16327 ( .A(j202_soc_core_qspi_wb_addr[2]), .Y(
        n28116) );
  sky130_fd_sc_hd__clkinv_1 U16328 ( .A(j202_soc_core_j22_cpu_ml_macl[4]), .Y(
        n19428) );
  sky130_fd_sc_hd__clkinv_1 U16329 ( .A(j202_soc_core_j22_cpu_ml_macl[20]), 
        .Y(n22141) );
  sky130_fd_sc_hd__clkinv_1 U16330 ( .A(j202_soc_core_intc_core_00_rg_itgt[52]), .Y(n25721) );
  sky130_fd_sc_hd__clkinv_1 U16331 ( .A(j202_soc_core_j22_cpu_rf_gpr[6]), .Y(
        n13944) );
  sky130_fd_sc_hd__clkinv_1 U16332 ( .A(j202_soc_core_intc_core_00_rg_itgt[24]), .Y(n27756) );
  sky130_fd_sc_hd__clkinv_1 U16333 ( .A(j202_soc_core_j22_cpu_id_opn_v_), .Y(
        n16048) );
  sky130_fd_sc_hd__clkinv_1 U16334 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__2_), 
        .Y(n21553) );
  sky130_fd_sc_hd__clkinv_1 U16335 ( .A(j202_soc_core_intc_core_00_rg_itgt[92]), .Y(n28531) );
  sky130_fd_sc_hd__clkinv_1 U16336 ( .A(j202_soc_core_j22_cpu_regop_We__3_), 
        .Y(n23555) );
  sky130_fd_sc_hd__clkinv_1 U16337 ( .A(j202_soc_core_intc_core_00_rg_itgt[44]), .Y(n25730) );
  sky130_fd_sc_hd__clkinv_1 U16338 ( .A(j202_soc_core_intr_level__2_), .Y(
        n16042) );
  sky130_fd_sc_hd__clkinv_1 U16339 ( .A(j202_soc_core_j22_cpu_ml_macl[3]), .Y(
        n17808) );
  sky130_fd_sc_hd__clkinv_1 U16340 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd), .Y(n28109) );
  sky130_fd_sc_hd__clkinv_1 U16341 ( .A(j202_soc_core_j22_cpu_ml_macl[19]), 
        .Y(n22953) );
  sky130_fd_sc_hd__clkinv_1 U16342 ( .A(j202_soc_core_intc_core_00_rg_ipr[117]), .Y(n25379) );
  sky130_fd_sc_hd__clkinv_1 U16343 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[3]), .Y(n26210) );
  sky130_fd_sc_hd__clkinv_1 U16344 ( .A(j202_soc_core_j22_cpu_rf_gbr[6]), .Y(
        n21554) );
  sky130_fd_sc_hd__clkinv_1 U16345 ( .A(j202_soc_core_intr_level__1_), .Y(
        n16041) );
  sky130_fd_sc_hd__clkinv_1 U16346 ( .A(j202_soc_core_intc_core_00_rg_itgt[36]), .Y(n28530) );
  sky130_fd_sc_hd__clkinv_1 U16347 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[123]), .Y(n27511) );
  sky130_fd_sc_hd__clkinv_1 U16348 ( .A(j202_soc_core_intc_core_00_rg_itgt[91]), .Y(n27707) );
  sky130_fd_sc_hd__clkinv_1 U16349 ( .A(j202_soc_core_intc_core_00_rg_ipr[113]), .Y(n25722) );
  sky130_fd_sc_hd__clkinv_1 U16350 ( .A(j202_soc_core_intr_level__3_), .Y(
        n16038) );
  sky130_fd_sc_hd__clkinv_1 U16351 ( .A(j202_soc_core_bldc_core_00_pwm_duty[7]), .Y(n25701) );
  sky130_fd_sc_hd__clkinv_1 U16352 ( .A(j202_soc_core_intc_core_00_rg_itgt[26]), .Y(n27155) );
  sky130_fd_sc_hd__clkinv_1 U16353 ( .A(j202_soc_core_intc_core_00_rg_itgt[59]), .Y(n27807) );
  sky130_fd_sc_hd__clkinv_1 U16354 ( .A(j202_soc_core_intc_core_00_rg_itgt[28]), .Y(n27052) );
  sky130_fd_sc_hd__clkinv_1 U16355 ( .A(j202_soc_core_j22_cpu_ml_macl[2]), .Y(
        n19186) );
  sky130_fd_sc_hd__clkinv_1 U16356 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[23]), .Y(n28722) );
  sky130_fd_sc_hd__clkinv_1 U16357 ( .A(j202_soc_core_j22_cpu_opst[0]), .Y(
        n27978) );
  sky130_fd_sc_hd__clkinv_1 U16358 ( .A(j202_soc_core_j22_cpu_ml_macl[18]), 
        .Y(n22198) );
  sky130_fd_sc_hd__clkinv_1 U16359 ( .A(j202_soc_core_intc_core_00_rg_ipr[116]), .Y(n27584) );
  sky130_fd_sc_hd__clkinv_1 U16360 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[1]), .Y(n17183) );
  sky130_fd_sc_hd__clkinv_1 U16361 ( .A(j202_soc_core_intc_core_00_rg_ipr[81]), 
        .Y(n25719) );
  sky130_fd_sc_hd__clkinv_1 U16362 ( .A(j202_soc_core_intc_core_00_rg_itgt[90]), .Y(n27285) );
  sky130_fd_sc_hd__clkinv_1 U16363 ( .A(j202_soc_core_j22_cpu_rf_pr[9]), .Y(
        n22855) );
  sky130_fd_sc_hd__clkinv_1 U16364 ( .A(j202_soc_core_intc_core_00_rg_ipr[106]), .Y(n27287) );
  sky130_fd_sc_hd__clkinv_1 U16365 ( .A(j202_soc_core_intc_core_00_bs_addr[9]), 
        .Y(n24970) );
  sky130_fd_sc_hd__clkinv_1 U16366 ( .A(j202_soc_core_j22_cpu_ml_macl[1]), .Y(
        n22724) );
  sky130_fd_sc_hd__clkinv_1 U16367 ( .A(j202_soc_core_intc_core_00_rg_ipr[114]), .Y(n28540) );
  sky130_fd_sc_hd__clkinv_1 U16368 ( .A(j202_soc_core_intc_core_00_rg_ipr[108]), .Y(n26266) );
  sky130_fd_sc_hd__clkinv_1 U16369 ( .A(j202_soc_core_j22_cpu_ml_macl[17]), 
        .Y(n22806) );
  sky130_fd_sc_hd__clkinv_1 U16370 ( .A(j202_soc_core_intc_core_00_rg_ipr[109]), .Y(n28529) );
  sky130_fd_sc_hd__clkinv_1 U16371 ( .A(j202_soc_core_intc_core_00_rg_ie[17]), 
        .Y(n25729) );
  sky130_fd_sc_hd__clkinv_1 U16372 ( .A(j202_soc_core_intc_core_00_rg_itgt[30]), .Y(n25855) );
  sky130_fd_sc_hd__clkinv_1 U16373 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[13]), .Y(n28366) );
  sky130_fd_sc_hd__clkinv_1 U16374 ( .A(j202_soc_core_j22_cpu_rf_gpr[505]), 
        .Y(n22876) );
  sky130_fd_sc_hd__clkinv_1 U16375 ( .A(j202_soc_core_intc_core_00_rg_ipr[110]), .Y(n27709) );
  sky130_fd_sc_hd__clkinv_1 U16376 ( .A(j202_soc_core_intc_core_00_rg_ipr[112]), .Y(n27053) );
  sky130_fd_sc_hd__clkinv_1 U16377 ( .A(j202_soc_core_intc_core_00_rg_ipr[111]), .Y(n27513) );
  sky130_fd_sc_hd__clkinv_1 U16378 ( .A(j202_soc_core_j22_cpu_rf_vbr[25]), .Y(
        n22878) );
  sky130_fd_sc_hd__clkinv_1 U16379 ( .A(j202_soc_core_j22_cpu_pc_hold), .Y(
        n23861) );
  sky130_fd_sc_hd__clkinv_1 U16380 ( .A(
        j202_soc_core_wbqspiflash_00_spi_len[0]), .Y(n23333) );
  sky130_fd_sc_hd__clkinv_1 U16381 ( .A(j202_soc_core_intc_core_00_rg_itgt[31]), .Y(n26453) );
  sky130_fd_sc_hd__clkinv_1 U16382 ( .A(j202_soc_core_qspi_wb_wdat[13]), .Y(
        n28360) );
  sky130_fd_sc_hd__clkinv_1 U16383 ( .A(j202_soc_core_j22_cpu_ml_mach[24]), 
        .Y(n22386) );
  sky130_fd_sc_hd__clkinv_1 U16384 ( .A(
        j202_soc_core_wbqspiflash_00_spi_len[1]), .Y(n26226) );
  sky130_fd_sc_hd__clkinv_1 U16385 ( .A(j202_soc_core_qspi_wb_wdat[19]), .Y(
        n25699) );
  sky130_fd_sc_hd__clkinv_1 U16386 ( .A(j202_soc_core_qspi_wb_addr[3]), .Y(
        n28106) );
  sky130_fd_sc_hd__clkinv_1 U16387 ( .A(j202_soc_core_intc_core_00_rg_itgt[88]), .Y(n24976) );
  sky130_fd_sc_hd__clkinv_1 U16388 ( .A(j202_soc_core_wbqspiflash_00_spi_spd), 
        .Y(n28110) );
  sky130_fd_sc_hd__clkinv_1 U16389 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[120]), .Y(n27847) );
  sky130_fd_sc_hd__clkinv_1 U16390 ( .A(j202_soc_core_intc_core_00_rg_itgt[57]), .Y(n26932) );
  sky130_fd_sc_hd__clkinv_1 U16391 ( .A(j202_soc_core_wbqspiflash_00_spi_in[1]), .Y(n28655) );
  sky130_fd_sc_hd__clkinv_1 U16392 ( .A(j202_soc_core_intc_core_00_rg_itgt[89]), .Y(n27535) );
  sky130_fd_sc_hd__clkinv_1 U16393 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[2]), .Y(n24948) );
  sky130_fd_sc_hd__clkinv_1 U16394 ( .A(j202_soc_core_j22_cpu_ml_mach[5]), .Y(
        n17490) );
  sky130_fd_sc_hd__clkinv_1 U16395 ( .A(j202_soc_core_intc_core_00_rg_ipr[28]), 
        .Y(n24029) );
  sky130_fd_sc_hd__clkinv_1 U16396 ( .A(j202_soc_core_intc_core_00_rg_ipr[88]), 
        .Y(n25862) );
  sky130_fd_sc_hd__clkinv_1 U16397 ( .A(j202_soc_core_uart_sio_ce), .Y(n28564)
         );
  sky130_fd_sc_hd__clkinv_1 U16398 ( .A(j202_soc_core_cmt_core_00_reg_addr[0]), 
        .Y(n23666) );
  sky130_fd_sc_hd__clkinv_1 U16399 ( .A(j202_soc_core_intc_core_00_rg_ipr[90]), 
        .Y(n25089) );
  sky130_fd_sc_hd__clkinv_1 U16400 ( .A(j202_soc_core_j22_cpu_ml_mach[4]), .Y(
        n17389) );
  sky130_fd_sc_hd__clkinv_1 U16401 ( .A(j202_soc_core_j22_cpu_ml_macl[22]), 
        .Y(n22337) );
  sky130_fd_sc_hd__clkinv_1 U16402 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[124]), .Y(n28546) );
  sky130_fd_sc_hd__clkinv_1 U16403 ( .A(j202_soc_core_bldc_core_00_comm[1]), 
        .Y(n28583) );
  sky130_fd_sc_hd__clkinv_1 U16404 ( .A(j202_soc_core_intc_core_00_rg_ipr[91]), 
        .Y(n25643) );
  sky130_fd_sc_hd__clkinv_1 U16405 ( .A(j202_soc_core_cmt_core_00_reg_addr[2]), 
        .Y(n24842) );
  sky130_fd_sc_hd__clkinv_1 U16406 ( .A(j202_soc_core_intc_core_00_rg_ipr[92]), 
        .Y(n26452) );
  sky130_fd_sc_hd__clkinv_1 U16407 ( .A(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[1]), .Y(n19859) );
  sky130_fd_sc_hd__clkinv_1 U16408 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[20]), .Y(n28712) );
  sky130_fd_sc_hd__clkinv_1 U16409 ( .A(j202_soc_core_intc_core_00_rg_ipr[93]), 
        .Y(n26953) );
  sky130_fd_sc_hd__clkinv_1 U16410 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[19]), .Y(n28188) );
  sky130_fd_sc_hd__clkinv_1 U16411 ( .A(j202_soc_core_intc_core_00_rg_ipr[94]), 
        .Y(n27100) );
  sky130_fd_sc_hd__clkinv_1 U16412 ( .A(j202_soc_core_intc_core_00_rg_ipr[95]), 
        .Y(n27075) );
  sky130_fd_sc_hd__clkinv_1 U16413 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[0]), .Y(n27731) );
  sky130_fd_sc_hd__clkinv_1 U16414 ( .A(j202_soc_core_intc_core_00_rg_itgt[46]), .Y(n25201) );
  sky130_fd_sc_hd__clkinv_1 U16415 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[3]), .Y(n28297) );
  sky130_fd_sc_hd__clkinv_1 U16416 ( .A(j202_soc_core_intc_core_00_rg_itgt[63]), .Y(n26955) );
  sky130_fd_sc_hd__clkinv_1 U16417 ( .A(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled), .Y(n25973) );
  sky130_fd_sc_hd__clkinv_1 U16418 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[2]), .Y(n17182) );
  sky130_fd_sc_hd__clkinv_1 U16419 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[126]), .Y(n25645) );
  sky130_fd_sc_hd__clkinv_1 U16420 ( .A(j202_soc_core_wbqspiflash_00_spi_in[0]), .Y(n28652) );
  sky130_fd_sc_hd__clkinv_1 U16421 ( .A(j202_soc_core_pwrite[0]), .Y(n24820)
         );
  sky130_fd_sc_hd__clkinv_1 U16422 ( .A(j202_soc_core_intc_core_00_rg_ie[12]), 
        .Y(n25507) );
  sky130_fd_sc_hd__clkinv_1 U16423 ( .A(j202_soc_core_intc_core_00_rg_itgt[94]), .Y(n25091) );
  sky130_fd_sc_hd__nor2_4 U16424 ( .A(j202_soc_core_j22_cpu_ma_M_area[1]), .B(
        j202_soc_core_j22_cpu_ma_M_area[0]), .Y(n21771) );
  sky130_fd_sc_hd__clkinv_1 U16425 ( .A(j202_soc_core_intc_core_00_rg_ipr[120]), .Y(n25856) );
  sky130_fd_sc_hd__clkinv_1 U16426 ( .A(j202_soc_core_j22_cpu_ml_mach[9]), .Y(
        n18044) );
  sky130_fd_sc_hd__clkinv_1 U16427 ( .A(j202_soc_core_j22_cpu_ml_macl[5]), .Y(
        n17769) );
  sky130_fd_sc_hd__clkinv_1 U16428 ( .A(j202_soc_core_qspi_wb_addr[24]), .Y(
        n26153) );
  sky130_fd_sc_hd__clkinv_1 U16429 ( .A(j202_soc_core_j22_cpu_ml_mach[25]), 
        .Y(n22383) );
  sky130_fd_sc_hd__clkinv_1 U16430 ( .A(j202_soc_core_ahb2apb_02_state[2]), 
        .Y(n24316) );
  sky130_fd_sc_hd__clkinv_1 U16431 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[0]), .Y(n28095) );
  sky130_fd_sc_hd__clkinv_1 U16432 ( .A(j202_soc_core_j22_cpu_ml_macl[21]), 
        .Y(n22113) );
  sky130_fd_sc_hd__clkinv_1 U16433 ( .A(j202_soc_core_intc_core_00_rg_ipr[98]), 
        .Y(n24980) );
  sky130_fd_sc_hd__clkinv_1 U16434 ( .A(j202_soc_core_ahb2apb_00_state[0]), 
        .Y(n20986) );
  sky130_fd_sc_hd__clkinv_1 U16435 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[21]), .Y(n28715) );
  sky130_fd_sc_hd__clkinv_1 U16436 ( .A(j202_soc_core_wbqspiflash_00_spif_ctrl), .Y(n26134) );
  sky130_fd_sc_hd__clkinv_1 U16437 ( .A(j202_soc_core_intc_core_00_rg_ipr[99]), 
        .Y(n27848) );
  sky130_fd_sc_hd__clkinv_1 U16438 ( .A(j202_soc_core_cmt_core_00_cks0[0]), 
        .Y(n24846) );
  sky130_fd_sc_hd__clkinv_1 U16439 ( .A(j202_soc_core_intc_core_00_rg_itgt[54]), .Y(n25205) );
  sky130_fd_sc_hd__clkinv_1 U16440 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[1]), 
        .Y(n24378) );
  sky130_fd_sc_hd__clkinv_1 U16441 ( .A(j202_soc_core_ahb2apb_02_state[0]), 
        .Y(n23312) );
  sky130_fd_sc_hd__clkinv_1 U16442 ( .A(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[1]), .Y(n24817) );
  sky130_fd_sc_hd__clkinv_1 U16443 ( .A(j202_soc_core_intc_core_00_rg_ipr[100]), .Y(n26995) );
  sky130_fd_sc_hd__clkinv_1 U16444 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[28]), .Y(n28726) );
  sky130_fd_sc_hd__clkinv_1 U16445 ( .A(j202_soc_core_intc_core_00_rg_itgt[29]), .Y(n27580) );
  sky130_fd_sc_hd__clkinv_1 U16446 ( .A(j202_soc_core_ahb2apb_00_state[1]), 
        .Y(n24812) );
  sky130_fd_sc_hd__clkinv_1 U16447 ( .A(j202_soc_core_wbqspiflash_00_spif_cmd), 
        .Y(n26135) );
  sky130_fd_sc_hd__clkinv_1 U16448 ( .A(j202_soc_core_intc_core_00_rg_ipr[101]), .Y(n26934) );
  sky130_fd_sc_hd__clkinv_1 U16449 ( .A(j202_soc_core_intc_core_00_rg_ipr[119]), .Y(n27025) );
  sky130_fd_sc_hd__clkinv_1 U16450 ( .A(j202_soc_core_uart_div0[7]), .Y(n27043) );
  sky130_fd_sc_hd__clkinv_1 U16451 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[125]), .Y(n27024) );
  sky130_fd_sc_hd__clkinv_1 U16452 ( .A(j202_soc_core_intc_core_00_rg_ipr[102]), .Y(n27537) );
  sky130_fd_sc_hd__clkinv_1 U16453 ( .A(j202_soc_core_intc_core_00_rg_itgt[60]), .Y(n25720) );
  sky130_fd_sc_hd__clkinv_1 U16454 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[2]), .Y(n20982) );
  sky130_fd_sc_hd__clkinv_1 U16455 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[0]), .Y(n28148) );
  sky130_fd_sc_hd__clkinv_1 U16456 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[22]), .Y(n28718) );
  sky130_fd_sc_hd__clkinv_1 U16457 ( .A(j202_soc_core_j22_cpu_ml_mach[6]), .Y(
        n17983) );
  sky130_fd_sc_hd__clkinv_1 U16458 ( .A(j202_soc_core_intc_core_00_rg_itgt[62]), .Y(n25199) );
  sky130_fd_sc_hd__clkinv_1 U16459 ( .A(j202_soc_core_intc_core_00_rg_ipr[103]), .Y(n27305) );
  sky130_fd_sc_hd__clkinv_1 U16460 ( .A(j202_soc_core_intc_core_00_rg_ipr[104]), .Y(n27156) );
  sky130_fd_sc_hd__clkinv_1 U16461 ( .A(j202_soc_core_qspi_wb_wdat[2]), .Y(
        n28283) );
  sky130_fd_sc_hd__clkinv_1 U16462 ( .A(j202_soc_core_intc_core_00_rg_itgt[93]), .Y(n26490) );
  sky130_fd_sc_hd__clkinv_1 U16463 ( .A(j202_soc_core_intc_core_00_rg_ipr[118]), .Y(n26491) );
  sky130_fd_sc_hd__clkinv_1 U16464 ( .A(j202_soc_core_intc_core_00_rg_itgt[61]), .Y(n25378) );
  sky130_fd_sc_hd__clkinv_1 U16465 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[121]), .Y(n27303) );
  sky130_fd_sc_hd__clkinv_1 U16466 ( .A(j202_soc_core_intc_core_00_rg_itgt[64]), .Y(n24983) );
  sky130_fd_sc_hd__clkinv_1 U16467 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[1]), 
        .Y(n23664) );
  sky130_fd_sc_hd__clkinv_1 U16468 ( .A(j202_soc_core_j22_cpu_pc[21]), .Y(
        n15655) );
  sky130_fd_sc_hd__clkinv_1 U16469 ( .A(j202_soc_core_intc_core_00_rg_itgt[78]), .Y(n25093) );
  sky130_fd_sc_hd__clkinv_1 U16470 ( .A(j202_soc_core_intc_core_00_rg_ie[4]), 
        .Y(n25371) );
  sky130_fd_sc_hd__clkinv_1 U16471 ( .A(j202_soc_core_intc_core_00_rg_itgt[96]), .Y(n28523) );
  sky130_fd_sc_hd__clkinv_1 U16472 ( .A(j202_soc_core_j22_cpu_rf_pr[8]), .Y(
        n21991) );
  sky130_fd_sc_hd__clkinv_1 U16473 ( .A(j202_soc_core_j22_cpu_rf_tmp[6]), .Y(
        n13940) );
  sky130_fd_sc_hd__clkinv_1 U16474 ( .A(j202_soc_core_cmt_core_00_cks1[1]), 
        .Y(n23679) );
  sky130_fd_sc_hd__clkinv_1 U16475 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[110]), .Y(n25647) );
  sky130_fd_sc_hd__clkinv_1 U16476 ( .A(j202_soc_core_j22_cpu_ml_mach[10]), 
        .Y(n18152) );
  sky130_fd_sc_hd__clkinv_1 U16477 ( .A(j202_soc_core_intc_core_00_rg_itgt[34]), .Y(n25626) );
  sky130_fd_sc_hd__clkinv_1 U16478 ( .A(j202_soc_core_intc_core_00_rg_itgt[47]), .Y(n26957) );
  sky130_fd_sc_hd__clkinv_1 U16479 ( .A(j202_soc_core_intc_core_00_rg_itgt[56]), .Y(n27667) );
  sky130_fd_sc_hd__clkinv_1 U16480 ( .A(j202_soc_core_intc_core_00_rg_ie[3]), 
        .Y(n25283) );
  sky130_fd_sc_hd__clkinv_1 U16481 ( .A(j202_soc_core_intc_core_00_rg_ipr[16]), 
        .Y(n25429) );
  sky130_fd_sc_hd__clkinv_1 U16482 ( .A(j202_soc_core_intc_core_00_rg_itgt[16]), .Y(n25768) );
  sky130_fd_sc_hd__clkinv_1 U16483 ( .A(j202_soc_core_intc_core_00_rg_itgt[79]), .Y(n27093) );
  sky130_fd_sc_hd__clkinv_1 U16484 ( .A(j202_soc_core_intc_core_00_rg_eimk[0]), 
        .Y(n27753) );
  sky130_fd_sc_hd__clkinv_1 U16485 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[8]), .Y(n23624) );
  sky130_fd_sc_hd__clkinv_1 U16486 ( .A(j202_soc_core_j22_cpu_rf_tmp[26]), .Y(
        n16006) );
  sky130_fd_sc_hd__clkinv_1 U16487 ( .A(j202_soc_core_intc_core_00_rg_itgt[42]), .Y(n25630) );
  sky130_fd_sc_hd__clkinv_1 U16488 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[5]), .Y(n24894) );
  sky130_fd_sc_hd__and2_0 U16489 ( .A(j202_soc_core_ahb2wbqspi_00_stb_o), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .X(n23476) );
  sky130_fd_sc_hd__clkinv_1 U16490 ( .A(j202_soc_core_j22_cpu_rf_pr[26]), .Y(
        n16011) );
  sky130_fd_sc_hd__clkinv_1 U16491 ( .A(j202_soc_core_intc_core_00_rg_itgt[33]), .Y(n26937) );
  sky130_fd_sc_hd__clkinv_1 U16492 ( .A(j202_soc_core_intc_core_00_rg_itgt[48]), .Y(n27668) );
  sky130_fd_sc_hd__clkinv_1 U16493 ( .A(j202_soc_core_intc_core_00_rg_itgt[68]), .Y(n28534) );
  sky130_fd_sc_hd__clkinv_1 U16494 ( .A(j202_soc_core_j22_cpu_pc[26]), .Y(
        n16009) );
  sky130_fd_sc_hd__clkinv_1 U16495 ( .A(j202_soc_core_qspi_wb_wdat[25]), .Y(
        n25213) );
  sky130_fd_sc_hd__clkinv_1 U16496 ( .A(j202_soc_core_j22_cpu_rf_gpr[26]), .Y(
        n16015) );
  sky130_fd_sc_hd__clkinv_1 U16497 ( .A(j202_soc_core_j22_cpu_rf_gpr[2]), .Y(
        n14107) );
  sky130_fd_sc_hd__clkinv_1 U16498 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[3]), .Y(n24891) );
  sky130_fd_sc_hd__clkinv_1 U16499 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[25]), .Y(n28455) );
  sky130_fd_sc_hd__clkinv_1 U16500 ( .A(j202_soc_core_j22_cpu_rf_gpr[8]), .Y(
        n21998) );
  sky130_fd_sc_hd__clkinv_1 U16501 ( .A(j202_soc_core_intc_core_00_rg_ipr[17]), 
        .Y(n25428) );
  sky130_fd_sc_hd__clkinv_1 U16502 ( .A(j202_soc_core_intc_core_00_rg_itgt[50]), .Y(n25628) );
  sky130_fd_sc_hd__clkinv_1 U16503 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[15]), .Y(n23629) );
  sky130_fd_sc_hd__clkinv_1 U16504 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[111]), .Y(n27079) );
  sky130_fd_sc_hd__clkinv_1 U16505 ( .A(j202_soc_core_cmt_core_00_cnt0[13]), 
        .Y(n27475) );
  sky130_fd_sc_hd__clkinv_1 U16506 ( .A(j202_soc_core_j22_cpu_rf_gbr[26]), .Y(
        n16013) );
  sky130_fd_sc_hd__clkinv_1 U16507 ( .A(j202_soc_core_intc_core_00_rg_itgt[40]), .Y(n27670) );
  sky130_fd_sc_hd__clkinv_1 U16508 ( .A(j202_soc_core_intc_core_00_rg_ipr[11]), 
        .Y(n25278) );
  sky130_fd_sc_hd__clkinv_1 U16509 ( .A(j202_soc_core_intc_core_00_rg_itgt[17]), .Y(n25761) );
  sky130_fd_sc_hd__clkinv_1 U16510 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[13]), .Y(n23632) );
  sky130_fd_sc_hd__clkinv_1 U16511 ( .A(j202_soc_core_intc_core_00_rg_itgt[65]), .Y(n27540) );
  sky130_fd_sc_hd__clkinv_1 U16512 ( .A(j202_soc_core_intc_core_00_rg_ipr[31]), 
        .Y(n25447) );
  sky130_fd_sc_hd__clkinv_1 U16513 ( .A(j202_soc_core_intc_core_00_rg_itgt[19]), .Y(n26265) );
  sky130_fd_sc_hd__clkinv_1 U16514 ( .A(j202_soc_core_intc_core_00_rg_itgt[67]), .Y(n27706) );
  sky130_fd_sc_hd__clkinv_1 U16515 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[9]), .Y(n23634) );
  sky130_fd_sc_hd__clkinv_1 U16516 ( .A(j202_soc_core_intc_core_00_rg_ipr[27]), 
        .Y(n25448) );
  sky130_fd_sc_hd__clkinv_1 U16517 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[7]), .Y(n24900) );
  sky130_fd_sc_hd__clkinv_1 U16518 ( .A(j202_soc_core_qspi_wb_wdat[5]), .Y(
        n28304) );
  sky130_fd_sc_hd__clkinv_1 U16519 ( .A(j202_soc_core_intc_core_00_rg_itgt[21]), .Y(n27582) );
  sky130_fd_sc_hd__clkinv_1 U16520 ( .A(j202_soc_core_j22_cpu_ml_mach[0]), .Y(
        n17529) );
  sky130_fd_sc_hd__clkinv_1 U16521 ( .A(j202_soc_core_j22_cpu_ml_macl[16]), 
        .Y(n22530) );
  sky130_fd_sc_hd__clkinv_1 U16522 ( .A(j202_soc_core_intc_core_00_rg_itgt[97]), .Y(n27302) );
  sky130_fd_sc_hd__clkinv_1 U16523 ( .A(j202_soc_core_intc_core_00_rg_itgt[58]), .Y(n25627) );
  sky130_fd_sc_hd__clkinv_1 U16524 ( .A(j202_soc_core_intc_core_00_rg_ie[2]), 
        .Y(n27201) );
  sky130_fd_sc_hd__clkinv_1 U16525 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[0]), 
        .Y(n24694) );
  sky130_fd_sc_hd__clkinv_1 U16526 ( .A(j202_soc_core_j22_cpu_ml_macl[15]), 
        .Y(n17589) );
  sky130_fd_sc_hd__clkinv_1 U16527 ( .A(j202_soc_core_j22_cpu_rf_tmp[3]), .Y(
        n21413) );
  sky130_fd_sc_hd__clkinv_1 U16528 ( .A(j202_soc_core_intc_core_00_rg_ie[0]), 
        .Y(n25357) );
  sky130_fd_sc_hd__clkinv_1 U16529 ( .A(j202_soc_core_j22_cpu_rfuo_sr__q_), 
        .Y(n21992) );
  sky130_fd_sc_hd__clkinv_1 U16530 ( .A(j202_soc_core_intc_core_00_rg_ipr[24]), 
        .Y(n25863) );
  sky130_fd_sc_hd__clkinv_1 U16531 ( .A(j202_soc_core_intc_core_00_rg_itgt[32]), .Y(n27672) );
  sky130_fd_sc_hd__clkinv_1 U16532 ( .A(j202_soc_core_cmt_core_00_cnt0[15]), 
        .Y(n27480) );
  sky130_fd_sc_hd__clkinv_1 U16533 ( .A(j202_soc_core_intc_core_00_rg_itgt[99]), .Y(n27510) );
  sky130_fd_sc_hd__clkinv_1 U16534 ( .A(j202_soc_core_intc_core_00_rg_itgt[39]), .Y(n26954) );
  sky130_fd_sc_hd__clkinv_1 U16535 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[1]), .Y(n27682) );
  sky130_fd_sc_hd__clkinv_1 U16536 ( .A(j202_soc_core_cmt_core_00_reg_addr[5]), 
        .Y(n23665) );
  sky130_fd_sc_hd__clkinv_1 U16537 ( .A(j202_soc_core_intc_core_00_rg_itgt[18]), .Y(n26816) );
  sky130_fd_sc_hd__clkinv_1 U16538 ( .A(j202_soc_core_intc_core_00_rg_itgt[66]), .Y(n27284) );
  sky130_fd_sc_hd__clkinv_1 U16539 ( .A(j202_soc_core_j22_cpu_ml_mach[29]), 
        .Y(n22417) );
  sky130_fd_sc_hd__clkinv_1 U16540 ( .A(j202_soc_core_j22_cpu_rf_pr[1]), .Y(
        n22780) );
  sky130_fd_sc_hd__clkinv_1 U16541 ( .A(j202_soc_core_intc_core_00_rg_ipr[29]), 
        .Y(n25446) );
  sky130_fd_sc_hd__clkinv_1 U16542 ( .A(j202_soc_core_j22_cpu_ml_macl[28]), 
        .Y(n22638) );
  sky130_fd_sc_hd__clkinv_1 U16543 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[9]), .Y(n25022) );
  sky130_fd_sc_hd__buf_4 U16544 ( .A(j202_soc_core_bootrom_00_address_w[3]), 
        .X(n20788) );
  sky130_fd_sc_hd__clkinv_1 U16545 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[31]), .Y(n28268) );
  sky130_fd_sc_hd__clkinv_1 U16546 ( .A(j202_soc_core_j22_cpu_rf_gbr[8]), .Y(
        n21993) );
  sky130_fd_sc_hd__clkinv_1 U16547 ( .A(j202_soc_core_j22_cpu_ml_macl[31]), 
        .Y(n18295) );
  sky130_fd_sc_hd__clkinv_1 U16548 ( .A(j202_soc_core_qspi_wb_wdat[7]), .Y(
        n28318) );
  sky130_fd_sc_hd__clkinv_1 U16549 ( .A(j202_soc_core_j22_cpu_ml_mach[12]), 
        .Y(n18238) );
  sky130_fd_sc_hd__clkinv_1 U16550 ( .A(j202_soc_core_j22_cpu_ml_mach[20]), 
        .Y(n22072) );
  sky130_fd_sc_hd__clkinv_1 U16551 ( .A(j202_soc_core_intc_core_00_rg_itgt[25]), .Y(n26994) );
  sky130_fd_sc_hd__clkinv_1 U16552 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[103]), .Y(n27076) );
  sky130_fd_sc_hd__clkinv_1 U16553 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[9]), .Y(n24902) );
  sky130_fd_sc_hd__clkinv_1 U16554 ( .A(j202_soc_core_intc_core_00_rg_itgt[35]), .Y(n27806) );
  sky130_fd_sc_hd__clkinv_1 U16555 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[8]), .Y(n23319) );
  sky130_fd_sc_hd__clkinv_1 U16556 ( .A(j202_soc_core_qspi_wb_wdat[6]), .Y(
        n28311) );
  sky130_fd_sc_hd__clkinv_1 U16557 ( .A(j202_soc_core_intc_core_00_rg_ipr[97]), 
        .Y(n27669) );
  sky130_fd_sc_hd__clkinv_1 U16558 ( .A(j202_soc_core_intc_core_00_rg_ie[1]), 
        .Y(n25752) );
  sky130_fd_sc_hd__clkinv_1 U16559 ( .A(j202_soc_core_intc_core_00_rg_ie[20]), 
        .Y(n26485) );
  sky130_fd_sc_hd__clkinv_1 U16560 ( .A(j202_soc_core_j22_cpu_ma_M_address[1]), 
        .Y(n22999) );
  sky130_fd_sc_hd__clkinv_1 U16561 ( .A(j202_soc_core_intc_core_00_rg_ie[18]), 
        .Y(n26822) );
  sky130_fd_sc_hd__clkinv_1 U16562 ( .A(j202_soc_core_j22_cpu_rf_gbr[5]), .Y(
        n21857) );
  sky130_fd_sc_hd__clkinv_1 U16563 ( .A(j202_soc_core_j22_cpu_rf_gbr[2]), .Y(
        n14108) );
  sky130_fd_sc_hd__clkinv_1 U16564 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[1]), 
        .Y(n18920) );
  sky130_fd_sc_hd__clkinv_1 U16565 ( .A(j202_soc_core_intc_core_00_rg_eimk[1]), 
        .Y(n27666) );
  sky130_fd_sc_hd__clkinv_1 U16566 ( .A(j202_soc_core_intc_core_00_rg_itgt[77]), .Y(n26492) );
  sky130_fd_sc_hd__clkinv_1 U16567 ( .A(j202_soc_core_j22_cpu_ml_mach[18]), 
        .Y(n22062) );
  sky130_fd_sc_hd__clkinv_1 U16568 ( .A(j202_soc_core_intc_core_00_rg_eimk[4]), 
        .Y(n26993) );
  sky130_fd_sc_hd__clkinv_1 U16569 ( .A(j202_soc_core_j22_cpu_ml_mach[16]), 
        .Y(n22056) );
  sky130_fd_sc_hd__clkinv_1 U16570 ( .A(j202_soc_core_wbqspiflash_00_spi_in[3]), .Y(n28661) );
  sky130_fd_sc_hd__clkinv_1 U16571 ( .A(j202_soc_core_j22_cpu_ma_M_address[0]), 
        .Y(n18979) );
  sky130_fd_sc_hd__clkinv_1 U16572 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[101]), .Y(n27023) );
  sky130_fd_sc_hd__clkinv_1 U16573 ( .A(j202_soc_core_intc_core_00_rg_eimk[5]), 
        .Y(n26931) );
  sky130_fd_sc_hd__clkinv_1 U16574 ( .A(j202_soc_core_intc_core_00_rg_ie[15]), 
        .Y(n25489) );
  sky130_fd_sc_hd__clkinv_1 U16575 ( .A(j202_soc_core_qspi_wb_wdat[26]), .Y(
        n25114) );
  sky130_fd_sc_hd__clkinv_1 U16576 ( .A(j202_soc_core_j22_cpu_pc[24]), .Y(
        n16028) );
  sky130_fd_sc_hd__clkinv_1 U16577 ( .A(j202_soc_core_j22_cpu_ml_macl[27]), 
        .Y(n18106) );
  sky130_fd_sc_hd__clkinv_1 U16578 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[17]), .Y(n28703) );
  sky130_fd_sc_hd__clkinv_1 U16579 ( .A(j202_soc_core_j22_cpu_ml_mach[30]), 
        .Y(n22465) );
  sky130_fd_sc_hd__clkinv_1 U16580 ( .A(j202_soc_core_aquc_SEL__0_), .Y(n22297) );
  sky130_fd_sc_hd__clkinv_1 U16581 ( .A(j202_soc_core_qspi_wb_wdat[3]), .Y(
        n28291) );
  sky130_fd_sc_hd__clkinv_1 U16582 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[1]), 
        .Y(n28752) );
  sky130_fd_sc_hd__clkinv_1 U16583 ( .A(j202_soc_core_j22_cpu_pc[23]), .Y(
        n15301) );
  sky130_fd_sc_hd__clkinv_1 U16584 ( .A(j202_soc_core_intc_core_00_rg_ie[10]), 
        .Y(n25455) );
  sky130_fd_sc_hd__clkinv_1 U16585 ( .A(j202_soc_core_intc_core_00_rg_itgt[69]), .Y(n26489) );
  sky130_fd_sc_hd__clkinv_1 U16586 ( .A(j202_soc_core_intc_core_00_rg_eimk[6]), 
        .Y(n27534) );
  sky130_fd_sc_hd__clkinv_1 U16587 ( .A(j202_soc_core_j22_cpu_ml_macl[11]), 
        .Y(n23972) );
  sky130_fd_sc_hd__clkinv_1 U16588 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[3]), .Y(n25023) );
  sky130_fd_sc_hd__clkinv_1 U16589 ( .A(j202_soc_core_qspi_wb_wdat[29]), .Y(
        n26969) );
  sky130_fd_sc_hd__clkinv_1 U16590 ( .A(
        j202_soc_core_memory0_ram_dout0_sel[11]), .Y(n13502) );
  sky130_fd_sc_hd__clkinv_1 U16591 ( .A(j202_soc_core_intc_core_00_rg_ipr[26]), 
        .Y(n25088) );
  sky130_fd_sc_hd__clkinv_1 U16592 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[14]), .Y(n23635) );
  sky130_fd_sc_hd__clkinv_1 U16593 ( .A(j202_soc_core_intc_core_00_rg_itgt[70]), .Y(n25090) );
  sky130_fd_sc_hd__clkinv_1 U16594 ( .A(j202_soc_core_intc_core_00_rg_ie[7]), 
        .Y(n25444) );
  sky130_fd_sc_hd__clkinv_1 U16595 ( .A(j202_soc_core_j22_cpu_ml_mach[14]), 
        .Y(n18308) );
  sky130_fd_sc_hd__clkinv_1 U16596 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .Y(n26261) );
  sky130_fd_sc_hd__clkinv_1 U16597 ( .A(j202_soc_core_j22_cpu_ml_macl[0]), .Y(
        n21931) );
  sky130_fd_sc_hd__clkinv_1 U16598 ( .A(j202_soc_core_intc_core_00_rg_ipr[19]), 
        .Y(n25431) );
  sky130_fd_sc_hd__clkinv_1 U16599 ( .A(j202_soc_core_cmt_core_00_cnt0[12]), 
        .Y(n26291) );
  sky130_fd_sc_hd__clkinv_1 U16600 ( .A(j202_soc_core_wbqspiflash_00_spi_valid), .Y(n26476) );
  sky130_fd_sc_hd__clkinv_1 U16601 ( .A(j202_soc_core_qspi_wb_wdat[4]), .Y(
        n28277) );
  sky130_fd_sc_hd__clkinv_1 U16602 ( .A(j202_soc_core_j22_cpu_ml_mach[17]), 
        .Y(n22063) );
  sky130_fd_sc_hd__clkinv_1 U16603 ( .A(j202_soc_core_intc_core_00_rg_ie[6]), 
        .Y(n25437) );
  sky130_fd_sc_hd__clkinv_1 U16604 ( .A(j202_soc_core_j22_cpu_ml_mach[15]), 
        .Y(n18296) );
  sky130_fd_sc_hd__clkinv_1 U16605 ( .A(j202_soc_core_intc_core_00_rg_eimk[2]), 
        .Y(n24974) );
  sky130_fd_sc_hd__clkinv_1 U16606 ( .A(j202_soc_core_j22_cpu_ml_mach[11]), 
        .Y(n18107) );
  sky130_fd_sc_hd__clkinv_1 U16607 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[18]), .Y(n28706) );
  sky130_fd_sc_hd__clkinv_1 U16608 ( .A(j202_soc_core_j22_cpu_pc[18]), .Y(
        n15518) );
  sky130_fd_sc_hd__clkinv_1 U16609 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[2]), .Y(n23317) );
  sky130_fd_sc_hd__clkinv_1 U16610 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[109]), .Y(n27026) );
  sky130_fd_sc_hd__clkinv_1 U16611 ( .A(j202_soc_core_j22_cpu_ml_mach[19]), 
        .Y(n22070) );
  sky130_fd_sc_hd__clkinv_1 U16612 ( .A(j202_soc_core_intc_core_00_rg_itgt[27]), .Y(n26264) );
  sky130_fd_sc_hd__clkinv_1 U16613 ( .A(j202_soc_core_qspi_wb_wdat[22]), .Y(
        n26506) );
  sky130_fd_sc_hd__clkinv_1 U16614 ( .A(j202_soc_core_j22_cpu_ml_mach[21]), 
        .Y(n22073) );
  sky130_fd_sc_hd__clkinv_1 U16615 ( .A(j202_soc_core_j22_cpu_rf_pr[2]), .Y(
        n19202) );
  sky130_fd_sc_hd__clkinv_1 U16616 ( .A(j202_soc_core_intc_core_00_rg_ie[9]), 
        .Y(n25469) );
  sky130_fd_sc_hd__clkinv_1 U16617 ( .A(j202_soc_core_cmt_core_00_cks1[0]), 
        .Y(n23671) );
  sky130_fd_sc_hd__clkinv_1 U16618 ( .A(j202_soc_core_cmt_core_00_cnt1[3]), 
        .Y(n25592) );
  sky130_fd_sc_hd__clkinv_1 U16619 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[102]), .Y(n25644) );
  sky130_fd_sc_hd__clkinv_1 U16620 ( .A(j202_soc_core_intc_core_00_rg_ipr[105]), .Y(n25629) );
  sky130_fd_sc_hd__clkinv_1 U16621 ( .A(j202_soc_core_intc_core_00_rg_itgt[37]), .Y(n25377) );
  sky130_fd_sc_hd__clkinv_1 U16622 ( .A(j202_soc_core_j22_cpu_pc[17]), .Y(
        n21008) );
  sky130_fd_sc_hd__clkinv_1 U16623 ( .A(j202_soc_core_intc_core_00_rg_ie[5]), 
        .Y(n25365) );
  sky130_fd_sc_hd__clkinv_1 U16624 ( .A(j202_soc_core_intc_core_00_rg_itgt[71]), .Y(n27090) );
  sky130_fd_sc_hd__clkinv_1 U16625 ( .A(j202_soc_core_intc_core_00_rg_eimk[3]), 
        .Y(n28521) );
  sky130_fd_sc_hd__clkinv_1 U16626 ( .A(j202_soc_core_intc_core_00_rg_eimk[7]), 
        .Y(n28525) );
  sky130_fd_sc_hd__clkinv_1 U16627 ( .A(j202_soc_core_intc_core_00_rg_ipr[73]), 
        .Y(n25625) );
  sky130_fd_sc_hd__clkinv_1 U16628 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[7]), .Y(n23623) );
  sky130_fd_sc_hd__or2_0 U16629 ( .A(io_in[37]), .B(wb_rst_i), .X(n3) );
  sky130_fd_sc_hd__nand2_1 U16756 ( .A(n13054), .B(n11293), .Y(n27881) );
  sky130_fd_sc_hd__nand2_2 U16757 ( .A(n12732), .B(n12731), .Y(n11293) );
  sky130_fd_sc_hd__nor2_1 U16758 ( .A(n13260), .B(n11294), .Y(n12503) );
  sky130_fd_sc_hd__nand4_1 U16759 ( .A(n20409), .B(n20408), .C(n20407), .D(
        n20404), .Y(n11294) );
  sky130_fd_sc_hd__nand3_1 U16760 ( .A(n13009), .B(n11296), .C(n24253), .Y(
        n23166) );
  sky130_fd_sc_hd__nand2_1 U16761 ( .A(n12475), .B(n27683), .Y(n11296) );
  sky130_fd_sc_hd__nand2b_1 U16762 ( .A_N(n11295), .B(n27552), .Y(n27554) );
  sky130_fd_sc_hd__o21ai_0 U16763 ( .A1(n27553), .A2(n27892), .B1(n11296), .Y(
        n11295) );
  sky130_fd_sc_hd__nor2_1 U16765 ( .A(n11299), .B(n11298), .Y(n11297) );
  sky130_fd_sc_hd__nand4_1 U16766 ( .A(n11304), .B(n11308), .C(n11305), .D(
        n11309), .Y(n11298) );
  sky130_fd_sc_hd__nand4_1 U16767 ( .A(n11306), .B(n11310), .C(n11303), .D(
        n11307), .Y(n11299) );
  sky130_fd_sc_hd__nand4_1 U16769 ( .A(n12014), .B(n12016), .C(n12015), .D(
        n13154), .Y(n11302) );
  sky130_fd_sc_hd__nand2_1 U16770 ( .A(j202_soc_core_memory0_ram_dout0[210]), 
        .B(n21732), .Y(n11303) );
  sky130_fd_sc_hd__nand2_1 U16771 ( .A(j202_soc_core_memory0_ram_dout0[114]), 
        .B(n21591), .Y(n11304) );
  sky130_fd_sc_hd__nand2_1 U16772 ( .A(j202_soc_core_memory0_ram_dout0[370]), 
        .B(n21596), .Y(n11305) );
  sky130_fd_sc_hd__nand2_1 U16773 ( .A(j202_soc_core_memory0_ram_dout0[434]), 
        .B(n21598), .Y(n11306) );
  sky130_fd_sc_hd__nand2_1 U16774 ( .A(j202_soc_core_memory0_ram_dout0[242]), 
        .B(n21735), .Y(n11307) );
  sky130_fd_sc_hd__nand2_1 U16775 ( .A(j202_soc_core_memory0_ram_dout0[18]), 
        .B(n21733), .Y(n11308) );
  sky130_fd_sc_hd__nand2_1 U16776 ( .A(j202_soc_core_memory0_ram_dout0[50]), 
        .B(n21604), .Y(n11309) );
  sky130_fd_sc_hd__nand2_1 U16777 ( .A(j202_soc_core_memory0_ram_dout0[178]), 
        .B(n21590), .Y(n11310) );
  sky130_fd_sc_hd__inv_1 U16778 ( .A(n20031), .Y(n11311) );
  sky130_fd_sc_hd__inv_1 U16779 ( .A(n11340), .Y(n11312) );
  sky130_fd_sc_hd__nand2_1 U16782 ( .A(n20715), .B(n29572), .Y(n11314) );
  sky130_fd_sc_hd__inv_1 U16784 ( .A(n12889), .Y(n11316) );
  sky130_fd_sc_hd__nand2_1 U16785 ( .A(n20718), .B(n11056), .Y(n11317) );
  sky130_fd_sc_hd__nand2_1 U16788 ( .A(n13157), .B(n13156), .Y(n11318) );
  sky130_fd_sc_hd__nand4_1 U16789 ( .A(n19934), .B(n19933), .C(n19932), .D(
        n19931), .Y(n13157) );
  sky130_fd_sc_hd__nand2_1 U16791 ( .A(n13155), .B(n20708), .Y(n11320) );
  sky130_fd_sc_hd__nand4_1 U16792 ( .A(n11643), .B(n19930), .C(n19929), .D(
        n19927), .Y(n11321) );
  sky130_fd_sc_hd__nand2_1 U16793 ( .A(n21007), .B(n12282), .Y(n11322) );
  sky130_fd_sc_hd__nand3_4 U16795 ( .A(n11324), .B(n20561), .C(n11323), .Y(
        n22278) );
  sky130_fd_sc_hd__nand2_1 U16797 ( .A(n11345), .B(n11348), .Y(n20988) );
  sky130_fd_sc_hd__nand2_1 U16798 ( .A(n11378), .B(n11387), .Y(n13008) );
  sky130_fd_sc_hd__nand3_1 U16799 ( .A(n27893), .B(n23208), .C(n24388), .Y(
        n23206) );
  sky130_fd_sc_hd__nand2_1 U16800 ( .A(n12732), .B(n11626), .Y(n27893) );
  sky130_fd_sc_hd__nor2_1 U16802 ( .A(n24265), .B(n27556), .Y(n11325) );
  sky130_fd_sc_hd__nand2_1 U16804 ( .A(n27556), .B(n24350), .Y(n12046) );
  sky130_fd_sc_hd__nand2_1 U16805 ( .A(n11326), .B(n23606), .Y(n11818) );
  sky130_fd_sc_hd__nand2_1 U16807 ( .A(n11337), .B(n11327), .Y(n20712) );
  sky130_fd_sc_hd__nand4_1 U16808 ( .A(n11332), .B(n11331), .C(n11330), .D(
        n11329), .Y(n11328) );
  sky130_fd_sc_hd__nand2_1 U16809 ( .A(j202_soc_core_memory0_ram_dout0[162]), 
        .B(n21590), .Y(n11329) );
  sky130_fd_sc_hd__nand2_1 U16810 ( .A(j202_soc_core_memory0_ram_dout0[34]), 
        .B(n21604), .Y(n11330) );
  sky130_fd_sc_hd__nand2_1 U16811 ( .A(j202_soc_core_memory0_ram_dout0[2]), 
        .B(n21733), .Y(n11331) );
  sky130_fd_sc_hd__nand2_1 U16812 ( .A(j202_soc_core_memory0_ram_dout0[130]), 
        .B(n21592), .Y(n11332) );
  sky130_fd_sc_hd__nand4_1 U16813 ( .A(n17241), .B(n11336), .C(n11335), .D(
        n11334), .Y(n11333) );
  sky130_fd_sc_hd__nand2_1 U16814 ( .A(j202_soc_core_memory0_ram_dout0[66]), 
        .B(n21734), .Y(n11334) );
  sky130_fd_sc_hd__nand2_1 U16815 ( .A(j202_soc_core_memory0_ram_dout0[98]), 
        .B(n21591), .Y(n11335) );
  sky130_fd_sc_hd__nand2_1 U16816 ( .A(j202_soc_core_memory0_ram_dout0[194]), 
        .B(n21732), .Y(n11336) );
  sky130_fd_sc_hd__nand4_1 U16817 ( .A(n13183), .B(n13184), .C(n17239), .D(
        n17240), .Y(n11338) );
  sky130_fd_sc_hd__nand4_1 U16818 ( .A(n13010), .B(n12620), .C(n13185), .D(
        n17238), .Y(n11339) );
  sky130_fd_sc_hd__nand4_1 U16819 ( .A(n11343), .B(n11342), .C(n11341), .D(
        n20027), .Y(n11340) );
  sky130_fd_sc_hd__nand2_1 U16820 ( .A(j202_soc_core_memory0_ram_dout0[419]), 
        .B(n21598), .Y(n11341) );
  sky130_fd_sc_hd__nand2_1 U16821 ( .A(j202_soc_core_memory0_ram_dout0[355]), 
        .B(n21596), .Y(n11342) );
  sky130_fd_sc_hd__nand2_1 U16822 ( .A(j202_soc_core_memory0_ram_dout0[451]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11343) );
  sky130_fd_sc_hd__nor2_1 U16824 ( .A(n29071), .B(n12692), .Y(n22279) );
  sky130_fd_sc_hd__nand2_4 U16825 ( .A(n29070), .B(n13180), .Y(n12692) );
  sky130_fd_sc_hd__nand2_1 U16826 ( .A(n22102), .B(n11478), .Y(n11473) );
  sky130_fd_sc_hd__nand2_1 U16827 ( .A(n11344), .B(n22100), .Y(n22102) );
  sky130_fd_sc_hd__nand2_1 U16828 ( .A(n22130), .B(n22101), .Y(n11344) );
  sky130_fd_sc_hd__nand4_1 U16830 ( .A(n11358), .B(n11354), .C(n11356), .D(
        n11355), .Y(n11346) );
  sky130_fd_sc_hd__nor2_1 U16832 ( .A(n11350), .B(n11349), .Y(n11348) );
  sky130_fd_sc_hd__nand4_1 U16833 ( .A(n20545), .B(n20433), .C(n20544), .D(
        n20546), .Y(n11349) );
  sky130_fd_sc_hd__nand4_1 U16834 ( .A(n11702), .B(n20431), .C(n20432), .D(
        n12803), .Y(n11350) );
  sky130_fd_sc_hd__nand2_1 U16836 ( .A(j202_soc_core_memory0_ram_dout0[432]), 
        .B(n21598), .Y(n11352) );
  sky130_fd_sc_hd__nand2_1 U16837 ( .A(j202_soc_core_memory0_ram_dout0[80]), 
        .B(n21734), .Y(n11353) );
  sky130_fd_sc_hd__nand2_1 U16838 ( .A(j202_soc_core_memory0_ram_dout0[272]), 
        .B(n21605), .Y(n11355) );
  sky130_fd_sc_hd__nand2_1 U16839 ( .A(j202_soc_core_memory0_ram_dout0[336]), 
        .B(n21593), .Y(n11356) );
  sky130_fd_sc_hd__nand2_1 U16840 ( .A(j202_soc_core_memory0_ram_dout0[176]), 
        .B(n21590), .Y(n11357) );
  sky130_fd_sc_hd__nand2_1 U16841 ( .A(j202_soc_core_memory0_ram_dout0[464]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11358) );
  sky130_fd_sc_hd__nand2_1 U16842 ( .A(n26400), .B(n29496), .Y(n26404) );
  sky130_fd_sc_hd__nand2_1 U16844 ( .A(n11361), .B(n26863), .Y(n26399) );
  sky130_fd_sc_hd__xnor2_1 U16845 ( .A(n22664), .B(n22663), .Y(n11361) );
  sky130_fd_sc_hd__nand2_1 U16846 ( .A(n22399), .B(n12928), .Y(n12927) );
  sky130_fd_sc_hd__nand2_1 U16847 ( .A(n22399), .B(n22421), .Y(n12926) );
  sky130_fd_sc_hd__nand2_1 U16848 ( .A(n11362), .B(n22428), .Y(n22430) );
  sky130_fd_sc_hd__nand2_1 U16849 ( .A(n22399), .B(n22469), .Y(n11362) );
  sky130_fd_sc_hd__nand2_1 U16850 ( .A(n22478), .B(n11363), .Y(n22399) );
  sky130_fd_sc_hd__nand2_1 U16851 ( .A(n22398), .B(n22470), .Y(n11363) );
  sky130_fd_sc_hd__nand2_1 U16852 ( .A(n11366), .B(n11364), .Y(n18911) );
  sky130_fd_sc_hd__nand2_1 U16853 ( .A(n11365), .B(n21430), .Y(n19444) );
  sky130_fd_sc_hd__nand2_1 U16854 ( .A(n11142), .B(n21431), .Y(n11365) );
  sky130_fd_sc_hd__inv_1 U16855 ( .A(n11368), .Y(n11367) );
  sky130_fd_sc_hd__nand2_1 U16856 ( .A(n21802), .B(n11493), .Y(n11368) );
  sky130_fd_sc_hd__o21a_1 U16857 ( .A1(n21504), .A2(n17897), .B1(n18888), .X(
        n11494) );
  sky130_fd_sc_hd__nand2_1 U16859 ( .A(n11371), .B(n24771), .Y(n11370) );
  sky130_fd_sc_hd__nand2_1 U16860 ( .A(n25250), .B(n12699), .Y(n11371) );
  sky130_fd_sc_hd__o21a_1 U16861 ( .A1(n24798), .A2(n25251), .B1(n11373), .X(
        n11372) );
  sky130_fd_sc_hd__nand2_1 U16862 ( .A(n23237), .B(n24499), .Y(n25251) );
  sky130_fd_sc_hd__nand2_1 U16863 ( .A(n11375), .B(n11374), .Y(n17959) );
  sky130_fd_sc_hd__nand2_1 U16864 ( .A(n17485), .B(n17486), .Y(n11374) );
  sky130_fd_sc_hd__xnor2_1 U16866 ( .A(n17485), .B(n11376), .Y(n17517) );
  sky130_fd_sc_hd__xnor2_1 U16867 ( .A(n17486), .B(n17484), .Y(n11376) );
  sky130_fd_sc_hd__nor2_1 U16868 ( .A(n29546), .B(n27298), .Y(n22281) );
  sky130_fd_sc_hd__nand2_1 U16870 ( .A(n13272), .B(n27556), .Y(n13274) );
  sky130_fd_sc_hd__nand2_1 U16872 ( .A(n13056), .B(n29546), .Y(n13055) );
  sky130_fd_sc_hd__nand2_1 U16873 ( .A(n11849), .B(n29546), .Y(n11867) );
  sky130_fd_sc_hd__nor2_2 U16874 ( .A(n17928), .B(n17929), .Y(n21808) );
  sky130_fd_sc_hd__nor2_1 U16875 ( .A(n11384), .B(n11379), .Y(n11378) );
  sky130_fd_sc_hd__nand4_1 U16876 ( .A(n11383), .B(n11382), .C(n11381), .D(
        n11380), .Y(n11379) );
  sky130_fd_sc_hd__nand2_1 U16877 ( .A(j202_soc_core_memory0_ram_dout0[32]), 
        .B(n21604), .Y(n11380) );
  sky130_fd_sc_hd__nand2_1 U16878 ( .A(j202_soc_core_memory0_ram_dout0[64]), 
        .B(n21734), .Y(n11381) );
  sky130_fd_sc_hd__nand2_2 U16880 ( .A(j202_soc_core_memory0_ram_dout0[256]), 
        .B(n21605), .Y(n11383) );
  sky130_fd_sc_hd__nand4_1 U16881 ( .A(n12002), .B(n12003), .C(n11386), .D(
        n11385), .Y(n11384) );
  sky130_fd_sc_hd__nand2_1 U16882 ( .A(j202_soc_core_memory0_ram_dout0[192]), 
        .B(n21732), .Y(n11385) );
  sky130_fd_sc_hd__nand2_1 U16883 ( .A(j202_soc_core_memory0_ram_dout0[352]), 
        .B(n21596), .Y(n11386) );
  sky130_fd_sc_hd__nor2_1 U16884 ( .A(n11389), .B(n11388), .Y(n11387) );
  sky130_fd_sc_hd__nand4_1 U16885 ( .A(n12808), .B(n12807), .C(n12806), .D(
        n12805), .Y(n11388) );
  sky130_fd_sc_hd__nand4_1 U16886 ( .A(n13117), .B(n13118), .C(n13119), .D(
        n12241), .Y(n11389) );
  sky130_fd_sc_hd__nand2b_4 U16888 ( .A_N(n11390), .B(n20977), .Y(n12501) );
  sky130_fd_sc_hd__nand2_1 U16889 ( .A(n11794), .B(n11827), .Y(n11390) );
  sky130_fd_sc_hd__nand3_2 U16890 ( .A(n11891), .B(n22674), .C(n12898), .Y(
        n11391) );
  sky130_fd_sc_hd__nand2_1 U16891 ( .A(n11391), .B(n29594), .Y(n12492) );
  sky130_fd_sc_hd__nand3_2 U16893 ( .A(n11133), .B(n11392), .C(n29077), .Y(
        n27957) );
  sky130_fd_sc_hd__o21a_1 U16894 ( .A1(n11133), .A2(n23589), .B1(n11392), .X(
        n24108) );
  sky130_fd_sc_hd__inv_2 U16896 ( .A(n11842), .Y(n11392) );
  sky130_fd_sc_hd__nand3_1 U16897 ( .A(n28924), .B(n28957), .C(n29518), .Y(
        n12626) );
  sky130_fd_sc_hd__nand3_2 U16898 ( .A(n11395), .B(n15214), .C(n15213), .Y(
        n28924) );
  sky130_fd_sc_hd__inv_2 U16899 ( .A(n21916), .Y(n23731) );
  sky130_fd_sc_hd__inv_1 U16900 ( .A(n11396), .Y(n27558) );
  sky130_fd_sc_hd__nor2_1 U16901 ( .A(n23161), .B(n11396), .Y(n27561) );
  sky130_fd_sc_hd__o2bb2ai_1 U16902 ( .B1(n11396), .B2(n27685), .A1_N(n12742), 
        .A2_N(n27683), .Y(n27689) );
  sky130_fd_sc_hd__nand2_1 U16903 ( .A(n12394), .B(n23143), .Y(n11396) );
  sky130_fd_sc_hd__nand4_1 U16904 ( .A(n11402), .B(n11401), .C(n11400), .D(
        n11399), .Y(n11398) );
  sky130_fd_sc_hd__nand2_1 U16905 ( .A(j202_soc_core_memory0_ram_dout0[120]), 
        .B(n21591), .Y(n11399) );
  sky130_fd_sc_hd__nand2_1 U16906 ( .A(j202_soc_core_memory0_ram_dout0[184]), 
        .B(n21590), .Y(n11400) );
  sky130_fd_sc_hd__nand2_1 U16907 ( .A(j202_soc_core_memory0_ram_dout0[472]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11401) );
  sky130_fd_sc_hd__nand2_1 U16908 ( .A(j202_soc_core_memory0_ram_dout0[344]), 
        .B(n21593), .Y(n11402) );
  sky130_fd_sc_hd__nand4_1 U16909 ( .A(n13106), .B(n13111), .C(n11405), .D(
        n11404), .Y(n11403) );
  sky130_fd_sc_hd__nand2_1 U16910 ( .A(j202_soc_core_memory0_ram_dout0[152]), 
        .B(n21592), .Y(n11404) );
  sky130_fd_sc_hd__nand2_1 U16911 ( .A(j202_soc_core_memory0_ram_dout0[312]), 
        .B(n21603), .Y(n11405) );
  sky130_fd_sc_hd__nand4_1 U16912 ( .A(n13108), .B(n13114), .C(n13113), .D(
        n13112), .Y(n11407) );
  sky130_fd_sc_hd__nand4_1 U16913 ( .A(n13110), .B(n13109), .C(n13107), .D(
        n14970), .Y(n11408) );
  sky130_fd_sc_hd__nor2_1 U16915 ( .A(n11555), .B(n11661), .Y(n11409) );
  sky130_fd_sc_hd__nand2_2 U16916 ( .A(n23797), .B(n12352), .Y(n11661) );
  sky130_fd_sc_hd__nand2_1 U16918 ( .A(n11410), .B(n26323), .Y(n18991) );
  sky130_fd_sc_hd__nand2_1 U16919 ( .A(n11410), .B(n26729), .Y(n26601) );
  sky130_fd_sc_hd__o21a_1 U16920 ( .A1(n26729), .A2(n11410), .B1(n24481), .X(
        n12454) );
  sky130_fd_sc_hd__nand2_2 U16921 ( .A(n26552), .B(n23045), .Y(n11410) );
  sky130_fd_sc_hd__nand2_1 U16922 ( .A(n11411), .B(n26443), .Y(n26444) );
  sky130_fd_sc_hd__xnor2_1 U16923 ( .A(n26705), .B(n26557), .Y(n11411) );
  sky130_fd_sc_hd__nand2_1 U16924 ( .A(n11412), .B(n11414), .Y(n18808) );
  sky130_fd_sc_hd__nand2b_1 U16925 ( .A_N(n11417), .B(n11421), .Y(n11413) );
  sky130_fd_sc_hd__nand3_1 U16926 ( .A(n11421), .B(n18593), .C(n11420), .Y(
        n11414) );
  sky130_fd_sc_hd__xor2_1 U16928 ( .A(n11416), .B(n18562), .X(n11419) );
  sky130_fd_sc_hd__nand2_1 U16929 ( .A(n11419), .B(n11418), .Y(n11420) );
  sky130_fd_sc_hd__nand2_1 U16930 ( .A(n12947), .B(n12946), .Y(n11418) );
  sky130_fd_sc_hd__nand2_1 U16931 ( .A(n11422), .B(n18595), .Y(n11421) );
  sky130_fd_sc_hd__nand2_1 U16932 ( .A(n12947), .B(n12946), .Y(n18594) );
  sky130_fd_sc_hd__xnor2_1 U16933 ( .A(n18247), .B(n11423), .Y(n18249) );
  sky130_fd_sc_hd__xnor2_1 U16934 ( .A(n18246), .B(n18245), .Y(n11423) );
  sky130_fd_sc_hd__xor2_1 U16935 ( .A(n25403), .B(n24087), .X(n24089) );
  sky130_fd_sc_hd__nor2_1 U16936 ( .A(n11424), .B(n12353), .Y(n24087) );
  sky130_fd_sc_hd__xnor2_1 U16937 ( .A(n18746), .B(n18745), .Y(n11585) );
  sky130_fd_sc_hd__nand2_1 U16938 ( .A(n11426), .B(n11425), .Y(n18690) );
  sky130_fd_sc_hd__nand2_1 U16939 ( .A(n18677), .B(n11428), .Y(n11425) );
  sky130_fd_sc_hd__xnor2_1 U16941 ( .A(n18676), .B(n11427), .Y(n18739) );
  sky130_fd_sc_hd__xnor2_1 U16942 ( .A(n11428), .B(n18677), .Y(n11427) );
  sky130_fd_sc_hd__o22ai_2 U16943 ( .A1(n18719), .A2(n18666), .B1(n18665), 
        .B2(n11514), .Y(n11428) );
  sky130_fd_sc_hd__o21ai_2 U16944 ( .A1(n22907), .A2(n18848), .B1(n18847), .Y(
        n22398) );
  sky130_fd_sc_hd__inv_2 U16945 ( .A(n22398), .Y(n22619) );
  sky130_fd_sc_hd__nand2_1 U16946 ( .A(n18846), .B(n19227), .Y(n18848) );
  sky130_fd_sc_hd__nand2_1 U16947 ( .A(n22480), .B(n22398), .Y(n12713) );
  sky130_fd_sc_hd__nand2_1 U16948 ( .A(n11431), .B(n11430), .Y(n12166) );
  sky130_fd_sc_hd__xnor2_1 U16949 ( .A(n18596), .B(n11432), .Y(n18614) );
  sky130_fd_sc_hd__xnor2_1 U16950 ( .A(n18597), .B(n18598), .Y(n11432) );
  sky130_fd_sc_hd__xor2_1 U16951 ( .A(n18395), .B(n11433), .X(n18596) );
  sky130_fd_sc_hd__xor2_1 U16952 ( .A(n18394), .B(n18393), .X(n11433) );
  sky130_fd_sc_hd__nand2_1 U16953 ( .A(n11435), .B(n11434), .Y(n18778) );
  sky130_fd_sc_hd__nand2_1 U16954 ( .A(n18773), .B(n18772), .Y(n11434) );
  sky130_fd_sc_hd__o21ai_1 U16955 ( .A1(n18772), .A2(n18773), .B1(n18771), .Y(
        n11435) );
  sky130_fd_sc_hd__xor2_1 U16956 ( .A(n11437), .B(n11436), .X(n18781) );
  sky130_fd_sc_hd__xnor2_1 U16957 ( .A(n18772), .B(n18771), .Y(n11436) );
  sky130_fd_sc_hd__nand2_1 U16958 ( .A(n22949), .B(n26863), .Y(n25663) );
  sky130_fd_sc_hd__nand2_1 U16959 ( .A(n21798), .B(n11438), .Y(n21800) );
  sky130_fd_sc_hd__nand2_1 U16960 ( .A(n19249), .B(n21799), .Y(n11438) );
  sky130_fd_sc_hd__o21ai_1 U16961 ( .A1(n18906), .A2(n11439), .B1(n18905), .Y(
        n18907) );
  sky130_fd_sc_hd__o21ai_1 U16962 ( .A1(n22527), .A2(n11439), .B1(n22526), .Y(
        n22528) );
  sky130_fd_sc_hd__o21ai_1 U16964 ( .A1(n18858), .A2(n11439), .B1(n18857), .Y(
        n18859) );
  sky130_fd_sc_hd__inv_2 U16965 ( .A(n19249), .Y(n11439) );
  sky130_fd_sc_hd__inv_2 U16966 ( .A(n11440), .Y(n17772) );
  sky130_fd_sc_hd__xnor2_1 U16967 ( .A(n11440), .B(n18511), .Y(n17709) );
  sky130_fd_sc_hd__xnor2_1 U16968 ( .A(n11440), .B(n18667), .Y(n17698) );
  sky130_fd_sc_hd__xnor2_1 U16969 ( .A(n11440), .B(n18226), .Y(n17767) );
  sky130_fd_sc_hd__xnor2_1 U16970 ( .A(n11440), .B(n18466), .Y(n17751) );
  sky130_fd_sc_hd__xnor2_1 U16971 ( .A(n11440), .B(n18673), .Y(n17537) );
  sky130_fd_sc_hd__xnor2_1 U16972 ( .A(n11440), .B(n18426), .Y(n17765) );
  sky130_fd_sc_hd__xnor2_1 U16973 ( .A(n11440), .B(n18685), .Y(n17538) );
  sky130_fd_sc_hd__xnor2_1 U16974 ( .A(n11440), .B(n22052), .Y(n17504) );
  sky130_fd_sc_hd__xnor2_1 U16975 ( .A(n11440), .B(n18651), .Y(n17472) );
  sky130_fd_sc_hd__xnor2_1 U16976 ( .A(n11440), .B(n18479), .Y(n17716) );
  sky130_fd_sc_hd__xnor2_1 U16977 ( .A(n11440), .B(n18661), .Y(n17579) );
  sky130_fd_sc_hd__xnor2_1 U16978 ( .A(n11440), .B(n18708), .Y(n17657) );
  sky130_fd_sc_hd__xnor2_1 U16979 ( .A(n11440), .B(n18654), .Y(n17656) );
  sky130_fd_sc_hd__xnor2_1 U16980 ( .A(n11440), .B(n18649), .Y(n17644) );
  sky130_fd_sc_hd__xnor2_1 U16981 ( .A(n11440), .B(n18721), .Y(n17464) );
  sky130_fd_sc_hd__xnor2_1 U16982 ( .A(n11440), .B(n18687), .Y(n17452) );
  sky130_fd_sc_hd__xnor2_1 U16983 ( .A(n11440), .B(n18367), .Y(n17768) );
  sky130_fd_sc_hd__nand2_1 U16984 ( .A(n27187), .B(n11440), .Y(n12783) );
  sky130_fd_sc_hd__nor2b_1 U16985 ( .B_N(n11440), .A(n21972), .Y(n11442) );
  sky130_fd_sc_hd__nand2_4 U16986 ( .A(n11444), .B(n27047), .Y(n27189) );
  sky130_fd_sc_hd__inv_2 U16987 ( .A(n23256), .Y(n11444) );
  sky130_fd_sc_hd__nand3_2 U16988 ( .A(n23269), .B(n23267), .C(n12990), .Y(
        n23256) );
  sky130_fd_sc_hd__nand3_2 U16989 ( .A(n12680), .B(n23251), .C(n23250), .Y(
        n12990) );
  sky130_fd_sc_hd__nand2_1 U16990 ( .A(n11446), .B(n11445), .Y(n18027) );
  sky130_fd_sc_hd__nand2_1 U16991 ( .A(n17994), .B(n17993), .Y(n11445) );
  sky130_fd_sc_hd__o21ai_1 U16992 ( .A1(n17994), .A2(n17993), .B1(n17992), .Y(
        n11446) );
  sky130_fd_sc_hd__xor2_1 U16993 ( .A(n17994), .B(n11447), .X(n18081) );
  sky130_fd_sc_hd__xor2_1 U16994 ( .A(n17993), .B(n17992), .X(n11447) );
  sky130_fd_sc_hd__nand2_1 U16995 ( .A(n11450), .B(n11449), .Y(n11448) );
  sky130_fd_sc_hd__nand2_1 U16996 ( .A(n11456), .B(n22619), .Y(n11450) );
  sky130_fd_sc_hd__nand2_1 U16997 ( .A(n11453), .B(n11457), .Y(n11452) );
  sky130_fd_sc_hd__inv_6 U16998 ( .A(n19249), .Y(n22897) );
  sky130_fd_sc_hd__nand3_1 U16999 ( .A(n19249), .B(n22471), .C(n12321), .Y(
        n11456) );
  sky130_fd_sc_hd__nand2_1 U17000 ( .A(n22661), .B(n22471), .Y(n11457) );
  sky130_fd_sc_hd__nand2_1 U17001 ( .A(n24806), .B(n11458), .Y(
        j202_soc_core_j22_cpu_ml_maclj[2]) );
  sky130_fd_sc_hd__nand3_1 U17002 ( .A(n11461), .B(n11460), .C(n25822), .Y(
        n11459) );
  sky130_fd_sc_hd__nand3_4 U17003 ( .A(n12487), .B(n23254), .C(n23268), .Y(
        n25822) );
  sky130_fd_sc_hd__nand2_1 U17004 ( .A(n12357), .B(n11462), .Y(n11461) );
  sky130_fd_sc_hd__nand3_2 U17005 ( .A(n12990), .B(n26878), .C(n23269), .Y(
        n12357) );
  sky130_fd_sc_hd__nand3_4 U17006 ( .A(n23227), .B(n23229), .C(n23228), .Y(
        n23269) );
  sky130_fd_sc_hd__inv_1 U17007 ( .A(n11463), .Y(n25116) );
  sky130_fd_sc_hd__nand2_2 U17008 ( .A(n11546), .B(n26548), .Y(n12352) );
  sky130_fd_sc_hd__nand2_1 U17010 ( .A(n26100), .B(n26443), .Y(n11465) );
  sky130_fd_sc_hd__nand2_1 U17011 ( .A(n11466), .B(n26859), .Y(n11485) );
  sky130_fd_sc_hd__nand2_1 U17012 ( .A(n11467), .B(n12596), .Y(n11466) );
  sky130_fd_sc_hd__nand2_1 U17013 ( .A(n27340), .B(n26323), .Y(n11467) );
  sky130_fd_sc_hd__nand3_2 U17014 ( .A(n11471), .B(n11483), .C(n11468), .Y(
        n26881) );
  sky130_fd_sc_hd__nand2_1 U17015 ( .A(n24997), .B(n26329), .Y(n11468) );
  sky130_fd_sc_hd__nand2_1 U17016 ( .A(n26864), .B(n22627), .Y(n11469) );
  sky130_fd_sc_hd__nand2_1 U17017 ( .A(n12706), .B(n24478), .Y(n11470) );
  sky130_fd_sc_hd__nand2_1 U17018 ( .A(n11485), .B(n11484), .Y(n11472) );
  sky130_fd_sc_hd__nand3_1 U17019 ( .A(n12713), .B(n11477), .C(n22616), .Y(
        n22481) );
  sky130_fd_sc_hd__nand2b_1 U17020 ( .A_N(n22618), .B(n11147), .Y(n11477) );
  sky130_fd_sc_hd__nand2_1 U17021 ( .A(n11480), .B(n11479), .Y(n22066) );
  sky130_fd_sc_hd__nand2_1 U17022 ( .A(n22058), .B(n11481), .Y(n11479) );
  sky130_fd_sc_hd__o21ai_1 U17023 ( .A1(n11481), .A2(n22058), .B1(n22057), .Y(
        n11480) );
  sky130_fd_sc_hd__xor2_1 U17024 ( .A(n22058), .B(n11482), .X(n22059) );
  sky130_fd_sc_hd__xnor2_1 U17025 ( .A(n22057), .B(n17376), .Y(n11482) );
  sky130_fd_sc_hd__nand3_1 U17026 ( .A(n11483), .B(n11484), .C(n11485), .Y(
        n25000) );
  sky130_fd_sc_hd__a21oi_1 U17027 ( .A1(n27340), .A2(n26406), .B1(n23939), .Y(
        n11484) );
  sky130_fd_sc_hd__nand3_1 U17028 ( .A(n11486), .B(n12352), .C(n11547), .Y(
        n11520) );
  sky130_fd_sc_hd__nand2_1 U17029 ( .A(n11487), .B(n11054), .Y(n11488) );
  sky130_fd_sc_hd__nand2_1 U17030 ( .A(n19463), .B(n17892), .Y(n11487) );
  sky130_fd_sc_hd__o21ai_1 U17031 ( .A1(n21803), .A2(n21808), .B1(n21809), .Y(
        n11492) );
  sky130_fd_sc_hd__inv_2 U17032 ( .A(n12317), .Y(n21802) );
  sky130_fd_sc_hd__inv_2 U17033 ( .A(n21462), .Y(n11496) );
  sky130_fd_sc_hd__nand2_1 U17034 ( .A(n17866), .B(n17867), .Y(n21462) );
  sky130_fd_sc_hd__nand2_1 U17036 ( .A(n17865), .B(n17864), .Y(n19240) );
  sky130_fd_sc_hd__clkinv_1 U17037 ( .A(n17866), .Y(n11497) );
  sky130_fd_sc_hd__xor2_1 U17038 ( .A(n11499), .B(n17781), .X(n17849) );
  sky130_fd_sc_hd__nand2_1 U17039 ( .A(n11501), .B(n11500), .Y(n17762) );
  sky130_fd_sc_hd__nand2_1 U17040 ( .A(n17759), .B(n17760), .Y(n11500) );
  sky130_fd_sc_hd__xnor2_1 U17042 ( .A(n17758), .B(n11502), .Y(n17857) );
  sky130_fd_sc_hd__xnor2_1 U17043 ( .A(n17760), .B(n17759), .Y(n11502) );
  sky130_fd_sc_hd__xnor2_1 U17044 ( .A(j202_soc_core_j22_cpu_ml_bufa[5]), .B(
        j202_soc_core_j22_cpu_ml_bufa[6]), .Y(n17387) );
  sky130_fd_sc_hd__o21a_2 U17045 ( .A1(n18916), .A2(n25193), .B1(n25140), .X(
        n25222) );
  sky130_fd_sc_hd__inv_2 U17046 ( .A(n11504), .Y(n25156) );
  sky130_fd_sc_hd__nand2_1 U17047 ( .A(n23010), .B(n23009), .Y(n11791) );
  sky130_fd_sc_hd__nand2_1 U17048 ( .A(n11505), .B(n26863), .Y(n25143) );
  sky130_fd_sc_hd__xnor2_1 U17049 ( .A(n22684), .B(n11506), .Y(n11505) );
  sky130_fd_sc_hd__nand3_1 U17050 ( .A(n22683), .B(n12321), .C(n19249), .Y(
        n11507) );
  sky130_fd_sc_hd__nand2_1 U17051 ( .A(n22683), .B(n22944), .Y(n11508) );
  sky130_fd_sc_hd__nand2_1 U17052 ( .A(n22131), .B(n22101), .Y(n22389) );
  sky130_fd_sc_hd__nor2_4 U17053 ( .A(n18848), .B(n22905), .Y(n22471) );
  sky130_fd_sc_hd__nand2_1 U17054 ( .A(n22965), .B(
        j202_soc_core_j22_cpu_ml_bufa[28]), .Y(n26396) );
  sky130_fd_sc_hd__a22oi_1 U17055 ( .A1(j202_soc_core_j22_cpu_ml_bufa[28]), 
        .A2(n27187), .B1(n24548), .B2(n27047), .Y(n24549) );
  sky130_fd_sc_hd__nand2_1 U17056 ( .A(n11509), .B(n29495), .Y(n11532) );
  sky130_fd_sc_hd__nand2_1 U17057 ( .A(n11104), .B(n12495), .Y(n11509) );
  sky130_fd_sc_hd__o22ai_1 U17058 ( .A1(n18719), .A2(n18303), .B1(n18302), 
        .B2(n11514), .Y(n18349) );
  sky130_fd_sc_hd__nand2_1 U17059 ( .A(n17369), .B(n11510), .Y(n22057) );
  sky130_fd_sc_hd__nand2_1 U17060 ( .A(n11514), .B(n18719), .Y(n11510) );
  sky130_fd_sc_hd__o22ai_1 U17061 ( .A1(n18719), .A2(n18446), .B1(n18423), 
        .B2(n11514), .Y(n18453) );
  sky130_fd_sc_hd__o22ai_1 U17062 ( .A1(n18719), .A2(n18423), .B1(n18374), 
        .B2(n11514), .Y(n18409) );
  sky130_fd_sc_hd__o22ai_1 U17063 ( .A1(n18719), .A2(n18717), .B1(n18653), 
        .B2(n11514), .Y(n18704) );
  sky130_fd_sc_hd__o22ai_1 U17064 ( .A1(n18719), .A2(n18631), .B1(n18718), 
        .B2(n11514), .Y(n18764) );
  sky130_fd_sc_hd__o22ai_1 U17066 ( .A1(n18719), .A2(n18623), .B1(n18631), 
        .B2(n11514), .Y(n18637) );
  sky130_fd_sc_hd__o22ai_1 U17067 ( .A1(n18719), .A2(n17380), .B1(n18623), 
        .B2(n11514), .Y(n18630) );
  sky130_fd_sc_hd__o22ai_1 U17068 ( .A1(n18719), .A2(n18718), .B1(n18717), 
        .B2(n11514), .Y(n18760) );
  sky130_fd_sc_hd__o22ai_1 U17069 ( .A1(n18719), .A2(n18653), .B1(n18666), 
        .B2(n11514), .Y(n18696) );
  sky130_fd_sc_hd__o22ai_1 U17070 ( .A1(n18719), .A2(n17378), .B1(n17380), 
        .B2(n11514), .Y(n18627) );
  sky130_fd_sc_hd__o22ai_1 U17071 ( .A1(n18719), .A2(n18665), .B1(n11514), 
        .B2(n18538), .Y(n18683) );
  sky130_fd_sc_hd__o22ai_1 U17072 ( .A1(n11514), .A2(n18446), .B1(n18719), 
        .B2(n18505), .Y(n18499) );
  sky130_fd_sc_hd__nand2_1 U17073 ( .A(n11512), .B(n11511), .Y(n18535) );
  sky130_fd_sc_hd__nand2b_1 U17074 ( .A_N(n18538), .B(n11162), .Y(n11511) );
  sky130_fd_sc_hd__nand2b_1 U17075 ( .A_N(n18505), .B(n11513), .Y(n11512) );
  sky130_fd_sc_hd__nand2_4 U17076 ( .A(n18719), .B(n17364), .Y(n11514) );
  sky130_fd_sc_hd__nand3_2 U17077 ( .A(n11515), .B(n11139), .C(n11140), .Y(
        n18826) );
  sky130_fd_sc_hd__nor2_2 U17078 ( .A(n18820), .B(n12320), .Y(n21794) );
  sky130_fd_sc_hd__nor2_2 U17080 ( .A(n18826), .B(n19246), .Y(n18903) );
  sky130_fd_sc_hd__nor2_2 U17081 ( .A(n18810), .B(n18811), .Y(n18872) );
  sky130_fd_sc_hd__xnor2_1 U17084 ( .A(n18490), .B(n11516), .Y(n18545) );
  sky130_fd_sc_hd__xnor2_1 U17085 ( .A(n18491), .B(n18492), .Y(n11516) );
  sky130_fd_sc_hd__xnor3_1 U17086 ( .A(n12776), .B(n18482), .C(n18483), .X(
        n18490) );
  sky130_fd_sc_hd__nand2_1 U17087 ( .A(n11519), .B(n29513), .Y(n23002) );
  sky130_fd_sc_hd__nand2_1 U17088 ( .A(n11519), .B(n12024), .Y(n12940) );
  sky130_fd_sc_hd__nand2_1 U17089 ( .A(n11519), .B(n12689), .Y(n26970) );
  sky130_fd_sc_hd__inv_1 U17090 ( .A(n25191), .Y(n25140) );
  sky130_fd_sc_hd__nand3_1 U17091 ( .A(n11769), .B(n24781), .C(n26691), .Y(
        n24782) );
  sky130_fd_sc_hd__nand2_1 U17092 ( .A(n11521), .B(n26535), .Y(n23797) );
  sky130_fd_sc_hd__nand4_1 U17095 ( .A(n11526), .B(n11525), .C(n11524), .D(
        n11523), .Y(n11522) );
  sky130_fd_sc_hd__nand2_1 U17096 ( .A(j202_soc_core_memory0_ram_dout0[113]), 
        .B(n21591), .Y(n11523) );
  sky130_fd_sc_hd__nand2_1 U17097 ( .A(j202_soc_core_memory0_ram_dout0[209]), 
        .B(n21732), .Y(n11524) );
  sky130_fd_sc_hd__nand2_1 U17098 ( .A(j202_soc_core_memory0_ram_dout0[433]), 
        .B(n21598), .Y(n11525) );
  sky130_fd_sc_hd__nand2_1 U17099 ( .A(j202_soc_core_memory0_ram_dout0[465]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11526) );
  sky130_fd_sc_hd__nand4_1 U17100 ( .A(n11531), .B(n11530), .C(n11529), .D(
        n11528), .Y(n11527) );
  sky130_fd_sc_hd__nand2_1 U17101 ( .A(j202_soc_core_memory0_ram_dout0[369]), 
        .B(n21596), .Y(n11528) );
  sky130_fd_sc_hd__nand2_1 U17102 ( .A(j202_soc_core_memory0_ram_dout0[241]), 
        .B(n21735), .Y(n11529) );
  sky130_fd_sc_hd__nand2_1 U17103 ( .A(j202_soc_core_memory0_ram_dout0[145]), 
        .B(n21592), .Y(n11530) );
  sky130_fd_sc_hd__nand2_1 U17104 ( .A(j202_soc_core_memory0_ram_dout0[17]), 
        .B(n21733), .Y(n11531) );
  sky130_fd_sc_hd__nor2_1 U17105 ( .A(n12153), .B(n11532), .Y(n12488) );
  sky130_fd_sc_hd__nand2_1 U17106 ( .A(n24263), .B(n11071), .Y(n24269) );
  sky130_fd_sc_hd__nand2_1 U17107 ( .A(n23164), .B(n23586), .Y(n11533) );
  sky130_fd_sc_hd__nand2_1 U17108 ( .A(n23079), .B(n11534), .Y(n29317) );
  sky130_fd_sc_hd__nand2b_1 U17109 ( .A_N(n23537), .B(n23536), .Y(n11534) );
  sky130_fd_sc_hd__clkinv_1 U17111 ( .A(n13525), .Y(n11537) );
  sky130_fd_sc_hd__nand2_1 U17112 ( .A(n13525), .B(n12200), .Y(n24430) );
  sky130_fd_sc_hd__inv_2 U17113 ( .A(n11540), .Y(n26512) );
  sky130_fd_sc_hd__nand2_1 U17114 ( .A(n11542), .B(n26716), .Y(n11541) );
  sky130_fd_sc_hd__nand2_1 U17115 ( .A(n12769), .B(n12768), .Y(n11542) );
  sky130_fd_sc_hd__o21ai_1 U17116 ( .A1(n26716), .A2(n26519), .B1(n24481), .Y(
        n11544) );
  sky130_fd_sc_hd__nand2_2 U17117 ( .A(n11546), .B(n11545), .Y(n26519) );
  sky130_fd_sc_hd__nand2_1 U17118 ( .A(n25119), .B(n25120), .Y(n11547) );
  sky130_fd_sc_hd__and2_0 U17119 ( .A(n25137), .B(n26443), .X(n11548) );
  sky130_fd_sc_hd__nand2_1 U17120 ( .A(n11550), .B(n11549), .Y(
        j202_soc_core_j22_cpu_rf_N323) );
  sky130_fd_sc_hd__and2_0 U17121 ( .A(n23791), .B(n23790), .X(n11549) );
  sky130_fd_sc_hd__nand2_1 U17122 ( .A(n25116), .B(n11157), .Y(n11550) );
  sky130_fd_sc_hd__o22ai_1 U17123 ( .A1(n25189), .A2(n26070), .B1(n25714), 
        .B2(n11551), .Y(n25190) );
  sky130_fd_sc_hd__o22ai_1 U17124 ( .A1(n27575), .A2(n11551), .B1(n27574), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N3113) );
  sky130_fd_sc_hd__o22ai_1 U17125 ( .A1(n26899), .A2(n11551), .B1(n26898), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N3337) );
  sky130_fd_sc_hd__o22ai_1 U17126 ( .A1(n27225), .A2(n11551), .B1(n27224), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N2965) );
  sky130_fd_sc_hd__o22ai_1 U17127 ( .A1(n27223), .A2(n11551), .B1(n27222), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N3039) );
  sky130_fd_sc_hd__o22ai_1 U17128 ( .A1(n27211), .A2(n11551), .B1(n27210), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N3224) );
  sky130_fd_sc_hd__o22ai_1 U17129 ( .A1(n27228), .A2(n11551), .B1(n27227), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N3187) );
  sky130_fd_sc_hd__o22ai_1 U17130 ( .A1(n27215), .A2(n11551), .B1(n27214), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N2928) );
  sky130_fd_sc_hd__o22ai_1 U17131 ( .A1(n26378), .A2(n11551), .B1(n26449), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N3261) );
  sky130_fd_sc_hd__o22ai_1 U17132 ( .A1(n11141), .A2(n11551), .B1(n27124), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N2706) );
  sky130_fd_sc_hd__o22ai_1 U17133 ( .A1(n27466), .A2(n11551), .B1(n27465), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N2780) );
  sky130_fd_sc_hd__o22ai_1 U17134 ( .A1(n27226), .A2(n11551), .B1(n23079), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N3150) );
  sky130_fd_sc_hd__o22ai_1 U17135 ( .A1(n27217), .A2(n11551), .B1(n27216), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N2854) );
  sky130_fd_sc_hd__o22ai_1 U17136 ( .A1(n27221), .A2(n11551), .B1(n27220), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N2891) );
  sky130_fd_sc_hd__o22ai_1 U17137 ( .A1(n27219), .A2(n11551), .B1(n27218), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N3002) );
  sky130_fd_sc_hd__o22ai_1 U17138 ( .A1(n27209), .A2(n11551), .B1(n23039), 
        .B2(n25222), .Y(j202_soc_core_j22_cpu_rf_N2743) );
  sky130_fd_sc_hd__o21a_1 U17139 ( .A1(n11153), .A2(n23847), .B1(n11552), .X(
        n12477) );
  sky130_fd_sc_hd__a21oi_1 U17140 ( .A1(n26550), .A2(n26406), .B1(n11624), .Y(
        n11552) );
  sky130_fd_sc_hd__nand2_1 U17141 ( .A(n26550), .B(n25871), .Y(n23847) );
  sky130_fd_sc_hd__nand2_1 U17142 ( .A(n11556), .B(n11553), .Y(n25073) );
  sky130_fd_sc_hd__and2_0 U17143 ( .A(n25069), .B(n26351), .X(n11555) );
  sky130_fd_sc_hd__nand2_1 U17144 ( .A(n12740), .B(n11153), .Y(n11558) );
  sky130_fd_sc_hd__o21ai_1 U17145 ( .A1(n25807), .A2(n11561), .B1(n27395), .Y(
        n11560) );
  sky130_fd_sc_hd__and2_1 U17146 ( .A(n26710), .B(n26323), .X(n11561) );
  sky130_fd_sc_hd__nand2b_1 U17147 ( .A_N(n26352), .B(n26710), .Y(n11564) );
  sky130_fd_sc_hd__o21ai_1 U17148 ( .A1(n25809), .A2(n18916), .B1(n25808), .Y(
        n11565) );
  sky130_fd_sc_hd__clkinv_1 U17149 ( .A(n11566), .Y(n25557) );
  sky130_fd_sc_hd__nand2_1 U17151 ( .A(n27388), .B(n24730), .Y(n11567) );
  sky130_fd_sc_hd__nand2_1 U17152 ( .A(n11569), .B(n26721), .Y(n11568) );
  sky130_fd_sc_hd__o21a_1 U17153 ( .A1(n11572), .A2(n24633), .B1(n24631), .X(
        n11571) );
  sky130_fd_sc_hd__and2_0 U17154 ( .A(n24630), .B(n26351), .X(n11572) );
  sky130_fd_sc_hd__xnor2_1 U17155 ( .A(n25128), .B(n24633), .Y(n11573) );
  sky130_fd_sc_hd__nand2_1 U17157 ( .A(n26315), .B(n12078), .Y(n27360) );
  sky130_fd_sc_hd__nand2_1 U17158 ( .A(n12079), .B(n11153), .Y(n11575) );
  sky130_fd_sc_hd__nand3_1 U17159 ( .A(n26315), .B(n12078), .C(n26352), .Y(
        n11576) );
  sky130_fd_sc_hd__nand2_1 U17160 ( .A(n11578), .B(n11153), .Y(n11577) );
  sky130_fd_sc_hd__nand2_1 U17161 ( .A(n18082), .B(n11579), .Y(n18086) );
  sky130_fd_sc_hd__nand2_1 U17162 ( .A(n11581), .B(n11580), .Y(n11579) );
  sky130_fd_sc_hd__nand2_1 U17163 ( .A(n22901), .B(n26863), .Y(n25217) );
  sky130_fd_sc_hd__inv_2 U17164 ( .A(n23236), .Y(n25218) );
  sky130_fd_sc_hd__buf_6 U17165 ( .A(n23045), .X(n26315) );
  sky130_fd_sc_hd__nand3_2 U17166 ( .A(n23177), .B(n23176), .C(n23175), .Y(
        n23178) );
  sky130_fd_sc_hd__o21a_1 U17167 ( .A1(n24732), .A2(n18916), .B1(n24731), .X(
        n11582) );
  sky130_fd_sc_hd__nand3_2 U17168 ( .A(n11131), .B(n11583), .C(n11590), .Y(
        n11778) );
  sky130_fd_sc_hd__xnor2_1 U17169 ( .A(n18744), .B(n11585), .Y(n12207) );
  sky130_fd_sc_hd__o2bb2ai_1 U17170 ( .B1(n27276), .B2(n27575), .A1_N(n11586), 
        .A2_N(n11109), .Y(j202_soc_core_j22_cpu_rf_N3096) );
  sky130_fd_sc_hd__nand2_1 U17171 ( .A(n11588), .B(n11587), .Y(n25046) );
  sky130_fd_sc_hd__o21a_1 U17172 ( .A1(n18916), .A2(n25045), .B1(n25044), .X(
        n11587) );
  sky130_fd_sc_hd__nand2_1 U17173 ( .A(n27382), .B(n25043), .Y(n11588) );
  sky130_fd_sc_hd__clkbuf_1 U17174 ( .A(n26064), .X(n11589) );
  sky130_fd_sc_hd__a21oi_2 U17175 ( .A1(n26802), .A2(n26068), .B1(n26073), .Y(
        n25186) );
  sky130_fd_sc_hd__xor2_1 U17178 ( .A(n11591), .B(n18387), .X(n18569) );
  sky130_fd_sc_hd__xor2_1 U17179 ( .A(n18389), .B(n18388), .X(n11591) );
  sky130_fd_sc_hd__nand2_1 U17180 ( .A(n11593), .B(n11592), .Y(n18597) );
  sky130_fd_sc_hd__nand2_1 U17181 ( .A(n18582), .B(n11597), .Y(n11592) );
  sky130_fd_sc_hd__nand2_1 U17182 ( .A(n18581), .B(n11594), .Y(n11593) );
  sky130_fd_sc_hd__nand2b_1 U17183 ( .A_N(n18582), .B(n11595), .Y(n11594) );
  sky130_fd_sc_hd__xnor2_1 U17184 ( .A(n18581), .B(n11596), .Y(n18604) );
  sky130_fd_sc_hd__xnor2_1 U17185 ( .A(n11597), .B(n18582), .Y(n11596) );
  sky130_fd_sc_hd__nand2_1 U17186 ( .A(n11599), .B(n11598), .Y(n11597) );
  sky130_fd_sc_hd__nand2_1 U17187 ( .A(n18388), .B(n18389), .Y(n11598) );
  sky130_fd_sc_hd__nand2_4 U17189 ( .A(n11601), .B(n11600), .Y(n27127) );
  sky130_fd_sc_hd__nand2_1 U17190 ( .A(n25326), .B(n25334), .Y(n11601) );
  sky130_fd_sc_hd__nand2_1 U17191 ( .A(n11603), .B(n11602), .Y(n18832) );
  sky130_fd_sc_hd__nand2_1 U17192 ( .A(n11605), .B(n18806), .Y(n11602) );
  sky130_fd_sc_hd__xor2_1 U17194 ( .A(n11605), .B(n11604), .X(n18829) );
  sky130_fd_sc_hd__xor2_1 U17195 ( .A(n18806), .B(n18805), .X(n11604) );
  sky130_fd_sc_hd__nand2_1 U17196 ( .A(n12696), .B(n12695), .Y(n11605) );
  sky130_fd_sc_hd__inv_2 U17197 ( .A(n21510), .Y(n18904) );
  sky130_fd_sc_hd__nand2_1 U17198 ( .A(n11606), .B(n24047), .Y(n11609) );
  sky130_fd_sc_hd__o21ai_1 U17199 ( .A1(n12929), .A2(n24371), .B1(n12240), .Y(
        n11606) );
  sky130_fd_sc_hd__nand2_1 U17200 ( .A(n11607), .B(n12664), .Y(n13328) );
  sky130_fd_sc_hd__nand2_1 U17201 ( .A(n18602), .B(n18339), .Y(n11607) );
  sky130_fd_sc_hd__o21ai_1 U17202 ( .A1(n18577), .A2(n18578), .B1(n18579), .Y(
        n18336) );
  sky130_fd_sc_hd__inv_1 U17203 ( .A(n26804), .Y(n13065) );
  sky130_fd_sc_hd__nand3_2 U17204 ( .A(n21949), .B(n21947), .C(n21948), .Y(
        n26804) );
  sky130_fd_sc_hd__clkbuf_1 U17206 ( .A(n27364), .X(n11611) );
  sky130_fd_sc_hd__clkbuf_1 U17207 ( .A(n26970), .X(n11612) );
  sky130_fd_sc_hd__inv_2 U17208 ( .A(n24186), .Y(n24187) );
  sky130_fd_sc_hd__nor2_1 U17209 ( .A(n17895), .B(n17896), .Y(n17897) );
  sky130_fd_sc_hd__nand2_1 U17210 ( .A(n12318), .B(n12319), .Y(n21431) );
  sky130_fd_sc_hd__clkbuf_1 U17211 ( .A(n23253), .X(n11614) );
  sky130_fd_sc_hd__xnor2_1 U17212 ( .A(n12569), .B(n25830), .Y(n17386) );
  sky130_fd_sc_hd__nand2_1 U17213 ( .A(n11616), .B(n11615), .Y(n17622) );
  sky130_fd_sc_hd__nand2_1 U17214 ( .A(n17620), .B(n11618), .Y(n11615) );
  sky130_fd_sc_hd__o21ai_1 U17215 ( .A1(n11618), .A2(n17620), .B1(n17619), .Y(
        n11616) );
  sky130_fd_sc_hd__xnor2_1 U17216 ( .A(n17619), .B(n11617), .Y(n17913) );
  sky130_fd_sc_hd__xnor2_1 U17217 ( .A(n11618), .B(n17620), .Y(n11617) );
  sky130_fd_sc_hd__xor2_1 U17218 ( .A(n17572), .B(n11619), .X(n11618) );
  sky130_fd_sc_hd__xnor2_1 U17219 ( .A(n12575), .B(n17573), .Y(n11619) );
  sky130_fd_sc_hd__nand2_1 U17220 ( .A(n25833), .B(n11620), .Y(
        j202_soc_core_j22_cpu_rf_N3279) );
  sky130_fd_sc_hd__nand2_1 U17221 ( .A(n27395), .B(n27460), .Y(n11620) );
  sky130_fd_sc_hd__nand2_4 U17222 ( .A(n23045), .B(n23001), .Y(n12353) );
  sky130_fd_sc_hd__nand2_1 U17223 ( .A(n11622), .B(n11621), .Y(n17879) );
  sky130_fd_sc_hd__nand2_1 U17224 ( .A(n17734), .B(n17735), .Y(n11621) );
  sky130_fd_sc_hd__xnor3_1 U17226 ( .A(n11623), .B(n17734), .C(n17733), .X(
        n17872) );
  sky130_fd_sc_hd__inv_2 U17227 ( .A(n18911), .Y(n22837) );
  sky130_fd_sc_hd__nand2b_1 U17228 ( .A_N(n23845), .B(n23846), .Y(n11624) );
  sky130_fd_sc_hd__nand2_1 U17229 ( .A(n22306), .B(n11625), .Y(n22307) );
  sky130_fd_sc_hd__inv_2 U17231 ( .A(n11628), .Y(n13276) );
  sky130_fd_sc_hd__nand2_1 U17232 ( .A(n28977), .B(n11129), .Y(n11628) );
  sky130_fd_sc_hd__xnor2_1 U17234 ( .A(n17551), .B(n11629), .Y(n17576) );
  sky130_fd_sc_hd__xnor2_1 U17235 ( .A(n17549), .B(n17550), .Y(n11629) );
  sky130_fd_sc_hd__nand2_1 U17236 ( .A(n11631), .B(n11630), .Y(n17522) );
  sky130_fd_sc_hd__nand2_1 U17237 ( .A(n17457), .B(n11635), .Y(n11630) );
  sky130_fd_sc_hd__nand2_1 U17238 ( .A(n17456), .B(n11632), .Y(n11631) );
  sky130_fd_sc_hd__nand2b_1 U17239 ( .A_N(n17457), .B(n11633), .Y(n11632) );
  sky130_fd_sc_hd__xnor2_1 U17240 ( .A(n11634), .B(n17456), .Y(n17569) );
  sky130_fd_sc_hd__xnor2_1 U17241 ( .A(n11635), .B(n17457), .Y(n11634) );
  sky130_fd_sc_hd__nand2_1 U17242 ( .A(n11637), .B(n11636), .Y(n11635) );
  sky130_fd_sc_hd__nand2_1 U17243 ( .A(n17551), .B(n17550), .Y(n11636) );
  sky130_fd_sc_hd__inv_2 U17245 ( .A(n23603), .Y(n23144) );
  sky130_fd_sc_hd__inv_1 U17246 ( .A(n17925), .Y(n12319) );
  sky130_fd_sc_hd__nand4_1 U17247 ( .A(n13095), .B(n13094), .C(n13096), .D(
        n11638), .Y(n13093) );
  sky130_fd_sc_hd__nand2_1 U17248 ( .A(j202_soc_core_memory0_ram_dout0[404]), 
        .B(n21597), .Y(n11638) );
  sky130_fd_sc_hd__inv_2 U17249 ( .A(n13011), .Y(n13272) );
  sky130_fd_sc_hd__nor2b_1 U17250 ( .B_N(n11138), .A(n11847), .Y(n24409) );
  sky130_fd_sc_hd__inv_1 U17251 ( .A(n11805), .Y(n12875) );
  sky130_fd_sc_hd__nor2_2 U17252 ( .A(n13377), .B(n13496), .Y(n21735) );
  sky130_fd_sc_hd__nand4_1 U17255 ( .A(n12818), .B(n12816), .C(n12817), .D(
        n12815), .Y(n12814) );
  sky130_fd_sc_hd__nand3b_1 U17257 ( .A_N(n23821), .B(n24456), .C(n12744), .Y(
        n11810) );
  sky130_fd_sc_hd__nand4_1 U17258 ( .A(n11639), .B(n12715), .C(n24458), .D(
        n13046), .Y(n13045) );
  sky130_fd_sc_hd__nor2_1 U17259 ( .A(n13048), .B(n13047), .Y(n11639) );
  sky130_fd_sc_hd__nand4_1 U17260 ( .A(n12093), .B(n11640), .C(n27785), .D(
        n11074), .Y(n27795) );
  sky130_fd_sc_hd__nand2_1 U17261 ( .A(n11888), .B(n17138), .Y(n17149) );
  sky130_fd_sc_hd__clkbuf_1 U17264 ( .A(n27964), .X(n11642) );
  sky130_fd_sc_hd__nand2_1 U17267 ( .A(n11698), .B(n24310), .Y(n13054) );
  sky130_fd_sc_hd__nand4_1 U17268 ( .A(n12971), .B(n11724), .C(n16832), .D(
        n11645), .Y(n12970) );
  sky130_fd_sc_hd__nand2_1 U17269 ( .A(j202_soc_core_memory0_ram_dout0[93]), 
        .B(n21734), .Y(n11645) );
  sky130_fd_sc_hd__clkbuf_1 U17270 ( .A(n28972), .X(n11646) );
  sky130_fd_sc_hd__nand2_2 U17271 ( .A(n12486), .B(n11996), .Y(n27566) );
  sky130_fd_sc_hd__nor2_2 U17272 ( .A(n23148), .B(n12501), .Y(n12486) );
  sky130_fd_sc_hd__nand4_1 U17273 ( .A(n16631), .B(n16630), .C(n20968), .D(
        n16633), .Y(n13245) );
  sky130_fd_sc_hd__nand2_1 U17274 ( .A(j202_soc_core_memory0_ram_dout0[220]), 
        .B(n21732), .Y(n16630) );
  sky130_fd_sc_hd__nand2_1 U17275 ( .A(n24559), .B(n11647), .Y(
        j202_soc_core_j22_cpu_rf_N2692) );
  sky130_fd_sc_hd__nand3_2 U17276 ( .A(n12489), .B(n12460), .C(n20975), .Y(
        n22019) );
  sky130_fd_sc_hd__inv_1 U17277 ( .A(n11648), .Y(n13087) );
  sky130_fd_sc_hd__nand4_1 U17278 ( .A(n13088), .B(n13089), .C(n13090), .D(
        n13091), .Y(n11648) );
  sky130_fd_sc_hd__nand4_1 U17279 ( .A(n19253), .B(n19252), .C(n11649), .D(
        n19306), .Y(n12958) );
  sky130_fd_sc_hd__nand2_1 U17280 ( .A(j202_soc_core_memory0_ram_dout0[236]), 
        .B(n21735), .Y(n11649) );
  sky130_fd_sc_hd__nand3_2 U17281 ( .A(n23951), .B(n12501), .C(n10974), .Y(
        n11842) );
  sky130_fd_sc_hd__inv_2 U17282 ( .A(n11650), .Y(n23951) );
  sky130_fd_sc_hd__o21a_1 U17285 ( .A1(n11651), .A2(n27795), .B1(n12129), .X(
        n10573) );
  sky130_fd_sc_hd__nand4_1 U17286 ( .A(n12327), .B(n27939), .C(n27794), .D(
        n27793), .Y(n11651) );
  sky130_fd_sc_hd__nand4_1 U17287 ( .A(n12962), .B(n12961), .C(n12963), .D(
        n11652), .Y(n12960) );
  sky130_fd_sc_hd__nand2_1 U17288 ( .A(j202_soc_core_memory0_ram_dout0[381]), 
        .B(n21596), .Y(n11652) );
  sky130_fd_sc_hd__nand2_1 U17289 ( .A(n12355), .B(n27215), .Y(n24555) );
  sky130_fd_sc_hd__inv_2 U17290 ( .A(n23585), .Y(n23160) );
  sky130_fd_sc_hd__o31a_1 U17291 ( .A1(n13259), .A2(n21778), .A3(n12503), .B1(
        n13261), .X(n20835) );
  sky130_fd_sc_hd__nand2_1 U17292 ( .A(n12884), .B(n29534), .Y(n12614) );
  sky130_fd_sc_hd__nor2_1 U17293 ( .A(n23211), .B(n23157), .Y(n11698) );
  sky130_fd_sc_hd__o22a_1 U17294 ( .A1(n26312), .A2(n12359), .B1(n26314), .B2(
        n23694), .X(n26551) );
  sky130_fd_sc_hd__nand2_1 U17295 ( .A(n12111), .B(n26443), .Y(n11653) );
  sky130_fd_sc_hd__nor2_1 U17296 ( .A(n11654), .B(n11999), .Y(n11998) );
  sky130_fd_sc_hd__nand4_1 U17297 ( .A(n21148), .B(n21144), .C(n21143), .D(
        n21036), .Y(n11654) );
  sky130_fd_sc_hd__nand2_1 U17305 ( .A(j202_soc_core_memory0_ram_dout0[92]), 
        .B(n21734), .Y(n16631) );
  sky130_fd_sc_hd__nand2_1 U17306 ( .A(n11657), .B(n27980), .Y(n27903) );
  sky130_fd_sc_hd__nand2_1 U17307 ( .A(n12393), .B(n11658), .Y(n11657) );
  sky130_fd_sc_hd__nand2_1 U17308 ( .A(n11105), .B(n11659), .Y(n11658) );
  sky130_fd_sc_hd__nand2_1 U17309 ( .A(n11660), .B(n29077), .Y(n27782) );
  sky130_fd_sc_hd__inv_1 U17310 ( .A(n27878), .Y(n11660) );
  sky130_fd_sc_hd__nand3_2 U17311 ( .A(n12261), .B(n12477), .C(n23855), .Y(
        n25878) );
  sky130_fd_sc_hd__nand3b_1 U17312 ( .A_N(n27566), .B(n12482), .C(n13269), .Y(
        n23146) );
  sky130_fd_sc_hd__nand3_2 U17313 ( .A(n22935), .B(n22916), .C(n22917), .Y(
        n28994) );
  sky130_fd_sc_hd__nand2_1 U17315 ( .A(n22718), .B(n26603), .Y(n11662) );
  sky130_fd_sc_hd__nor2_1 U17316 ( .A(n11663), .B(n13031), .Y(n12657) );
  sky130_fd_sc_hd__nand4_1 U17317 ( .A(n13034), .B(n13038), .C(n13033), .D(
        n13223), .Y(n11663) );
  sky130_fd_sc_hd__o21ai_1 U17319 ( .A1(n18127), .A2(n18128), .B1(n18126), .Y(
        n18130) );
  sky130_fd_sc_hd__nand2_1 U17320 ( .A(n11666), .B(n11665), .Y(n18040) );
  sky130_fd_sc_hd__nand2_1 U17321 ( .A(n18003), .B(n11668), .Y(n11665) );
  sky130_fd_sc_hd__o21ai_1 U17322 ( .A1(n11668), .A2(n18003), .B1(n18002), .Y(
        n11666) );
  sky130_fd_sc_hd__xnor2_1 U17323 ( .A(n18003), .B(n11667), .Y(n17999) );
  sky130_fd_sc_hd__xnor2_1 U17324 ( .A(n11668), .B(n18002), .Y(n11667) );
  sky130_fd_sc_hd__nand2b_4 U17325 ( .A_N(n23167), .B(n29595), .Y(
        j202_soc_core_ahb2apb_01_N22) );
  sky130_fd_sc_hd__nor2_1 U17326 ( .A(n22675), .B(n12085), .Y(n23167) );
  sky130_fd_sc_hd__nor2_2 U17327 ( .A(n13489), .B(n13499), .Y(n21603) );
  sky130_fd_sc_hd__nor2b_1 U17328 ( .B_N(n17101), .A(n11678), .Y(n13126) );
  sky130_fd_sc_hd__nor2_4 U17330 ( .A(n11900), .B(n12346), .Y(n13236) );
  sky130_fd_sc_hd__nand3_2 U17331 ( .A(n13191), .B(n13192), .C(n13190), .Y(
        n13189) );
  sky130_fd_sc_hd__inv_2 U17332 ( .A(n11682), .Y(n26529) );
  sky130_fd_sc_hd__inv_2 U17336 ( .A(n24659), .Y(n23803) );
  sky130_fd_sc_hd__nand3_2 U17337 ( .A(n13162), .B(n24452), .C(n23802), .Y(
        n24659) );
  sky130_fd_sc_hd__nand2_1 U17339 ( .A(n17054), .B(n11671), .Y(n11670) );
  sky130_fd_sc_hd__nor2b_1 U17340 ( .B_N(n17302), .A(n17056), .Y(n11672) );
  sky130_fd_sc_hd__nand2_1 U17341 ( .A(n17053), .B(n20787), .Y(n11674) );
  sky130_fd_sc_hd__clkbuf_1 U17342 ( .A(n12656), .X(n11675) );
  sky130_fd_sc_hd__nand2_1 U17343 ( .A(n11677), .B(n11676), .Y(n17099) );
  sky130_fd_sc_hd__nand2_1 U17344 ( .A(n17062), .B(n17061), .Y(n11677) );
  sky130_fd_sc_hd__nand2_1 U17345 ( .A(n13128), .B(n13127), .Y(n11678) );
  sky130_fd_sc_hd__nand2_1 U17346 ( .A(n11680), .B(n27980), .Y(n27573) );
  sky130_fd_sc_hd__nand4_1 U17347 ( .A(n27569), .B(n27597), .C(n27570), .D(
        n11681), .Y(n11680) );
  sky130_fd_sc_hd__nand2_1 U17348 ( .A(n13084), .B(n13517), .Y(n11682) );
  sky130_fd_sc_hd__nand2_1 U17349 ( .A(n13140), .B(n29077), .Y(n27258) );
  sky130_fd_sc_hd__nand3_1 U17351 ( .A(n11812), .B(n11813), .C(n27776), .Y(
        n11869) );
  sky130_fd_sc_hd__inv_1 U17352 ( .A(n11691), .Y(n12988) );
  sky130_fd_sc_hd__nand3_1 U17353 ( .A(n13230), .B(n13231), .C(n20834), .Y(
        n29053) );
  sky130_fd_sc_hd__nand2_1 U17354 ( .A(n21519), .B(n12235), .Y(n13230) );
  sky130_fd_sc_hd__inv_2 U17355 ( .A(n11683), .Y(n24203) );
  sky130_fd_sc_hd__nand2_1 U17356 ( .A(n28994), .B(n27824), .Y(n11683) );
  sky130_fd_sc_hd__nor2_1 U17357 ( .A(n29009), .B(n29014), .Y(n13116) );
  sky130_fd_sc_hd__nand3_2 U17358 ( .A(n18880), .B(n11614), .C(n18870), .Y(
        n22936) );
  sky130_fd_sc_hd__nand2_1 U17359 ( .A(n24112), .B(n11684), .Y(n18880) );
  sky130_fd_sc_hd__inv_2 U17360 ( .A(n22028), .Y(n26872) );
  sky130_fd_sc_hd__nand3_1 U17361 ( .A(n11685), .B(n25045), .C(n25030), .Y(
        n19243) );
  sky130_fd_sc_hd__nand2_1 U17362 ( .A(n12348), .B(n19237), .Y(n11685) );
  sky130_fd_sc_hd__nand4_1 U17363 ( .A(n12857), .B(n12856), .C(n12858), .D(
        n12855), .Y(n12854) );
  sky130_fd_sc_hd__inv_2 U17364 ( .A(n11686), .Y(n22935) );
  sky130_fd_sc_hd__nand3_2 U17366 ( .A(n11690), .B(n22767), .C(n22768), .Y(
        n22827) );
  sky130_fd_sc_hd__nand2_1 U17367 ( .A(n22414), .B(n11060), .Y(n28978) );
  sky130_fd_sc_hd__a211o_1 U17368 ( .A1(n24119), .A2(n25108), .B1(n24118), 
        .C1(n12457), .X(n29114) );
  sky130_fd_sc_hd__xnor2_1 U17369 ( .A(n17628), .B(n11687), .Y(n17679) );
  sky130_fd_sc_hd__xnor2_1 U17370 ( .A(n17627), .B(n17629), .Y(n11687) );
  sky130_fd_sc_hd__xnor2_1 U17371 ( .A(n17676), .B(n17677), .Y(n12316) );
  sky130_fd_sc_hd__nand2_1 U17372 ( .A(n11689), .B(n11688), .Y(n17676) );
  sky130_fd_sc_hd__nand2_1 U17373 ( .A(n17628), .B(n17629), .Y(n11688) );
  sky130_fd_sc_hd__o21ai_1 U17374 ( .A1(n17629), .A2(n17628), .B1(n17627), .Y(
        n11689) );
  sky130_fd_sc_hd__nand3_2 U17375 ( .A(n22766), .B(n13318), .C(n24700), .Y(
        n11690) );
  sky130_fd_sc_hd__a22oi_2 U17376 ( .A1(j202_soc_core_memory0_ram_dout0[353]), 
        .A2(n21596), .B1(n21597), .B2(j202_soc_core_memory0_ram_dout0[385]), 
        .Y(n19930) );
  sky130_fd_sc_hd__nand2_1 U17377 ( .A(n12013), .B(n22716), .Y(n11691) );
  sky130_fd_sc_hd__nand2_1 U17378 ( .A(n11718), .B(n16144), .Y(n11692) );
  sky130_fd_sc_hd__o22ai_1 U17379 ( .A1(n18224), .A2(n17586), .B1(n17585), 
        .B2(n18225), .Y(n17633) );
  sky130_fd_sc_hd__xor2_1 U17380 ( .A(n17521), .B(n11693), .X(n17568) );
  sky130_fd_sc_hd__xnor2_1 U17381 ( .A(n12572), .B(n17522), .Y(n11693) );
  sky130_fd_sc_hd__nor2_2 U17382 ( .A(n17926), .B(n17927), .Y(n21805) );
  sky130_fd_sc_hd__inv_2 U17383 ( .A(n25046), .Y(n11694) );
  sky130_fd_sc_hd__inv_2 U17384 ( .A(n11695), .Y(n13192) );
  sky130_fd_sc_hd__nand2_1 U17385 ( .A(n13080), .B(n13187), .Y(n11695) );
  sky130_fd_sc_hd__nand3_2 U17386 ( .A(n12587), .B(n20835), .C(n12347), .Y(
        n12346) );
  sky130_fd_sc_hd__inv_2 U17387 ( .A(n11696), .Y(n12587) );
  sky130_fd_sc_hd__nand2_1 U17388 ( .A(n20957), .B(n20959), .Y(n11696) );
  sky130_fd_sc_hd__inv_2 U17389 ( .A(j202_soc_core_intc_core_00_rg_ipr[5]), 
        .Y(n24056) );
  sky130_fd_sc_hd__mux2i_1 U17390 ( .A0(n11699), .A1(n19648), .S(n26840), .Y(
        n19775) );
  sky130_fd_sc_hd__clkbuf_1 U17391 ( .A(n27202), .X(n11700) );
  sky130_fd_sc_hd__nand3_1 U17392 ( .A(n22285), .B(n12515), .C(n22284), .Y(
        n13228) );
  sky130_fd_sc_hd__nand4_1 U17393 ( .A(n11852), .B(n11851), .C(n11853), .D(
        n11701), .Y(n11850) );
  sky130_fd_sc_hd__nand2_1 U17394 ( .A(j202_soc_core_memory0_ram_dout0[282]), 
        .B(n21605), .Y(n11701) );
  sky130_fd_sc_hd__nand2_1 U17395 ( .A(j202_soc_core_memory0_ram_dout0[240]), 
        .B(n21735), .Y(n11702) );
  sky130_fd_sc_hd__inv_1 U17396 ( .A(n11703), .Y(n19448) );
  sky130_fd_sc_hd__clkbuf_1 U17397 ( .A(n27421), .X(n11704) );
  sky130_fd_sc_hd__clkbuf_1 U17398 ( .A(n12840), .X(n11705) );
  sky130_fd_sc_hd__inv_1 U17399 ( .A(n11707), .Y(n22667) );
  sky130_fd_sc_hd__nand2_1 U17400 ( .A(n22270), .B(n12296), .Y(n11707) );
  sky130_fd_sc_hd__nand3_2 U17401 ( .A(n24591), .B(n24590), .C(n22768), .Y(
        n22270) );
  sky130_fd_sc_hd__inv_2 U17402 ( .A(n24189), .Y(n24190) );
  sky130_fd_sc_hd__nor2_2 U17403 ( .A(n13491), .B(n13496), .Y(n21590) );
  sky130_fd_sc_hd__nand4_1 U17404 ( .A(n12623), .B(n12801), .C(n12800), .D(
        n12589), .Y(n12799) );
  sky130_fd_sc_hd__a21oi_2 U17405 ( .A1(n12510), .A2(n17004), .B1(n17003), .Y(
        n12400) );
  sky130_fd_sc_hd__nand2_1 U17406 ( .A(n11708), .B(n27980), .Y(n24302) );
  sky130_fd_sc_hd__nand3_1 U17407 ( .A(n11826), .B(n11825), .C(n12764), .Y(
        n11708) );
  sky130_fd_sc_hd__nand4_2 U17408 ( .A(n11898), .B(n17126), .C(n17130), .D(
        n11897), .Y(n27823) );
  sky130_fd_sc_hd__nand3_1 U17409 ( .A(n27300), .B(n13303), .C(n11709), .Y(
        n10579) );
  sky130_fd_sc_hd__o21ai_1 U17410 ( .A1(n24107), .A2(n12361), .B1(n27980), .Y(
        n11709) );
  sky130_fd_sc_hd__inv_2 U17411 ( .A(n27686), .Y(n27687) );
  sky130_fd_sc_hd__nand2_1 U17412 ( .A(n11906), .B(n11710), .Y(n18982) );
  sky130_fd_sc_hd__nand2_1 U17413 ( .A(n22236), .B(n11712), .Y(n11711) );
  sky130_fd_sc_hd__nand2b_1 U17414 ( .A_N(n22237), .B(n11713), .Y(n11712) );
  sky130_fd_sc_hd__nand2_1 U17415 ( .A(n29005), .B(n27824), .Y(n24221) );
  sky130_fd_sc_hd__nor2b_1 U17416 ( .B_N(n11158), .A(n22352), .Y(n11715) );
  sky130_fd_sc_hd__o21ai_2 U17417 ( .A1(n21385), .A2(n21388), .B1(n21386), .Y(
        n19423) );
  sky130_fd_sc_hd__clkbuf_1 U17418 ( .A(j202_soc_core_j22_cpu_ml_bufa[2]), .X(
        n11716) );
  sky130_fd_sc_hd__inv_2 U17421 ( .A(n12714), .Y(n12641) );
  sky130_fd_sc_hd__nor2_1 U17423 ( .A(n27791), .B(n23967), .Y(n23964) );
  sky130_fd_sc_hd__nand4_1 U17424 ( .A(n12859), .B(n12869), .C(n12853), .D(
        n12863), .Y(n11718) );
  sky130_fd_sc_hd__inv_2 U17426 ( .A(n13236), .Y(n23953) );
  sky130_fd_sc_hd__nand2_1 U17427 ( .A(n11719), .B(n11965), .Y(n27792) );
  sky130_fd_sc_hd__nand2_1 U17428 ( .A(n11721), .B(n11720), .Y(n11719) );
  sky130_fd_sc_hd__nand2_1 U17429 ( .A(n27789), .B(n29548), .Y(n11720) );
  sky130_fd_sc_hd__inv_2 U17430 ( .A(n12467), .Y(n11721) );
  sky130_fd_sc_hd__nand3_1 U17431 ( .A(n24589), .B(n24587), .C(n24588), .Y(
        j202_soc_core_j22_cpu_ml_maclj[4]) );
  sky130_fd_sc_hd__nand3_1 U17432 ( .A(n25052), .B(n25050), .C(n25051), .Y(
        j202_soc_core_j22_cpu_ml_maclj[10]) );
  sky130_fd_sc_hd__nand3_1 U17433 ( .A(n24059), .B(n24058), .C(n24057), .Y(
        j202_soc_core_j22_cpu_ml_maclj[1]) );
  sky130_fd_sc_hd__nand3_1 U17434 ( .A(n24065), .B(n24063), .C(n24064), .Y(
        j202_soc_core_j22_cpu_ml_maclj[5]) );
  sky130_fd_sc_hd__nand3_1 U17435 ( .A(n24605), .B(n24604), .C(n24603), .Y(
        j202_soc_core_j22_cpu_ml_maclj[0]) );
  sky130_fd_sc_hd__a2bb2oi_2 U17436 ( .B1(n23777), .B2(n12727), .A1_N(n26312), 
        .A2_N(n23753), .Y(n26552) );
  sky130_fd_sc_hd__nand2_1 U17437 ( .A(n28921), .B(n22712), .Y(n21378) );
  sky130_fd_sc_hd__o21a_1 U17438 ( .A1(n20719), .A2(n20718), .B1(n20717), .X(
        n28921) );
  sky130_fd_sc_hd__nand4_1 U17440 ( .A(n12860), .B(n12862), .C(n12861), .D(
        n11722), .Y(n11757) );
  sky130_fd_sc_hd__nand2_1 U17441 ( .A(j202_soc_core_memory0_ram_dout0[25]), 
        .B(n21733), .Y(n11722) );
  sky130_fd_sc_hd__nand2_1 U17444 ( .A(j202_soc_core_memory0_ram_dout0[349]), 
        .B(n21593), .Y(n11724) );
  sky130_fd_sc_hd__nand2_1 U17446 ( .A(n11906), .B(n11726), .Y(n11944) );
  sky130_fd_sc_hd__nand2_1 U17449 ( .A(n11728), .B(n11727), .Y(n26799) );
  sky130_fd_sc_hd__nand2_1 U17450 ( .A(n11729), .B(n26775), .Y(n11728) );
  sky130_fd_sc_hd__nor2_2 U17452 ( .A(n23211), .B(n12467), .Y(n12511) );
  sky130_fd_sc_hd__nand3_1 U17454 ( .A(n13186), .B(n13321), .C(n25816), .Y(
        n13007) );
  sky130_fd_sc_hd__nand2_1 U17455 ( .A(n20972), .B(n12229), .Y(n12489) );
  sky130_fd_sc_hd__nand3_1 U17456 ( .A(n20966), .B(n13243), .C(n13246), .Y(
        n20972) );
  sky130_fd_sc_hd__nand2_1 U17457 ( .A(n11730), .B(n12955), .Y(n20974) );
  sky130_fd_sc_hd__nor2_1 U17458 ( .A(n12814), .B(n12809), .Y(n11730) );
  sky130_fd_sc_hd__nand2_1 U17460 ( .A(n24557), .B(n11732), .Y(
        j202_soc_core_j22_cpu_rf_N2951) );
  sky130_fd_sc_hd__nand2_1 U17461 ( .A(n11611), .B(n27224), .Y(n11732) );
  sky130_fd_sc_hd__nand2_1 U17462 ( .A(n24556), .B(n11733), .Y(
        j202_soc_core_j22_cpu_rf_N3025) );
  sky130_fd_sc_hd__nand2_1 U17463 ( .A(n11611), .B(n27222), .Y(n11733) );
  sky130_fd_sc_hd__nand2_1 U17464 ( .A(n24099), .B(n11735), .Y(n11734) );
  sky130_fd_sc_hd__or3_1 U17465 ( .A(n24100), .B(n24254), .C(n27980), .X(
        n11735) );
  sky130_fd_sc_hd__nand2_1 U17469 ( .A(n11739), .B(n11738), .Y(n10496) );
  sky130_fd_sc_hd__nand2_1 U17470 ( .A(n24111), .B(n11138), .Y(n11738) );
  sky130_fd_sc_hd__nand2_1 U17471 ( .A(n13239), .B(n13237), .Y(n11739) );
  sky130_fd_sc_hd__inv_1 U17473 ( .A(n23223), .Y(n23240) );
  sky130_fd_sc_hd__nand2_1 U17474 ( .A(n11741), .B(n11740), .Y(n18419) );
  sky130_fd_sc_hd__nand2_1 U17475 ( .A(n18395), .B(n18394), .Y(n11740) );
  sky130_fd_sc_hd__nand2_1 U17479 ( .A(n11745), .B(n11744), .Y(n18439) );
  sky130_fd_sc_hd__nand2_1 U17480 ( .A(n18400), .B(n18401), .Y(n11744) );
  sky130_fd_sc_hd__nand2_4 U17482 ( .A(n12134), .B(n23253), .Y(n18183) );
  sky130_fd_sc_hd__clkbuf_1 U17484 ( .A(n21791), .X(n11747) );
  sky130_fd_sc_hd__inv_2 U17485 ( .A(n18434), .Y(n12701) );
  sky130_fd_sc_hd__nand2_1 U17486 ( .A(n26375), .B(n11748), .Y(
        j202_soc_core_j22_cpu_rf_N2876) );
  sky130_fd_sc_hd__nand2_1 U17487 ( .A(n27371), .B(n11136), .Y(n11748) );
  sky130_fd_sc_hd__clkbuf_1 U17488 ( .A(j202_soc_core_j22_cpu_ml_bufa[1]), .X(
        n11749) );
  sky130_fd_sc_hd__nand2_1 U17489 ( .A(n26372), .B(n11750), .Y(
        j202_soc_core_j22_cpu_rf_N3061) );
  sky130_fd_sc_hd__nand2_1 U17490 ( .A(n27371), .B(n11137), .Y(n11750) );
  sky130_fd_sc_hd__nand3_4 U17491 ( .A(n11751), .B(n26359), .C(n26357), .Y(
        n26393) );
  sky130_fd_sc_hd__nand2_1 U17492 ( .A(n26358), .B(n26709), .Y(n11751) );
  sky130_fd_sc_hd__o21ai_1 U17493 ( .A1(n26443), .A2(n27371), .B1(n11752), .Y(
        n26324) );
  sky130_fd_sc_hd__nand2_1 U17494 ( .A(n27371), .B(n11153), .Y(n11752) );
  sky130_fd_sc_hd__o21a_1 U17495 ( .A1(n19173), .A2(n17818), .B1(n19176), .X(
        n21388) );
  sky130_fd_sc_hd__nor2_1 U17496 ( .A(n12086), .B(n11753), .Y(n12087) );
  sky130_fd_sc_hd__nand4_1 U17497 ( .A(n16670), .B(n16668), .C(n13059), .D(
        n13063), .Y(n11753) );
  sky130_fd_sc_hd__nand3_2 U17499 ( .A(n27780), .B(n22022), .C(n22023), .Y(
        n12728) );
  sky130_fd_sc_hd__nand2_1 U17500 ( .A(n12642), .B(n23951), .Y(n11874) );
  sky130_fd_sc_hd__nand2_1 U17501 ( .A(n11868), .B(n12476), .Y(n22020) );
  sky130_fd_sc_hd__nor2_1 U17502 ( .A(n12728), .B(n24451), .Y(n24461) );
  sky130_fd_sc_hd__nand2_1 U17504 ( .A(n27978), .B(n27979), .Y(n11755) );
  sky130_fd_sc_hd__nand2_2 U17505 ( .A(n11626), .B(n12004), .Y(n23184) );
  sky130_fd_sc_hd__inv_1 U17506 ( .A(n11757), .Y(n12859) );
  sky130_fd_sc_hd__nand2_1 U17507 ( .A(n19407), .B(n19406), .Y(n11758) );
  sky130_fd_sc_hd__nand2_1 U17508 ( .A(n28980), .B(n27824), .Y(n24178) );
  sky130_fd_sc_hd__nand3_1 U17509 ( .A(n22667), .B(n12671), .C(n19503), .Y(
        n28980) );
  sky130_fd_sc_hd__inv_2 U17512 ( .A(n11760), .Y(n24094) );
  sky130_fd_sc_hd__nand2_1 U17513 ( .A(n11761), .B(n29524), .Y(n11760) );
  sky130_fd_sc_hd__inv_2 U17514 ( .A(n28972), .Y(n11761) );
  sky130_fd_sc_hd__nand4_1 U17516 ( .A(n12332), .B(n12331), .C(n11762), .D(
        n13485), .Y(n13086) );
  sky130_fd_sc_hd__nand2_1 U17517 ( .A(j202_soc_core_memory0_ram_dout0[308]), 
        .B(n21603), .Y(n11762) );
  sky130_fd_sc_hd__nor2_1 U17519 ( .A(n12712), .B(n12008), .Y(n12007) );
  sky130_fd_sc_hd__inv_1 U17522 ( .A(n11763), .Y(n12470) );
  sky130_fd_sc_hd__nor2_4 U17526 ( .A(n23081), .B(n23169), .Y(n27226) );
  sky130_fd_sc_hd__nand2_1 U17527 ( .A(n27382), .B(n26323), .Y(n11765) );
  sky130_fd_sc_hd__nand2_1 U17528 ( .A(n11055), .B(n25230), .Y(n25233) );
  sky130_fd_sc_hd__clkbuf_1 U17529 ( .A(n12374), .X(n11766) );
  sky130_fd_sc_hd__o2bb2ai_1 U17530 ( .B1(n27333), .B2(n25157), .A1_N(n26371), 
        .A2_N(n25158), .Y(j202_soc_core_j22_cpu_rf_N3078) );
  sky130_fd_sc_hd__nand2_4 U17531 ( .A(n11559), .B(n25845), .Y(n25810) );
  sky130_fd_sc_hd__and2_0 U17534 ( .A(n24158), .B(n12592), .X(n11772) );
  sky130_fd_sc_hd__clkbuf_1 U17535 ( .A(n23248), .X(n11774) );
  sky130_fd_sc_hd__xnor2_1 U17536 ( .A(n18524), .B(n18525), .Y(n18507) );
  sky130_fd_sc_hd__nand2_1 U17537 ( .A(n11777), .B(n11775), .Y(
        j202_soc_core_j22_cpu_rf_N3102) );
  sky130_fd_sc_hd__nand2_1 U17538 ( .A(n24163), .B(n11108), .Y(n11775) );
  sky130_fd_sc_hd__nand2_1 U17540 ( .A(n11778), .B(n11109), .Y(n11777) );
  sky130_fd_sc_hd__nand2_1 U17541 ( .A(n11780), .B(n11779), .Y(
        j202_soc_core_j22_cpu_rf_N3115) );
  sky130_fd_sc_hd__nand2_1 U17542 ( .A(n11104), .B(n11108), .Y(n11779) );
  sky130_fd_sc_hd__nand2_1 U17543 ( .A(n12385), .B(n11109), .Y(n11780) );
  sky130_fd_sc_hd__nand2_1 U17544 ( .A(n11782), .B(n11781), .Y(n18787) );
  sky130_fd_sc_hd__nand2_1 U17545 ( .A(n18757), .B(n18758), .Y(n11781) );
  sky130_fd_sc_hd__nand2_1 U17546 ( .A(n18756), .B(n11783), .Y(n11782) );
  sky130_fd_sc_hd__nand2b_1 U17547 ( .A_N(n18757), .B(n11784), .Y(n11783) );
  sky130_fd_sc_hd__xnor2_1 U17548 ( .A(n11785), .B(n18756), .Y(n18784) );
  sky130_fd_sc_hd__xnor2_1 U17549 ( .A(n18758), .B(n18757), .Y(n11785) );
  sky130_fd_sc_hd__nand2_1 U17550 ( .A(n11787), .B(n11786), .Y(n18724) );
  sky130_fd_sc_hd__nand2_1 U17551 ( .A(n18697), .B(n11789), .Y(n11786) );
  sky130_fd_sc_hd__o21ai_1 U17552 ( .A1(n11789), .A2(n18697), .B1(n18696), .Y(
        n11787) );
  sky130_fd_sc_hd__xnor2_1 U17553 ( .A(n18696), .B(n11788), .Y(n18730) );
  sky130_fd_sc_hd__xnor2_1 U17554 ( .A(n11789), .B(n18697), .Y(n11788) );
  sky130_fd_sc_hd__and2_0 U17555 ( .A(n24002), .B(n24003), .X(n11790) );
  sky130_fd_sc_hd__clkbuf_1 U17556 ( .A(n13140), .X(n11792) );
  sky130_fd_sc_hd__inv_2 U17557 ( .A(n29015), .Y(n13140) );
  sky130_fd_sc_hd__nand2_1 U17559 ( .A(n11906), .B(n29586), .Y(n11794) );
  sky130_fd_sc_hd__inv_1 U17564 ( .A(n23165), .Y(n11797) );
  sky130_fd_sc_hd__nand2b_1 U17567 ( .A_N(n24448), .B(n27948), .Y(n13048) );
  sky130_fd_sc_hd__nand2_1 U17568 ( .A(n24264), .B(n11799), .Y(n24448) );
  sky130_fd_sc_hd__nand2_1 U17569 ( .A(n11801), .B(n27683), .Y(n11799) );
  sky130_fd_sc_hd__inv_2 U17570 ( .A(n11800), .Y(n12512) );
  sky130_fd_sc_hd__nor2_1 U17571 ( .A(n12692), .B(n12362), .Y(n11800) );
  sky130_fd_sc_hd__nand3b_4 U17572 ( .A_N(n12362), .B(n11626), .C(n24399), .Y(
        n12665) );
  sky130_fd_sc_hd__nand3_2 U17573 ( .A(n11801), .B(n12461), .C(n24257), .Y(
        n23582) );
  sky130_fd_sc_hd__nand2_1 U17574 ( .A(n13079), .B(n11801), .Y(n13187) );
  sky130_fd_sc_hd__nand3_1 U17575 ( .A(n12286), .B(n23953), .C(n11801), .Y(
        n13270) );
  sky130_fd_sc_hd__nand2_1 U17576 ( .A(n23151), .B(n11801), .Y(n23152) );
  sky130_fd_sc_hd__inv_2 U17577 ( .A(n12362), .Y(n11801) );
  sky130_fd_sc_hd__nand2_1 U17578 ( .A(n23964), .B(n27782), .Y(n11802) );
  sky130_fd_sc_hd__nor2_2 U17580 ( .A(n27687), .B(n11804), .Y(n13043) );
  sky130_fd_sc_hd__inv_1 U17581 ( .A(n24402), .Y(n11804) );
  sky130_fd_sc_hd__inv_1 U17582 ( .A(n12485), .Y(n11806) );
  sky130_fd_sc_hd__inv_1 U17583 ( .A(n11810), .Y(n11807) );
  sky130_fd_sc_hd__nand2_1 U17585 ( .A(n23819), .B(n11867), .Y(n11809) );
  sky130_fd_sc_hd__nand3_2 U17587 ( .A(n12011), .B(n21316), .C(n11811), .Y(
        n28972) );
  sky130_fd_sc_hd__inv_2 U17588 ( .A(n12238), .Y(n11812) );
  sky130_fd_sc_hd__inv_1 U17589 ( .A(n13233), .Y(n11813) );
  sky130_fd_sc_hd__nand2_1 U17590 ( .A(n11132), .B(n11134), .Y(n11814) );
  sky130_fd_sc_hd__inv_2 U17593 ( .A(n27551), .Y(n24353) );
  sky130_fd_sc_hd__nand2_1 U17595 ( .A(n29532), .B(n23158), .Y(n11816) );
  sky130_fd_sc_hd__nand2_1 U17596 ( .A(n27691), .B(n24262), .Y(n24402) );
  sky130_fd_sc_hd__nand2_1 U17598 ( .A(n12665), .B(n24307), .Y(n24308) );
  sky130_fd_sc_hd__nand2_2 U17599 ( .A(n11873), .B(n29522), .Y(n12362) );
  sky130_fd_sc_hd__nor2_1 U17600 ( .A(n11819), .B(n11817), .Y(n23965) );
  sky130_fd_sc_hd__nand2_1 U17603 ( .A(n20976), .B(n12460), .Y(n11821) );
  sky130_fd_sc_hd__nand4_1 U17604 ( .A(n13251), .B(n16629), .C(n11822), .D(
        n13254), .Y(n13249) );
  sky130_fd_sc_hd__nand2_1 U17605 ( .A(j202_soc_core_memory0_ram_dout0[380]), 
        .B(n21596), .Y(n13254) );
  sky130_fd_sc_hd__nand2_1 U17606 ( .A(j202_soc_core_memory0_ram_dout0[476]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11822) );
  sky130_fd_sc_hd__nand2_1 U17607 ( .A(j202_soc_core_memory0_ram_dout0[284]), 
        .B(n21605), .Y(n16629) );
  sky130_fd_sc_hd__nand2_1 U17608 ( .A(j202_soc_core_memory0_ram_dout0[348]), 
        .B(n21593), .Y(n13251) );
  sky130_fd_sc_hd__inv_1 U17609 ( .A(n24298), .Y(n11826) );
  sky130_fd_sc_hd__nand2_1 U17610 ( .A(n29490), .B(n24296), .Y(n24298) );
  sky130_fd_sc_hd__inv_1 U17613 ( .A(n10926), .Y(n11825) );
  sky130_fd_sc_hd__nand2_1 U17614 ( .A(n20146), .B(n12230), .Y(n11827) );
  sky130_fd_sc_hd__nand2_1 U17615 ( .A(n12770), .B(n12657), .Y(n20146) );
  sky130_fd_sc_hd__nand2_1 U17616 ( .A(n12978), .B(n12979), .Y(n11906) );
  sky130_fd_sc_hd__inv_1 U17617 ( .A(n11828), .Y(n11830) );
  sky130_fd_sc_hd__inv_1 U17618 ( .A(n11829), .Y(n11834) );
  sky130_fd_sc_hd__nand4_1 U17619 ( .A(n11831), .B(n24338), .C(n11077), .D(
        n11830), .Y(n11829) );
  sky130_fd_sc_hd__nand2b_1 U17620 ( .A_N(n11832), .B(n27563), .Y(n11828) );
  sky130_fd_sc_hd__inv_2 U17621 ( .A(n24339), .Y(n11831) );
  sky130_fd_sc_hd__nand2_1 U17622 ( .A(n24337), .B(n24456), .Y(n11832) );
  sky130_fd_sc_hd__clkbuf_1 U17623 ( .A(n23582), .X(n11833) );
  sky130_fd_sc_hd__nor2_1 U17624 ( .A(n11838), .B(n11837), .Y(n11836) );
  sky130_fd_sc_hd__nand2_1 U17625 ( .A(n23582), .B(n24334), .Y(n11837) );
  sky130_fd_sc_hd__nand2_1 U17626 ( .A(n24333), .B(n27550), .Y(n11838) );
  sky130_fd_sc_hd__nand2_1 U17627 ( .A(n11840), .B(n12393), .Y(n13232) );
  sky130_fd_sc_hd__nor2_1 U17628 ( .A(n11841), .B(n13189), .Y(n11840) );
  sky130_fd_sc_hd__nand2_1 U17629 ( .A(n27948), .B(n27947), .Y(n11841) );
  sky130_fd_sc_hd__nand2_2 U17631 ( .A(n27790), .B(n11843), .Y(n23154) );
  sky130_fd_sc_hd__inv_2 U17632 ( .A(n24360), .Y(n11843) );
  sky130_fd_sc_hd__nor2_2 U17633 ( .A(n12378), .B(n12879), .Y(n24360) );
  sky130_fd_sc_hd__nand3_1 U17634 ( .A(n12082), .B(n12081), .C(n13198), .Y(
        n12879) );
  sky130_fd_sc_hd__nand3_2 U17635 ( .A(n11844), .B(n27230), .C(n22272), .Y(
        n27790) );
  sky130_fd_sc_hd__inv_2 U17636 ( .A(n13103), .Y(n27230) );
  sky130_fd_sc_hd__nand3_2 U17637 ( .A(n21783), .B(n21782), .C(n12297), .Y(
        n13103) );
  sky130_fd_sc_hd__inv_2 U17638 ( .A(n12378), .Y(n22272) );
  sky130_fd_sc_hd__nand3_2 U17639 ( .A(n13070), .B(n13071), .C(n12293), .Y(
        n12378) );
  sky130_fd_sc_hd__inv_2 U17640 ( .A(n12615), .Y(n11844) );
  sky130_fd_sc_hd__nand2_1 U17641 ( .A(n22273), .B(n29072), .Y(n12615) );
  sky130_fd_sc_hd__inv_2 U17642 ( .A(n11845), .Y(n12436) );
  sky130_fd_sc_hd__nand2_1 U17643 ( .A(n11845), .B(n24094), .Y(n24095) );
  sky130_fd_sc_hd__nor2_2 U17644 ( .A(n12745), .B(n11845), .Y(n12515) );
  sky130_fd_sc_hd__nand2_1 U17646 ( .A(n13270), .B(n11847), .Y(n11846) );
  sky130_fd_sc_hd__nand2_1 U17647 ( .A(n13226), .B(n22282), .Y(n11847) );
  sky130_fd_sc_hd__nor2_1 U17648 ( .A(n11848), .B(n23166), .Y(n12326) );
  sky130_fd_sc_hd__nor2_1 U17649 ( .A(n11848), .B(n27172), .Y(n27173) );
  sky130_fd_sc_hd__nor3_1 U17650 ( .A(n11848), .B(n23166), .C(n23137), .Y(
        n13046) );
  sky130_fd_sc_hd__inv_1 U17652 ( .A(n11849), .Y(n11868) );
  sky130_fd_sc_hd__nor2_1 U17654 ( .A(n11854), .B(n11850), .Y(n11876) );
  sky130_fd_sc_hd__nand2_1 U17655 ( .A(j202_soc_core_memory0_ram_dout0[250]), 
        .B(n21735), .Y(n11851) );
  sky130_fd_sc_hd__nand2_1 U17656 ( .A(j202_soc_core_memory0_ram_dout0[186]), 
        .B(n21590), .Y(n11852) );
  sky130_fd_sc_hd__nand2_1 U17657 ( .A(j202_soc_core_memory0_ram_dout0[58]), 
        .B(n21604), .Y(n11853) );
  sky130_fd_sc_hd__nand4_1 U17658 ( .A(n11858), .B(n11857), .C(n11856), .D(
        n11855), .Y(n11854) );
  sky130_fd_sc_hd__nand2_1 U17659 ( .A(j202_soc_core_memory0_ram_dout0[314]), 
        .B(n21603), .Y(n11855) );
  sky130_fd_sc_hd__nand2_1 U17660 ( .A(j202_soc_core_memory0_ram_dout0[442]), 
        .B(n21598), .Y(n11856) );
  sky130_fd_sc_hd__nand2_1 U17661 ( .A(j202_soc_core_memory0_ram_dout0[410]), 
        .B(n21597), .Y(n11857) );
  sky130_fd_sc_hd__nand2_1 U17662 ( .A(j202_soc_core_memory0_ram_dout0[346]), 
        .B(n21593), .Y(n11858) );
  sky130_fd_sc_hd__nand2_1 U17663 ( .A(n11859), .B(n27980), .Y(n27181) );
  sky130_fd_sc_hd__nand3_1 U17664 ( .A(n11860), .B(n12395), .C(n27169), .Y(
        n11859) );
  sky130_fd_sc_hd__nor2_1 U17665 ( .A(n11862), .B(n11861), .Y(n11860) );
  sky130_fd_sc_hd__nand2_1 U17666 ( .A(n11076), .B(n11130), .Y(n11861) );
  sky130_fd_sc_hd__nand2_1 U17667 ( .A(n27168), .B(n27563), .Y(n11862) );
  sky130_fd_sc_hd__nand2_1 U17670 ( .A(n11866), .B(n23586), .Y(n27259) );
  sky130_fd_sc_hd__nand2_1 U17671 ( .A(n11865), .B(n11864), .Y(n12238) );
  sky130_fd_sc_hd__nand2_1 U17672 ( .A(n13056), .B(n11798), .Y(n11864) );
  sky130_fd_sc_hd__nand3_1 U17673 ( .A(n11866), .B(n11798), .C(n23586), .Y(
        n11865) );
  sky130_fd_sc_hd__inv_1 U17675 ( .A(n11874), .Y(n12598) );
  sky130_fd_sc_hd__nand2_2 U17677 ( .A(n23213), .B(n12376), .Y(n23185) );
  sky130_fd_sc_hd__inv_1 U17678 ( .A(n11871), .Y(n23213) );
  sky130_fd_sc_hd__nand3_1 U17679 ( .A(n23951), .B(n11872), .C(n12501), .Y(
        n11871) );
  sky130_fd_sc_hd__nor2_1 U17680 ( .A(n11107), .B(n29009), .Y(n11872) );
  sky130_fd_sc_hd__nor2_1 U17681 ( .A(n27258), .B(n23185), .Y(n27774) );
  sky130_fd_sc_hd__buf_6 U17682 ( .A(n23951), .X(n11873) );
  sky130_fd_sc_hd__inv_1 U17683 ( .A(n11875), .Y(n12009) );
  sky130_fd_sc_hd__nand2_1 U17686 ( .A(n11877), .B(n11876), .Y(n12911) );
  sky130_fd_sc_hd__nor2_1 U17687 ( .A(n11880), .B(n11878), .Y(n11877) );
  sky130_fd_sc_hd__nand4_1 U17688 ( .A(n15785), .B(n15784), .C(n15781), .D(
        n11879), .Y(n11878) );
  sky130_fd_sc_hd__nand2_1 U17689 ( .A(j202_soc_core_memory0_ram_dout0[474]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11879) );
  sky130_fd_sc_hd__nand4_1 U17690 ( .A(n11896), .B(n15782), .C(n15783), .D(
        n15890), .Y(n11880) );
  sky130_fd_sc_hd__inv_2 U17691 ( .A(n11881), .Y(n24204) );
  sky130_fd_sc_hd__nand2_1 U17692 ( .A(n28995), .B(n24225), .Y(n11881) );
  sky130_fd_sc_hd__nand3_1 U17693 ( .A(n22414), .B(n22413), .C(n22412), .Y(
        n28995) );
  sky130_fd_sc_hd__nand2_1 U17694 ( .A(n12329), .B(n12330), .Y(n22414) );
  sky130_fd_sc_hd__inv_2 U17695 ( .A(n11882), .Y(n23045) );
  sky130_fd_sc_hd__nand4_1 U17696 ( .A(n18985), .B(n18983), .C(n18984), .D(
        n18982), .Y(n11882) );
  sky130_fd_sc_hd__nand2_1 U17697 ( .A(n11884), .B(n11883), .Y(n23173) );
  sky130_fd_sc_hd__nand2_1 U17698 ( .A(n12426), .B(n12427), .Y(n13688) );
  sky130_fd_sc_hd__nand2_1 U17699 ( .A(n12432), .B(n12429), .Y(n13687) );
  sky130_fd_sc_hd__nand3_1 U17700 ( .A(n11963), .B(n26610), .C(n16555), .Y(
        n11959) );
  sky130_fd_sc_hd__nand2_1 U17701 ( .A(n16556), .B(n22513), .Y(n11963) );
  sky130_fd_sc_hd__nand2_1 U17702 ( .A(n14060), .B(n11885), .Y(n14062) );
  sky130_fd_sc_hd__mux2i_1 U17703 ( .A0(n11146), .A1(n11887), .S(n27455), .Y(
        n11885) );
  sky130_fd_sc_hd__nand3_2 U17704 ( .A(n11886), .B(n14057), .C(n14058), .Y(
        n27455) );
  sky130_fd_sc_hd__nand2_1 U17705 ( .A(n21960), .B(n16513), .Y(n11886) );
  sky130_fd_sc_hd__nand2_1 U17706 ( .A(n17149), .B(n12073), .Y(n11899) );
  sky130_fd_sc_hd__nor2_1 U17707 ( .A(n11890), .B(n11889), .Y(n11888) );
  sky130_fd_sc_hd__inv_2 U17711 ( .A(n12464), .Y(n11892) );
  sky130_fd_sc_hd__nand2_1 U17713 ( .A(j202_soc_core_memory0_ram_dout0[378]), 
        .B(n21596), .Y(n11896) );
  sky130_fd_sc_hd__inv_1 U17715 ( .A(n11946), .Y(n11897) );
  sky130_fd_sc_hd__nand3_1 U17716 ( .A(n12911), .B(n15898), .C(n22581), .Y(
        n12628) );
  sky130_fd_sc_hd__nand2_1 U17717 ( .A(n12911), .B(n15898), .Y(n26535) );
  sky130_fd_sc_hd__inv_1 U17718 ( .A(n12346), .Y(n23589) );
  sky130_fd_sc_hd__nand3_2 U17719 ( .A(n12880), .B(n12482), .C(n13236), .Y(
        n27890) );
  sky130_fd_sc_hd__nand3_1 U17721 ( .A(n11873), .B(n27556), .C(n10973), .Y(
        n11901) );
  sky130_fd_sc_hd__inv_2 U17722 ( .A(n11902), .Y(n24091) );
  sky130_fd_sc_hd__nor2_1 U17723 ( .A(n11903), .B(n27566), .Y(n11902) );
  sky130_fd_sc_hd__inv_2 U17724 ( .A(n11904), .Y(n24456) );
  sky130_fd_sc_hd__nor2_1 U17725 ( .A(n11905), .B(n27566), .Y(n11904) );
  sky130_fd_sc_hd__nand2_1 U17726 ( .A(n27260), .B(n11767), .Y(n11905) );
  sky130_fd_sc_hd__nand2_1 U17727 ( .A(n11906), .B(n18981), .Y(n26531) );
  sky130_fd_sc_hd__o22ai_2 U17728 ( .A1(n13602), .A2(n24430), .B1(n11908), 
        .B2(n11907), .Y(n13603) );
  sky130_fd_sc_hd__nand2_1 U17729 ( .A(n11913), .B(n13601), .Y(n11908) );
  sky130_fd_sc_hd__nand2_1 U17730 ( .A(n13603), .B(n11909), .Y(n14847) );
  sky130_fd_sc_hd__inv_2 U17731 ( .A(n11910), .Y(n12158) );
  sky130_fd_sc_hd__nand2_1 U17732 ( .A(n13603), .B(n11911), .Y(n11910) );
  sky130_fd_sc_hd__nand2_1 U17733 ( .A(n13649), .B(n13656), .Y(n11912) );
  sky130_fd_sc_hd__nor2_1 U17734 ( .A(n11914), .B(n12085), .Y(n23288) );
  sky130_fd_sc_hd__nand2_1 U17735 ( .A(n17145), .B(n12416), .Y(n12085) );
  sky130_fd_sc_hd__nand2_1 U17736 ( .A(n24113), .B(n23525), .Y(n11916) );
  sky130_fd_sc_hd__nand2_1 U17737 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[6]), .B(j202_soc_core_bootrom_00_sel_w), .Y(n11917) );
  sky130_fd_sc_hd__nand2_1 U17738 ( .A(n13524), .B(n11919), .Y(n11918) );
  sky130_fd_sc_hd__o21ai_1 U17739 ( .A1(n11910), .A2(n11960), .B1(n11954), .Y(
        n11920) );
  sky130_fd_sc_hd__nand2_1 U17741 ( .A(j202_soc_core_memory0_ram_dout0[159]), 
        .B(n21592), .Y(n11921) );
  sky130_fd_sc_hd__nand2_1 U17742 ( .A(j202_soc_core_memory0_ram_dout0[31]), 
        .B(n21733), .Y(n11922) );
  sky130_fd_sc_hd__nand2_1 U17743 ( .A(j202_soc_core_memory0_ram_dout0[191]), 
        .B(n21590), .Y(n11923) );
  sky130_fd_sc_hd__nand2_1 U17744 ( .A(j202_soc_core_memory0_ram_dout0[287]), 
        .B(n21605), .Y(n11924) );
  sky130_fd_sc_hd__nand4_1 U17745 ( .A(n11927), .B(n11926), .C(n11925), .D(
        n12246), .Y(n11929) );
  sky130_fd_sc_hd__nand2_1 U17746 ( .A(j202_soc_core_memory0_ram_dout0[127]), 
        .B(n21591), .Y(n11925) );
  sky130_fd_sc_hd__nand2_1 U17747 ( .A(j202_soc_core_memory0_ram_dout0[383]), 
        .B(n21596), .Y(n11926) );
  sky130_fd_sc_hd__nand2_1 U17748 ( .A(j202_soc_core_memory0_ram_dout0[63]), 
        .B(n21604), .Y(n11927) );
  sky130_fd_sc_hd__nor2_1 U17749 ( .A(n11929), .B(n11928), .Y(n12979) );
  sky130_fd_sc_hd__nor2_1 U17750 ( .A(n11931), .B(n11930), .Y(n11935) );
  sky130_fd_sc_hd__nand2_1 U17751 ( .A(n17151), .B(n17134), .Y(n11931) );
  sky130_fd_sc_hd__nand4_1 U17752 ( .A(n17151), .B(n17132), .C(n17134), .D(
        n17133), .Y(n17141) );
  sky130_fd_sc_hd__nand3_2 U17753 ( .A(n17131), .B(n11974), .C(n17130), .Y(
        n21022) );
  sky130_fd_sc_hd__nand2_1 U17754 ( .A(n17139), .B(n13292), .Y(n17140) );
  sky130_fd_sc_hd__nand2_2 U17755 ( .A(n11934), .B(n11932), .Y(n11936) );
  sky130_fd_sc_hd__nand2_1 U17756 ( .A(n10934), .B(n11935), .Y(n11934) );
  sky130_fd_sc_hd__inv_1 U17757 ( .A(n11936), .Y(n24188) );
  sky130_fd_sc_hd__inv_1 U17758 ( .A(n11938), .Y(n11937) );
  sky130_fd_sc_hd__nand2_1 U17759 ( .A(n28918), .B(n24123), .Y(n11938) );
  sky130_fd_sc_hd__nand2_2 U17760 ( .A(n11939), .B(n11046), .Y(n28920) );
  sky130_fd_sc_hd__nand2b_1 U17761 ( .A_N(n12913), .B(n11940), .Y(n11939) );
  sky130_fd_sc_hd__nor2_1 U17762 ( .A(n12914), .B(n29521), .Y(n11941) );
  sky130_fd_sc_hd__nand2_1 U17763 ( .A(n26887), .B(n11144), .Y(n11943) );
  sky130_fd_sc_hd__nand2_1 U17769 ( .A(n11049), .B(n12628), .Y(n12073) );
  sky130_fd_sc_hd__nand3_1 U17770 ( .A(n28957), .B(n28960), .C(n28924), .Y(
        n11946) );
  sky130_fd_sc_hd__inv_2 U17771 ( .A(n11947), .Y(n15063) );
  sky130_fd_sc_hd__nor2_1 U17772 ( .A(n13638), .B(n23112), .Y(n11947) );
  sky130_fd_sc_hd__nand2_2 U17773 ( .A(n13751), .B(
        j202_soc_core_j22_cpu_regop_Ra__0_), .Y(n13638) );
  sky130_fd_sc_hd__nand3_1 U17774 ( .A(n13613), .B(n13604), .C(
        j202_soc_core_j22_cpu_regop_Rn__2_), .Y(n23112) );
  sky130_fd_sc_hd__nand2_1 U17775 ( .A(n14381), .B(n14383), .Y(n11949) );
  sky130_fd_sc_hd__xor2_1 U17776 ( .A(n15421), .B(n11950), .X(n26096) );
  sky130_fd_sc_hd__nand2_1 U17777 ( .A(n15416), .B(n11951), .Y(n11950) );
  sky130_fd_sc_hd__nand2_1 U17778 ( .A(n22513), .B(n15417), .Y(n11951) );
  sky130_fd_sc_hd__nand2b_1 U17779 ( .A_N(n23518), .B(n11163), .Y(n14143) );
  sky130_fd_sc_hd__nand2_1 U17780 ( .A(n13627), .B(
        j202_soc_core_j22_cpu_regop_Rn__0_), .Y(n23518) );
  sky130_fd_sc_hd__inv_2 U17781 ( .A(n26709), .Y(n26426) );
  sky130_fd_sc_hd__o2bb2ai_1 U17782 ( .B1(n13793), .B2(n26325), .A1_N(n26720), 
        .A2_N(n16289), .Y(n14558) );
  sky130_fd_sc_hd__nand2_1 U17783 ( .A(n11953), .B(n11952), .Y(n14560) );
  sky130_fd_sc_hd__nand2_1 U17784 ( .A(n26720), .B(n16261), .Y(n11952) );
  sky130_fd_sc_hd__nand2_1 U17785 ( .A(n26709), .B(n16289), .Y(n11953) );
  sky130_fd_sc_hd__nand3_1 U17786 ( .A(n11960), .B(n11959), .C(n11957), .Y(
        n26883) );
  sky130_fd_sc_hd__nand2_1 U17787 ( .A(n11955), .B(n12158), .Y(n11954) );
  sky130_fd_sc_hd__o21ai_1 U17788 ( .A1(n11910), .A2(n11957), .B1(n16557), .Y(
        n11956) );
  sky130_fd_sc_hd__nand2_1 U17789 ( .A(n11963), .B(n16555), .Y(n25838) );
  sky130_fd_sc_hd__nor2b_1 U17790 ( .B_N(n11961), .A(n16555), .Y(n11958) );
  sky130_fd_sc_hd__nand2_1 U17791 ( .A(n11962), .B(n11961), .Y(n11960) );
  sky130_fd_sc_hd__nand3_1 U17792 ( .A(n23608), .B(n24421), .C(n11965), .Y(
        n27875) );
  sky130_fd_sc_hd__nand3_1 U17793 ( .A(n13071), .B(n12293), .C(n13070), .Y(
        n28975) );
  sky130_fd_sc_hd__nand3_1 U17794 ( .A(n18923), .B(n18921), .C(n21776), .Y(
        n13070) );
  sky130_fd_sc_hd__nand2_1 U17795 ( .A(n28916), .B(n21750), .Y(n13071) );
  sky130_fd_sc_hd__nand4_1 U17796 ( .A(n11969), .B(n11968), .C(n11967), .D(
        n11966), .Y(n12625) );
  sky130_fd_sc_hd__nand2_1 U17797 ( .A(j202_soc_core_memory0_ram_dout0[279]), 
        .B(n21605), .Y(n11966) );
  sky130_fd_sc_hd__nand2_1 U17798 ( .A(j202_soc_core_memory0_ram_dout0[471]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n11967) );
  sky130_fd_sc_hd__nand2_1 U17799 ( .A(j202_soc_core_memory0_ram_dout0[247]), 
        .B(n21735), .Y(n11968) );
  sky130_fd_sc_hd__nand2_1 U17800 ( .A(j202_soc_core_memory0_ram_dout0[311]), 
        .B(n21603), .Y(n11969) );
  sky130_fd_sc_hd__nand2_1 U17801 ( .A(n18923), .B(n18921), .Y(n23753) );
  sky130_fd_sc_hd__nand3_1 U17802 ( .A(n18923), .B(n18921), .C(n22581), .Y(
        n12915) );
  sky130_fd_sc_hd__nand4_1 U17803 ( .A(n13151), .B(n29500), .C(n13150), .D(
        n13147), .Y(n18923) );
  sky130_fd_sc_hd__nand2b_1 U17804 ( .A_N(n23509), .B(n11163), .Y(n12170) );
  sky130_fd_sc_hd__nand2_1 U17805 ( .A(n13626), .B(
        j202_soc_core_j22_cpu_regop_Rn__2_), .Y(n23509) );
  sky130_fd_sc_hd__clkinv_1 U17806 ( .A(n23179), .Y(n22674) );
  sky130_fd_sc_hd__nand2_1 U17807 ( .A(n22670), .B(n11973), .Y(n11972) );
  sky130_fd_sc_hd__o22ai_1 U17809 ( .A1(n11145), .A2(n16492), .B1(n13793), 
        .B2(n26577), .Y(n14127) );
  sky130_fd_sc_hd__nand3_2 U17810 ( .A(n13897), .B(n12249), .C(n13896), .Y(
        n26600) );
  sky130_fd_sc_hd__nand2_1 U17811 ( .A(n11976), .B(n11975), .Y(n14128) );
  sky130_fd_sc_hd__nand2_1 U17812 ( .A(n27409), .B(n16529), .Y(n11975) );
  sky130_fd_sc_hd__nand2_1 U17813 ( .A(n11977), .B(n11146), .Y(n11976) );
  sky130_fd_sc_hd__nor2_1 U17814 ( .A(n21326), .B(n22586), .Y(n11979) );
  sky130_fd_sc_hd__inv_1 U17815 ( .A(n21325), .Y(n11980) );
  sky130_fd_sc_hd__o21a_1 U17816 ( .A1(n11161), .A2(n23697), .B1(n21522), .X(
        n12690) );
  sky130_fd_sc_hd__nand2_1 U17817 ( .A(n21318), .B(n21317), .Y(n23697) );
  sky130_fd_sc_hd__nand2_1 U17818 ( .A(n22242), .B(n22768), .Y(n21565) );
  sky130_fd_sc_hd__o21a_1 U17819 ( .A1(n11985), .A2(n27408), .B1(n11984), .X(
        n11982) );
  sky130_fd_sc_hd__nand2_1 U17820 ( .A(n11986), .B(n26600), .Y(n11983) );
  sky130_fd_sc_hd__o21a_1 U17821 ( .A1(n21525), .A2(n11145), .B1(n21551), .X(
        n11984) );
  sky130_fd_sc_hd__nand2b_1 U17822 ( .A_N(n26352), .B(n26600), .Y(n11985) );
  sky130_fd_sc_hd__nand4_1 U17823 ( .A(n21146), .B(n21147), .C(n21037), .D(
        n21149), .Y(n11987) );
  sky130_fd_sc_hd__and2_0 U17825 ( .A(n21161), .B(n21142), .X(n11989) );
  sky130_fd_sc_hd__nor2b_1 U17826 ( .B_N(n21580), .A(n21579), .Y(n11990) );
  sky130_fd_sc_hd__nand2b_1 U17831 ( .A_N(n21141), .B(n20908), .Y(n21161) );
  sky130_fd_sc_hd__nand2_1 U17833 ( .A(n19354), .B(n17302), .Y(n17278) );
  sky130_fd_sc_hd__nor2_2 U17834 ( .A(n11994), .B(n12136), .Y(n17302) );
  sky130_fd_sc_hd__inv_2 U17835 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .Y(n11994) );
  sky130_fd_sc_hd__inv_2 U17836 ( .A(n21130), .Y(n21274) );
  sky130_fd_sc_hd__nand2b_1 U17837 ( .A_N(n21096), .B(n11995), .Y(n21130) );
  sky130_fd_sc_hd__nand2_1 U17838 ( .A(n21187), .B(n21286), .Y(n21096) );
  sky130_fd_sc_hd__nor2_1 U17839 ( .A(n19298), .B(n19299), .Y(n21187) );
  sky130_fd_sc_hd__nor2_1 U17840 ( .A(n22287), .B(n11996), .Y(n23141) );
  sky130_fd_sc_hd__nor2_1 U17841 ( .A(n11996), .B(n12615), .Y(n13224) );
  sky130_fd_sc_hd__nand2_1 U17844 ( .A(n12000), .B(n11998), .Y(n21318) );
  sky130_fd_sc_hd__nand4_1 U17845 ( .A(n21033), .B(n21032), .C(n21038), .D(
        n21035), .Y(n11999) );
  sky130_fd_sc_hd__inv_2 U17846 ( .A(n13269), .Y(n27260) );
  sky130_fd_sc_hd__inv_2 U17848 ( .A(n22277), .Y(n13152) );
  sky130_fd_sc_hd__inv_2 U17849 ( .A(n22278), .Y(n12595) );
  sky130_fd_sc_hd__nand2_1 U17850 ( .A(j202_soc_core_memory0_ram_dout0[96]), 
        .B(n21591), .Y(n12002) );
  sky130_fd_sc_hd__nand2_1 U17851 ( .A(j202_soc_core_memory0_ram_dout0[128]), 
        .B(n21592), .Y(n12003) );
  sky130_fd_sc_hd__nand2_2 U17852 ( .A(n23184), .B(n24388), .Y(n12712) );
  sky130_fd_sc_hd__inv_1 U17853 ( .A(n12714), .Y(n12004) );
  sky130_fd_sc_hd__nand2_1 U17854 ( .A(n23184), .B(n24388), .Y(n12005) );
  sky130_fd_sc_hd__nand2_1 U17855 ( .A(n12009), .B(n12007), .Y(n12006) );
  sky130_fd_sc_hd__nand3_1 U17856 ( .A(n27261), .B(n24357), .C(n27877), .Y(
        n12008) );
  sky130_fd_sc_hd__nand2_1 U17858 ( .A(n22019), .B(n28972), .Y(n22287) );
  sky130_fd_sc_hd__nand2_1 U17859 ( .A(n12414), .B(n11061), .Y(n12011) );
  sky130_fd_sc_hd__inv_2 U17860 ( .A(n12012), .Y(n27551) );
  sky130_fd_sc_hd__nand2b_1 U17861 ( .A_N(n24353), .B(n24257), .Y(n12388) );
  sky130_fd_sc_hd__nand2_2 U17862 ( .A(n27684), .B(n10975), .Y(n12012) );
  sky130_fd_sc_hd__nand2_1 U17863 ( .A(n12496), .B(n22715), .Y(n22716) );
  sky130_fd_sc_hd__nand2_1 U17864 ( .A(j202_soc_core_memory0_ram_dout0[274]), 
        .B(n21605), .Y(n12014) );
  sky130_fd_sc_hd__nand2_1 U17865 ( .A(j202_soc_core_memory0_ram_dout0[402]), 
        .B(n21597), .Y(n12015) );
  sky130_fd_sc_hd__nand2_1 U17866 ( .A(j202_soc_core_memory0_ram_dout0[466]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12016) );
  sky130_fd_sc_hd__inv_1 U17868 ( .A(n12876), .Y(n12017) );
  sky130_fd_sc_hd__inv_1 U17869 ( .A(n24331), .Y(n12018) );
  sky130_fd_sc_hd__nand2_1 U17870 ( .A(n12019), .B(n12693), .Y(n10581) );
  sky130_fd_sc_hd__nand2_1 U17871 ( .A(n12020), .B(n27980), .Y(n12019) );
  sky130_fd_sc_hd__nor2_1 U17872 ( .A(n12022), .B(n12150), .Y(n12021) );
  sky130_fd_sc_hd__nand3_1 U17874 ( .A(n27558), .B(n12482), .C(n12023), .Y(
        n24337) );
  sky130_fd_sc_hd__inv_2 U17876 ( .A(n12150), .Y(n12023) );
  sky130_fd_sc_hd__nand2_1 U17877 ( .A(n28917), .B(n22581), .Y(n22518) );
  sky130_fd_sc_hd__nand3_1 U17878 ( .A(n26531), .B(n10967), .C(n12024), .Y(
        n26532) );
  sky130_fd_sc_hd__nor2_1 U17879 ( .A(n12030), .B(n12025), .Y(n12978) );
  sky130_fd_sc_hd__nand4_1 U17880 ( .A(n12029), .B(n12028), .C(n12027), .D(
        n12026), .Y(n12025) );
  sky130_fd_sc_hd__nand2_1 U17881 ( .A(j202_soc_core_memory0_ram_dout0[351]), 
        .B(n21593), .Y(n12026) );
  sky130_fd_sc_hd__nand2_1 U17882 ( .A(j202_soc_core_memory0_ram_dout0[255]), 
        .B(n21735), .Y(n12027) );
  sky130_fd_sc_hd__nand2_1 U17883 ( .A(j202_soc_core_memory0_ram_dout0[95]), 
        .B(n21734), .Y(n12028) );
  sky130_fd_sc_hd__nand2_1 U17884 ( .A(j202_soc_core_memory0_ram_dout0[319]), 
        .B(n21603), .Y(n12029) );
  sky130_fd_sc_hd__nand4_1 U17885 ( .A(n12033), .B(n12034), .C(n12032), .D(
        n12031), .Y(n12030) );
  sky130_fd_sc_hd__nand2_1 U17886 ( .A(j202_soc_core_memory0_ram_dout0[223]), 
        .B(n21732), .Y(n12031) );
  sky130_fd_sc_hd__nand2_1 U17887 ( .A(j202_soc_core_memory0_ram_dout0[447]), 
        .B(n21598), .Y(n12032) );
  sky130_fd_sc_hd__nand2_1 U17888 ( .A(j202_soc_core_memory0_ram_dout0[479]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12033) );
  sky130_fd_sc_hd__nand2_1 U17889 ( .A(j202_soc_core_memory0_ram_dout0[415]), 
        .B(n21597), .Y(n12034) );
  sky130_fd_sc_hd__clkbuf_1 U17890 ( .A(n12038), .X(n12035) );
  sky130_fd_sc_hd__nand2_1 U17891 ( .A(n12035), .B(n29075), .Y(n27296) );
  sky130_fd_sc_hd__nand2_1 U17892 ( .A(n12035), .B(n29072), .Y(n25341) );
  sky130_fd_sc_hd__inv_1 U17893 ( .A(n12038), .Y(n12036) );
  sky130_fd_sc_hd__nor2_1 U17894 ( .A(n12038), .B(n24325), .Y(n12423) );
  sky130_fd_sc_hd__nor2_1 U17895 ( .A(n12037), .B(n25814), .Y(n25817) );
  sky130_fd_sc_hd__nand2_1 U17896 ( .A(n27878), .B(n23601), .Y(n12038) );
  sky130_fd_sc_hd__nand3_4 U17897 ( .A(n12041), .B(n12040), .C(n20713), .Y(
        n13180) );
  sky130_fd_sc_hd__nand2_1 U17898 ( .A(n20710), .B(n12289), .Y(n12040) );
  sky130_fd_sc_hd__nor2_1 U17899 ( .A(n27722), .B(n12042), .Y(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_N497) );
  sky130_fd_sc_hd__xnor2_1 U17901 ( .A(n12761), .B(n12760), .Y(n12045) );
  sky130_fd_sc_hd__nand2_1 U17902 ( .A(n12045), .B(n18812), .Y(n22751) );
  sky130_fd_sc_hd__inv_2 U17903 ( .A(n12046), .Y(n27683) );
  sky130_fd_sc_hd__nand4_1 U17904 ( .A(n12049), .B(n12048), .C(n12047), .D(
        n16971), .Y(n12972) );
  sky130_fd_sc_hd__nand2_1 U17905 ( .A(j202_soc_core_memory0_ram_dout0[125]), 
        .B(n21591), .Y(n12047) );
  sky130_fd_sc_hd__nand2_1 U17906 ( .A(j202_soc_core_memory0_ram_dout0[29]), 
        .B(n21733), .Y(n12048) );
  sky130_fd_sc_hd__nand2_1 U17907 ( .A(j202_soc_core_memory0_ram_dout0[157]), 
        .B(n21592), .Y(n12049) );
  sky130_fd_sc_hd__nand3_1 U17909 ( .A(n12894), .B(n15765), .C(n15764), .Y(
        n20714) );
  sky130_fd_sc_hd__nand2_1 U17910 ( .A(n20044), .B(n12287), .Y(n20717) );
  sky130_fd_sc_hd__nand3_1 U17911 ( .A(n12051), .B(n25826), .C(
        j202_soc_core_j22_cpu_ml_macl[5]), .Y(n24063) );
  sky130_fd_sc_hd__nand3_1 U17912 ( .A(n12051), .B(n25826), .C(
        j202_soc_core_j22_cpu_ml_macl[2]), .Y(n24806) );
  sky130_fd_sc_hd__o21ai_1 U17913 ( .A1(n24369), .A2(n24368), .B1(n12051), .Y(
        n24370) );
  sky130_fd_sc_hd__nand2_1 U17914 ( .A(n12051), .B(n25233), .Y(n12785) );
  sky130_fd_sc_hd__nand2_2 U17915 ( .A(n12052), .B(n23257), .Y(n12917) );
  sky130_fd_sc_hd__nand2_1 U17916 ( .A(n12052), .B(n25826), .Y(n12918) );
  sky130_fd_sc_hd__nand3_2 U17917 ( .A(n23269), .B(n12990), .C(n23267), .Y(
        n12052) );
  sky130_fd_sc_hd__nand2_1 U17918 ( .A(n12054), .B(n12053), .Y(n18613) );
  sky130_fd_sc_hd__nand2_1 U17919 ( .A(n18603), .B(n18604), .Y(n12053) );
  sky130_fd_sc_hd__xor2_1 U17921 ( .A(n12057), .B(n12055), .X(n18610) );
  sky130_fd_sc_hd__xnor2_1 U17922 ( .A(n12056), .B(n18603), .Y(n12055) );
  sky130_fd_sc_hd__inv_2 U17923 ( .A(n18604), .Y(n12056) );
  sky130_fd_sc_hd__nand2_1 U17924 ( .A(n18589), .B(n12058), .Y(n12057) );
  sky130_fd_sc_hd__o21ai_1 U17925 ( .A1(n18587), .A2(n18588), .B1(n18586), .Y(
        n12058) );
  sky130_fd_sc_hd__nor2_1 U17926 ( .A(n10938), .B(n27875), .Y(n12288) );
  sky130_fd_sc_hd__nand2_1 U17928 ( .A(n12064), .B(n29077), .Y(n12290) );
  sky130_fd_sc_hd__nand2_1 U17929 ( .A(n12064), .B(n12376), .Y(n12291) );
  sky130_fd_sc_hd__inv_2 U17930 ( .A(n12064), .Y(n12062) );
  sky130_fd_sc_hd__nand2_1 U17931 ( .A(n27522), .B(n12063), .Y(n10491) );
  sky130_fd_sc_hd__nand2_1 U17932 ( .A(n12064), .B(n11133), .Y(n12063) );
  sky130_fd_sc_hd__inv_1 U17933 ( .A(n23605), .Y(n27934) );
  sky130_fd_sc_hd__nand2_1 U17934 ( .A(n12067), .B(n12066), .Y(n23605) );
  sky130_fd_sc_hd__inv_1 U17935 ( .A(n29548), .Y(n12066) );
  sky130_fd_sc_hd__inv_1 U17936 ( .A(n27890), .Y(n12067) );
  sky130_fd_sc_hd__nand2_1 U17937 ( .A(n12069), .B(n13544), .Y(n12068) );
  sky130_fd_sc_hd__nand2_1 U17938 ( .A(n12070), .B(n13542), .Y(n12069) );
  sky130_fd_sc_hd__nand2_1 U17939 ( .A(n13543), .B(n13638), .Y(n12070) );
  sky130_fd_sc_hd__nand2_1 U17940 ( .A(n12072), .B(n23861), .Y(n27928) );
  sky130_fd_sc_hd__nand2_1 U17941 ( .A(n12072), .B(
        j202_soc_core_j22_cpu_pc_hold), .Y(n27956) );
  sky130_fd_sc_hd__nand2b_1 U17942 ( .A_N(n12072), .B(n27176), .Y(n10607) );
  sky130_fd_sc_hd__nand2_1 U17943 ( .A(n29015), .B(n12072), .Y(n24303) );
  sky130_fd_sc_hd__nand3_1 U17944 ( .A(n12073), .B(n12279), .C(n28962), .Y(
        n17127) );
  sky130_fd_sc_hd__nand4_1 U17945 ( .A(n12075), .B(n12076), .C(n12074), .D(
        n12077), .Y(n12849) );
  sky130_fd_sc_hd__nand2_1 U17946 ( .A(j202_soc_core_memory0_ram_dout0[213]), 
        .B(n21732), .Y(n12074) );
  sky130_fd_sc_hd__nand2_1 U17947 ( .A(j202_soc_core_memory0_ram_dout0[21]), 
        .B(n21733), .Y(n12075) );
  sky130_fd_sc_hd__nand2_1 U17948 ( .A(j202_soc_core_memory0_ram_dout0[85]), 
        .B(n21734), .Y(n12076) );
  sky130_fd_sc_hd__nand2_1 U17949 ( .A(j202_soc_core_memory0_ram_dout0[245]), 
        .B(n21735), .Y(n12077) );
  sky130_fd_sc_hd__nand4b_1 U17950 ( .A_N(n12079), .B(n26552), .C(n26551), .D(
        n26553), .Y(n26554) );
  sky130_fd_sc_hd__nand3_1 U17951 ( .A(n13231), .B(n20834), .C(n21753), .Y(
        n12080) );
  sky130_fd_sc_hd__nand2_1 U17952 ( .A(n20833), .B(n13288), .Y(n13231) );
  sky130_fd_sc_hd__clkinv_1 U17953 ( .A(n12080), .Y(n12081) );
  sky130_fd_sc_hd__nand2_1 U17954 ( .A(n13230), .B(n13199), .Y(n12083) );
  sky130_fd_sc_hd__nand2_1 U17955 ( .A(n21752), .B(n12084), .Y(n13199) );
  sky130_fd_sc_hd__nand4_1 U17957 ( .A(n13061), .B(n16672), .C(n13060), .D(
        n16665), .Y(n12086) );
  sky130_fd_sc_hd__nor2_1 U17958 ( .A(n12090), .B(n12089), .Y(n12088) );
  sky130_fd_sc_hd__nand4_1 U17959 ( .A(n16671), .B(n13062), .C(n16666), .D(
        n16669), .Y(n12089) );
  sky130_fd_sc_hd__nand4_1 U17960 ( .A(n13057), .B(n13058), .C(n16667), .D(
        n16796), .Y(n12090) );
  sky130_fd_sc_hd__nand2_1 U17961 ( .A(n12091), .B(n12471), .Y(
        j202_soc_core_j22_cpu_id_idec_N937) );
  sky130_fd_sc_hd__nand2_1 U17962 ( .A(n12092), .B(n27980), .Y(n12091) );
  sky130_fd_sc_hd__nand4_1 U17963 ( .A(n12093), .B(n27939), .C(n12327), .D(
        n27938), .Y(n12092) );
  sky130_fd_sc_hd__nand2_1 U17964 ( .A(n12105), .B(n12094), .Y(n21755) );
  sky130_fd_sc_hd__nand4_1 U17965 ( .A(n12099), .B(n12098), .C(n12097), .D(
        n12096), .Y(n12095) );
  sky130_fd_sc_hd__nand2_1 U17966 ( .A(j202_soc_core_memory0_ram_dout0[101]), 
        .B(n21591), .Y(n12096) );
  sky130_fd_sc_hd__nand2_1 U17967 ( .A(j202_soc_core_memory0_ram_dout0[165]), 
        .B(n21590), .Y(n12097) );
  sky130_fd_sc_hd__nand2_1 U17968 ( .A(j202_soc_core_memory0_ram_dout0[5]), 
        .B(n21733), .Y(n12098) );
  sky130_fd_sc_hd__nand2_1 U17969 ( .A(j202_soc_core_memory0_ram_dout0[229]), 
        .B(n21735), .Y(n12099) );
  sky130_fd_sc_hd__nand4_1 U17970 ( .A(n12104), .B(n12103), .C(n12102), .D(
        n12101), .Y(n12100) );
  sky130_fd_sc_hd__nand2_1 U17971 ( .A(j202_soc_core_memory0_ram_dout0[69]), 
        .B(n21734), .Y(n12101) );
  sky130_fd_sc_hd__nand2_1 U17972 ( .A(j202_soc_core_memory0_ram_dout0[261]), 
        .B(n21605), .Y(n12102) );
  sky130_fd_sc_hd__nand2_1 U17973 ( .A(j202_soc_core_memory0_ram_dout0[37]), 
        .B(n21604), .Y(n12103) );
  sky130_fd_sc_hd__nand2_1 U17974 ( .A(j202_soc_core_memory0_ram_dout0[293]), 
        .B(n21603), .Y(n12104) );
  sky130_fd_sc_hd__nand4_1 U17975 ( .A(n21599), .B(n21600), .C(n21601), .D(
        n21602), .Y(n12106) );
  sky130_fd_sc_hd__nand4_1 U17976 ( .A(n13073), .B(n21594), .C(n21595), .D(
        n21731), .Y(n12107) );
  sky130_fd_sc_hd__a22oi_1 U17978 ( .A1(n11669), .A2(n23762), .B1(n12771), 
        .B2(n23777), .Y(n26543) );
  sky130_fd_sc_hd__inv_2 U17979 ( .A(n24226), .Y(n24227) );
  sky130_fd_sc_hd__nand4_1 U17980 ( .A(n12968), .B(n12967), .C(n12965), .D(
        n12966), .Y(n12109) );
  sky130_fd_sc_hd__inv_2 U17981 ( .A(n24195), .Y(n24196) );
  sky130_fd_sc_hd__inv_1 U17982 ( .A(n13121), .Y(n13120) );
  sky130_fd_sc_hd__or2_0 U17984 ( .A(n27228), .B(n27461), .X(n12110) );
  sky130_fd_sc_hd__nand2_1 U17985 ( .A(n12110), .B(n24560), .Y(
        j202_soc_core_j22_cpu_rf_N3173) );
  sky130_fd_sc_hd__nand2_1 U17986 ( .A(n26323), .B(n27364), .Y(n12112) );
  sky130_fd_sc_hd__inv_2 U17987 ( .A(n24217), .Y(n24218) );
  sky130_fd_sc_hd__nand2_1 U17988 ( .A(n23981), .B(n23980), .Y(n24001) );
  sky130_fd_sc_hd__inv_1 U17989 ( .A(n12842), .Y(n24106) );
  sky130_fd_sc_hd__nand2_1 U17990 ( .A(n24350), .B(n12150), .Y(n12115) );
  sky130_fd_sc_hd__nand2_1 U17991 ( .A(n11069), .B(n12116), .Y(n27773) );
  sky130_fd_sc_hd__inv_1 U17992 ( .A(n12115), .Y(n12116) );
  sky130_fd_sc_hd__nor2_1 U17993 ( .A(n24295), .B(n12114), .Y(n24296) );
  sky130_fd_sc_hd__inv_2 U17994 ( .A(n11771), .Y(n27359) );
  sky130_fd_sc_hd__nor2_1 U17995 ( .A(n13233), .B(n12238), .Y(n12117) );
  sky130_fd_sc_hd__a22oi_1 U17996 ( .A1(j202_soc_core_memory0_ram_dout0[457]), 
        .A2(j202_soc_core_memory0_ram_dout0_sel[14]), .B1(n21598), .B2(
        j202_soc_core_memory0_ram_dout0[425]), .Y(n20933) );
  sky130_fd_sc_hd__xnor2_1 U17997 ( .A(n17431), .B(n12711), .Y(n17560) );
  sky130_fd_sc_hd__buf_6 U18002 ( .A(n24216), .X(n12121) );
  sky130_fd_sc_hd__inv_2 U18003 ( .A(n24215), .Y(n24216) );
  sky130_fd_sc_hd__inv_2 U18004 ( .A(n24201), .Y(n24202) );
  sky130_fd_sc_hd__nand2_1 U18005 ( .A(n17145), .B(n12416), .Y(n24127) );
  sky130_fd_sc_hd__inv_2 U18006 ( .A(n18291), .Y(n18292) );
  sky130_fd_sc_hd__buf_6 U18007 ( .A(n24220), .X(n29305) );
  sky130_fd_sc_hd__inv_2 U18008 ( .A(n24219), .Y(n24220) );
  sky130_fd_sc_hd__nor2_1 U18009 ( .A(n27928), .B(n13187), .Y(n24410) );
  sky130_fd_sc_hd__nand3_1 U18010 ( .A(n27171), .B(n13083), .C(n24455), .Y(
        n23159) );
  sky130_fd_sc_hd__o21ai_2 U18012 ( .A1(n23539), .A2(n23543), .B1(n23178), .Y(
        j202_soc_core_j22_cpu_rf_N3079) );
  sky130_fd_sc_hd__inv_1 U18013 ( .A(n13008), .Y(n20560) );
  sky130_fd_sc_hd__nand2_1 U18014 ( .A(n22027), .B(n27947), .Y(n29079) );
  sky130_fd_sc_hd__inv_1 U18015 ( .A(n23161), .Y(n23139) );
  sky130_fd_sc_hd__mux2_2 U18016 ( .A0(n19777), .A1(n19776), .S(n11700), .X(
        n12126) );
  sky130_fd_sc_hd__o22ai_1 U18017 ( .A1(n19664), .A2(n19651), .B1(n13027), 
        .B2(n13024), .Y(n12127) );
  sky130_fd_sc_hd__mux2_2 U18018 ( .A0(n19646), .A1(n19645), .S(n25769), .X(
        n19776) );
  sky130_fd_sc_hd__inv_1 U18019 ( .A(n20714), .Y(n12914) );
  sky130_fd_sc_hd__nor2_1 U18020 ( .A(n29009), .B(n13140), .Y(n13115) );
  sky130_fd_sc_hd__inv_2 U18021 ( .A(n24211), .Y(n24212) );
  sky130_fd_sc_hd__o2bb2ai_1 U18022 ( .B1(n27467), .B2(n11141), .A1_N(n11141), 
        .A2_N(n12151), .Y(j202_soc_core_j22_cpu_rf_N2686) );
  sky130_fd_sc_hd__buf_6 U18024 ( .A(n24222), .X(n29307) );
  sky130_fd_sc_hd__inv_2 U18025 ( .A(n24221), .Y(n24222) );
  sky130_fd_sc_hd__nor2_1 U18026 ( .A(n12109), .B(n12960), .Y(n12130) );
  sky130_fd_sc_hd__o211ai_2 U18027 ( .A1(n26352), .A2(n26912), .B1(n21819), 
        .C1(n21818), .Y(n21820) );
  sky130_fd_sc_hd__inv_2 U18028 ( .A(n24182), .Y(n24183) );
  sky130_fd_sc_hd__a21oi_1 U18029 ( .A1(n20955), .A2(n20956), .B1(n12191), .Y(
        n28970) );
  sky130_fd_sc_hd__inv_2 U18030 ( .A(n24176), .Y(n24177) );
  sky130_fd_sc_hd__inv_4 U18031 ( .A(n19249), .Y(n22912) );
  sky130_fd_sc_hd__nand2_1 U18032 ( .A(n24109), .B(n13083), .Y(n27882) );
  sky130_fd_sc_hd__buf_2 U18034 ( .A(n18366), .X(n12131) );
  sky130_fd_sc_hd__xnor2_1 U18035 ( .A(j202_soc_core_j22_cpu_ml_bufa[24]), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .Y(n18366) );
  sky130_fd_sc_hd__nand3_1 U18036 ( .A(n24347), .B(n27877), .C(n24452), .Y(
        n23147) );
  sky130_fd_sc_hd__buf_6 U18037 ( .A(n24198), .X(n29278) );
  sky130_fd_sc_hd__inv_2 U18038 ( .A(n24197), .Y(n24198) );
  sky130_fd_sc_hd__inv_2 U18039 ( .A(n24180), .Y(n24181) );
  sky130_fd_sc_hd__inv_2 U18040 ( .A(n24199), .Y(n24200) );
  sky130_fd_sc_hd__o22a_1 U18041 ( .A1(n11161), .A2(n12877), .B1(n21915), .B2(
        n26535), .X(n19168) );
  sky130_fd_sc_hd__nand2_2 U18042 ( .A(n12436), .B(n11646), .Y(n24307) );
  sky130_fd_sc_hd__inv_2 U18043 ( .A(n24206), .Y(n24207) );
  sky130_fd_sc_hd__nand2_2 U18046 ( .A(n12641), .B(n27683), .Y(n13179) );
  sky130_fd_sc_hd__inv_2 U18047 ( .A(n12954), .Y(n24205) );
  sky130_fd_sc_hd__inv_2 U18048 ( .A(n24178), .Y(n24179) );
  sky130_fd_sc_hd__nand3_1 U18050 ( .A(n22257), .B(n22256), .C(n22255), .Y(
        n29004) );
  sky130_fd_sc_hd__a2bb2oi_2 U18051 ( .B1(n18978), .B2(n20830), .A1_N(n18977), 
        .A2_N(j202_soc_core_memory0_ram_dout0[495]), .Y(n20145) );
  sky130_fd_sc_hd__inv_1 U18053 ( .A(n12501), .Y(n24437) );
  sky130_fd_sc_hd__nand3_1 U18055 ( .A(n12313), .B(n23278), .C(n25336), .Y(
        n22245) );
  sky130_fd_sc_hd__nor2_1 U18056 ( .A(n23136), .B(n27876), .Y(n24458) );
  sky130_fd_sc_hd__inv_1 U18057 ( .A(n12483), .Y(n12139) );
  sky130_fd_sc_hd__inv_2 U18058 ( .A(n23973), .Y(n23974) );
  sky130_fd_sc_hd__buf_2 U18059 ( .A(n17426), .X(n12133) );
  sky130_fd_sc_hd__buf_4 U18060 ( .A(n17387), .X(n17972) );
  sky130_fd_sc_hd__a22oi_2 U18061 ( .A1(n13229), .A2(n27980), .B1(n12912), 
        .B2(n12227), .Y(n12377) );
  sky130_fd_sc_hd__o22ai_1 U18063 ( .A1(n18660), .A2(n18137), .B1(n18109), 
        .B2(n12991), .Y(n18134) );
  sky130_fd_sc_hd__nand2_1 U18064 ( .A(n24335), .B(n27556), .Y(n23210) );
  sky130_fd_sc_hd__and2_4 U18065 ( .A(n18871), .B(n17357), .X(n12134) );
  sky130_fd_sc_hd__inv_1 U18066 ( .A(n17815), .Y(n12790) );
  sky130_fd_sc_hd__clkbuf_1 U18068 ( .A(j202_soc_core_j22_cpu_ml_bufa[21]), 
        .X(n12138) );
  sky130_fd_sc_hd__nor2_4 U18069 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .B(n17175), .Y(n13388) );
  sky130_fd_sc_hd__xnor2_1 U18070 ( .A(n18523), .B(n18507), .Y(n18550) );
  sky130_fd_sc_hd__inv_1 U18071 ( .A(n12483), .Y(n12140) );
  sky130_fd_sc_hd__inv_1 U18072 ( .A(n12483), .Y(n18514) );
  sky130_fd_sc_hd__buf_4 U18073 ( .A(n12303), .X(n12141) );
  sky130_fd_sc_hd__o22a_4 U18075 ( .A1(n17142), .A2(n21022), .B1(n17140), .B2(
        n17141), .X(n12416) );
  sky130_fd_sc_hd__inv_2 U18076 ( .A(n23126), .Y(n23130) );
  sky130_fd_sc_hd__inv_2 U18077 ( .A(n13396), .Y(n17277) );
  sky130_fd_sc_hd__inv_2 U18078 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .Y(n13396) );
  sky130_fd_sc_hd__inv_6 U18079 ( .A(n29249), .Y(n12517) );
  sky130_fd_sc_hd__nand2_1 U18080 ( .A(n12146), .B(n27006), .Y(
        j202_soc_core_j22_cpu_ml_N323) );
  sky130_fd_sc_hd__nand2_1 U18081 ( .A(n11166), .B(n12147), .Y(n12146) );
  sky130_fd_sc_hd__inv_6 U18085 ( .A(n29248), .Y(n12531) );
  sky130_fd_sc_hd__inv_6 U18086 ( .A(n29248), .Y(n12524) );
  sky130_fd_sc_hd__nand2_1 U18087 ( .A(n17274), .B(n17289), .Y(n15423) );
  sky130_fd_sc_hd__clkinv_1 U18088 ( .A(n14884), .Y(n15425) );
  sky130_fd_sc_hd__nand2_1 U18089 ( .A(n18915), .B(n24279), .Y(n16054) );
  sky130_fd_sc_hd__and2_0 U18090 ( .A(n16782), .B(n16781), .X(n16784) );
  sky130_fd_sc_hd__inv_2 U18092 ( .A(n14749), .Y(n13774) );
  sky130_fd_sc_hd__nor2_1 U18093 ( .A(n18830), .B(n18829), .Y(n18807) );
  sky130_fd_sc_hd__and2_0 U18094 ( .A(n20908), .B(n21251), .X(n13275) );
  sky130_fd_sc_hd__clkinv_1 U18095 ( .A(n20873), .Y(n20892) );
  sky130_fd_sc_hd__nand3_1 U18096 ( .A(n23770), .B(n26443), .C(n26717), .Y(
        n24537) );
  sky130_fd_sc_hd__nor2_1 U18097 ( .A(n12505), .B(n13702), .Y(n13706) );
  sky130_fd_sc_hd__and2_0 U18098 ( .A(n19516), .B(n19517), .X(n19529) );
  sky130_fd_sc_hd__clkinv_1 U18099 ( .A(n27914), .Y(n13602) );
  sky130_fd_sc_hd__nand2_1 U18100 ( .A(n26260), .B(n26202), .Y(n28743) );
  sky130_fd_sc_hd__inv_2 U18101 ( .A(n25219), .Y(n24499) );
  sky130_fd_sc_hd__clkinv_1 U18102 ( .A(j202_soc_core_j22_cpu_memop_MEM__0_), 
        .Y(n27721) );
  sky130_fd_sc_hd__clkinv_1 U18103 ( .A(j202_soc_core_j22_cpu_memop_MEM__2_), 
        .Y(n24279) );
  sky130_fd_sc_hd__nand2_1 U18104 ( .A(n27232), .B(n29514), .Y(n27794) );
  sky130_fd_sc_hd__nor2_1 U18105 ( .A(n12141), .B(n18467), .Y(n18488) );
  sky130_fd_sc_hd__nor2_1 U18106 ( .A(n12141), .B(n18368), .Y(n18406) );
  sky130_fd_sc_hd__o22ai_1 U18107 ( .A1(n18224), .A2(n18105), .B1(n18064), 
        .B2(n18225), .Y(n18100) );
  sky130_fd_sc_hd__o22ai_1 U18108 ( .A1(n18514), .A2(n18377), .B1(n18376), 
        .B2(n18424), .Y(n18383) );
  sky130_fd_sc_hd__o22ai_1 U18109 ( .A1(n18067), .A2(n17978), .B1(n17944), 
        .B2(n18068), .Y(n17964) );
  sky130_fd_sc_hd__and2_0 U18110 ( .A(n15615), .B(n15593), .X(n15344) );
  sky130_fd_sc_hd__buf_2 U18111 ( .A(j202_soc_core_j22_cpu_ml_bufb[6]), .X(
        n18667) );
  sky130_fd_sc_hd__o21ai_1 U18112 ( .A1(n19222), .A2(n21437), .B1(n21438), .Y(
        n21875) );
  sky130_fd_sc_hd__and2_0 U18113 ( .A(n20532), .B(n20502), .X(n20516) );
  sky130_fd_sc_hd__and2_0 U18115 ( .A(n20574), .B(n20571), .X(n20584) );
  sky130_fd_sc_hd__clkinv_1 U18116 ( .A(n20885), .Y(n20245) );
  sky130_fd_sc_hd__and2_0 U18117 ( .A(n20741), .B(n20772), .X(n21191) );
  sky130_fd_sc_hd__clkinv_1 U18118 ( .A(n21077), .Y(n21042) );
  sky130_fd_sc_hd__clkinv_1 U18119 ( .A(n17279), .Y(n19355) );
  sky130_fd_sc_hd__and2_0 U18120 ( .A(n21706), .B(n21186), .X(n21680) );
  sky130_fd_sc_hd__and2_0 U18121 ( .A(n20118), .B(n20843), .X(n20003) );
  sky130_fd_sc_hd__clkinv_1 U18122 ( .A(n17169), .Y(n17301) );
  sky130_fd_sc_hd__inv_2 U18123 ( .A(n20221), .Y(n20059) );
  sky130_fd_sc_hd__clkinv_1 U18124 ( .A(n18267), .Y(n12444) );
  sky130_fd_sc_hd__nand2_1 U18125 ( .A(n25259), .B(n24793), .Y(n24794) );
  sky130_fd_sc_hd__and2_0 U18126 ( .A(n22469), .B(n22474), .X(n22477) );
  sky130_fd_sc_hd__clkinv_1 U18127 ( .A(n22907), .Y(n21974) );
  sky130_fd_sc_hd__inv_2 U18128 ( .A(n22065), .Y(n22068) );
  sky130_fd_sc_hd__clkinv_1 U18129 ( .A(n21491), .Y(n21868) );
  sky130_fd_sc_hd__nor4_1 U18131 ( .A(n21043), .B(n21042), .C(n21176), .D(
        n21227), .Y(n21136) );
  sky130_fd_sc_hd__clkinv_1 U18132 ( .A(n16596), .Y(n16945) );
  sky130_fd_sc_hd__and2_0 U18133 ( .A(n13481), .B(n16919), .X(n16937) );
  sky130_fd_sc_hd__and2_0 U18134 ( .A(j202_soc_core_j22_cpu_ma_M_area[1]), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[6]), .X(n13409) );
  sky130_fd_sc_hd__and2_0 U18135 ( .A(n20908), .B(n21235), .X(n21063) );
  sky130_fd_sc_hd__clkinv_1 U18136 ( .A(n21722), .Y(n21251) );
  sky130_fd_sc_hd__nand2_1 U18137 ( .A(n20778), .B(n17314), .Y(n21221) );
  sky130_fd_sc_hd__and2_0 U18138 ( .A(n21613), .B(n20772), .X(n17328) );
  sky130_fd_sc_hd__clkinv_1 U18139 ( .A(n20860), .Y(n21675) );
  sky130_fd_sc_hd__buf_2 U18141 ( .A(j202_soc_core_bootrom_00_address_w[7]), 
        .X(n17289) );
  sky130_fd_sc_hd__nor2_1 U18142 ( .A(j202_soc_core_memory0_ram_dout0_sel[11]), 
        .B(n13501), .Y(n13487) );
  sky130_fd_sc_hd__nand3_1 U18143 ( .A(n19666), .B(n25461), .C(
        j202_soc_core_intc_core_00_rg_ipr[40]), .Y(n19667) );
  sky130_fd_sc_hd__nor2_1 U18144 ( .A(n24792), .B(n12983), .Y(n12982) );
  sky130_fd_sc_hd__inv_2 U18145 ( .A(n26333), .Y(n26077) );
  sky130_fd_sc_hd__o22ai_1 U18146 ( .A1(n18882), .A2(n22806), .B1(n22724), 
        .B2(n18307), .Y(n17815) );
  sky130_fd_sc_hd__clkinv_1 U18147 ( .A(j202_soc_core_j22_cpu_rfuo_sr__t_), 
        .Y(n23928) );
  sky130_fd_sc_hd__and2_0 U18148 ( .A(n19196), .B(n19195), .X(n13338) );
  sky130_fd_sc_hd__clkinv_1 U18149 ( .A(j202_soc_core_bootrom_00_address_w[7]), 
        .Y(n17293) );
  sky130_fd_sc_hd__clkinv_1 U18150 ( .A(n21705), .Y(n21235) );
  sky130_fd_sc_hd__clkinv_1 U18151 ( .A(n21720), .Y(n21288) );
  sky130_fd_sc_hd__a21boi_0 U18152 ( .A1(j202_soc_core_memory0_ram_dout0[361]), 
        .A2(n21596), .B1_N(n20932), .Y(n20934) );
  sky130_fd_sc_hd__nor2_1 U18153 ( .A(n24778), .B(n13142), .Y(n13141) );
  sky130_fd_sc_hd__nand2_1 U18154 ( .A(n13068), .B(n21813), .Y(n13067) );
  sky130_fd_sc_hd__nand4bb_1 U18155 ( .A_N(n26643), .B_N(n26642), .C(n26641), 
        .D(n26640), .Y(n26753) );
  sky130_fd_sc_hd__nand4bb_1 U18156 ( .A_N(n26678), .B_N(n26677), .C(n26676), 
        .D(n26675), .Y(n26754) );
  sky130_fd_sc_hd__inv_2 U18157 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(
        n26690) );
  sky130_fd_sc_hd__and2_0 U18158 ( .A(n25836), .B(n25835), .X(n13342) );
  sky130_fd_sc_hd__nor2_1 U18159 ( .A(n12345), .B(n12344), .Y(n12343) );
  sky130_fd_sc_hd__nor2_1 U18160 ( .A(n12334), .B(n12339), .Y(n12333) );
  sky130_fd_sc_hd__a21oi_1 U18162 ( .A1(n29075), .A2(n29036), .B1(n11793), .Y(
        n13076) );
  sky130_fd_sc_hd__clkinv_1 U18163 ( .A(n17171), .Y(n20378) );
  sky130_fd_sc_hd__clkinv_1 U18164 ( .A(n19856), .Y(n21727) );
  sky130_fd_sc_hd__clkinv_1 U18165 ( .A(
        j202_soc_core_memory0_ram_dout0_sel[10]), .Y(n13500) );
  sky130_fd_sc_hd__nor2_1 U18167 ( .A(j202_soc_core_memory0_ram_dout0_sel[10]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[9]), .Y(n13486) );
  sky130_fd_sc_hd__inv_2 U18168 ( .A(n13481), .Y(n21179) );
  sky130_fd_sc_hd__clkinv_1 U18170 ( .A(j202_soc_core_memory0_ram_dout0_sel[8]), .Y(n13371) );
  sky130_fd_sc_hd__mux2_2 U18171 ( .A0(n19650), .A1(n19649), .S(n25769), .X(
        n19770) );
  sky130_fd_sc_hd__clkinv_1 U18172 ( .A(n19825), .Y(n13023) );
  sky130_fd_sc_hd__nand2_1 U18173 ( .A(n19577), .B(n19576), .Y(n26839) );
  sky130_fd_sc_hd__a21oi_1 U18174 ( .A1(n19707), .A2(n19706), .B1(n19705), .Y(
        n19720) );
  sky130_fd_sc_hd__a2bb2oi_1 U18175 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[59]), .B2(n25501), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[62]), .A2_N(n25087), .Y(n19702) );
  sky130_fd_sc_hd__and2_0 U18177 ( .A(n29056), .B(
        j202_soc_core_wbqspiflash_00_spi_spd), .X(n26203) );
  sky130_fd_sc_hd__and2_0 U18178 ( .A(n24865), .B(n24864), .X(n24869) );
  sky130_fd_sc_hd__and2_0 U18179 ( .A(n23681), .B(n23680), .X(n23682) );
  sky130_fd_sc_hd__clkinv_1 U18181 ( .A(n20152), .Y(n27603) );
  sky130_fd_sc_hd__nand2_1 U18182 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[0]), .Y(n23012) );
  sky130_fd_sc_hd__inv_2 U18183 ( .A(n21926), .Y(n22721) );
  sky130_fd_sc_hd__clkinv_1 U18184 ( .A(n24168), .Y(n13064) );
  sky130_fd_sc_hd__nor2_1 U18186 ( .A(n23212), .B(n12511), .Y(n27169) );
  sky130_fd_sc_hd__clkinv_1 U18187 ( .A(n13549), .Y(n23493) );
  sky130_fd_sc_hd__nand3_1 U18188 ( .A(n11521), .B(n24785), .C(n12152), .Y(
        n23915) );
  sky130_fd_sc_hd__inv_2 U18190 ( .A(n13051), .Y(n12482) );
  sky130_fd_sc_hd__clkinv_1 U18191 ( .A(n22545), .Y(n23574) );
  sky130_fd_sc_hd__o21ai_1 U18192 ( .A1(n16991), .A2(n17110), .B1(n16990), .Y(
        n16992) );
  sky130_fd_sc_hd__clkinv_1 U18193 ( .A(n24046), .Y(n12688) );
  sky130_fd_sc_hd__nor2_1 U18194 ( .A(n13262), .B(n13263), .Y(n13264) );
  sky130_fd_sc_hd__nand3_1 U18195 ( .A(n19327), .B(n12206), .C(n19326), .Y(
        n13262) );
  sky130_fd_sc_hd__nor2_1 U18196 ( .A(n22923), .B(n22965), .Y(n21972) );
  sky130_fd_sc_hd__nand2_1 U18197 ( .A(n25826), .B(n11713), .Y(n22925) );
  sky130_fd_sc_hd__and2_0 U18198 ( .A(n21312), .B(n21311), .X(n21314) );
  sky130_fd_sc_hd__clkinv_1 U18199 ( .A(j202_soc_core_wbqspiflash_00_state[3]), 
        .Y(n26042) );
  sky130_fd_sc_hd__nand2_1 U18201 ( .A(j202_soc_core_memory0_ram_dout0[288]), 
        .B(n21603), .Y(n12808) );
  sky130_fd_sc_hd__nor2_1 U18202 ( .A(n28590), .B(n19828), .Y(n13020) );
  sky130_fd_sc_hd__inv_2 U18203 ( .A(n19620), .Y(n26838) );
  sky130_fd_sc_hd__clkinv_1 U18204 ( .A(n19720), .Y(n26829) );
  sky130_fd_sc_hd__nor2_1 U18205 ( .A(n13561), .B(n13560), .Y(n23485) );
  sky130_fd_sc_hd__nand3_1 U18206 ( .A(n27650), .B(n29593), .C(n27649), .Y(
        n27660) );
  sky130_fd_sc_hd__nand2_1 U18207 ( .A(n27823), .B(n12691), .Y(n17144) );
  sky130_fd_sc_hd__clkinv_1 U18208 ( .A(j202_soc_core_qspi_wb_addr[20]), .Y(
        n28068) );
  sky130_fd_sc_hd__clkinv_1 U18210 ( .A(n28740), .Y(n28719) );
  sky130_fd_sc_hd__clkinv_1 U18211 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[0]), 
        .Y(n28753) );
  sky130_fd_sc_hd__and2_0 U18212 ( .A(n28230), .B(n25955), .X(n28260) );
  sky130_fd_sc_hd__clkinv_1 U18213 ( .A(n27473), .Y(n27482) );
  sky130_fd_sc_hd__clkinv_1 U18214 ( .A(n24478), .Y(n12618) );
  sky130_fd_sc_hd__clkinv_1 U18215 ( .A(n27489), .Y(n26301) );
  sky130_fd_sc_hd__clkinv_1 U18216 ( .A(n26284), .Y(n28619) );
  sky130_fd_sc_hd__clkinv_1 U18217 ( .A(n27676), .Y(n27851) );
  sky130_fd_sc_hd__clkinv_1 U18218 ( .A(n27581), .Y(n28536) );
  sky130_fd_sc_hd__clkinv_1 U18219 ( .A(n27583), .Y(n28538) );
  sky130_fd_sc_hd__nor2_1 U18220 ( .A(n28590), .B(n27583), .Y(n27581) );
  sky130_fd_sc_hd__clkinv_1 U18221 ( .A(n27008), .Y(n28542) );
  sky130_fd_sc_hd__clkinv_1 U18222 ( .A(n27010), .Y(n28544) );
  sky130_fd_sc_hd__nor2_1 U18223 ( .A(n28590), .B(n27010), .Y(n27008) );
  sky130_fd_sc_hd__clkinv_1 U18224 ( .A(n27754), .Y(n28545) );
  sky130_fd_sc_hd__clkinv_1 U18225 ( .A(n27757), .Y(n28547) );
  sky130_fd_sc_hd__nor2_1 U18226 ( .A(n28590), .B(n27757), .Y(n27754) );
  sky130_fd_sc_hd__clkinv_1 U18227 ( .A(n27152), .Y(n28533) );
  sky130_fd_sc_hd__clkinv_1 U18228 ( .A(n27154), .Y(n28535) );
  sky130_fd_sc_hd__nor2_1 U18229 ( .A(n28590), .B(n27154), .Y(n27152) );
  sky130_fd_sc_hd__nand2_1 U18230 ( .A(n28526), .B(n29594), .Y(n28524) );
  sky130_fd_sc_hd__a21oi_1 U18231 ( .A1(n27641), .A2(n27656), .B1(n28590), .Y(
        n28476) );
  sky130_fd_sc_hd__nand2_1 U18232 ( .A(j202_soc_core_qspi_wb_wdat[2]), .B(
        n29594), .Y(n28615) );
  sky130_fd_sc_hd__nand2_1 U18233 ( .A(j202_soc_core_qspi_wb_wdat[16]), .B(
        n29594), .Y(n28606) );
  sky130_fd_sc_hd__clkinv_1 U18234 ( .A(n12162), .Y(n12898) );
  sky130_fd_sc_hd__nor2_1 U18235 ( .A(n26014), .B(n25993), .Y(n28215) );
  sky130_fd_sc_hd__nand2_1 U18236 ( .A(n28737), .B(
        j202_soc_core_wbqspiflash_00_spi_spd), .Y(n28723) );
  sky130_fd_sc_hd__clkinv_1 U18237 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .Y(n28058) );
  sky130_fd_sc_hd__and2_0 U18238 ( .A(n12726), .B(n22502), .X(n12295) );
  sky130_fd_sc_hd__inv_2 U18239 ( .A(n27047), .Y(n26865) );
  sky130_fd_sc_hd__and2_0 U18240 ( .A(n25081), .B(n22406), .X(n13319) );
  sky130_fd_sc_hd__clkinv_1 U18241 ( .A(n18883), .Y(n25264) );
  sky130_fd_sc_hd__inv_2 U18242 ( .A(n26507), .Y(n27407) );
  sky130_fd_sc_hd__inv_2 U18243 ( .A(n19012), .Y(n17718) );
  sky130_fd_sc_hd__clkinv_1 U18244 ( .A(n25824), .Y(n25344) );
  sky130_fd_sc_hd__clkinv_1 U18245 ( .A(j202_soc_core_j22_cpu_macop_MAC_[0]), 
        .Y(n26398) );
  sky130_fd_sc_hd__and2_0 U18246 ( .A(n16030), .B(n16029), .X(n16145) );
  sky130_fd_sc_hd__clkinv_1 U18247 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[0]), 
        .Y(n27137) );
  sky130_fd_sc_hd__inv_1 U18248 ( .A(n23039), .Y(n26360) );
  sky130_fd_sc_hd__clkinv_1 U18249 ( .A(n26516), .Y(n26951) );
  sky130_fd_sc_hd__nand2b_2 U18250 ( .A_N(n23856), .B(n12366), .Y(n26898) );
  sky130_fd_sc_hd__clkinv_1 U18251 ( .A(n22929), .Y(n22978) );
  sky130_fd_sc_hd__clkinv_1 U18252 ( .A(n22654), .Y(n22980) );
  sky130_fd_sc_hd__nand2_2 U18253 ( .A(n19535), .B(n19534), .Y(n26847) );
  sky130_fd_sc_hd__o21a_1 U18254 ( .A1(n22456), .A2(n24166), .B1(n21966), .X(
        n22580) );
  sky130_fd_sc_hd__a21oi_1 U18255 ( .A1(n26804), .A2(n22768), .B1(n21965), .Y(
        n21966) );
  sky130_fd_sc_hd__inv_2 U18256 ( .A(n24593), .Y(n26891) );
  sky130_fd_sc_hd__and2_0 U18257 ( .A(n24920), .B(n24919), .X(n24930) );
  sky130_fd_sc_hd__clkinv_1 U18258 ( .A(n26300), .Y(n28622) );
  sky130_fd_sc_hd__nor2_1 U18259 ( .A(n28947), .B(n28948), .Y(n24565) );
  sky130_fd_sc_hd__nor4_1 U18260 ( .A(n23907), .B(n23546), .C(n28642), .D(
        n28640), .Y(n28647) );
  sky130_fd_sc_hd__clkinv_1 U18261 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[0]), .Y(n20984) );
  sky130_fd_sc_hd__clkinv_1 U18262 ( .A(n28108), .Y(n28259) );
  sky130_fd_sc_hd__clkinv_1 U18263 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .Y(n28727) );
  sky130_fd_sc_hd__clkinv_1 U18264 ( .A(n23784), .Y(n26895) );
  sky130_fd_sc_hd__nor2_1 U18265 ( .A(n23706), .B(n23705), .Y(n24593) );
  sky130_fd_sc_hd__nand2_1 U18266 ( .A(n23485), .B(n29594), .Y(n26897) );
  sky130_fd_sc_hd__clkinv_1 U18267 ( .A(n24534), .Y(n24546) );
  sky130_fd_sc_hd__nor2_1 U18269 ( .A(n12328), .B(n23569), .Y(n12327) );
  sky130_fd_sc_hd__clkinv_1 U18270 ( .A(n13240), .Y(n13238) );
  sky130_fd_sc_hd__and2_0 U18271 ( .A(j202_soc_core_j22_cpu_memop_MEM__2_), 
        .B(j202_soc_core_j22_cpu_memop_MEM__0_), .X(n23300) );
  sky130_fd_sc_hd__and2_1 U18272 ( .A(n18899), .B(n23300), .X(n22929) );
  sky130_fd_sc_hd__o21a_1 U18274 ( .A1(n13599), .A2(n27914), .B1(n13598), .X(
        n27919) );
  sky130_fd_sc_hd__clkinv_1 U18275 ( .A(n27919), .Y(n27176) );
  sky130_fd_sc_hd__and2_0 U18276 ( .A(n13367), .B(n13366), .X(n13368) );
  sky130_fd_sc_hd__and2_0 U18277 ( .A(n13365), .B(n13364), .X(n13369) );
  sky130_fd_sc_hd__clkinv_1 U18279 ( .A(gpio_en_o[1]), .Y(io_oeb[1]) );
  sky130_fd_sc_hd__clkinv_1 U18280 ( .A(gpio_en_o[2]), .Y(io_oeb[2]) );
  sky130_fd_sc_hd__clkinv_1 U18281 ( .A(gpio_en_o[3]), .Y(io_oeb[3]) );
  sky130_fd_sc_hd__clkinv_1 U18282 ( .A(gpio_en_o[5]), .Y(io_oeb[7]) );
  sky130_fd_sc_hd__clkinv_1 U18283 ( .A(gpio_en_o[6]), .Y(io_oeb[26]) );
  sky130_fd_sc_hd__clkinv_1 U18284 ( .A(gpio_en_o[7]), .Y(io_oeb[27]) );
  sky130_fd_sc_hd__clkinv_1 U18285 ( .A(gpio_en_o[9]), .Y(io_oeb[29]) );
  sky130_fd_sc_hd__clkinv_1 U18286 ( .A(gpio_en_o[10]), .Y(io_oeb[30]) );
  sky130_fd_sc_hd__clkinv_1 U18287 ( .A(gpio_en_o[11]), .Y(io_oeb[31]) );
  sky130_fd_sc_hd__clkinv_1 U18288 ( .A(gpio_en_o[13]), .Y(io_oeb[33]) );
  sky130_fd_sc_hd__clkinv_1 U18289 ( .A(gpio_en_o[14]), .Y(io_oeb[34]) );
  sky130_fd_sc_hd__clkinv_1 U18290 ( .A(gpio_en_o[15]), .Y(io_oeb[35]) );
  sky130_fd_sc_hd__nand2b_1 U18291 ( .A_N(n18353), .B(n18656), .Y(n18058) );
  sky130_fd_sc_hd__clkinv_1 U18292 ( .A(n18309), .Y(n12304) );
  sky130_fd_sc_hd__o22ai_1 U18293 ( .A1(n18750), .A2(n18304), .B1(n18320), 
        .B2(n18747), .Y(n18348) );
  sky130_fd_sc_hd__clkinv_1 U18294 ( .A(n18353), .Y(n12302) );
  sky130_fd_sc_hd__nand2b_1 U18295 ( .A_N(n18353), .B(n22112), .Y(n17512) );
  sky130_fd_sc_hd__and2_0 U18296 ( .A(n15614), .B(n15558), .X(n13419) );
  sky130_fd_sc_hd__o22ai_1 U18297 ( .A1(n18344), .A2(n18343), .B1(n18294), 
        .B2(n17402), .Y(n12305) );
  sky130_fd_sc_hd__clkinv_1 U18298 ( .A(n18253), .Y(n12721) );
  sky130_fd_sc_hd__clkinv_1 U18299 ( .A(n18254), .Y(n12720) );
  sky130_fd_sc_hd__xor2_1 U18300 ( .A(n12138), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n17506) );
  sky130_fd_sc_hd__o22ai_1 U18301 ( .A1(n18660), .A2(n18658), .B1(n18516), 
        .B2(n12991), .Y(n18671) );
  sky130_fd_sc_hd__clkinv_1 U18302 ( .A(n17604), .Y(n12749) );
  sky130_fd_sc_hd__clkinv_1 U18303 ( .A(j202_soc_core_j22_cpu_ml_bufa[11]), 
        .Y(n17688) );
  sky130_fd_sc_hd__clkinv_1 U18304 ( .A(n18576), .Y(n12611) );
  sky130_fd_sc_hd__o22ai_1 U18305 ( .A1(n18750), .A2(n18447), .B1(n18428), 
        .B2(n18747), .Y(n18450) );
  sky130_fd_sc_hd__fa_1 U18306 ( .A(n18533), .B(n18532), .CIN(n18531), .COUT(
        n18734), .SUM(n18542) );
  sky130_fd_sc_hd__o22ai_1 U18307 ( .A1(n18660), .A2(n18516), .B1(n18485), 
        .B2(n12991), .Y(n18522) );
  sky130_fd_sc_hd__clkinv_1 U18308 ( .A(n18804), .Y(n12634) );
  sky130_fd_sc_hd__or2_0 U18309 ( .A(n17985), .B(n17984), .X(n18016) );
  sky130_fd_sc_hd__clkinv_1 U18310 ( .A(n26757), .Y(n21932) );
  sky130_fd_sc_hd__and2_0 U18311 ( .A(n15227), .B(n15593), .X(n12192) );
  sky130_fd_sc_hd__and2_0 U18312 ( .A(n18927), .B(n21186), .X(n21082) );
  sky130_fd_sc_hd__clkinv_1 U18313 ( .A(n15580), .Y(n15227) );
  sky130_fd_sc_hd__clkinv_1 U18314 ( .A(n18266), .Y(n12445) );
  sky130_fd_sc_hd__clkinv_1 U18315 ( .A(n18563), .Y(n12950) );
  sky130_fd_sc_hd__clkinv_1 U18316 ( .A(n18154), .Y(n12565) );
  sky130_fd_sc_hd__nor2_1 U18317 ( .A(n12141), .B(n18650), .Y(n18699) );
  sky130_fd_sc_hd__and2_0 U18318 ( .A(n22129), .B(n22357), .X(n22101) );
  sky130_fd_sc_hd__clkinv_1 U18319 ( .A(n18074), .Y(n12994) );
  sky130_fd_sc_hd__clkinv_1 U18320 ( .A(n18011), .Y(n12684) );
  sky130_fd_sc_hd__nor2b_1 U18321 ( .B_N(n18353), .A(n18344), .Y(n17626) );
  sky130_fd_sc_hd__clkinv_1 U18322 ( .A(j202_soc_core_j22_cpu_ml_bufa[9]), .Y(
        n12569) );
  sky130_fd_sc_hd__buf_2 U18323 ( .A(j202_soc_core_j22_cpu_ml_bufb[5]), .X(
        n18511) );
  sky130_fd_sc_hd__clkinv_1 U18324 ( .A(n18476), .Y(n12925) );
  sky130_fd_sc_hd__clkinv_1 U18325 ( .A(n17523), .Y(n12572) );
  sky130_fd_sc_hd__clkinv_1 U18326 ( .A(n15593), .Y(n13478) );
  sky130_fd_sc_hd__and2_0 U18328 ( .A(n21078), .B(n20772), .X(n21607) );
  sky130_fd_sc_hd__and2_0 U18329 ( .A(n21648), .B(n21094), .X(n21172) );
  sky130_fd_sc_hd__and2_0 U18330 ( .A(n20532), .B(n20648), .X(n15682) );
  sky130_fd_sc_hd__nand2_1 U18331 ( .A(n17293), .B(
        j202_soc_core_bootrom_00_address_w[11]), .Y(n16845) );
  sky130_fd_sc_hd__clkinv_1 U18332 ( .A(n16773), .Y(n16579) );
  sky130_fd_sc_hd__and2_0 U18333 ( .A(n21253), .B(n20772), .X(n21229) );
  sky130_fd_sc_hd__nand4bb_1 U18334 ( .A_N(n16111), .B_N(n15803), .C(n15802), 
        .D(n15801), .Y(n15804) );
  sky130_fd_sc_hd__inv_2 U18335 ( .A(n21053), .Y(n21608) );
  sky130_fd_sc_hd__nor4_1 U18336 ( .A(n20079), .B(n20082), .C(n20348), .D(
        n20078), .Y(n20086) );
  sky130_fd_sc_hd__and2_0 U18339 ( .A(n16689), .B(n16880), .X(n16965) );
  sky130_fd_sc_hd__and2_0 U18340 ( .A(n20054), .B(n20885), .X(n20352) );
  sky130_fd_sc_hd__clkinv_1 U18341 ( .A(n15708), .Y(n17163) );
  sky130_fd_sc_hd__o2bb2ai_1 U18342 ( .B1(n15708), .B2(n15368), .A1_N(n15584), 
        .A2_N(n15259), .Y(n15260) );
  sky130_fd_sc_hd__nor2_1 U18343 ( .A(n11153), .B(n21915), .Y(n12981) );
  sky130_fd_sc_hd__clkinv_1 U18344 ( .A(n17747), .Y(n12653) );
  sky130_fd_sc_hd__clkinv_1 U18345 ( .A(n17702), .Y(n12607) );
  sky130_fd_sc_hd__and2_0 U18346 ( .A(n24785), .B(n24774), .X(n25308) );
  sky130_fd_sc_hd__a21oi_1 U18347 ( .A1(n18288), .A2(n21875), .B1(n18287), .Y(
        n18289) );
  sky130_fd_sc_hd__inv_2 U18348 ( .A(n21253), .Y(n19351) );
  sky130_fd_sc_hd__a31o_1 U18349 ( .A1(n15611), .A2(n15610), .A3(n15609), .B1(
        n15708), .X(n15634) );
  sky130_fd_sc_hd__and2_0 U18350 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_duty[9]), .X(n15647) );
  sky130_fd_sc_hd__and2_0 U18351 ( .A(n15359), .B(n15558), .X(n15551) );
  sky130_fd_sc_hd__a21boi_0 U18352 ( .A1(n13304), .A2(n21064), .B1_N(n21063), 
        .Y(n21153) );
  sky130_fd_sc_hd__clkinv_1 U18353 ( .A(n21648), .Y(n21054) );
  sky130_fd_sc_hd__clkinv_1 U18354 ( .A(n21201), .Y(n19279) );
  sky130_fd_sc_hd__inv_2 U18355 ( .A(n20659), .Y(n20439) );
  sky130_fd_sc_hd__clkinv_1 U18356 ( .A(n20849), .Y(n20172) );
  sky130_fd_sc_hd__inv_2 U18357 ( .A(n20919), .Y(n20180) );
  sky130_fd_sc_hd__a31o_1 U18358 ( .A1(n20051), .A2(n20050), .A3(n20075), .B1(
        n20906), .X(n20071) );
  sky130_fd_sc_hd__clkinv_1 U18359 ( .A(n17166), .Y(n17193) );
  sky130_fd_sc_hd__inv_2 U18360 ( .A(n20047), .Y(n20871) );
  sky130_fd_sc_hd__inv_2 U18361 ( .A(n21697), .Y(n21124) );
  sky130_fd_sc_hd__inv_2 U18362 ( .A(n21244), .Y(n21178) );
  sky130_fd_sc_hd__and2_0 U18363 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[1]), 
        .B(j202_soc_core_uart_TOP_rx_fifo_rp[0]), .X(n21668) );
  sky130_fd_sc_hd__nor2_1 U18364 ( .A(n13383), .B(n17184), .Y(n21666) );
  sky130_fd_sc_hd__nor2_1 U18365 ( .A(n17182), .B(n17184), .Y(n21699) );
  sky130_fd_sc_hd__inv_2 U18366 ( .A(n20384), .Y(n19834) );
  sky130_fd_sc_hd__inv_2 U18367 ( .A(n20074), .Y(n20918) );
  sky130_fd_sc_hd__a21oi_1 U18368 ( .A1(n18856), .A2(n22944), .B1(n18855), .Y(
        n18857) );
  sky130_fd_sc_hd__and2_0 U18369 ( .A(n15274), .B(n15294), .X(n12285) );
  sky130_fd_sc_hd__nor2_1 U18370 ( .A(n12700), .B(n24770), .Y(n12699) );
  sky130_fd_sc_hd__clkinv_1 U18371 ( .A(n24797), .Y(n12694) );
  sky130_fd_sc_hd__clkinv_1 U18373 ( .A(j202_soc_core_j22_cpu_rf_vbr[29]), .Y(
        n22441) );
  sky130_fd_sc_hd__clkinv_1 U18374 ( .A(j202_soc_core_j22_cpu_rf_gpr[509]), 
        .Y(n22442) );
  sky130_fd_sc_hd__and2_0 U18375 ( .A(n12927), .B(n22658), .X(n12280) );
  sky130_fd_sc_hd__clkinv_1 U18376 ( .A(n22659), .Y(n12928) );
  sky130_fd_sc_hd__clkinv_1 U18377 ( .A(n18901), .Y(n18831) );
  sky130_fd_sc_hd__nor2_1 U18378 ( .A(n12207), .B(n18832), .Y(n22908) );
  sky130_fd_sc_hd__clkinv_1 U18380 ( .A(n19164), .Y(n12399) );
  sky130_fd_sc_hd__a21boi_0 U18381 ( .A1(n26077), .A2(n26724), .B1_N(n24715), 
        .Y(n24716) );
  sky130_fd_sc_hd__nand2_1 U18382 ( .A(n24265), .B(n23603), .Y(n23606) );
  sky130_fd_sc_hd__nand3_1 U18383 ( .A(n18988), .B(n18987), .C(n26780), .Y(
        n23922) );
  sky130_fd_sc_hd__inv_1 U18384 ( .A(n26526), .Y(n19164) );
  sky130_fd_sc_hd__clkinv_1 U18385 ( .A(n21790), .Y(n12368) );
  sky130_fd_sc_hd__and2_0 U18386 ( .A(n21677), .B(n21773), .X(n12206) );
  sky130_fd_sc_hd__and2_0 U18387 ( .A(n21632), .B(n21706), .X(n21079) );
  sky130_fd_sc_hd__clkinv_1 U18388 ( .A(n21709), .Y(n21636) );
  sky130_fd_sc_hd__nor2_1 U18389 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .B(n14965), .Y(n20626) );
  sky130_fd_sc_hd__and2_0 U18390 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_duty[5]), .X(n20703) );
  sky130_fd_sc_hd__clkinv_1 U18391 ( .A(n14724), .Y(n13986) );
  sky130_fd_sc_hd__clkinv_1 U18392 ( .A(n26755), .Y(n26758) );
  sky130_fd_sc_hd__clkinv_1 U18393 ( .A(n27368), .Y(n26568) );
  sky130_fd_sc_hd__clkinv_1 U18394 ( .A(n26539), .Y(n26548) );
  sky130_fd_sc_hd__and2_0 U18395 ( .A(n21317), .B(n21750), .X(n12231) );
  sky130_fd_sc_hd__nand2_1 U18396 ( .A(n12628), .B(n11049), .Y(n12421) );
  sky130_fd_sc_hd__clkinv_1 U18397 ( .A(n24607), .Y(n24755) );
  sky130_fd_sc_hd__and2_0 U18398 ( .A(n28888), .B(
        j202_soc_core_intc_core_00_bs_addr[8]), .X(n24749) );
  sky130_fd_sc_hd__clkinv_1 U18399 ( .A(j202_soc_core_intc_core_00_bs_addr[6]), 
        .Y(n28884) );
  sky130_fd_sc_hd__clkinv_1 U18400 ( .A(n15496), .Y(n13153) );
  sky130_fd_sc_hd__clkinv_1 U18401 ( .A(n16134), .Y(n12855) );
  sky130_fd_sc_hd__a21boi_0 U18403 ( .A1(n17315), .A2(n20801), .B1_N(n17303), 
        .Y(n19398) );
  sky130_fd_sc_hd__clkinv_1 U18404 ( .A(
        j202_soc_core_memory0_ram_dout0_sel[12]), .Y(n13505) );
  sky130_fd_sc_hd__clkinv_1 U18405 ( .A(n20864), .Y(n20927) );
  sky130_fd_sc_hd__and2_0 U18406 ( .A(n26529), .B(n26539), .X(n23769) );
  sky130_fd_sc_hd__o21ai_1 U18407 ( .A1(n23144), .A2(n12012), .B1(n27259), .Y(
        n23604) );
  sky130_fd_sc_hd__clkbuf_1 U18408 ( .A(n23213), .X(n23954) );
  sky130_fd_sc_hd__and2_0 U18409 ( .A(n27912), .B(n27909), .X(n13654) );
  sky130_fd_sc_hd__clkinv_1 U18410 ( .A(n24658), .Y(n24093) );
  sky130_fd_sc_hd__inv_2 U18411 ( .A(n27789), .Y(n24386) );
  sky130_fd_sc_hd__clkinv_1 U18412 ( .A(j202_soc_core_gpio_core_00_reg_addr[1]), .Y(n27629) );
  sky130_fd_sc_hd__clkinv_1 U18413 ( .A(j202_soc_core_pwrite[1]), .Y(n28882)
         );
  sky130_fd_sc_hd__clkinv_1 U18414 ( .A(j202_soc_core_intc_core_00_bs_addr[3]), 
        .Y(n28886) );
  sky130_fd_sc_hd__and2_0 U18415 ( .A(n25916), .B(n28058), .X(n26189) );
  sky130_fd_sc_hd__a21oi_1 U18416 ( .A1(n22944), .A2(n21493), .B1(n21492), .Y(
        n21494) );
  sky130_fd_sc_hd__nand2b_1 U18419 ( .A_N(n12399), .B(n26539), .Y(n24781) );
  sky130_fd_sc_hd__inv_2 U18420 ( .A(n17706), .Y(n21505) );
  sky130_fd_sc_hd__a21boi_0 U18421 ( .A1(n26077), .A2(n26728), .B1_N(n25028), 
        .Y(n25029) );
  sky130_fd_sc_hd__nand3_1 U18422 ( .A(n23014), .B(n26443), .C(n25130), .Y(
        n23034) );
  sky130_fd_sc_hd__and2_0 U18423 ( .A(n22769), .B(n22770), .X(n13318) );
  sky130_fd_sc_hd__clkinv_1 U18424 ( .A(n17816), .Y(n12791) );
  sky130_fd_sc_hd__and2_0 U18425 ( .A(n24954), .B(n24957), .X(n27732) );
  sky130_fd_sc_hd__nor2_1 U18426 ( .A(n18893), .B(n26863), .Y(n22028) );
  sky130_fd_sc_hd__inv_2 U18427 ( .A(j202_soc_core_j22_cpu_regop_We__2_), .Y(
        n23279) );
  sky130_fd_sc_hd__nand3_2 U18428 ( .A(n14034), .B(n14033), .C(n14032), .Y(
        n26723) );
  sky130_fd_sc_hd__nor2_2 U18429 ( .A(n13659), .B(n13682), .Y(n13794) );
  sky130_fd_sc_hd__inv_2 U18430 ( .A(n29568), .Y(n23089) );
  sky130_fd_sc_hd__and2_0 U18431 ( .A(n26863), .B(n26398), .X(n22627) );
  sky130_fd_sc_hd__nand2b_1 U18432 ( .A_N(n23693), .B(n22712), .Y(n21523) );
  sky130_fd_sc_hd__nand3_1 U18433 ( .A(n19197), .B(n29535), .C(n13338), .Y(
        n12325) );
  sky130_fd_sc_hd__nor2_1 U18434 ( .A(n13103), .B(n12378), .Y(n12733) );
  sky130_fd_sc_hd__nor2_1 U18435 ( .A(n23144), .B(n24705), .Y(n23821) );
  sky130_fd_sc_hd__and2_0 U18436 ( .A(n27914), .B(n27913), .X(n27917) );
  sky130_fd_sc_hd__clkinv_1 U18437 ( .A(n24049), .Y(n12929) );
  sky130_fd_sc_hd__and2_0 U18438 ( .A(n25056), .B(n26329), .X(n25074) );
  sky130_fd_sc_hd__and2_0 U18439 ( .A(n24896), .B(n24950), .X(n24946) );
  sky130_fd_sc_hd__clkinv_1 U18440 ( .A(j202_soc_core_j22_cpu_rf_pr[13]), .Y(
        n21845) );
  sky130_fd_sc_hd__and2_0 U18441 ( .A(n21780), .B(n21779), .X(n13343) );
  sky130_fd_sc_hd__nor2_1 U18442 ( .A(n17300), .B(n20804), .Y(n21207) );
  sky130_fd_sc_hd__nand2_1 U18443 ( .A(n17293), .B(n20687), .Y(n21705) );
  sky130_fd_sc_hd__nand2_1 U18444 ( .A(n20626), .B(
        j202_soc_core_bootrom_00_address_w[9]), .Y(n19856) );
  sky130_fd_sc_hd__clkinv_1 U18445 ( .A(n13004), .Y(n19327) );
  sky130_fd_sc_hd__clkinv_1 U18446 ( .A(n23172), .Y(n23520) );
  sky130_fd_sc_hd__clkinv_1 U18447 ( .A(n20989), .Y(n22321) );
  sky130_fd_sc_hd__and2_0 U18448 ( .A(n24910), .B(n24909), .X(n24917) );
  sky130_fd_sc_hd__and2_0 U18449 ( .A(n24908), .B(n24907), .X(n24918) );
  sky130_fd_sc_hd__and2_0 U18450 ( .A(n24914), .B(n24913), .X(n24915) );
  sky130_fd_sc_hd__and2_0 U18451 ( .A(n24926), .B(n24925), .X(n24927) );
  sky130_fd_sc_hd__and2_0 U18452 ( .A(n24922), .B(n24921), .X(n24929) );
  sky130_fd_sc_hd__and2_0 U18453 ( .A(n24924), .B(n24923), .X(n24928) );
  sky130_fd_sc_hd__clkinv_1 U18454 ( .A(n23669), .Y(n24896) );
  sky130_fd_sc_hd__nor2_1 U18455 ( .A(n21427), .B(n13146), .Y(n13144) );
  sky130_fd_sc_hd__clkinv_1 U18456 ( .A(n26805), .Y(n26801) );
  sky130_fd_sc_hd__clkinv_1 U18457 ( .A(n26780), .Y(n26693) );
  sky130_fd_sc_hd__a22oi_1 U18458 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__14_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__14_), .Y(n21166) );
  sky130_fd_sc_hd__clkinv_1 U18459 ( .A(j202_soc_core_ahb2apb_01_state[0]), 
        .Y(n24005) );
  sky130_fd_sc_hd__clkinv_1 U18460 ( .A(j202_soc_core_ahb2apb_01_state[2]), 
        .Y(n24319) );
  sky130_fd_sc_hd__clkinv_1 U18461 ( .A(j202_soc_core_wbqspiflash_00_state[2]), 
        .Y(n23467) );
  sky130_fd_sc_hd__clkinv_1 U18462 ( .A(n26029), .Y(n26030) );
  sky130_fd_sc_hd__clkinv_1 U18463 ( .A(n25953), .Y(n26035) );
  sky130_fd_sc_hd__inv_2 U18464 ( .A(n26728), .Y(n26571) );
  sky130_fd_sc_hd__nor2_1 U18466 ( .A(n13380), .B(n13496), .Y(n21604) );
  sky130_fd_sc_hd__buf_2 U18467 ( .A(n24417), .X(n12729) );
  sky130_fd_sc_hd__nand2_1 U18468 ( .A(j202_soc_core_memory0_ram_dout0[459]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n13178) );
  sky130_fd_sc_hd__nand2_1 U18469 ( .A(n12830), .B(n12819), .Y(n12878) );
  sky130_fd_sc_hd__nor2_2 U18470 ( .A(n13493), .B(n13496), .Y(n21591) );
  sky130_fd_sc_hd__nor2_1 U18471 ( .A(n13500), .B(n13499), .Y(n21593) );
  sky130_fd_sc_hd__nor2_1 U18472 ( .A(n13502), .B(n13501), .Y(n21596) );
  sky130_fd_sc_hd__nor2_1 U18473 ( .A(n13505), .B(n13504), .Y(n21597) );
  sky130_fd_sc_hd__clkinv_1 U18474 ( .A(
        j202_soc_core_memory0_ram_dout0_sel[13]), .Y(n13498) );
  sky130_fd_sc_hd__nor2_1 U18475 ( .A(n13488), .B(n13499), .Y(n21605) );
  sky130_fd_sc_hd__nor2_1 U18476 ( .A(n13376), .B(n13496), .Y(n21733) );
  sky130_fd_sc_hd__nor2_2 U18478 ( .A(n13378), .B(n13496), .Y(n21732) );
  sky130_fd_sc_hd__and2_0 U18479 ( .A(j202_soc_core_intc_core_00_in_intreq[20]), .B(j202_soc_core_intc_core_00_rg_itgt[20]), .X(n19562) );
  sky130_fd_sc_hd__o22ai_1 U18480 ( .A1(n19664), .A2(n19651), .B1(n13027), 
        .B2(n13024), .Y(n19658) );
  sky130_fd_sc_hd__clkinv_1 U18481 ( .A(n26839), .Y(n26841) );
  sky130_fd_sc_hd__buf_2 U18482 ( .A(n13700), .X(n16513) );
  sky130_fd_sc_hd__clkinv_1 U18483 ( .A(n26863), .Y(n26318) );
  sky130_fd_sc_hd__nand2_1 U18484 ( .A(n23237), .B(n26863), .Y(n22311) );
  sky130_fd_sc_hd__clkinv_1 U18485 ( .A(n14846), .Y(n23706) );
  sky130_fd_sc_hd__clkinv_1 U18486 ( .A(j202_soc_core_j22_cpu_regop_Rs__1_), 
        .Y(n22873) );
  sky130_fd_sc_hd__clkinv_1 U18487 ( .A(n22034), .Y(n22866) );
  sky130_fd_sc_hd__clkinv_1 U18488 ( .A(n24159), .Y(n18894) );
  sky130_fd_sc_hd__nand2_1 U18489 ( .A(n12560), .B(n27980), .Y(n22289) );
  sky130_fd_sc_hd__and2_1 U18490 ( .A(n20428), .B(
        j202_soc_core_j22_cpu_id_opn_v_), .X(n21775) );
  sky130_fd_sc_hd__and2_0 U18491 ( .A(n20711), .B(n21750), .X(n12232) );
  sky130_fd_sc_hd__inv_2 U18493 ( .A(n27889), .Y(n27958) );
  sky130_fd_sc_hd__clkinv_1 U18495 ( .A(j202_soc_core_intc_core_00_bs_addr[0]), 
        .Y(n27074) );
  sky130_fd_sc_hd__clkinv_1 U18496 ( .A(j202_soc_core_intc_core_00_bs_addr[1]), 
        .Y(n27070) );
  sky130_fd_sc_hd__inv_2 U18497 ( .A(j202_soc_core_intc_core_00_rg_ipr[41]), 
        .Y(n24027) );
  sky130_fd_sc_hd__clkinv_1 U18498 ( .A(j202_soc_core_intc_core_00_rg_ipr[22]), 
        .Y(n26499) );
  sky130_fd_sc_hd__and2_0 U18499 ( .A(n28743), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[2]), .X(n29118) );
  sky130_fd_sc_hd__clkinv_1 U18500 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[11]), .Y(n28347) );
  sky130_fd_sc_hd__clkinv_1 U18501 ( .A(
        j202_soc_core_intc_core_00_in_intreq[11]), .Y(n27011) );
  sky130_fd_sc_hd__clkinv_1 U18502 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[14]), .Y(n28368) );
  sky130_fd_sc_hd__clkinv_1 U18503 ( .A(
        j202_soc_core_intc_core_00_in_intreq[14]), .Y(n25496) );
  sky130_fd_sc_hd__and2_0 U18504 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[0]), 
        .B(j202_soc_core_uart_TOP_tx_fifo_rp[1]), .X(n28777) );
  sky130_fd_sc_hd__clkinv_1 U18505 ( .A(
        j202_soc_core_intc_core_00_in_intreq[13]), .Y(n25512) );
  sky130_fd_sc_hd__clkinv_1 U18506 ( .A(
        j202_soc_core_intc_core_00_in_intreq[8]), .Y(n25473) );
  sky130_fd_sc_hd__clkinv_1 U18507 ( .A(n28222), .Y(n28223) );
  sky130_fd_sc_hd__clkinv_1 U18508 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[19]), .Y(n28404) );
  sky130_fd_sc_hd__clkinv_1 U18509 ( .A(
        j202_soc_core_intc_core_00_in_intreq[9]), .Y(n25467) );
  sky130_fd_sc_hd__and2_0 U18510 ( .A(n24849), .B(n24848), .X(n24859) );
  sky130_fd_sc_hd__and2_0 U18511 ( .A(n24851), .B(n24850), .X(n24858) );
  sky130_fd_sc_hd__and2_0 U18512 ( .A(n24855), .B(n24854), .X(n24856) );
  sky130_fd_sc_hd__and2_0 U18513 ( .A(n24861), .B(n24860), .X(n24871) );
  sky130_fd_sc_hd__and2_0 U18514 ( .A(n24867), .B(n24866), .X(n24868) );
  sky130_fd_sc_hd__and2_0 U18515 ( .A(n24863), .B(n24862), .X(n24870) );
  sky130_fd_sc_hd__clkinv_1 U18516 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[25]), .Y(n28451) );
  sky130_fd_sc_hd__clkinv_1 U18517 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[1]), .Y(n27642) );
  sky130_fd_sc_hd__clkinv_1 U18518 ( .A(j202_soc_core_intc_core_00_rg_ipr[1]), 
        .Y(n27677) );
  sky130_fd_sc_hd__clkinv_1 U18519 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[1]), .Y(n27611) );
  sky130_fd_sc_hd__clkinv_1 U18520 ( .A(n27312), .Y(n27852) );
  sky130_fd_sc_hd__nor2_1 U18521 ( .A(n28590), .B(n27306), .Y(n27869) );
  sky130_fd_sc_hd__inv_2 U18522 ( .A(j202_soc_core_intc_core_00_rg_ipr[61]), 
        .Y(n26952) );
  sky130_fd_sc_hd__inv_2 U18523 ( .A(j202_soc_core_intc_core_00_rg_ipr[48]), 
        .Y(n25519) );
  sky130_fd_sc_hd__inv_2 U18524 ( .A(j202_soc_core_intc_core_00_rg_ipr[46]), 
        .Y(n25450) );
  sky130_fd_sc_hd__inv_2 U18525 ( .A(j202_soc_core_intc_core_00_rg_ipr[45]), 
        .Y(n25460) );
  sky130_fd_sc_hd__inv_2 U18527 ( .A(j202_soc_core_intc_core_00_rg_ipr[42]), 
        .Y(n25449) );
  sky130_fd_sc_hd__inv_2 U18528 ( .A(j202_soc_core_intc_core_00_rg_ipr[39]), 
        .Y(n25485) );
  sky130_fd_sc_hd__inv_2 U18529 ( .A(j202_soc_core_intc_core_00_rg_ipr[38]), 
        .Y(n25464) );
  sky130_fd_sc_hd__inv_2 U18530 ( .A(j202_soc_core_intc_core_00_rg_ipr[36]), 
        .Y(n25483) );
  sky130_fd_sc_hd__clkinv_1 U18531 ( .A(n25481), .Y(n27019) );
  sky130_fd_sc_hd__clkinv_1 U18532 ( .A(n25482), .Y(n27021) );
  sky130_fd_sc_hd__clkinv_1 U18533 ( .A(n28520), .Y(n28541) );
  sky130_fd_sc_hd__inv_2 U18534 ( .A(j202_soc_core_intc_core_00_rg_ipr[77]), 
        .Y(n27805) );
  sky130_fd_sc_hd__inv_2 U18535 ( .A(j202_soc_core_intc_core_00_rg_ipr[76]), 
        .Y(n26263) );
  sky130_fd_sc_hd__clkinv_1 U18537 ( .A(n27752), .Y(n27990) );
  sky130_fd_sc_hd__clkinv_1 U18538 ( .A(j202_soc_core_intc_core_00_rg_ipr[15]), 
        .Y(n25277) );
  sky130_fd_sc_hd__clkinv_1 U18539 ( .A(
        j202_soc_core_intc_core_00_in_intreq[15]), .Y(n25487) );
  sky130_fd_sc_hd__clkinv_1 U18540 ( .A(
        j202_soc_core_intc_core_00_in_intreq[10]), .Y(n25453) );
  sky130_fd_sc_hd__clkinv_1 U18541 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[27]), .Y(n28467) );
  sky130_fd_sc_hd__and2_0 U18542 ( .A(n28904), .B(n28903), .X(n28914) );
  sky130_fd_sc_hd__clkinv_1 U18543 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[2]), .Y(n28284) );
  sky130_fd_sc_hd__clkinv_1 U18544 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[5]), .Y(n28305) );
  sky130_fd_sc_hd__clkinv_1 U18545 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[6]), .Y(n28312) );
  sky130_fd_sc_hd__clkinv_1 U18546 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[7]), .Y(n28319) );
  sky130_fd_sc_hd__clkinv_1 U18547 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[12]), .Y(n28354) );
  sky130_fd_sc_hd__clkinv_1 U18548 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[18]), .Y(n28396) );
  sky130_fd_sc_hd__clkinv_1 U18549 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[22]), .Y(n28429) );
  sky130_fd_sc_hd__clkinv_1 U18550 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[23]), .Y(n28438) );
  sky130_fd_sc_hd__clkinv_1 U18551 ( .A(gpio_en_o[24]), .Y(n28445) );
  sky130_fd_sc_hd__clkinv_1 U18552 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[26]), .Y(n28459) );
  sky130_fd_sc_hd__clkinv_1 U18553 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[28]), .Y(n28479) );
  sky130_fd_sc_hd__clkinv_1 U18554 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[29]), .Y(n28485) );
  sky130_fd_sc_hd__clkinv_1 U18555 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[30]), .Y(n28493) );
  sky130_fd_sc_hd__clkinv_1 U18556 ( .A(n28476), .Y(n28506) );
  sky130_fd_sc_hd__clkinv_1 U18557 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[15]), .Y(n28375) );
  sky130_fd_sc_hd__clkinv_1 U18558 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[10]), .Y(n28340) );
  sky130_fd_sc_hd__and2_0 U18559 ( .A(n22039), .B(n22873), .X(n22969) );
  sky130_fd_sc_hd__clkinv_1 U18560 ( .A(n22611), .Y(n12499) );
  sky130_fd_sc_hd__clkinv_1 U18561 ( .A(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_), .Y(n25680) );
  sky130_fd_sc_hd__and2_0 U18562 ( .A(j202_soc_core_aquc_STB_), .B(
        j202_soc_core_aquc_CE__0_), .X(n23909) );
  sky130_fd_sc_hd__clkinv_1 U18563 ( .A(
        j202_soc_core_wbqspiflash_00_write_in_progress), .Y(n26171) );
  sky130_fd_sc_hd__clkinv_1 U18564 ( .A(n26859), .Y(n27341) );
  sky130_fd_sc_hd__clkinv_1 U18565 ( .A(n25215), .Y(n27184) );
  sky130_fd_sc_hd__clkinv_1 U18566 ( .A(n26861), .Y(n27339) );
  sky130_fd_sc_hd__inv_2 U18567 ( .A(n12645), .Y(n27276) );
  sky130_fd_sc_hd__clkinv_1 U18569 ( .A(n12647), .Y(n27394) );
  sky130_fd_sc_hd__nand2_1 U18570 ( .A(n29517), .B(n26539), .Y(n12619) );
  sky130_fd_sc_hd__clkinv_1 U18571 ( .A(n25332), .Y(n25326) );
  sky130_fd_sc_hd__inv_2 U18572 ( .A(n27371), .Y(n26395) );
  sky130_fd_sc_hd__inv_2 U18573 ( .A(n11766), .Y(n27464) );
  sky130_fd_sc_hd__clkinv_1 U18574 ( .A(n25259), .Y(n27434) );
  sky130_fd_sc_hd__clkinv_1 U18575 ( .A(n27418), .Y(n27452) );
  sky130_fd_sc_hd__clkinv_1 U18576 ( .A(n27456), .Y(n24112) );
  sky130_fd_sc_hd__nand2_1 U18577 ( .A(n13580), .B(n13579), .Y(n27450) );
  sky130_fd_sc_hd__clkinv_1 U18578 ( .A(n27438), .Y(n27446) );
  sky130_fd_sc_hd__nand2_1 U18579 ( .A(n26861), .B(n24023), .Y(n27343) );
  sky130_fd_sc_hd__or2_0 U18580 ( .A(n18993), .B(n18992), .X(n18995) );
  sky130_fd_sc_hd__clkinv_1 U18581 ( .A(j202_soc_core_j22_cpu_macop_MAC_[1]), 
        .Y(n24288) );
  sky130_fd_sc_hd__clkinv_1 U18582 ( .A(n27442), .Y(n27335) );
  sky130_fd_sc_hd__nand2_1 U18583 ( .A(n26528), .B(n26539), .Y(n12593) );
  sky130_fd_sc_hd__nand3_1 U18584 ( .A(n12326), .B(n24449), .C(n24450), .Y(
        n24451) );
  sky130_fd_sc_hd__and2_0 U18585 ( .A(n27265), .B(n24364), .X(n27177) );
  sky130_fd_sc_hd__nand3_2 U18586 ( .A(n23177), .B(n23078), .C(n23077), .Y(
        n23079) );
  sky130_fd_sc_hd__clkinv_1 U18587 ( .A(n27467), .Y(n12455) );
  sky130_fd_sc_hd__nand3_2 U18588 ( .A(n19168), .B(n19166), .C(n19167), .Y(
        n12840) );
  sky130_fd_sc_hd__clkinv_1 U18589 ( .A(n26557), .Y(n27370) );
  sky130_fd_sc_hd__clkinv_1 U18590 ( .A(n12120), .Y(n27576) );
  sky130_fd_sc_hd__clkinv_1 U18591 ( .A(n26898), .Y(n26383) );
  sky130_fd_sc_hd__nor2_1 U18592 ( .A(n13082), .B(n11070), .Y(n13081) );
  sky130_fd_sc_hd__clkinv_1 U18593 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[4]), .Y(n26986) );
  sky130_fd_sc_hd__clkinv_1 U18594 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[5]), .Y(n26924) );
  sky130_fd_sc_hd__a21oi_1 U18595 ( .A1(n22513), .A2(n16993), .B1(n16992), .Y(
        n16998) );
  sky130_fd_sc_hd__clkinv_1 U18596 ( .A(n27343), .Y(n27006) );
  sky130_fd_sc_hd__clkinv_1 U18597 ( .A(n26946), .Y(n26450) );
  sky130_fd_sc_hd__clkinv_1 U18598 ( .A(n27340), .Y(n27349) );
  sky130_fd_sc_hd__nand2_1 U18599 ( .A(n24012), .B(j202_soc_core_pwrite[1]), 
        .Y(n25534) );
  sky130_fd_sc_hd__clkinv_1 U18600 ( .A(n24753), .Y(n24012) );
  sky130_fd_sc_hd__clkinv_1 U18602 ( .A(n27491), .Y(n27498) );
  sky130_fd_sc_hd__clkinv_1 U18603 ( .A(n12417), .Y(n27064) );
  sky130_fd_sc_hd__inv_2 U18604 ( .A(n24565), .Y(n22711) );
  sky130_fd_sc_hd__nor2_1 U18605 ( .A(n28590), .B(n24979), .Y(n27860) );
  sky130_fd_sc_hd__nor2_1 U18606 ( .A(n28590), .B(n24977), .Y(n27856) );
  sky130_fd_sc_hd__nor2_1 U18607 ( .A(n28590), .B(n24762), .Y(n27850) );
  sky130_fd_sc_hd__nor2_1 U18608 ( .A(n28590), .B(n24754), .Y(n27862) );
  sky130_fd_sc_hd__clkinv_1 U18609 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[6]), .Y(n27527) );
  sky130_fd_sc_hd__clkinv_1 U18610 ( .A(j202_soc_core_ahb2apb_00_state[2]), 
        .Y(n24814) );
  sky130_fd_sc_hd__nand3_1 U18611 ( .A(n20983), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_sck), .C(n20982), .Y(n24575) );
  sky130_fd_sc_hd__clkinv_1 U18612 ( .A(n25928), .Y(n26161) );
  sky130_fd_sc_hd__clkinv_1 U18613 ( .A(j202_soc_core_wbqspiflash_00_state[4]), 
        .Y(n26255) );
  sky130_fd_sc_hd__and2_0 U18614 ( .A(n25226), .B(n25224), .X(n20980) );
  sky130_fd_sc_hd__nor2_1 U18615 ( .A(n13248), .B(n13247), .Y(n13246) );
  sky130_fd_sc_hd__and2_0 U18616 ( .A(n20144), .B(n21750), .X(n12234) );
  sky130_fd_sc_hd__clkinv_1 U18617 ( .A(j202_soc_core_j22_cpu_id_op2_v_), .Y(
        n20428) );
  sky130_fd_sc_hd__nand3_1 U18618 ( .A(n27560), .B(n13160), .C(n11833), .Y(
        n27562) );
  sky130_fd_sc_hd__clkinv_1 U18619 ( .A(n20427), .Y(n13259) );
  sky130_fd_sc_hd__a21oi_1 U18620 ( .A1(j202_soc_core_memory0_ram_dout0[480]), 
        .A2(n21771), .B1(n20260), .Y(n20430) );
  sky130_fd_sc_hd__nand2_1 U18621 ( .A(n12878), .B(n19158), .Y(n12877) );
  sky130_fd_sc_hd__inv_2 U18622 ( .A(n19685), .Y(n26823) );
  sky130_fd_sc_hd__nand3_1 U18623 ( .A(n13018), .B(n13016), .C(n13015), .Y(
        n13014) );
  sky130_fd_sc_hd__clkinv_1 U18624 ( .A(n13020), .Y(n13017) );
  sky130_fd_sc_hd__inv_1 U18625 ( .A(n26904), .Y(n26834) );
  sky130_fd_sc_hd__clkinv_1 U18626 ( .A(
        j202_soc_core_intc_core_00_in_intreq[12]), .Y(n25504) );
  sky130_fd_sc_hd__clkinv_1 U18627 ( .A(n25351), .Y(n27194) );
  sky130_fd_sc_hd__clkinv_1 U18628 ( .A(n13007), .Y(n27522) );
  sky130_fd_sc_hd__clkinv_1 U18630 ( .A(n26790), .Y(n27402) );
  sky130_fd_sc_hd__clkinv_1 U18631 ( .A(n27654), .Y(n27656) );
  sky130_fd_sc_hd__clkinv_1 U18632 ( .A(n25237), .Y(n27435) );
  sky130_fd_sc_hd__clkinv_1 U18633 ( .A(n24208), .Y(n24209) );
  sky130_fd_sc_hd__clkinv_1 U18634 ( .A(n24193), .Y(n24194) );
  sky130_fd_sc_hd__clkinv_1 U18635 ( .A(n24174), .Y(n24175) );
  sky130_fd_sc_hd__clkinv_1 U18636 ( .A(gpio_en_o[0]), .Y(io_oeb[0]) );
  sky130_fd_sc_hd__clkinv_1 U18637 ( .A(gpio_en_o[4]), .Y(io_oeb[4]) );
  sky130_fd_sc_hd__clkinv_1 U18638 ( .A(gpio_en_o[8]), .Y(io_oeb[28]) );
  sky130_fd_sc_hd__clkinv_1 U18639 ( .A(gpio_en_o[16]), .Y(io_oeb[36]) );
  sky130_fd_sc_hd__nand2_1 U18640 ( .A(n23457), .B(n23456), .Y(io_out[8]) );
  sky130_fd_sc_hd__nor2b_1 U18641 ( .B_N(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[0]), .A(
        j202_soc_core_wbqspiflash_00_spif_override), .Y(io_out[10]) );
  sky130_fd_sc_hd__nor2b_1 U18642 ( .B_N(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[1]), .A(
        j202_soc_core_wbqspiflash_00_spif_override), .Y(io_out[11]) );
  sky130_fd_sc_hd__nor2_1 U18643 ( .A(n12766), .B(n12765), .Y(n12764) );
  sky130_fd_sc_hd__clkinv_1 U18644 ( .A(j202_soc_core_uart_TOP_tx_fifo_gb), 
        .Y(n27992) );
  sky130_fd_sc_hd__and2_0 U18645 ( .A(n27719), .B(
        j202_soc_core_wbqspiflash_00_spi_out[8]), .X(n29155) );
  sky130_fd_sc_hd__and2_0 U18646 ( .A(n27719), .B(
        j202_soc_core_wbqspiflash_00_spi_out[9]), .X(n29156) );
  sky130_fd_sc_hd__and2_0 U18647 ( .A(n27719), .B(
        j202_soc_core_wbqspiflash_00_spi_out[10]), .X(n29157) );
  sky130_fd_sc_hd__and2_0 U18648 ( .A(n27719), .B(
        j202_soc_core_wbqspiflash_00_spi_out[11]), .X(n29158) );
  sky130_fd_sc_hd__and2_0 U18649 ( .A(n27719), .B(
        j202_soc_core_wbqspiflash_00_spi_out[12]), .X(n29159) );
  sky130_fd_sc_hd__and2_0 U18650 ( .A(n27719), .B(
        j202_soc_core_wbqspiflash_00_spi_out[13]), .X(n29160) );
  sky130_fd_sc_hd__and2_0 U18651 ( .A(n27719), .B(
        j202_soc_core_wbqspiflash_00_spi_out[22]), .X(n29161) );
  sky130_fd_sc_hd__and2_0 U18652 ( .A(n27719), .B(
        j202_soc_core_wbqspiflash_00_spi_out[23]), .X(n29162) );
  sky130_fd_sc_hd__and2_0 U18653 ( .A(n27719), .B(
        j202_soc_core_wbqspiflash_00_spi_out[24]), .X(n29163) );
  sky130_fd_sc_hd__and2_0 U18654 ( .A(n27719), .B(
        j202_soc_core_wbqspiflash_00_spi_out[25]), .X(n29164) );
  sky130_fd_sc_hd__clkinv_1 U18656 ( .A(n28014), .Y(n28017) );
  sky130_fd_sc_hd__nor2_1 U18657 ( .A(n23972), .B(n12918), .Y(n12583) );
  sky130_fd_sc_hd__nand2b_1 U18658 ( .A_N(n26313), .B(n22581), .Y(n21366) );
  sky130_fd_sc_hd__and2_1 U18659 ( .A(n29067), .B(n29012), .X(n12244) );
  sky130_fd_sc_hd__and2_1 U18660 ( .A(n29067), .B(n29013), .X(n12260) );
  sky130_fd_sc_hd__and2_1 U18661 ( .A(n29067), .B(n29034), .X(n12263) );
  sky130_fd_sc_hd__and2_1 U18662 ( .A(n29067), .B(n29035), .X(n12245) );
  sky130_fd_sc_hd__and2_1 U18663 ( .A(n29067), .B(n29011), .X(n12242) );
  sky130_fd_sc_hd__and2_1 U18665 ( .A(n29067), .B(n29064), .X(n12239) );
  sky130_fd_sc_hd__and2_1 U18666 ( .A(n29067), .B(n29032), .X(n12255) );
  sky130_fd_sc_hd__and2_1 U18667 ( .A(n29067), .B(n29063), .X(n12254) );
  sky130_fd_sc_hd__o31ai_1 U18668 ( .A1(j202_soc_core_gpio_core_00_reg_addr[3]), .A2(n23454), .A3(n27658), .B1(n29594), .Y(n10676) );
  sky130_fd_sc_hd__clkbuf_1 U18669 ( .A(n10676), .X(n29315) );
  sky130_fd_sc_hd__clkinv_1 U18670 ( .A(n28881), .Y(n29086) );
  sky130_fd_sc_hd__nor2_1 U18671 ( .A(n23947), .B(n12918), .Y(n12582) );
  sky130_fd_sc_hd__clkinv_1 U18672 ( .A(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_wen), .Y(
        n25682) );
  sky130_fd_sc_hd__nand3_1 U18673 ( .A(n12916), .B(n25826), .C(
        j202_soc_core_j22_cpu_ml_macl[8]), .Y(n25827) );
  sky130_fd_sc_hd__clkinv_1 U18674 ( .A(n23442), .Y(n29239) );
  sky130_fd_sc_hd__and2_0 U18675 ( .A(n23907), .B(n23881), .X(n29166) );
  sky130_fd_sc_hd__and2_0 U18676 ( .A(n29056), .B(n23881), .X(n29203) );
  sky130_fd_sc_hd__and2_0 U18677 ( .A(n23907), .B(n23882), .X(n29167) );
  sky130_fd_sc_hd__and2_0 U18678 ( .A(n29056), .B(n23882), .X(n29204) );
  sky130_fd_sc_hd__and2_0 U18679 ( .A(n23907), .B(n23883), .X(n29168) );
  sky130_fd_sc_hd__and2_0 U18680 ( .A(n29056), .B(n23883), .X(n29206) );
  sky130_fd_sc_hd__and2_0 U18681 ( .A(n23907), .B(n23884), .X(n29169) );
  sky130_fd_sc_hd__and2_0 U18682 ( .A(n29056), .B(n23884), .X(n29207) );
  sky130_fd_sc_hd__and2_0 U18683 ( .A(n23907), .B(n23885), .X(n29170) );
  sky130_fd_sc_hd__and2_0 U18684 ( .A(n29056), .B(n23885), .X(n29208) );
  sky130_fd_sc_hd__and2_0 U18685 ( .A(n23907), .B(n23886), .X(n29171) );
  sky130_fd_sc_hd__and2_0 U18686 ( .A(n29056), .B(n23886), .X(n29209) );
  sky130_fd_sc_hd__and2_0 U18687 ( .A(n23900), .B(n23907), .X(n29185) );
  sky130_fd_sc_hd__and2_0 U18688 ( .A(n29056), .B(n23900), .X(n29193) );
  sky130_fd_sc_hd__and2_0 U18689 ( .A(n23907), .B(n23887), .X(n29172) );
  sky130_fd_sc_hd__and2_0 U18690 ( .A(n29056), .B(n23887), .X(n29217) );
  sky130_fd_sc_hd__and2_0 U18691 ( .A(n23901), .B(n23907), .X(n29186) );
  sky130_fd_sc_hd__and2_0 U18692 ( .A(n29056), .B(n23901), .X(n29210) );
  sky130_fd_sc_hd__and2_0 U18693 ( .A(n23907), .B(n23888), .X(n29173) );
  sky130_fd_sc_hd__and2_0 U18694 ( .A(n29056), .B(n23888), .X(n29194) );
  sky130_fd_sc_hd__and2_0 U18695 ( .A(n23902), .B(n23907), .X(n29187) );
  sky130_fd_sc_hd__and2_0 U18696 ( .A(n29056), .B(n23902), .X(n29211) );
  sky130_fd_sc_hd__and2_0 U18697 ( .A(n23907), .B(n23889), .X(n29174) );
  sky130_fd_sc_hd__and2_0 U18698 ( .A(n29056), .B(n23889), .X(n29212) );
  sky130_fd_sc_hd__and2_0 U18699 ( .A(n23907), .B(n23890), .X(n29175) );
  sky130_fd_sc_hd__and2_0 U18700 ( .A(n29056), .B(n23890), .X(n29195) );
  sky130_fd_sc_hd__and2_0 U18701 ( .A(n23907), .B(n23891), .X(n29176) );
  sky130_fd_sc_hd__and2_0 U18702 ( .A(n29056), .B(n23891), .X(n29213) );
  sky130_fd_sc_hd__and2_0 U18703 ( .A(n23903), .B(n23907), .X(n29188) );
  sky130_fd_sc_hd__and2_0 U18704 ( .A(n29056), .B(n23903), .X(n29196) );
  sky130_fd_sc_hd__and2_0 U18705 ( .A(n23904), .B(n23907), .X(n29189) );
  sky130_fd_sc_hd__and2_0 U18706 ( .A(n29056), .B(n23904), .X(n29200) );
  sky130_fd_sc_hd__and2_0 U18707 ( .A(n23905), .B(n23907), .X(n29190) );
  sky130_fd_sc_hd__and2_0 U18708 ( .A(n29056), .B(n23905), .X(n29214) );
  sky130_fd_sc_hd__and2_0 U18709 ( .A(n23907), .B(n23892), .X(n29177) );
  sky130_fd_sc_hd__and2_0 U18710 ( .A(n29056), .B(n23892), .X(n29219) );
  sky130_fd_sc_hd__and2_0 U18711 ( .A(n23907), .B(n23893), .X(n29178) );
  sky130_fd_sc_hd__and2_0 U18712 ( .A(n29056), .B(n23893), .X(n29218) );
  sky130_fd_sc_hd__and2_0 U18713 ( .A(n23907), .B(n23894), .X(n29179) );
  sky130_fd_sc_hd__and2_0 U18714 ( .A(n29056), .B(n23894), .X(n29201) );
  sky130_fd_sc_hd__and2_0 U18715 ( .A(n23907), .B(n23895), .X(n29180) );
  sky130_fd_sc_hd__and2_0 U18716 ( .A(n29056), .B(n23895), .X(n29197) );
  sky130_fd_sc_hd__and2_0 U18717 ( .A(n23907), .B(n23896), .X(n29181) );
  sky130_fd_sc_hd__and2_0 U18718 ( .A(n29056), .B(n23896), .X(n29202) );
  sky130_fd_sc_hd__and2_0 U18719 ( .A(n23907), .B(n23897), .X(n29182) );
  sky130_fd_sc_hd__and2_0 U18720 ( .A(n29056), .B(n23897), .X(n29198) );
  sky130_fd_sc_hd__and2_0 U18721 ( .A(n23906), .B(n23907), .X(n29191) );
  sky130_fd_sc_hd__and2_0 U18722 ( .A(n29056), .B(n23906), .X(n29199) );
  sky130_fd_sc_hd__and2_0 U18723 ( .A(n23908), .B(n23907), .X(n29192) );
  sky130_fd_sc_hd__and2_0 U18724 ( .A(n29056), .B(n23908), .X(n29215) );
  sky130_fd_sc_hd__and2_0 U18725 ( .A(n23907), .B(n23898), .X(n29183) );
  sky130_fd_sc_hd__and2_0 U18726 ( .A(n29056), .B(n23898), .X(n29205) );
  sky130_fd_sc_hd__and2_0 U18727 ( .A(n23907), .B(n23899), .X(n29184) );
  sky130_fd_sc_hd__and2_0 U18728 ( .A(n29056), .B(n23899), .X(n29216) );
  sky130_fd_sc_hd__nand3_1 U18729 ( .A(n22506), .B(n22507), .C(n11062), .Y(
        n29001) );
  sky130_fd_sc_hd__nand3_1 U18730 ( .A(n12916), .B(n26977), .C(n26871), .Y(
        n26880) );
  sky130_fd_sc_hd__nand3_1 U18731 ( .A(n12916), .B(n25826), .C(
        j202_soc_core_j22_cpu_ml_macl[15]), .Y(n25266) );
  sky130_fd_sc_hd__nand3_1 U18732 ( .A(n12916), .B(n25826), .C(
        j202_soc_core_j22_cpu_ml_macl[10]), .Y(n25050) );
  sky130_fd_sc_hd__o21a_1 U18733 ( .A1(n26951), .A2(n12420), .B1(n25054), .X(
        n25055) );
  sky130_fd_sc_hd__o22ai_1 U18734 ( .A1(n27226), .A2(n27427), .B1(n23079), 
        .B2(n12474), .Y(j202_soc_core_j22_cpu_rf_N3143) );
  sky130_fd_sc_hd__clkbuf_1 U18735 ( .A(n23325), .X(n29242) );
  sky130_fd_sc_hd__nand3_1 U18737 ( .A(n12916), .B(n25826), .C(
        j202_soc_core_j22_cpu_ml_macl[4]), .Y(n24587) );
  sky130_fd_sc_hd__nand3_1 U18738 ( .A(n12916), .B(n25826), .C(
        j202_soc_core_j22_cpu_ml_macl[1]), .Y(n24058) );
  sky130_fd_sc_hd__nand3_1 U18739 ( .A(n12916), .B(n25826), .C(
        j202_soc_core_j22_cpu_ml_macl[0]), .Y(n24604) );
  sky130_fd_sc_hd__o22ai_1 U18740 ( .A1(n27226), .A2(n24055), .B1(n23079), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N3155) );
  sky130_fd_sc_hd__clkinv_1 U18741 ( .A(n26899), .Y(n12469) );
  sky130_fd_sc_hd__nor2_1 U18742 ( .A(n27298), .B(n11130), .Y(n13193) );
  sky130_fd_sc_hd__nand3_1 U18743 ( .A(n21351), .B(n21350), .C(n21349), .Y(
        n28947) );
  sky130_fd_sc_hd__and2_0 U18744 ( .A(n27719), .B(
        j202_soc_core_wbqspiflash_00_spi_out[26]), .X(n29165) );
  sky130_fd_sc_hd__and2_0 U18745 ( .A(n27996), .B(n28624), .X(n10911) );
  sky130_fd_sc_hd__and2_0 U18746 ( .A(n23911), .B(n28623), .X(n29232) );
  sky130_fd_sc_hd__clkinv_1 U18747 ( .A(n28000), .Y(j202_soc_core_uart_TOP_N95) );
  sky130_fd_sc_hd__nand2b_1 U18748 ( .A_N(n23697), .B(n22581), .Y(n21338) );
  sky130_fd_sc_hd__nand2_1 U18749 ( .A(n23338), .B(n26159), .Y(
        j202_soc_core_wbqspiflash_00_N755) );
  sky130_fd_sc_hd__and2_0 U18750 ( .A(n28640), .B(n28639), .X(n28644) );
  sky130_fd_sc_hd__nand2b_1 U18751 ( .A_N(n26526), .B(n22581), .Y(n15525) );
  sky130_fd_sc_hd__nand2_1 U18752 ( .A(n11126), .B(n25108), .Y(n25109) );
  sky130_fd_sc_hd__nor2_1 U18753 ( .A(n28590), .B(n12200), .Y(n29347) );
  sky130_fd_sc_hd__o211ai_1 U18754 ( .A1(n11793), .A2(n24704), .B1(n24706), 
        .C1(n12226), .Y(n24707) );
  sky130_fd_sc_hd__clkinv_1 U18755 ( .A(n27167), .Y(n29357) );
  sky130_fd_sc_hd__nor2_1 U18756 ( .A(n13158), .B(n13157), .Y(n20707) );
  sky130_fd_sc_hd__nand2_1 U18757 ( .A(n23492), .B(n23704), .Y(n29236) );
  sky130_fd_sc_hd__nand2_1 U18758 ( .A(n24110), .B(n13238), .Y(n13237) );
  sky130_fd_sc_hd__a31o_1 U18759 ( .A1(n27657), .A2(n27656), .A3(n24173), .B1(
        n28590), .X(n29243) );
  sky130_fd_sc_hd__and2_0 U18760 ( .A(j202_soc_core_j22_cpu_memop_MEM__2_), 
        .B(j202_soc_core_j22_cpu_memop_MEM__1_), .X(n15778) );
  sky130_fd_sc_hd__nand3_1 U18761 ( .A(n19075), .B(n22234), .C(n19074), .Y(
        n28983) );
  sky130_fd_sc_hd__and2_0 U18762 ( .A(n22503), .B(n19073), .X(n19074) );
  sky130_fd_sc_hd__clkinv_1 U18763 ( .A(n12200), .Y(
        j202_soc_core_ahbcs_6__HREADY_) );
  sky130_fd_sc_hd__clkinv_1 U18764 ( .A(la_oenb[31]), .Y(n23866) );
  sky130_fd_sc_hd__clkinv_1 U18765 ( .A(la_oenb[30]), .Y(n23867) );
  sky130_fd_sc_hd__clkinv_1 U18766 ( .A(la_oenb[29]), .Y(n23868) );
  sky130_fd_sc_hd__clkinv_1 U18767 ( .A(la_oenb[28]), .Y(n23869) );
  sky130_fd_sc_hd__clkinv_1 U18768 ( .A(la_oenb[27]), .Y(n23870) );
  sky130_fd_sc_hd__clkinv_1 U18769 ( .A(la_oenb[26]), .Y(n23871) );
  sky130_fd_sc_hd__clkinv_1 U18770 ( .A(la_oenb[25]), .Y(n23872) );
  sky130_fd_sc_hd__clkinv_1 U18771 ( .A(la_oenb[24]), .Y(n23873) );
  sky130_fd_sc_hd__clkinv_1 U18772 ( .A(la_oenb[23]), .Y(n23874) );
  sky130_fd_sc_hd__clkinv_1 U18773 ( .A(la_oenb[22]), .Y(n23875) );
  sky130_fd_sc_hd__clkinv_1 U18774 ( .A(la_oenb[21]), .Y(n23876) );
  sky130_fd_sc_hd__clkinv_1 U18775 ( .A(la_oenb[20]), .Y(n23877) );
  sky130_fd_sc_hd__clkinv_1 U18776 ( .A(la_oenb[19]), .Y(n23878) );
  sky130_fd_sc_hd__clkinv_1 U18777 ( .A(la_oenb[18]), .Y(n23879) );
  sky130_fd_sc_hd__clkinv_1 U18778 ( .A(la_oenb[17]), .Y(n23880) );
  sky130_fd_sc_hd__and2_0 U18779 ( .A(n29092), .B(wbs_dat_i[1]), .X(n13) );
  sky130_fd_sc_hd__and2_0 U18780 ( .A(n29092), .B(wbs_dat_i[2]), .X(n14) );
  sky130_fd_sc_hd__and2_0 U18781 ( .A(n29092), .B(wbs_dat_i[3]), .X(n15) );
  sky130_fd_sc_hd__and2_0 U18782 ( .A(n29092), .B(wbs_dat_i[4]), .X(n16) );
  sky130_fd_sc_hd__and2_0 U18783 ( .A(n29092), .B(wbs_dat_i[5]), .X(n17) );
  sky130_fd_sc_hd__and2_0 U18784 ( .A(n29092), .B(wbs_dat_i[6]), .X(n18) );
  sky130_fd_sc_hd__and2_0 U18785 ( .A(n29092), .B(wbs_dat_i[7]), .X(n19) );
  sky130_fd_sc_hd__and2_0 U18786 ( .A(n29092), .B(wbs_dat_i[8]), .X(n21) );
  sky130_fd_sc_hd__and2_0 U18787 ( .A(n23690), .B(wbs_dat_i[9]), .X(n220) );
  sky130_fd_sc_hd__and2_0 U18788 ( .A(n23690), .B(wbs_dat_i[10]), .X(n230) );
  sky130_fd_sc_hd__and2_0 U18789 ( .A(n23690), .B(wbs_dat_i[11]), .X(n240) );
  sky130_fd_sc_hd__and2_0 U18790 ( .A(n23690), .B(wbs_dat_i[12]), .X(n250) );
  sky130_fd_sc_hd__and2_0 U18791 ( .A(n23690), .B(wbs_dat_i[13]), .X(n260) );
  sky130_fd_sc_hd__and2_0 U18792 ( .A(n23690), .B(wbs_dat_i[14]), .X(n270) );
  sky130_fd_sc_hd__a31o_1 U18793 ( .A1(n29092), .A2(wbs_we_i), .A3(
        wbs_sel_i[1]), .B1(wb_rst_i), .X(n20) );
  sky130_fd_sc_hd__and2_0 U18794 ( .A(n23690), .B(wbs_dat_i[15]), .X(n280) );
  sky130_fd_sc_hd__and2_0 U18795 ( .A(n23690), .B(wbs_dat_i[16]), .X(n300) );
  sky130_fd_sc_hd__and2_0 U18796 ( .A(n23690), .B(wbs_dat_i[17]), .X(n310) );
  sky130_fd_sc_hd__and2_0 U18797 ( .A(n23690), .B(wbs_dat_i[18]), .X(n320) );
  sky130_fd_sc_hd__and2_0 U18798 ( .A(n23690), .B(wbs_dat_i[19]), .X(n330) );
  sky130_fd_sc_hd__and2_0 U18799 ( .A(n23690), .B(wbs_dat_i[20]), .X(n340) );
  sky130_fd_sc_hd__and2_0 U18800 ( .A(n29092), .B(wbs_dat_i[21]), .X(n350) );
  sky130_fd_sc_hd__and2_0 U18801 ( .A(n29092), .B(wbs_dat_i[22]), .X(n360) );
  sky130_fd_sc_hd__a31o_1 U18802 ( .A1(n29092), .A2(wbs_we_i), .A3(
        wbs_sel_i[2]), .B1(wb_rst_i), .X(n290) );
  sky130_fd_sc_hd__and2_0 U18803 ( .A(n29092), .B(wbs_dat_i[23]), .X(n370) );
  sky130_fd_sc_hd__and2_0 U18804 ( .A(n29092), .B(wbs_dat_i[24]), .X(n390) );
  sky130_fd_sc_hd__and2_0 U18805 ( .A(n23690), .B(wbs_dat_i[25]), .X(n400) );
  sky130_fd_sc_hd__and2_0 U18806 ( .A(n29092), .B(wbs_dat_i[26]), .X(n410) );
  sky130_fd_sc_hd__and2_0 U18807 ( .A(n29092), .B(wbs_dat_i[27]), .X(n420) );
  sky130_fd_sc_hd__and2_0 U18808 ( .A(n29092), .B(wbs_dat_i[28]), .X(n430) );
  sky130_fd_sc_hd__and2_0 U18809 ( .A(n29092), .B(wbs_dat_i[29]), .X(n440) );
  sky130_fd_sc_hd__and2_0 U18810 ( .A(n29092), .B(wbs_dat_i[30]), .X(n450) );
  sky130_fd_sc_hd__a31o_1 U18811 ( .A1(n29092), .A2(wbs_we_i), .A3(
        wbs_sel_i[3]), .B1(wb_rst_i), .X(n380) );
  sky130_fd_sc_hd__and2_0 U18812 ( .A(n29092), .B(wbs_dat_i[31]), .X(n460) );
  sky130_fd_sc_hd__clkbuf_1 U18813 ( .A(n23690), .X(n29092) );
  sky130_fd_sc_hd__and4_1 U18814 ( .A(n13173), .B(n13178), .C(n13165), .D(
        n13177), .X(n12148) );
  sky130_fd_sc_hd__inv_2 U18815 ( .A(n12187), .Y(n15128) );
  sky130_fd_sc_hd__inv_2 U18816 ( .A(n12187), .Y(n16278) );
  sky130_fd_sc_hd__and2_4 U18818 ( .A(n22278), .B(n13152), .X(n12150) );
  sky130_fd_sc_hd__and4_1 U18820 ( .A(n13167), .B(n13175), .C(n13171), .D(
        n13172), .X(n12155) );
  sky130_fd_sc_hd__clkinv_1 U18821 ( .A(n25338), .Y(n27187) );
  sky130_fd_sc_hd__inv_2 U18822 ( .A(n16261), .Y(n13793) );
  sky130_fd_sc_hd__clkinv_1 U18823 ( .A(n18916), .Y(n26329) );
  sky130_fd_sc_hd__nand2b_1 U18824 ( .A_N(n12353), .B(n24781), .Y(n25259) );
  sky130_fd_sc_hd__nand2_2 U18825 ( .A(n17391), .B(n17390), .Y(n17392) );
  sky130_fd_sc_hd__and2_4 U18826 ( .A(n18871), .B(n17357), .X(n12159) );
  sky130_fd_sc_hd__buf_4 U18827 ( .A(j202_soc_core_j22_cpu_ml_bufa[17]), .X(
        n18300) );
  sky130_fd_sc_hd__and2_1 U18830 ( .A(n20308), .B(n20842), .X(n12165) );
  sky130_fd_sc_hd__buf_6 U18831 ( .A(n23256), .X(n12916) );
  sky130_fd_sc_hd__buf_2 U18832 ( .A(n13396), .X(n17314) );
  sky130_fd_sc_hd__clkinv_1 U18833 ( .A(n23530), .Y(n27192) );
  sky130_fd_sc_hd__clkinv_1 U18834 ( .A(n27192), .Y(n27460) );
  sky130_fd_sc_hd__nand3_2 U18836 ( .A(n18865), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .C(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .Y(n17357) );
  sky130_fd_sc_hd__clkinv_1 U18838 ( .A(n13986), .Y(n23502) );
  sky130_fd_sc_hd__or2_1 U18839 ( .A(n17839), .B(n17840), .X(n12173) );
  sky130_fd_sc_hd__or2_2 U18841 ( .A(n13675), .B(n13659), .X(n12176) );
  sky130_fd_sc_hd__nand2_2 U18842 ( .A(n24591), .B(n24590), .Y(n27208) );
  sky130_fd_sc_hd__xor2_1 U18843 ( .A(j202_soc_core_j22_cpu_ml_bufa[20]), .B(
        j202_soc_core_j22_cpu_ml_bufa[19]), .X(n12483) );
  sky130_fd_sc_hd__or2_2 U18844 ( .A(n18827), .B(n18828), .X(n12178) );
  sky130_fd_sc_hd__and2_1 U18846 ( .A(n20736), .B(n21685), .X(n12180) );
  sky130_fd_sc_hd__clkinv_1 U18847 ( .A(n17217), .Y(n20387) );
  sky130_fd_sc_hd__inv_2 U18848 ( .A(n14668), .Y(n14204) );
  sky130_fd_sc_hd__and4_1 U18849 ( .A(n14585), .B(n14584), .C(n14583), .D(
        n14582), .X(n12188) );
  sky130_fd_sc_hd__and4_1 U18850 ( .A(n13970), .B(n13969), .C(n13968), .D(
        n13967), .X(n12189) );
  sky130_fd_sc_hd__and4_1 U18851 ( .A(n13631), .B(n13630), .C(n13629), .D(
        n13628), .X(n12190) );
  sky130_fd_sc_hd__clkinv_1 U18852 ( .A(j202_soc_core_intc_core_00_rg_ipr[10]), 
        .Y(n25349) );
  sky130_fd_sc_hd__clkinv_1 U18853 ( .A(j202_soc_core_intc_core_00_rg_ipr[25]), 
        .Y(n25196) );
  sky130_fd_sc_hd__inv_2 U18854 ( .A(j202_soc_core_intc_core_00_rg_ipr[21]), 
        .Y(n19623) );
  sky130_fd_sc_hd__and4_1 U18855 ( .A(n14646), .B(n14645), .C(n14644), .D(
        n14643), .X(n12195) );
  sky130_fd_sc_hd__inv_2 U18856 ( .A(n14465), .Y(n16369) );
  sky130_fd_sc_hd__inv_2 U18857 ( .A(n14465), .Y(n16285) );
  sky130_fd_sc_hd__o211a_2 U18858 ( .A1(n26565), .A2(n11143), .B1(n21323), 
        .C1(n21322), .X(n12196) );
  sky130_fd_sc_hd__o211a_2 U18860 ( .A1(n26570), .A2(n11143), .B1(n15658), 
        .C1(n15657), .X(n12198) );
  sky130_fd_sc_hd__o211a_2 U18861 ( .A1(n25403), .A2(n11143), .B1(n15769), 
        .C1(n15768), .X(n12199) );
  sky130_fd_sc_hd__and4_1 U18862 ( .A(n13834), .B(n13833), .C(n13832), .D(
        n13831), .X(n12201) );
  sky130_fd_sc_hd__and4_1 U18863 ( .A(n14607), .B(n14606), .C(n14605), .D(
        n14604), .X(n12202) );
  sky130_fd_sc_hd__and4_1 U18864 ( .A(n13746), .B(n13745), .C(n13744), .D(
        n13743), .X(n12203) );
  sky130_fd_sc_hd__o21a_1 U18866 ( .A1(n19815), .A2(n19796), .B1(n19795), .X(
        n12205) );
  sky130_fd_sc_hd__nor2_1 U18867 ( .A(n23769), .B(n12353), .Y(n23770) );
  sky130_fd_sc_hd__clkinv_1 U18868 ( .A(n24768), .Y(n24770) );
  sky130_fd_sc_hd__inv_2 U18869 ( .A(n11104), .Y(n25157) );
  sky130_fd_sc_hd__clkbuf_1 U18870 ( .A(n12502), .X(n12757) );
  sky130_fd_sc_hd__a22o_1 U18871 ( .A1(n17497), .A2(n17496), .B1(n17495), .B2(
        n17494), .X(n12209) );
  sky130_fd_sc_hd__and4_1 U18872 ( .A(n14160), .B(n14159), .C(n14158), .D(
        n14157), .X(n12210) );
  sky130_fd_sc_hd__and4_1 U18873 ( .A(n14748), .B(n14747), .C(n14746), .D(
        n14745), .X(n12211) );
  sky130_fd_sc_hd__and4_1 U18874 ( .A(n25395), .B(n26398), .C(n25394), .D(
        n25393), .X(n12212) );
  sky130_fd_sc_hd__and4_1 U18875 ( .A(n14392), .B(n14391), .C(n14390), .D(
        n14389), .X(n12214) );
  sky130_fd_sc_hd__and4_1 U18876 ( .A(n13910), .B(n13909), .C(n13908), .D(
        n13907), .X(n12215) );
  sky130_fd_sc_hd__o211a_2 U18877 ( .A1(n26704), .A2(n11143), .B1(n15303), 
        .C1(n15302), .X(n12216) );
  sky130_fd_sc_hd__and4_1 U18878 ( .A(n14147), .B(n14146), .C(n14145), .D(
        n14144), .X(n12217) );
  sky130_fd_sc_hd__and4_1 U18879 ( .A(n13819), .B(n13818), .C(n13817), .D(
        n13816), .X(n12218) );
  sky130_fd_sc_hd__and4_1 U18880 ( .A(n15110), .B(n15109), .C(n15108), .D(
        n15107), .X(n12219) );
  sky130_fd_sc_hd__and4_1 U18881 ( .A(n13808), .B(n13807), .C(n13806), .D(
        n13805), .X(n12221) );
  sky130_fd_sc_hd__and4_1 U18882 ( .A(n13963), .B(n13962), .C(n13961), .D(
        n13960), .X(n12222) );
  sky130_fd_sc_hd__and4_1 U18883 ( .A(n14048), .B(n14047), .C(n14046), .D(
        n14045), .X(n12223) );
  sky130_fd_sc_hd__and4_1 U18884 ( .A(n14729), .B(n14728), .C(n14727), .D(
        n14726), .X(n12224) );
  sky130_fd_sc_hd__inv_2 U18885 ( .A(n23163), .Y(n23164) );
  sky130_fd_sc_hd__and3_1 U18886 ( .A(n20960), .B(n13235), .C(n20962), .X(
        n12225) );
  sky130_fd_sc_hd__o21a_1 U18887 ( .A1(n11106), .A2(n24705), .B1(n27785), .X(
        n12226) );
  sky130_fd_sc_hd__buf_4 U18888 ( .A(n18903), .X(n12321) );
  sky130_fd_sc_hd__buf_2 U18889 ( .A(n18903), .X(n22521) );
  sky130_fd_sc_hd__nand3_1 U18891 ( .A(n20283), .B(n20282), .C(n20281), .Y(
        n29033) );
  sky130_fd_sc_hd__and2_1 U18892 ( .A(n29067), .B(n27621), .X(n12228) );
  sky130_fd_sc_hd__and2_1 U18893 ( .A(n12792), .B(n20971), .X(n12229) );
  sky130_fd_sc_hd__and2_1 U18894 ( .A(n29067), .B(n29066), .X(n12236) );
  sky130_fd_sc_hd__nand2_1 U18895 ( .A(n13011), .B(n29070), .Y(n12450) );
  sky130_fd_sc_hd__and4_1 U18896 ( .A(n20272), .B(n20271), .C(n20270), .D(
        n20269), .X(n12241) );
  sky130_fd_sc_hd__and4_1 U18897 ( .A(n16235), .B(n16226), .C(n16234), .D(
        n16232), .X(n12246) );
  sky130_fd_sc_hd__and4_1 U18898 ( .A(n20825), .B(n20824), .C(n20823), .D(
        n20822), .X(n12248) );
  sky130_fd_sc_hd__and4_1 U18899 ( .A(n13886), .B(n13885), .C(n13884), .D(
        n13883), .X(n12249) );
  sky130_fd_sc_hd__nor2_1 U18900 ( .A(n21778), .B(n20430), .Y(n12250) );
  sky130_fd_sc_hd__and4_1 U18901 ( .A(n13164), .B(n13176), .C(n13168), .D(
        n13169), .X(n12257) );
  sky130_fd_sc_hd__and4_1 U18902 ( .A(n14362), .B(n14361), .C(n14360), .D(
        n14359), .X(n12258) );
  sky130_fd_sc_hd__and4_1 U18903 ( .A(n14260), .B(n14259), .C(n14258), .D(
        n14257), .X(n12259) );
  sky130_fd_sc_hd__o211ai_1 U18904 ( .A1(n25871), .A2(n26550), .B1(n24481), 
        .C1(n23849), .Y(n12261) );
  sky130_fd_sc_hd__and2_1 U18905 ( .A(n29067), .B(n27620), .X(n12265) );
  sky130_fd_sc_hd__and2_1 U18906 ( .A(n29067), .B(n29061), .X(n12266) );
  sky130_fd_sc_hd__and2_1 U18909 ( .A(n29067), .B(n24322), .X(n12274) );
  sky130_fd_sc_hd__clkinv_1 U18910 ( .A(n29035), .Y(n27639) );
  sky130_fd_sc_hd__clkinv_1 U18911 ( .A(n29011), .Y(n27638) );
  sky130_fd_sc_hd__clkinv_1 U18912 ( .A(n29010), .Y(n27637) );
  sky130_fd_sc_hd__clkinv_1 U18913 ( .A(n29012), .Y(n27636) );
  sky130_fd_sc_hd__clkinv_1 U18914 ( .A(n29013), .Y(n27635) );
  sky130_fd_sc_hd__clkinv_1 U18916 ( .A(n29061), .Y(n27622) );
  sky130_fd_sc_hd__nand3_1 U18917 ( .A(n22295), .B(n22294), .C(n22293), .Y(
        n29061) );
  sky130_fd_sc_hd__clkinv_1 U18919 ( .A(n27224), .Y(n27225) );
  sky130_fd_sc_hd__clkinv_1 U18920 ( .A(n27227), .Y(n27228) );
  sky130_fd_sc_hd__clkinv_1 U18921 ( .A(n27214), .Y(n27215) );
  sky130_fd_sc_hd__clkinv_1 U18922 ( .A(n27210), .Y(n27211) );
  sky130_fd_sc_hd__inv_1 U18923 ( .A(n23178), .Y(n26371) );
  sky130_fd_sc_hd__nand3_1 U18924 ( .A(n23177), .B(n23120), .C(n23119), .Y(
        n27574) );
  sky130_fd_sc_hd__nor2_1 U18925 ( .A(n23481), .B(n13552), .Y(n23174) );
  sky130_fd_sc_hd__a21o_2 U18926 ( .A1(n23517), .A2(n23516), .B1(n14849), .X(
        n27214) );
  sky130_fd_sc_hd__a21o_2 U18927 ( .A1(n23527), .A2(n23526), .B1(n14849), .X(
        n27124) );
  sky130_fd_sc_hd__xor2_1 U18928 ( .A(j202_soc_core_qspi_wb_addr[8]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[8]), .X(n12292) );
  sky130_fd_sc_hd__nor2_1 U18929 ( .A(n20429), .B(n20547), .Y(n21750) );
  sky130_fd_sc_hd__clkinv_1 U18930 ( .A(n21750), .Y(n21778) );
  sky130_fd_sc_hd__clkinv_1 U18931 ( .A(n24778), .Y(n24785) );
  sky130_fd_sc_hd__clkinv_1 U18933 ( .A(n22682), .Y(n22421) );
  sky130_fd_sc_hd__a22oi_1 U18934 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__7_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__7_), .Y(n12293) );
  sky130_fd_sc_hd__clkinv_1 U18935 ( .A(n20967), .Y(n21776) );
  sky130_fd_sc_hd__and3_1 U18936 ( .A(n26396), .B(n26397), .C(n26398), .X(
        n12294) );
  sky130_fd_sc_hd__buf_4 U18937 ( .A(j202_soc_core_j22_cpu_ml_bufa[23]), .X(
        n22029) );
  sky130_fd_sc_hd__clkinv_1 U18938 ( .A(n18656), .Y(n18057) );
  sky130_fd_sc_hd__clkinv_1 U18939 ( .A(n23296), .Y(n22702) );
  sky130_fd_sc_hd__nor2_1 U18940 ( .A(n11713), .B(n18916), .Y(n26802) );
  sky130_fd_sc_hd__clkinv_1 U18942 ( .A(n21813), .Y(n22713) );
  sky130_fd_sc_hd__a22oi_1 U18943 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__4_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__4_), .Y(n12297) );
  sky130_fd_sc_hd__nand2_1 U18944 ( .A(n23573), .B(n23297), .Y(n23293) );
  sky130_fd_sc_hd__clkinv_1 U18945 ( .A(n23293), .Y(n22768) );
  sky130_fd_sc_hd__clkinv_1 U18946 ( .A(n22450), .Y(n24061) );
  sky130_fd_sc_hd__clkinv_1 U18947 ( .A(n19828), .Y(n13022) );
  sky130_fd_sc_hd__clkinv_1 U18948 ( .A(n18882), .Y(n23257) );
  sky130_fd_sc_hd__nor2_1 U18949 ( .A(n12302), .B(n12141), .Y(n18379) );
  sky130_fd_sc_hd__nor2_1 U18950 ( .A(n12141), .B(n18375), .Y(n18408) );
  sky130_fd_sc_hd__nor2_1 U18951 ( .A(n12141), .B(n18427), .Y(n18451) );
  sky130_fd_sc_hd__nor2_1 U18952 ( .A(n12141), .B(n18709), .Y(n18754) );
  sky130_fd_sc_hd__nor2_1 U18953 ( .A(n12141), .B(n18668), .Y(n18677) );
  sky130_fd_sc_hd__nor2_1 U18954 ( .A(n12141), .B(n18480), .Y(n18532) );
  sky130_fd_sc_hd__nor2_1 U18955 ( .A(n12141), .B(n18655), .Y(n18703) );
  sky130_fd_sc_hd__nor2_1 U18956 ( .A(n12141), .B(n17381), .Y(n18629) );
  sky130_fd_sc_hd__nor2_1 U18957 ( .A(n12141), .B(n18632), .Y(n18763) );
  sky130_fd_sc_hd__nor2_1 U18958 ( .A(n12141), .B(n18620), .Y(n18634) );
  sky130_fd_sc_hd__nor2_1 U18959 ( .A(n12141), .B(n18512), .Y(n18680) );
  sky130_fd_sc_hd__nor2_1 U18960 ( .A(n12141), .B(n17368), .Y(n22058) );
  sky130_fd_sc_hd__nor2_1 U18961 ( .A(n12141), .B(n17362), .Y(n17377) );
  sky130_fd_sc_hd__nor2_1 U18962 ( .A(n12141), .B(n17373), .Y(n18616) );
  sky130_fd_sc_hd__nor2_1 U18963 ( .A(n12141), .B(n22053), .Y(n22065) );
  sky130_fd_sc_hd__nand2b_1 U18964 ( .A_N(n12305), .B(n12304), .Y(n18325) );
  sky130_fd_sc_hd__xnor2_1 U18965 ( .A(n18309), .B(n12305), .Y(n18555) );
  sky130_fd_sc_hd__nand2_1 U18966 ( .A(n12307), .B(n12306), .Y(n18417) );
  sky130_fd_sc_hd__nand2_1 U18967 ( .A(n18357), .B(n18356), .Y(n12306) );
  sky130_fd_sc_hd__o21ai_1 U18968 ( .A1(n18356), .A2(n18357), .B1(n18355), .Y(
        n12307) );
  sky130_fd_sc_hd__xnor2_1 U18969 ( .A(n18355), .B(n12308), .Y(n18599) );
  sky130_fd_sc_hd__xnor2_1 U18970 ( .A(n18356), .B(n18357), .Y(n12308) );
  sky130_fd_sc_hd__nand2_1 U18971 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[23]), .Y(n12309) );
  sky130_fd_sc_hd__nand2_1 U18972 ( .A(n12311), .B(n26863), .Y(n12310) );
  sky130_fd_sc_hd__xnor2_1 U18973 ( .A(n22108), .B(n12312), .Y(n12311) );
  sky130_fd_sc_hd__o21ai_1 U18974 ( .A1(n22897), .A2(n22107), .B1(n22106), .Y(
        n12312) );
  sky130_fd_sc_hd__nand2_1 U18975 ( .A(n23275), .B(n23274), .Y(n25337) );
  sky130_fd_sc_hd__nand2_2 U18976 ( .A(n23234), .B(n26863), .Y(n23275) );
  sky130_fd_sc_hd__nand2_1 U18977 ( .A(n12315), .B(n12314), .Y(n17901) );
  sky130_fd_sc_hd__nand2_1 U18978 ( .A(n17676), .B(n17677), .Y(n12314) );
  sky130_fd_sc_hd__o21ai_1 U18979 ( .A1(n17677), .A2(n17676), .B1(n17675), .Y(
        n12315) );
  sky130_fd_sc_hd__xnor2_1 U18980 ( .A(n17675), .B(n12316), .Y(n17906) );
  sky130_fd_sc_hd__nand2_1 U18981 ( .A(n12320), .B(n18820), .Y(n21792) );
  sky130_fd_sc_hd__xnor2_1 U18982 ( .A(n18549), .B(n12921), .Y(n12320) );
  sky130_fd_sc_hd__inv_2 U18983 ( .A(n12321), .Y(n21512) );
  sky130_fd_sc_hd__nand2_1 U18984 ( .A(n12321), .B(n12178), .Y(n18906) );
  sky130_fd_sc_hd__nand2_1 U18985 ( .A(n19475), .B(n12321), .Y(n19477) );
  sky130_fd_sc_hd__nand2_1 U18986 ( .A(n22133), .B(n12321), .Y(n22135) );
  sky130_fd_sc_hd__nand2_1 U18987 ( .A(n22943), .B(n12321), .Y(n22946) );
  sky130_fd_sc_hd__nand2_1 U18988 ( .A(n22800), .B(n22521), .Y(n22802) );
  sky130_fd_sc_hd__nand2_1 U18989 ( .A(n22525), .B(n18903), .Y(n22527) );
  sky130_fd_sc_hd__nand2_1 U18990 ( .A(n22105), .B(n12321), .Y(n22107) );
  sky130_fd_sc_hd__nand2_1 U18991 ( .A(n18856), .B(n12321), .Y(n18858) );
  sky130_fd_sc_hd__nand2_1 U18992 ( .A(n21493), .B(n12321), .Y(n21495) );
  sky130_fd_sc_hd__nand2_1 U18993 ( .A(n22167), .B(n12321), .Y(n22169) );
  sky130_fd_sc_hd__nand2_1 U18994 ( .A(n22191), .B(n22521), .Y(n22193) );
  sky130_fd_sc_hd__nand2_1 U18995 ( .A(n22363), .B(n22521), .Y(n22365) );
  sky130_fd_sc_hd__nand2_1 U18996 ( .A(n22400), .B(n12321), .Y(n22402) );
  sky130_fd_sc_hd__nand2_1 U18997 ( .A(n22557), .B(n22521), .Y(n22559) );
  sky130_fd_sc_hd__nand2_1 U18998 ( .A(n22660), .B(n12321), .Y(n22662) );
  sky130_fd_sc_hd__nand2_1 U18999 ( .A(n22431), .B(n12321), .Y(n22433) );
  sky130_fd_sc_hd__nand2_1 U19000 ( .A(n22482), .B(n12321), .Y(n22484) );
  sky130_fd_sc_hd__nand2_1 U19001 ( .A(n12322), .B(n18819), .Y(n21419) );
  sky130_fd_sc_hd__xnor2_1 U19002 ( .A(n18546), .B(n18477), .Y(n12322) );
  sky130_fd_sc_hd__nor2_4 U19003 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]), .B(n12323), .Y(n17358) );
  sky130_fd_sc_hd__inv_2 U19004 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[4]), 
        .Y(n12323) );
  sky130_fd_sc_hd__nand2_1 U19005 ( .A(n12325), .B(n22768), .Y(n12324) );
  sky130_fd_sc_hd__nand2_1 U19006 ( .A(n19197), .B(n13338), .Y(n25232) );
  sky130_fd_sc_hd__nand2_1 U19007 ( .A(n12324), .B(n19211), .Y(n12329) );
  sky130_fd_sc_hd__nand2_1 U19009 ( .A(n27786), .B(n27787), .Y(n12328) );
  sky130_fd_sc_hd__nand2_1 U19010 ( .A(n12841), .B(n22218), .Y(n12330) );
  sky130_fd_sc_hd__nand2_1 U19011 ( .A(j202_soc_core_memory0_ram_dout0[52]), 
        .B(n21604), .Y(n12331) );
  sky130_fd_sc_hd__nand2_1 U19012 ( .A(j202_soc_core_memory0_ram_dout0[276]), 
        .B(n21605), .Y(n12332) );
  sky130_fd_sc_hd__nand2_1 U19013 ( .A(n12333), .B(n12343), .Y(n20833) );
  sky130_fd_sc_hd__nand4_1 U19014 ( .A(n12337), .B(n12336), .C(n12338), .D(
        n12335), .Y(n12334) );
  sky130_fd_sc_hd__nand2_1 U19015 ( .A(j202_soc_core_memory0_ram_dout0[310]), 
        .B(n21603), .Y(n12335) );
  sky130_fd_sc_hd__nand2_1 U19016 ( .A(j202_soc_core_memory0_ram_dout0[22]), 
        .B(n21733), .Y(n12336) );
  sky130_fd_sc_hd__nand2_1 U19017 ( .A(j202_soc_core_memory0_ram_dout0[54]), 
        .B(n21604), .Y(n12337) );
  sky130_fd_sc_hd__nand2_1 U19018 ( .A(j202_soc_core_memory0_ram_dout0[86]), 
        .B(n21734), .Y(n12338) );
  sky130_fd_sc_hd__nand4_1 U19019 ( .A(n15391), .B(n12342), .C(n12341), .D(
        n12340), .Y(n12339) );
  sky130_fd_sc_hd__nand2_1 U19020 ( .A(j202_soc_core_memory0_ram_dout0[118]), 
        .B(n21591), .Y(n12340) );
  sky130_fd_sc_hd__nand2_1 U19021 ( .A(j202_soc_core_memory0_ram_dout0[150]), 
        .B(n21592), .Y(n12341) );
  sky130_fd_sc_hd__nand2_1 U19022 ( .A(j202_soc_core_memory0_ram_dout0[214]), 
        .B(n21732), .Y(n12342) );
  sky130_fd_sc_hd__nand4_1 U19023 ( .A(n15394), .B(n15395), .C(n15389), .D(
        n15390), .Y(n12344) );
  sky130_fd_sc_hd__nand4_1 U19024 ( .A(n15393), .B(n15307), .C(n15392), .D(
        n15388), .Y(n12345) );
  sky130_fd_sc_hd__nand2_1 U19025 ( .A(n12641), .B(n24310), .Y(n24300) );
  sky130_fd_sc_hd__nand2_2 U19026 ( .A(n24400), .B(n12641), .Y(n27964) );
  sky130_fd_sc_hd__nand2_1 U19027 ( .A(n12731), .B(n12641), .Y(n24294) );
  sky130_fd_sc_hd__xnor2_1 U19028 ( .A(n18026), .B(n18027), .Y(n17950) );
  sky130_fd_sc_hd__nor2_2 U19029 ( .A(n22243), .B(n22242), .Y(n23278) );
  sky130_fd_sc_hd__and2_0 U19030 ( .A(n20958), .B(n20836), .X(n12347) );
  sky130_fd_sc_hd__nand2_1 U19031 ( .A(n23241), .B(n24499), .Y(n25083) );
  sky130_fd_sc_hd__nand2b_1 U19032 ( .A_N(n25027), .B(n12349), .Y(n12348) );
  sky130_fd_sc_hd__nor2_1 U19033 ( .A(n17146), .B(n12421), .Y(n17135) );
  sky130_fd_sc_hd__nor2_1 U19034 ( .A(n24061), .B(n22458), .Y(n24381) );
  sky130_fd_sc_hd__nand2b_1 U19035 ( .A_N(n21916), .B(n22714), .Y(n13066) );
  sky130_fd_sc_hd__nor2_1 U19036 ( .A(n29077), .B(n23185), .Y(n27880) );
  sky130_fd_sc_hd__or2_0 U19037 ( .A(n26378), .B(n27461), .X(n12354) );
  sky130_fd_sc_hd__nand2_1 U19038 ( .A(n12354), .B(n24558), .Y(
        j202_soc_core_j22_cpu_rf_N3247) );
  sky130_fd_sc_hd__nand3_1 U19039 ( .A(n12990), .B(n23269), .C(n26878), .Y(
        n12356) );
  sky130_fd_sc_hd__nand3_2 U19040 ( .A(n12990), .B(n23269), .C(n26878), .Y(
        n25875) );
  sky130_fd_sc_hd__nand2_1 U19041 ( .A(n10976), .B(n11124), .Y(n12358) );
  sky130_fd_sc_hd__nand2_1 U19042 ( .A(n10976), .B(n11124), .Y(n12497) );
  sky130_fd_sc_hd__nor2_1 U19043 ( .A(n12972), .B(n12970), .Y(n12360) );
  sky130_fd_sc_hd__nand4_1 U19044 ( .A(n13050), .B(n13043), .C(n13044), .D(
        n23160), .Y(n12361) );
  sky130_fd_sc_hd__buf_8 U19046 ( .A(n11122), .X(n12412) );
  sky130_fd_sc_hd__o2bb2ai_1 U19047 ( .B1(n23178), .B2(n12468), .A1_N(n11137), 
        .A2_N(n24629), .Y(j202_soc_core_j22_cpu_rf_N3067) );
  sky130_fd_sc_hd__buf_6 U19048 ( .A(n24175), .X(n29254) );
  sky130_fd_sc_hd__o2bb2ai_1 U19049 ( .B1(n27212), .B2(n25707), .A1_N(n23106), 
        .A2_N(n24629), .Y(j202_soc_core_j22_cpu_rf_N2808) );
  sky130_fd_sc_hd__o2bb2ai_1 U19050 ( .B1(n27220), .B2(n12468), .A1_N(n11136), 
        .A2_N(n24629), .Y(j202_soc_core_j22_cpu_rf_N2882) );
  sky130_fd_sc_hd__buf_4 U19051 ( .A(n17390), .X(n18370) );
  sky130_fd_sc_hd__nand2_1 U19052 ( .A(n17388), .B(n17387), .Y(n17973) );
  sky130_fd_sc_hd__buf_4 U19054 ( .A(n17406), .X(n12367) );
  sky130_fd_sc_hd__buf_4 U19055 ( .A(j202_soc_core_j22_cpu_ml_bufa[3]), .X(
        n24132) );
  sky130_fd_sc_hd__a21o_1 U19056 ( .A1(n18470), .A2(n12367), .B1(n18468), .X(
        n18487) );
  sky130_fd_sc_hd__nand2b_1 U19057 ( .A_N(n24353), .B(n27683), .Y(n24347) );
  sky130_fd_sc_hd__nand2_1 U19059 ( .A(j202_soc_core_memory0_ram_dout0[476]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12369) );
  sky130_fd_sc_hd__o211ai_1 U19060 ( .A1(n11153), .A2(n12988), .B1(n12987), 
        .C1(n12984), .Y(n22718) );
  sky130_fd_sc_hd__nor2_1 U19061 ( .A(n12985), .B(n12986), .Y(n12984) );
  sky130_fd_sc_hd__nand4_1 U19062 ( .A(n13254), .B(n16629), .C(n13251), .D(
        n12369), .Y(n12370) );
  sky130_fd_sc_hd__nand2_1 U19063 ( .A(n26443), .B(n12371), .Y(n12372) );
  sky130_fd_sc_hd__nand2_1 U19064 ( .A(n26323), .B(n12374), .Y(n12373) );
  sky130_fd_sc_hd__nand2_1 U19065 ( .A(n12622), .B(n11124), .Y(n12375) );
  sky130_fd_sc_hd__nor2_1 U19066 ( .A(n15278), .B(n15279), .Y(n12379) );
  sky130_fd_sc_hd__nor2_1 U19067 ( .A(n15278), .B(n15279), .Y(n13151) );
  sky130_fd_sc_hd__nor2_1 U19068 ( .A(n13161), .B(n27561), .Y(n13160) );
  sky130_fd_sc_hd__inv_2 U19069 ( .A(n13180), .Y(n13011) );
  sky130_fd_sc_hd__nand3_1 U19070 ( .A(n12940), .B(n12352), .C(n12937), .Y(
        n12936) );
  sky130_fd_sc_hd__nand2_1 U19071 ( .A(n12438), .B(n23803), .Y(n12380) );
  sky130_fd_sc_hd__nand2_2 U19072 ( .A(n26825), .B(n19697), .Y(n26824) );
  sky130_fd_sc_hd__fah_1 U19074 ( .A(n18051), .B(n18050), .CI(n18049), .COUT(
        n18160), .SUM(n18035) );
  sky130_fd_sc_hd__nand2_1 U19075 ( .A(n23233), .B(n26862), .Y(n25665) );
  sky130_fd_sc_hd__nand2_1 U19076 ( .A(n12840), .B(n23920), .Y(n26606) );
  sky130_fd_sc_hd__nand3_1 U19078 ( .A(n27779), .B(n27780), .C(n27778), .Y(
        n27784) );
  sky130_fd_sc_hd__nand3_1 U19079 ( .A(n24341), .B(n27892), .C(n24309), .Y(
        n27783) );
  sky130_fd_sc_hd__a21boi_1 U19080 ( .A1(n27558), .A2(n24355), .B1_N(n12388), 
        .Y(n24356) );
  sky130_fd_sc_hd__nand2_1 U19081 ( .A(n11135), .B(n21813), .Y(n21522) );
  sky130_fd_sc_hd__nor2_1 U19083 ( .A(n24446), .B(n12114), .Y(n12390) );
  sky130_fd_sc_hd__nor2_1 U19084 ( .A(n24446), .B(n12842), .Y(n27965) );
  sky130_fd_sc_hd__inv_2 U19086 ( .A(n26105), .Y(n12391) );
  sky130_fd_sc_hd__inv_2 U19087 ( .A(n26105), .Y(n12392) );
  sky130_fd_sc_hd__nand3_1 U19089 ( .A(n22706), .B(n22705), .C(n22704), .Y(
        n28996) );
  sky130_fd_sc_hd__nand3_1 U19090 ( .A(n27884), .B(n27885), .C(n12288), .Y(
        n12597) );
  sky130_fd_sc_hd__or2_0 U19091 ( .A(n27333), .B(n27461), .X(n12396) );
  sky130_fd_sc_hd__nand2_1 U19092 ( .A(n12396), .B(n24553), .Y(
        j202_soc_core_j22_cpu_rf_N3062) );
  sky130_fd_sc_hd__a22oi_2 U19093 ( .A1(j202_soc_core_memory0_ram_dout0[163]), 
        .A2(n21590), .B1(n21732), .B2(j202_soc_core_memory0_ram_dout0[195]), 
        .Y(n19936) );
  sky130_fd_sc_hd__nor2_1 U19094 ( .A(n12361), .B(n24298), .Y(n12397) );
  sky130_fd_sc_hd__fah_1 U19095 ( .A(n18350), .B(n18349), .CI(n18348), .COUT(
        n18393), .SUM(n18584) );
  sky130_fd_sc_hd__nor2_1 U19096 ( .A(n27791), .B(n27792), .Y(n27939) );
  sky130_fd_sc_hd__nand2_1 U19097 ( .A(n29328), .B(n22715), .Y(n19408) );
  sky130_fd_sc_hd__o21a_1 U19098 ( .A1(n24122), .A2(n12456), .B1(n24121), .X(
        n12398) );
  sky130_fd_sc_hd__nand2_1 U19099 ( .A(n12398), .B(n24120), .Y(
        j202_soc_core_ahb2aqu_00_N161) );
  sky130_fd_sc_hd__inv_1 U19100 ( .A(n12627), .Y(n12456) );
  sky130_fd_sc_hd__nand2_1 U19101 ( .A(n12959), .B(n12360), .Y(n12414) );
  sky130_fd_sc_hd__nand2_1 U19102 ( .A(n20710), .B(n20709), .Y(n26526) );
  sky130_fd_sc_hd__a21oi_1 U19103 ( .A1(n12510), .A2(n17004), .B1(n17003), .Y(
        n24124) );
  sky130_fd_sc_hd__nand2_1 U19104 ( .A(n11936), .B(n25108), .Y(n23305) );
  sky130_fd_sc_hd__a22oi_2 U19105 ( .A1(j202_soc_core_memory0_ram_dout0[83]), 
        .A2(n21734), .B1(n21732), .B2(j202_soc_core_memory0_ram_dout0[211]), 
        .Y(n15755) );
  sky130_fd_sc_hd__o31ai_2 U19106 ( .A1(n28590), .A2(n26242), .A3(n23441), 
        .B1(n23442), .Y(n29240) );
  sky130_fd_sc_hd__a22oi_2 U19107 ( .A1(j202_soc_core_memory0_ram_dout0[260]), 
        .A2(n21605), .B1(n21735), .B2(j202_soc_core_memory0_ram_dout0[228]), 
        .Y(n19333) );
  sky130_fd_sc_hd__a22oi_2 U19109 ( .A1(j202_soc_core_memory0_ram_dout0[4]), 
        .A2(n21733), .B1(n21592), .B2(j202_soc_core_memory0_ram_dout0[132]), 
        .Y(n19331) );
  sky130_fd_sc_hd__inv_2 U19110 ( .A(n12676), .Y(n12417) );
  sky130_fd_sc_hd__nand2_1 U19111 ( .A(n12624), .B(n11124), .Y(n12418) );
  sky130_fd_sc_hd__nand2_1 U19112 ( .A(n12624), .B(n11124), .Y(n29233) );
  sky130_fd_sc_hd__nand4_1 U19113 ( .A(n29500), .B(n12379), .C(n13147), .D(
        n13150), .Y(n12419) );
  sky130_fd_sc_hd__a21oi_1 U19114 ( .A1(n25047), .A2(n26722), .B1(n25046), .Y(
        n12420) );
  sky130_fd_sc_hd__nor2_1 U19115 ( .A(n25273), .B(n25269), .Y(n12422) );
  sky130_fd_sc_hd__nor2_1 U19116 ( .A(n24326), .B(n12424), .Y(n24330) );
  sky130_fd_sc_hd__nand2_1 U19117 ( .A(n19169), .B(n23011), .Y(n19170) );
  sky130_fd_sc_hd__inv_2 U19118 ( .A(n12435), .Y(n26470) );
  sky130_fd_sc_hd__nand4_1 U19119 ( .A(n23155), .B(n23156), .C(n22282), .D(
        n23154), .Y(n13083) );
  sky130_fd_sc_hd__nand3_1 U19120 ( .A(n23163), .B(n13078), .C(n13273), .Y(
        n12912) );
  sky130_fd_sc_hd__nand2_1 U19121 ( .A(n15275), .B(n12285), .Y(n15279) );
  sky130_fd_sc_hd__nand2_2 U19122 ( .A(n12915), .B(n12247), .Y(n28960) );
  sky130_fd_sc_hd__nand2_1 U19124 ( .A(n18256), .B(n18255), .Y(n12442) );
  sky130_fd_sc_hd__nand2_1 U19125 ( .A(n12440), .B(n12441), .Y(n12443) );
  sky130_fd_sc_hd__nand2_1 U19126 ( .A(n12442), .B(n12443), .Y(n18257) );
  sky130_fd_sc_hd__nand2_1 U19127 ( .A(n18267), .B(n18266), .Y(n12446) );
  sky130_fd_sc_hd__nand2_1 U19128 ( .A(n12444), .B(n12445), .Y(n12447) );
  sky130_fd_sc_hd__nand2_1 U19129 ( .A(n12446), .B(n12447), .Y(n18284) );
  sky130_fd_sc_hd__xnor2_1 U19130 ( .A(n18258), .B(n18257), .Y(n18264) );
  sky130_fd_sc_hd__nand2_1 U19131 ( .A(n20988), .B(n20987), .Y(n26536) );
  sky130_fd_sc_hd__nor2_1 U19132 ( .A(n13259), .B(n12503), .Y(n21914) );
  sky130_fd_sc_hd__nand3_1 U19133 ( .A(n12414), .B(n21814), .C(n21776), .Y(
        n12448) );
  sky130_fd_sc_hd__nand3_2 U19134 ( .A(n21817), .B(n21816), .C(n21815), .Y(
        n26912) );
  sky130_fd_sc_hd__inv_2 U19136 ( .A(n26912), .Y(n27417) );
  sky130_fd_sc_hd__mux2_2 U19137 ( .A0(n19756), .A1(n19755), .S(n26824), .X(
        n19788) );
  sky130_fd_sc_hd__mux2_2 U19138 ( .A0(n19699), .A1(n19698), .S(n26824), .X(
        n19743) );
  sky130_fd_sc_hd__nand2_1 U19139 ( .A(n23735), .B(n26539), .Y(n12689) );
  sky130_fd_sc_hd__nor2_1 U19140 ( .A(n13193), .B(n27231), .Y(n27233) );
  sky130_fd_sc_hd__clkbuf_1 U19141 ( .A(n27881), .X(n12679) );
  sky130_fd_sc_hd__nor2_1 U19142 ( .A(n24423), .B(n27881), .Y(n13049) );
  sky130_fd_sc_hd__nand2_1 U19143 ( .A(n13011), .B(n29070), .Y(n13051) );
  sky130_fd_sc_hd__o21a_1 U19144 ( .A1(n23920), .A2(n12840), .B1(n24785), .X(
        n12452) );
  sky130_fd_sc_hd__nand2_1 U19145 ( .A(n12452), .B(n19170), .Y(n19197) );
  sky130_fd_sc_hd__buf_6 U19147 ( .A(n12133), .X(n17786) );
  sky130_fd_sc_hd__nand2_1 U19148 ( .A(n12454), .B(n18990), .Y(n19039) );
  sky130_fd_sc_hd__nand3_1 U19149 ( .A(n12258), .B(n14380), .C(n14379), .Y(
        n26729) );
  sky130_fd_sc_hd__nand3_1 U19150 ( .A(n21366), .B(n21365), .C(n21364), .Y(
        n28948) );
  sky130_fd_sc_hd__clkbuf_1 U19151 ( .A(n24360), .X(n12461) );
  sky130_fd_sc_hd__nor2_2 U19152 ( .A(n28975), .B(n12879), .Y(n12462) );
  sky130_fd_sc_hd__nand3_1 U19153 ( .A(n24381), .B(n24382), .C(n24380), .Y(
        n24384) );
  sky130_fd_sc_hd__nand2_1 U19155 ( .A(n12640), .B(n23209), .Y(n12466) );
  sky130_fd_sc_hd__o2bb2ai_1 U19156 ( .B1(n23178), .B2(n11047), .A1_N(n11137), 
        .A2_N(n11612), .Y(j202_soc_core_j22_cpu_rf_N3081) );
  sky130_fd_sc_hd__o21ai_1 U19158 ( .A1(n17125), .A2(n26538), .B1(n16830), .Y(
        n12465) );
  sky130_fd_sc_hd__o2bb2ai_1 U19159 ( .B1(n27209), .B2(n27359), .A1_N(n26360), 
        .A2_N(n24497), .Y(j202_soc_core_j22_cpu_rf_N2749) );
  sky130_fd_sc_hd__nor2_1 U19160 ( .A(n12825), .B(n12820), .Y(n12819) );
  sky130_fd_sc_hd__nand3_1 U19161 ( .A(n12880), .B(n13236), .C(n12482), .Y(
        n12467) );
  sky130_fd_sc_hd__inv_2 U19162 ( .A(n25705), .Y(n12468) );
  sky130_fd_sc_hd__and2_1 U19164 ( .A(n25705), .B(n26450), .X(n13334) );
  sky130_fd_sc_hd__nor2_1 U19165 ( .A(n12836), .B(n12831), .Y(n12830) );
  sky130_fd_sc_hd__inv_2 U19166 ( .A(n23140), .Y(n12732) );
  sky130_fd_sc_hd__nand3_2 U19167 ( .A(n12436), .B(n11873), .C(n13116), .Y(
        n12744) );
  sky130_fd_sc_hd__o22ai_1 U19168 ( .A1(n18660), .A2(n17976), .B1(n17975), 
        .B2(n12991), .Y(n18005) );
  sky130_fd_sc_hd__o22ai_1 U19169 ( .A1(n18660), .A2(n18659), .B1(n12991), 
        .B2(n18658), .Y(n18695) );
  sky130_fd_sc_hd__o2bb2ai_1 U19170 ( .B1(n26898), .B2(n11047), .A1_N(n11612), 
        .A2_N(n12469), .Y(j202_soc_core_j22_cpu_rf_N3341) );
  sky130_fd_sc_hd__a21o_1 U19171 ( .A1(n17402), .A2(n18344), .B1(n18343), .X(
        n18390) );
  sky130_fd_sc_hd__inv_2 U19173 ( .A(n26881), .Y(n12478) );
  sky130_fd_sc_hd__inv_2 U19174 ( .A(n26881), .Y(n23944) );
  sky130_fd_sc_hd__clkbuf_1 U19175 ( .A(n21875), .X(n12578) );
  sky130_fd_sc_hd__buf_2 U19176 ( .A(j202_soc_core_j22_cpu_ml_bufa[13]), .X(
        n17400) );
  sky130_fd_sc_hd__nand3_2 U19178 ( .A(n13198), .B(n13199), .C(n21753), .Y(
        n29072) );
  sky130_fd_sc_hd__nor2_2 U19179 ( .A(n24447), .B(n23566), .Y(n13044) );
  sky130_fd_sc_hd__inv_1 U19180 ( .A(n12450), .Y(n24335) );
  sky130_fd_sc_hd__fah_1 U19181 ( .A(n18100), .B(n18099), .CI(n18098), .COUT(
        n18162), .SUM(n18121) );
  sky130_fd_sc_hd__nor2_2 U19182 ( .A(n17819), .B(n17820), .Y(n21385) );
  sky130_fd_sc_hd__nand2_1 U19183 ( .A(n20146), .B(n12220), .Y(n18983) );
  sky130_fd_sc_hd__and3_1 U19184 ( .A(n18979), .B(
        j202_soc_core_j22_cpu_ma_M_MEM[1]), .C(
        j202_soc_core_j22_cpu_ma_M_address[1]), .X(n22715) );
  sky130_fd_sc_hd__nand3_1 U19185 ( .A(n12675), .B(n26422), .C(n12674), .Y(
        n21918) );
  sky130_fd_sc_hd__nand3_1 U19186 ( .A(n23145), .B(n27564), .C(n23146), .Y(
        n24447) );
  sky130_fd_sc_hd__nand3_2 U19187 ( .A(n12670), .B(n19408), .C(n19409), .Y(
        n27421) );
  sky130_fd_sc_hd__nand2b_1 U19188 ( .A_N(n18353), .B(n21887), .Y(n17586) );
  sky130_fd_sc_hd__o211ai_1 U19189 ( .A1(n22662), .A2(n22897), .B1(n12773), 
        .C1(n12280), .Y(n22663) );
  sky130_fd_sc_hd__o21ai_1 U19190 ( .A1(n22193), .A2(n22897), .B1(n22192), .Y(
        n22194) );
  sky130_fd_sc_hd__nand3_1 U19191 ( .A(n23953), .B(n12598), .C(n13268), .Y(
        n13273) );
  sky130_fd_sc_hd__nor2_1 U19192 ( .A(n13250), .B(n12370), .Y(n12490) );
  sky130_fd_sc_hd__nor2_1 U19193 ( .A(n13250), .B(n13249), .Y(n20966) );
  sky130_fd_sc_hd__nand3_1 U19194 ( .A(n26315), .B(n23765), .C(n23764), .Y(
        n27382) );
  sky130_fd_sc_hd__nand2_2 U19195 ( .A(n26315), .B(n26555), .Y(n27371) );
  sky130_fd_sc_hd__nand2_2 U19196 ( .A(n26315), .B(n26551), .Y(n27364) );
  sky130_fd_sc_hd__nand3_1 U19197 ( .A(n25143), .B(n22686), .C(n25142), .Y(
        n23010) );
  sky130_fd_sc_hd__a21oi_1 U19198 ( .A1(n22398), .A2(n22189), .B1(n22188), .Y(
        n22798) );
  sky130_fd_sc_hd__o2bb2ai_1 U19199 ( .B1(n27575), .B2(n24546), .A1_N(n11109), 
        .A2_N(n12435), .Y(j202_soc_core_j22_cpu_rf_N3107) );
  sky130_fd_sc_hd__o21a_1 U19200 ( .A1(n26951), .A2(n25293), .B1(n25292), .X(
        n25294) );
  sky130_fd_sc_hd__clkbuf_1 U19201 ( .A(n12486), .X(n12742) );
  sky130_fd_sc_hd__nor2_1 U19202 ( .A(n12553), .B(n12552), .Y(n12551) );
  sky130_fd_sc_hd__nor2_1 U19203 ( .A(n13247), .B(n13244), .Y(n20965) );
  sky130_fd_sc_hd__nand2_1 U19204 ( .A(n13257), .B(n13256), .Y(n13244) );
  sky130_fd_sc_hd__inv_1 U19205 ( .A(n11124), .Y(n12494) );
  sky130_fd_sc_hd__nand2b_4 U19206 ( .A_N(n23157), .B(n27898), .Y(n24455) );
  sky130_fd_sc_hd__nand2_1 U19207 ( .A(n24417), .B(n12804), .Y(n23607) );
  sky130_fd_sc_hd__o21a_1 U19208 ( .A1(n26951), .A2(n24689), .B1(n24688), .X(
        n24690) );
  sky130_fd_sc_hd__nand2_1 U19209 ( .A(n21384), .B(n13141), .Y(n13145) );
  sky130_fd_sc_hd__fah_1 U19210 ( .A(n18193), .B(n18192), .CI(n18191), .COUT(
        n18245), .SUM(n18208) );
  sky130_fd_sc_hd__o22ai_1 U19211 ( .A1(n26707), .A2(n11153), .B1(n24778), 
        .B2(n23013), .Y(n12495) );
  sky130_fd_sc_hd__o21a_1 U19212 ( .A1(n26951), .A2(n25557), .B1(n25556), .X(
        n25558) );
  sky130_fd_sc_hd__inv_6 U19213 ( .A(n29249), .Y(n12537) );
  sky130_fd_sc_hd__a22oi_2 U19214 ( .A1(j202_soc_core_memory0_ram_dout0[100]), 
        .A2(n21591), .B1(n21590), .B2(j202_soc_core_memory0_ram_dout0[164]), 
        .Y(n19330) );
  sky130_fd_sc_hd__nor2_1 U19215 ( .A(n13267), .B(n13266), .Y(n21769) );
  sky130_fd_sc_hd__a21o_1 U19216 ( .A1(n22969), .A2(n22609), .B1(n22608), .X(
        n12500) );
  sky130_fd_sc_hd__o22ai_1 U19217 ( .A1(n25219), .A2(n17389), .B1(n22141), 
        .B2(n18307), .Y(n17514) );
  sky130_fd_sc_hd__o22ai_1 U19218 ( .A1(n25219), .A2(n18308), .B1(n22628), 
        .B2(n18307), .Y(n18556) );
  sky130_fd_sc_hd__nand2_2 U19220 ( .A(n17401), .B(n18112), .Y(n17402) );
  sky130_fd_sc_hd__o2bb2ai_1 U19221 ( .B1(n27224), .B2(n26915), .A1_N(n12504), 
        .A2_N(n27224), .Y(j202_soc_core_j22_cpu_rf_N2942) );
  sky130_fd_sc_hd__nand2b_1 U19222 ( .A_N(n24353), .B(n24351), .Y(n27171) );
  sky130_fd_sc_hd__o2bb2ai_1 U19223 ( .B1(n27210), .B2(n26915), .A1_N(n12504), 
        .A2_N(n27210), .Y(j202_soc_core_j22_cpu_rf_N3201) );
  sky130_fd_sc_hd__nor2_1 U19224 ( .A(n12548), .B(n12543), .Y(n12542) );
  sky130_fd_sc_hd__inv_6 U19226 ( .A(n12479), .Y(n12527) );
  sky130_fd_sc_hd__nand2_1 U19228 ( .A(n27888), .B(n12881), .Y(n12513) );
  sky130_fd_sc_hd__nand2_1 U19229 ( .A(n27888), .B(n12881), .Y(n12514) );
  sky130_fd_sc_hd__nand2_1 U19230 ( .A(n12466), .B(n12881), .Y(n10584) );
  sky130_fd_sc_hd__nand2_1 U19231 ( .A(n12729), .B(n27683), .Y(n27895) );
  sky130_fd_sc_hd__nand2_2 U19233 ( .A(n12515), .B(n23180), .Y(n27892) );
  sky130_fd_sc_hd__a22oi_1 U19234 ( .A1(j202_soc_core_memory0_ram_dout0[115]), 
        .A2(n21591), .B1(n21598), .B2(j202_soc_core_memory0_ram_dout0[435]), 
        .Y(n15754) );
  sky130_fd_sc_hd__inv_6 U19236 ( .A(n29249), .Y(n12535) );
  sky130_fd_sc_hd__inv_6 U19237 ( .A(n29249), .Y(n12536) );
  sky130_fd_sc_hd__inv_6 U19238 ( .A(n12479), .Y(n12528) );
  sky130_fd_sc_hd__inv_6 U19239 ( .A(n12479), .Y(n12526) );
  sky130_fd_sc_hd__inv_6 U19240 ( .A(n29248), .Y(n12522) );
  sky130_fd_sc_hd__inv_6 U19241 ( .A(n29248), .Y(n12523) );
  sky130_fd_sc_hd__inv_6 U19242 ( .A(n29248), .Y(n12529) );
  sky130_fd_sc_hd__inv_6 U19243 ( .A(n29248), .Y(n12530) );
  sky130_fd_sc_hd__nand2_1 U19244 ( .A(n20972), .B(n12229), .Y(n20976) );
  sky130_fd_sc_hd__nand2_1 U19245 ( .A(n12542), .B(n12551), .Y(n21340) );
  sky130_fd_sc_hd__nand4_1 U19246 ( .A(n12547), .B(n12546), .C(n12545), .D(
        n12544), .Y(n12543) );
  sky130_fd_sc_hd__nand2_1 U19247 ( .A(j202_soc_core_memory0_ram_dout0[205]), 
        .B(n21732), .Y(n12544) );
  sky130_fd_sc_hd__nand2_1 U19248 ( .A(j202_soc_core_memory0_ram_dout0[237]), 
        .B(n21735), .Y(n12545) );
  sky130_fd_sc_hd__nand2_1 U19249 ( .A(j202_soc_core_memory0_ram_dout0[141]), 
        .B(n21592), .Y(n12546) );
  sky130_fd_sc_hd__nand2_1 U19250 ( .A(j202_soc_core_memory0_ram_dout0[173]), 
        .B(n21590), .Y(n12547) );
  sky130_fd_sc_hd__nand4_1 U19251 ( .A(n21295), .B(n12550), .C(n21168), .D(
        n12549), .Y(n12548) );
  sky130_fd_sc_hd__nand2_1 U19252 ( .A(j202_soc_core_memory0_ram_dout0[109]), 
        .B(n21591), .Y(n12549) );
  sky130_fd_sc_hd__nand2_1 U19253 ( .A(j202_soc_core_memory0_ram_dout0[77]), 
        .B(n21734), .Y(n12550) );
  sky130_fd_sc_hd__nand4_1 U19254 ( .A(n21298), .B(n21296), .C(n21297), .D(
        n21167), .Y(n12552) );
  sky130_fd_sc_hd__nand4_1 U19255 ( .A(n13225), .B(n12648), .C(n12594), .D(
        n12554), .Y(n12553) );
  sky130_fd_sc_hd__and3_1 U19256 ( .A(n21294), .B(n21312), .C(n21313), .X(
        n12554) );
  sky130_fd_sc_hd__nor2_1 U19257 ( .A(n11105), .B(n12556), .Y(n12555) );
  sky130_fd_sc_hd__nand2_1 U19259 ( .A(n27553), .B(n29015), .Y(n12559) );
  sky130_fd_sc_hd__nand2_1 U19260 ( .A(n12562), .B(n12561), .Y(n18203) );
  sky130_fd_sc_hd__nand2_1 U19261 ( .A(n12564), .B(n18202), .Y(n12561) );
  sky130_fd_sc_hd__o21ai_1 U19262 ( .A1(n18202), .A2(n12564), .B1(n18201), .Y(
        n12562) );
  sky130_fd_sc_hd__xor2_1 U19263 ( .A(n12563), .B(n18201), .X(n18210) );
  sky130_fd_sc_hd__xor2_1 U19264 ( .A(n18202), .B(n12564), .X(n12563) );
  sky130_fd_sc_hd__nand2b_1 U19265 ( .A_N(n18153), .B(n12565), .Y(n12564) );
  sky130_fd_sc_hd__xnor2_1 U19266 ( .A(n12566), .B(n18571), .Y(n18592) );
  sky130_fd_sc_hd__xnor2_1 U19267 ( .A(n18572), .B(n18573), .Y(n12566) );
  sky130_fd_sc_hd__nand2_1 U19268 ( .A(n12610), .B(n18574), .Y(n12609) );
  sky130_fd_sc_hd__nand2_1 U19269 ( .A(n12568), .B(n12567), .Y(n18574) );
  sky130_fd_sc_hd__nand2_1 U19270 ( .A(n18572), .B(n18573), .Y(n12567) );
  sky130_fd_sc_hd__o21ai_1 U19271 ( .A1(n18572), .A2(n18573), .B1(n18571), .Y(
        n12568) );
  sky130_fd_sc_hd__inv_1 U19272 ( .A(n24308), .Y(n24341) );
  sky130_fd_sc_hd__nand2_1 U19273 ( .A(n12571), .B(n12570), .Y(n17495) );
  sky130_fd_sc_hd__nand2_1 U19274 ( .A(n17522), .B(n17523), .Y(n12570) );
  sky130_fd_sc_hd__nand2_1 U19276 ( .A(n12574), .B(n12573), .Y(n17570) );
  sky130_fd_sc_hd__nand2_1 U19277 ( .A(n17573), .B(n17574), .Y(n12573) );
  sky130_fd_sc_hd__o21ai_1 U19278 ( .A1(n17574), .A2(n17573), .B1(n17572), .Y(
        n12574) );
  sky130_fd_sc_hd__inv_2 U19279 ( .A(n17574), .Y(n12575) );
  sky130_fd_sc_hd__a22oi_2 U19280 ( .A1(j202_soc_core_memory0_ram_dout0[168]), 
        .A2(n21590), .B1(n21732), .B2(j202_soc_core_memory0_ram_dout0[200]), 
        .Y(n20406) );
  sky130_fd_sc_hd__xnor2_1 U19281 ( .A(n18610), .B(n12576), .Y(n18811) );
  sky130_fd_sc_hd__xnor2_1 U19282 ( .A(n18608), .B(n18609), .Y(n12576) );
  sky130_fd_sc_hd__clkbuf_1 U19283 ( .A(n22835), .X(n12579) );
  sky130_fd_sc_hd__nand3b_1 U19285 ( .A_N(n12582), .B(n23946), .C(n23945), .Y(
        j202_soc_core_j22_cpu_ml_maclj[12]) );
  sky130_fd_sc_hd__nand3b_1 U19286 ( .A_N(n12583), .B(n23971), .C(n23970), .Y(
        j202_soc_core_j22_cpu_ml_maclj[11]) );
  sky130_fd_sc_hd__nand2b_1 U19287 ( .A_N(n17454), .B(n12584), .Y(n17475) );
  sky130_fd_sc_hd__inv_1 U19288 ( .A(n17436), .Y(n12585) );
  sky130_fd_sc_hd__nand2b_1 U19289 ( .A_N(n17437), .B(n12585), .Y(n17434) );
  sky130_fd_sc_hd__nor2_1 U19290 ( .A(n18283), .B(n18284), .Y(n21878) );
  sky130_fd_sc_hd__nor2_1 U19291 ( .A(n12851), .B(n12852), .Y(n12850) );
  sky130_fd_sc_hd__a22oi_2 U19292 ( .A1(j202_soc_core_memory0_ram_dout0[360]), 
        .A2(n21596), .B1(j202_soc_core_memory0_ram_dout0_sel[14]), .B2(
        j202_soc_core_memory0_ram_dout0[456]), .Y(n20405) );
  sky130_fd_sc_hd__o22ai_1 U19293 ( .A1(n23144), .A2(n13076), .B1(n23210), 
        .B2(n13236), .Y(n13079) );
  sky130_fd_sc_hd__nand2_1 U19294 ( .A(j202_soc_core_memory0_ram_dout0[135]), 
        .B(n21592), .Y(n12589) );
  sky130_fd_sc_hd__nand2_1 U19295 ( .A(n12590), .B(n27970), .Y(n27923) );
  sky130_fd_sc_hd__nand2_1 U19296 ( .A(n27903), .B(n12284), .Y(n12590) );
  sky130_fd_sc_hd__inv_2 U19297 ( .A(n27045), .Y(n26581) );
  sky130_fd_sc_hd__o2bb2ai_1 U19298 ( .B1(n27333), .B2(n24546), .A1_N(n26371), 
        .A2_N(n12435), .Y(j202_soc_core_j22_cpu_rf_N3070) );
  sky130_fd_sc_hd__clkbuf_1 U19299 ( .A(j202_soc_core_j22_cpu_ml_bufa[24]), 
        .X(n24583) );
  sky130_fd_sc_hd__nor2_1 U19301 ( .A(n18290), .B(n19481), .Y(n18268) );
  sky130_fd_sc_hd__inv_1 U19302 ( .A(n13098), .Y(n13097) );
  sky130_fd_sc_hd__nand2_1 U19303 ( .A(n27522), .B(n12290), .Y(n10492) );
  sky130_fd_sc_hd__clkbuf_1 U19304 ( .A(n24712), .X(n12591) );
  sky130_fd_sc_hd__nand2_1 U19305 ( .A(n27964), .B(n24091), .Y(n24092) );
  sky130_fd_sc_hd__or2_0 U19306 ( .A(n18916), .B(n24159), .X(n12592) );
  sky130_fd_sc_hd__nor2_1 U19307 ( .A(n29577), .B(n12439), .Y(n12883) );
  sky130_fd_sc_hd__nand2_1 U19308 ( .A(j202_soc_core_memory0_ram_dout0[301]), 
        .B(n21603), .Y(n12594) );
  sky130_fd_sc_hd__a21oi_1 U19309 ( .A1(n13301), .A2(n22721), .B1(n17817), .Y(
        n19173) );
  sky130_fd_sc_hd__nand2_1 U19310 ( .A(n12790), .B(n12791), .Y(n13301) );
  sky130_fd_sc_hd__and2_0 U19311 ( .A(n23942), .B(n23941), .X(n12596) );
  sky130_fd_sc_hd__nand2_1 U19312 ( .A(n12597), .B(n27980), .Y(n27887) );
  sky130_fd_sc_hd__o21ai_2 U19313 ( .A1(n17869), .A2(n19241), .B1(n17868), .Y(
        n19463) );
  sky130_fd_sc_hd__clkbuf_1 U19314 ( .A(n21516), .X(n12599) );
  sky130_fd_sc_hd__nand3_2 U19315 ( .A(n22272), .B(n22273), .C(n27230), .Y(
        n23211) );
  sky130_fd_sc_hd__xnor2_1 U19316 ( .A(n18078), .B(n18079), .Y(n18080) );
  sky130_fd_sc_hd__nand3_1 U19317 ( .A(n23948), .B(n12602), .C(n12600), .Y(
        j202_soc_core_j22_cpu_ml_maclj[14]) );
  sky130_fd_sc_hd__inv_1 U19318 ( .A(n12601), .Y(n12600) );
  sky130_fd_sc_hd__nor2_1 U19319 ( .A(n23949), .B(n12918), .Y(n12601) );
  sky130_fd_sc_hd__nor2_1 U19320 ( .A(n12300), .B(n26976), .Y(n12602) );
  sky130_fd_sc_hd__nand2_1 U19321 ( .A(n12604), .B(n12603), .Y(n17704) );
  sky130_fd_sc_hd__nand2_1 U19322 ( .A(n17701), .B(n17702), .Y(n12603) );
  sky130_fd_sc_hd__nand2_1 U19323 ( .A(n17700), .B(n12605), .Y(n12604) );
  sky130_fd_sc_hd__nand2b_1 U19324 ( .A_N(n17701), .B(n12607), .Y(n12605) );
  sky130_fd_sc_hd__xor2_1 U19325 ( .A(n12606), .B(n17700), .X(n17885) );
  sky130_fd_sc_hd__xnor2_1 U19326 ( .A(n12607), .B(n17701), .Y(n12606) );
  sky130_fd_sc_hd__inv_1 U19327 ( .A(n13093), .Y(n13092) );
  sky130_fd_sc_hd__nand2_1 U19328 ( .A(n13205), .B(n13204), .Y(n18810) );
  sky130_fd_sc_hd__nand2_1 U19329 ( .A(n12609), .B(n12608), .Y(n18608) );
  sky130_fd_sc_hd__nand2_1 U19330 ( .A(n18575), .B(n18576), .Y(n12608) );
  sky130_fd_sc_hd__nand2b_1 U19331 ( .A_N(n18575), .B(n12611), .Y(n12610) );
  sky130_fd_sc_hd__xnor2_1 U19332 ( .A(n12612), .B(n18574), .Y(n18593) );
  sky130_fd_sc_hd__xnor2_1 U19333 ( .A(n18576), .B(n18575), .Y(n12612) );
  sky130_fd_sc_hd__a21oi_2 U19334 ( .A1(n18816), .A2(n22754), .B1(n18815), .Y(
        n19247) );
  sky130_fd_sc_hd__clkbuf_1 U19335 ( .A(j202_soc_core_j22_cpu_ml_bufa[0]), .X(
        n12613) );
  sky130_fd_sc_hd__nand3_2 U19336 ( .A(n22717), .B(n12989), .C(n12988), .Y(
        n27442) );
  sky130_fd_sc_hd__nor2_1 U19337 ( .A(n13135), .B(n13130), .Y(n13129) );
  sky130_fd_sc_hd__clkbuf_1 U19339 ( .A(n29053), .X(n12617) );
  sky130_fd_sc_hd__nand2_1 U19340 ( .A(n21447), .B(n12166), .Y(n18844) );
  sky130_fd_sc_hd__inv_1 U19341 ( .A(n18055), .Y(n18056) );
  sky130_fd_sc_hd__inv_1 U19342 ( .A(n13086), .Y(n13085) );
  sky130_fd_sc_hd__nand2_1 U19343 ( .A(j202_soc_core_memory0_ram_dout0[226]), 
        .B(n21735), .Y(n12620) );
  sky130_fd_sc_hd__nand2_2 U19345 ( .A(n12622), .B(n11124), .Y(n10585) );
  sky130_fd_sc_hd__nor2_4 U19346 ( .A(n22278), .B(n13152), .Y(n24265) );
  sky130_fd_sc_hd__inv_1 U19347 ( .A(n12864), .Y(n12863) );
  sky130_fd_sc_hd__nand2_1 U19348 ( .A(j202_soc_core_memory0_ram_dout0[71]), 
        .B(n21734), .Y(n12623) );
  sky130_fd_sc_hd__inv_1 U19349 ( .A(n12625), .Y(n13147) );
  sky130_fd_sc_hd__nand2_1 U19350 ( .A(n20833), .B(n20832), .Y(n23757) );
  sky130_fd_sc_hd__nor2_1 U19351 ( .A(n12849), .B(n12844), .Y(n12843) );
  sky130_fd_sc_hd__fah_1 U19352 ( .A(n18361), .B(n18360), .CI(n18359), .COUT(
        n18416), .SUM(n18356) );
  sky130_fd_sc_hd__clkbuf_1 U19353 ( .A(j202_soc_core_j22_cpu_ml_bufa[11]), 
        .X(n12630) );
  sky130_fd_sc_hd__nand2_1 U19354 ( .A(n12632), .B(n12631), .Y(n18830) );
  sky130_fd_sc_hd__nand2b_1 U19355 ( .A_N(n12636), .B(n18804), .Y(n12631) );
  sky130_fd_sc_hd__nand2_1 U19356 ( .A(n12633), .B(n18803), .Y(n12632) );
  sky130_fd_sc_hd__nand2_1 U19357 ( .A(n12636), .B(n12634), .Y(n12633) );
  sky130_fd_sc_hd__xor2_1 U19358 ( .A(n12636), .B(n12635), .X(n18828) );
  sky130_fd_sc_hd__xnor2_1 U19359 ( .A(n18804), .B(n18803), .Y(n12635) );
  sky130_fd_sc_hd__xor2_1 U19360 ( .A(n18799), .B(n12697), .X(n12636) );
  sky130_fd_sc_hd__nand2_1 U19361 ( .A(n12638), .B(n12637), .Y(n18741) );
  sky130_fd_sc_hd__nand2_1 U19362 ( .A(n18736), .B(n18737), .Y(n12637) );
  sky130_fd_sc_hd__o21ai_1 U19363 ( .A1(n18737), .A2(n18736), .B1(n18735), .Y(
        n12638) );
  sky130_fd_sc_hd__xnor2_1 U19364 ( .A(n18736), .B(n12639), .Y(n18798) );
  sky130_fd_sc_hd__xnor2_1 U19365 ( .A(n18737), .B(n18735), .Y(n12639) );
  sky130_fd_sc_hd__inv_1 U19366 ( .A(n12854), .Y(n12853) );
  sky130_fd_sc_hd__nand2_1 U19367 ( .A(n13068), .B(n26539), .Y(n12643) );
  sky130_fd_sc_hd__clkbuf_2 U19368 ( .A(n26550), .X(n12647) );
  sky130_fd_sc_hd__nand2_1 U19369 ( .A(j202_soc_core_memory0_ram_dout0[269]), 
        .B(n21605), .Y(n12648) );
  sky130_fd_sc_hd__nand2_1 U19370 ( .A(n12650), .B(n12649), .Y(n17876) );
  sky130_fd_sc_hd__nand2_1 U19371 ( .A(n17746), .B(n17747), .Y(n12649) );
  sky130_fd_sc_hd__nand2_1 U19372 ( .A(n17745), .B(n12651), .Y(n12650) );
  sky130_fd_sc_hd__nand2b_1 U19373 ( .A_N(n17746), .B(n12653), .Y(n12651) );
  sky130_fd_sc_hd__xor2_1 U19374 ( .A(n17745), .B(n12652), .X(n17763) );
  sky130_fd_sc_hd__xnor2_1 U19375 ( .A(n12653), .B(n17746), .Y(n12652) );
  sky130_fd_sc_hd__nand2_2 U19377 ( .A(n24094), .B(n12735), .Y(n27772) );
  sky130_fd_sc_hd__nand2_1 U19378 ( .A(n20719), .B(n11056), .Y(n20720) );
  sky130_fd_sc_hd__nand3_1 U19379 ( .A(n19937), .B(n19936), .C(n19935), .Y(
        n20719) );
  sky130_fd_sc_hd__nor2_1 U19380 ( .A(n12958), .B(n12956), .Y(n12955) );
  sky130_fd_sc_hd__nand3_2 U19381 ( .A(n23142), .B(n23586), .C(n29036), .Y(
        n27564) );
  sky130_fd_sc_hd__fah_1 U19382 ( .A(n17647), .B(n17646), .CI(n17645), .COUT(
        n17674), .SUM(n17701) );
  sky130_fd_sc_hd__nand2_1 U19384 ( .A(n12660), .B(n12659), .Y(n18560) );
  sky130_fd_sc_hd__nand2_1 U19385 ( .A(n18328), .B(n12661), .Y(n12659) );
  sky130_fd_sc_hd__o21ai_1 U19386 ( .A1(n12661), .A2(n18328), .B1(n18327), .Y(
        n12660) );
  sky130_fd_sc_hd__xor2_1 U19387 ( .A(n18328), .B(n12662), .X(n18552) );
  sky130_fd_sc_hd__xnor2_1 U19388 ( .A(n12663), .B(n18327), .Y(n12662) );
  sky130_fd_sc_hd__xnor2_1 U19389 ( .A(n18605), .B(n13328), .Y(n18607) );
  sky130_fd_sc_hd__nand2_1 U19390 ( .A(n18599), .B(n18600), .Y(n12664) );
  sky130_fd_sc_hd__nand2_1 U19391 ( .A(n22319), .B(n22320), .Y(n28999) );
  sky130_fd_sc_hd__nand2_1 U19392 ( .A(n23727), .B(n26539), .Y(n12666) );
  sky130_fd_sc_hd__nand3_1 U19393 ( .A(n12668), .B(n19414), .C(n12667), .Y(
        n19443) );
  sky130_fd_sc_hd__and2_1 U19394 ( .A(n26712), .B(n24785), .X(n12667) );
  sky130_fd_sc_hd__nand2_1 U19395 ( .A(n24592), .B(n12669), .Y(n12668) );
  sky130_fd_sc_hd__and3_1 U19396 ( .A(n26422), .B(n19412), .C(n19411), .X(
        n12669) );
  sky130_fd_sc_hd__nand2_1 U19398 ( .A(n19491), .B(n12672), .Y(n12671) );
  sky130_fd_sc_hd__o21a_1 U19399 ( .A1(n19492), .A2(n19493), .B1(n22929), .X(
        n12672) );
  sky130_fd_sc_hd__nand3_2 U19400 ( .A(n19448), .B(n24367), .C(n12673), .Y(
        n24591) );
  sky130_fd_sc_hd__nand2_1 U19401 ( .A(n27453), .B(n26323), .Y(n12674) );
  sky130_fd_sc_hd__nand2_1 U19402 ( .A(n12676), .B(n26443), .Y(n12675) );
  sky130_fd_sc_hd__inv_2 U19403 ( .A(n27453), .Y(n12676) );
  sky130_fd_sc_hd__o21ai_1 U19404 ( .A1(n19477), .A2(n22897), .B1(n19476), .Y(
        n19478) );
  sky130_fd_sc_hd__nor2_4 U19405 ( .A(n12745), .B(n12502), .Y(n22274) );
  sky130_fd_sc_hd__nor2_1 U19407 ( .A(n23239), .B(n23238), .Y(n12680) );
  sky130_fd_sc_hd__nand2_1 U19408 ( .A(n12682), .B(n12681), .Y(n18031) );
  sky130_fd_sc_hd__nand2_1 U19409 ( .A(n18010), .B(n18011), .Y(n12681) );
  sky130_fd_sc_hd__nand2_1 U19410 ( .A(n12687), .B(n12683), .Y(n12682) );
  sky130_fd_sc_hd__nand2_1 U19411 ( .A(n12685), .B(n12684), .Y(n12683) );
  sky130_fd_sc_hd__xnor2_1 U19412 ( .A(n12686), .B(n12687), .Y(n18075) );
  sky130_fd_sc_hd__xnor2_1 U19413 ( .A(n18011), .B(n18010), .Y(n12686) );
  sky130_fd_sc_hd__nand2_1 U19414 ( .A(n17996), .B(n17995), .Y(n12687) );
  sky130_fd_sc_hd__buf_4 U19416 ( .A(n12363), .X(n25223) );
  sky130_fd_sc_hd__nand2_1 U19417 ( .A(n24105), .B(n23210), .Y(n12884) );
  sky130_fd_sc_hd__and2_0 U19418 ( .A(n27602), .B(
        j202_soc_core_ahbcs_6__HREADY_), .X(n12691) );
  sky130_fd_sc_hd__nor2_1 U19419 ( .A(n13244), .B(n13245), .Y(n13243) );
  sky130_fd_sc_hd__nand2_2 U19420 ( .A(n23586), .B(n24265), .Y(n13194) );
  sky130_fd_sc_hd__o21a_1 U19421 ( .A1(n24332), .A2(n27956), .B1(n27176), .X(
        n12693) );
  sky130_fd_sc_hd__nand2_1 U19422 ( .A(n18799), .B(n18798), .Y(n12695) );
  sky130_fd_sc_hd__o21ai_1 U19423 ( .A1(n18798), .A2(n18799), .B1(n18797), .Y(
        n12696) );
  sky130_fd_sc_hd__xnor2_1 U19424 ( .A(n18798), .B(n18797), .Y(n12697) );
  sky130_fd_sc_hd__fah_1 U19425 ( .A(n18411), .B(n18412), .CI(n18413), .COUT(
        n18442), .SUM(n18435) );
  sky130_fd_sc_hd__xnor2_1 U19426 ( .A(n18439), .B(n12698), .Y(n18818) );
  sky130_fd_sc_hd__xnor2_1 U19427 ( .A(n18438), .B(n18437), .Y(n12698) );
  sky130_fd_sc_hd__nand2_1 U19428 ( .A(n25249), .B(n24767), .Y(n12700) );
  sky130_fd_sc_hd__xnor3_1 U19429 ( .A(n12701), .B(n18435), .C(n18433), .X(
        n18400) );
  sky130_fd_sc_hd__xnor2_1 U19430 ( .A(n18456), .B(n18457), .Y(n18436) );
  sky130_fd_sc_hd__nand2_1 U19431 ( .A(n12703), .B(n12702), .Y(n18456) );
  sky130_fd_sc_hd__nand2_1 U19432 ( .A(n18435), .B(n18434), .Y(n12702) );
  sky130_fd_sc_hd__o21ai_1 U19434 ( .A1(n22281), .A2(n23154), .B1(n22280), .Y(
        n13226) );
  sky130_fd_sc_hd__clkbuf_1 U19436 ( .A(n23242), .X(n12706) );
  sky130_fd_sc_hd__or2_0 U19437 ( .A(n26102), .B(n26101), .X(n12707) );
  sky130_fd_sc_hd__clkbuf_1 U19439 ( .A(j202_soc_core_j22_cpu_ml_bufa[10]), 
        .X(n12708) );
  sky130_fd_sc_hd__nand2_4 U19440 ( .A(n17427), .B(n12133), .Y(n17771) );
  sky130_fd_sc_hd__nand2_1 U19441 ( .A(n12710), .B(n12709), .Y(n17518) );
  sky130_fd_sc_hd__nand2_1 U19442 ( .A(n17431), .B(n17432), .Y(n12709) );
  sky130_fd_sc_hd__o21ai_1 U19443 ( .A1(n17432), .A2(n17431), .B1(n17430), .Y(
        n12710) );
  sky130_fd_sc_hd__xnor2_1 U19444 ( .A(n17432), .B(n17430), .Y(n12711) );
  sky130_fd_sc_hd__inv_2 U19445 ( .A(n22287), .Y(n23143) );
  sky130_fd_sc_hd__nor2_1 U19446 ( .A(n12972), .B(n12970), .Y(n12969) );
  sky130_fd_sc_hd__fah_1 U19447 ( .A(n18647), .B(n18646), .CI(n18645), .COUT(
        n18852), .SUM(n18849) );
  sky130_fd_sc_hd__inv_1 U19448 ( .A(n15219), .Y(n13150) );
  sky130_fd_sc_hd__nand2_1 U19449 ( .A(n12718), .B(n12717), .Y(n18267) );
  sky130_fd_sc_hd__nand2_1 U19450 ( .A(n18253), .B(n18254), .Y(n12717) );
  sky130_fd_sc_hd__nand2_1 U19451 ( .A(n12722), .B(n12719), .Y(n12718) );
  sky130_fd_sc_hd__nand2_1 U19452 ( .A(n12721), .B(n12720), .Y(n12719) );
  sky130_fd_sc_hd__xnor2_1 U19453 ( .A(n12723), .B(n12722), .Y(n18261) );
  sky130_fd_sc_hd__nand2_1 U19454 ( .A(n18165), .B(n18164), .Y(n12722) );
  sky130_fd_sc_hd__xnor2_1 U19455 ( .A(n18254), .B(n18253), .Y(n12723) );
  sky130_fd_sc_hd__fah_1 U19456 ( .A(n18097), .B(n18096), .CI(n18095), .COUT(
        n18163), .SUM(n18158) );
  sky130_fd_sc_hd__o21ai_2 U19457 ( .A1(n21498), .A2(n22897), .B1(n21499), .Y(
        n18875) );
  sky130_fd_sc_hd__nand2_1 U19458 ( .A(n27044), .B(n11153), .Y(n12724) );
  sky130_fd_sc_hd__clkbuf_1 U19459 ( .A(j202_soc_core_j22_cpu_ml_bufa[22]), 
        .X(n12725) );
  sky130_fd_sc_hd__and2_0 U19460 ( .A(n22503), .B(n22504), .X(n12726) );
  sky130_fd_sc_hd__inv_2 U19462 ( .A(n23210), .Y(n12731) );
  sky130_fd_sc_hd__nand2_1 U19463 ( .A(n12737), .B(n12736), .Y(
        j202_soc_core_j22_cpu_rf_N3082) );
  sky130_fd_sc_hd__nand2_1 U19464 ( .A(n11771), .B(n11137), .Y(n12736) );
  sky130_fd_sc_hd__nand2_1 U19465 ( .A(n24497), .B(n26371), .Y(n12737) );
  sky130_fd_sc_hd__nand2_4 U19466 ( .A(n26512), .B(n12738), .Y(n24497) );
  sky130_fd_sc_hd__a21o_1 U19468 ( .A1(n10971), .A2(n18067), .B1(n18066), .X(
        n18098) );
  sky130_fd_sc_hd__fah_1 U19469 ( .A(n18122), .B(n18121), .CI(n18120), .COUT(
        n18173), .SUM(n18175) );
  sky130_fd_sc_hd__clkbuf_1 U19470 ( .A(n21878), .X(n12741) );
  sky130_fd_sc_hd__nand4_1 U19471 ( .A(n12810), .B(n12811), .C(n12812), .D(
        n12813), .Y(n12809) );
  sky130_fd_sc_hd__nor2_1 U19472 ( .A(n12964), .B(n12960), .Y(n12959) );
  sky130_fd_sc_hd__nand2_1 U19473 ( .A(n12747), .B(n12746), .Y(n17600) );
  sky130_fd_sc_hd__nand2_1 U19474 ( .A(n17603), .B(n17604), .Y(n12746) );
  sky130_fd_sc_hd__nand2_1 U19475 ( .A(n17602), .B(n12748), .Y(n12747) );
  sky130_fd_sc_hd__nand2b_1 U19476 ( .A_N(n17603), .B(n12749), .Y(n12748) );
  sky130_fd_sc_hd__xnor2_1 U19477 ( .A(n12750), .B(n17602), .Y(n17915) );
  sky130_fd_sc_hd__xnor2_1 U19478 ( .A(n17604), .B(n17603), .Y(n12750) );
  sky130_fd_sc_hd__fah_1 U19479 ( .A(n17623), .B(n17622), .CI(n17621), .COUT(
        n17924), .SUM(n17923) );
  sky130_fd_sc_hd__nand2_1 U19480 ( .A(n17901), .B(n12751), .Y(n17597) );
  sky130_fd_sc_hd__nand2_1 U19481 ( .A(n12752), .B(n17595), .Y(n12751) );
  sky130_fd_sc_hd__nand2_1 U19482 ( .A(n12754), .B(n12753), .Y(n17610) );
  sky130_fd_sc_hd__nand2_1 U19483 ( .A(n17615), .B(n12756), .Y(n12753) );
  sky130_fd_sc_hd__xnor2_1 U19485 ( .A(n17614), .B(n12755), .Y(n17670) );
  sky130_fd_sc_hd__xnor2_1 U19486 ( .A(n12756), .B(n17615), .Y(n12755) );
  sky130_fd_sc_hd__o22ai_1 U19487 ( .A1(n17537), .A2(n17786), .B1(n17579), 
        .B2(n17771), .Y(n12756) );
  sky130_fd_sc_hd__nand2_1 U19488 ( .A(n12759), .B(n12758), .Y(n18813) );
  sky130_fd_sc_hd__nand2_1 U19489 ( .A(n12761), .B(n18614), .Y(n12758) );
  sky130_fd_sc_hd__o21ai_1 U19490 ( .A1(n18614), .A2(n12761), .B1(n18613), .Y(
        n12759) );
  sky130_fd_sc_hd__xnor2_1 U19491 ( .A(n18614), .B(n18613), .Y(n12760) );
  sky130_fd_sc_hd__xor2_1 U19492 ( .A(n12762), .B(n18601), .X(n12761) );
  sky130_fd_sc_hd__clkbuf_1 U19493 ( .A(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]), .X(n12763) );
  sky130_fd_sc_hd__nand2_1 U19494 ( .A(n24301), .B(n24300), .Y(n12766) );
  sky130_fd_sc_hd__clkbuf_1 U19495 ( .A(j202_soc_core_j22_cpu_ml_bufa[29]), 
        .X(n12767) );
  sky130_fd_sc_hd__o21a_1 U19496 ( .A1(n26579), .A2(n26432), .B1(n24494), .X(
        n12768) );
  sky130_fd_sc_hd__nand2_1 U19497 ( .A(n26519), .B(n26323), .Y(n12769) );
  sky130_fd_sc_hd__nand2_1 U19499 ( .A(n12415), .B(n18919), .Y(n18985) );
  sky130_fd_sc_hd__nand3_2 U19500 ( .A(n26444), .B(n12772), .C(n26445), .Y(
        n12802) );
  sky130_fd_sc_hd__nand2_1 U19501 ( .A(n26404), .B(n26403), .Y(n12772) );
  sky130_fd_sc_hd__nand2_1 U19502 ( .A(n22944), .B(n22660), .Y(n12773) );
  sky130_fd_sc_hd__nand2_1 U19503 ( .A(n12775), .B(n12774), .Y(n18541) );
  sky130_fd_sc_hd__nand2_1 U19504 ( .A(n18483), .B(n18484), .Y(n12774) );
  sky130_fd_sc_hd__o21ai_1 U19505 ( .A1(n18484), .A2(n18483), .B1(n18482), .Y(
        n12775) );
  sky130_fd_sc_hd__nand2_1 U19506 ( .A(n12778), .B(n12777), .Y(n18803) );
  sky130_fd_sc_hd__nand2_1 U19507 ( .A(n18802), .B(n18801), .Y(n12777) );
  sky130_fd_sc_hd__xnor2_1 U19509 ( .A(n12779), .B(n18800), .Y(n18791) );
  sky130_fd_sc_hd__xnor2_1 U19510 ( .A(n18801), .B(n18802), .Y(n12779) );
  sky130_fd_sc_hd__nand2_1 U19511 ( .A(n12782), .B(n12275), .Y(
        j202_soc_core_j22_cpu_ml_machj[7]) );
  sky130_fd_sc_hd__nand2_1 U19512 ( .A(n27187), .B(n19012), .Y(n12781) );
  sky130_fd_sc_hd__nand2_1 U19513 ( .A(n12916), .B(n24736), .Y(n12782) );
  sky130_fd_sc_hd__nand2_1 U19514 ( .A(n12784), .B(n12276), .Y(
        j202_soc_core_j22_cpu_ml_machj[5]) );
  sky130_fd_sc_hd__nand2_1 U19515 ( .A(n12916), .B(n12995), .Y(n12784) );
  sky130_fd_sc_hd__nand2_1 U19516 ( .A(n12785), .B(n12156), .Y(
        j202_soc_core_j22_cpu_ml_machj[2]) );
  sky130_fd_sc_hd__nand2_1 U19517 ( .A(n12786), .B(n12157), .Y(n29321) );
  sky130_fd_sc_hd__nand2_1 U19518 ( .A(n12916), .B(n12996), .Y(n12786) );
  sky130_fd_sc_hd__nand2_1 U19519 ( .A(n12788), .B(n12787), .Y(n18399) );
  sky130_fd_sc_hd__nand2_1 U19520 ( .A(n18597), .B(n18598), .Y(n12787) );
  sky130_fd_sc_hd__o21ai_1 U19521 ( .A1(n18598), .A2(n18597), .B1(n18596), .Y(
        n12788) );
  sky130_fd_sc_hd__clkbuf_1 U19522 ( .A(n18997), .X(n12789) );
  sky130_fd_sc_hd__nand2_1 U19523 ( .A(n20970), .B(n12793), .Y(n12792) );
  sky130_fd_sc_hd__and2_0 U19524 ( .A(n20968), .B(n20969), .X(n12793) );
  sky130_fd_sc_hd__nand4_1 U19525 ( .A(n12798), .B(n12797), .C(n12796), .D(
        n12795), .Y(n12794) );
  sky130_fd_sc_hd__nand2_1 U19526 ( .A(j202_soc_core_memory0_ram_dout0[423]), 
        .B(n21598), .Y(n12795) );
  sky130_fd_sc_hd__nand2_1 U19527 ( .A(j202_soc_core_memory0_ram_dout0[199]), 
        .B(n21732), .Y(n12796) );
  sky130_fd_sc_hd__nand2_1 U19528 ( .A(j202_soc_core_memory0_ram_dout0[263]), 
        .B(n21605), .Y(n12797) );
  sky130_fd_sc_hd__nand2_1 U19529 ( .A(j202_soc_core_memory0_ram_dout0[359]), 
        .B(n21596), .Y(n12798) );
  sky130_fd_sc_hd__nand2_1 U19530 ( .A(j202_soc_core_memory0_ram_dout0[103]), 
        .B(n21591), .Y(n12800) );
  sky130_fd_sc_hd__nand2_1 U19531 ( .A(j202_soc_core_memory0_ram_dout0[455]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12801) );
  sky130_fd_sc_hd__nand2_1 U19532 ( .A(n12802), .B(n27192), .Y(n26468) );
  sky130_fd_sc_hd__nand2_1 U19533 ( .A(n12802), .B(n26516), .Y(n26448) );
  sky130_fd_sc_hd__and3_1 U19534 ( .A(n20543), .B(n20556), .C(n20557), .X(
        n12803) );
  sky130_fd_sc_hd__nand2_1 U19535 ( .A(j202_soc_core_memory0_ram_dout0[384]), 
        .B(n21597), .Y(n12805) );
  sky130_fd_sc_hd__nand2_1 U19536 ( .A(j202_soc_core_memory0_ram_dout0[224]), 
        .B(n21735), .Y(n12806) );
  sky130_fd_sc_hd__nand2_1 U19537 ( .A(j202_soc_core_memory0_ram_dout0[0]), 
        .B(n21733), .Y(n12807) );
  sky130_fd_sc_hd__nand2_1 U19538 ( .A(j202_soc_core_memory0_ram_dout0[12]), 
        .B(n21733), .Y(n12810) );
  sky130_fd_sc_hd__nand2_1 U19539 ( .A(j202_soc_core_memory0_ram_dout0[364]), 
        .B(n21596), .Y(n12811) );
  sky130_fd_sc_hd__nand2_1 U19540 ( .A(j202_soc_core_memory0_ram_dout0[44]), 
        .B(n21604), .Y(n12812) );
  sky130_fd_sc_hd__nand2_1 U19541 ( .A(j202_soc_core_memory0_ram_dout0[332]), 
        .B(n21593), .Y(n12813) );
  sky130_fd_sc_hd__nand2_1 U19542 ( .A(j202_soc_core_memory0_ram_dout0[300]), 
        .B(n21603), .Y(n12815) );
  sky130_fd_sc_hd__nand2_1 U19543 ( .A(j202_soc_core_memory0_ram_dout0[108]), 
        .B(n21591), .Y(n12816) );
  sky130_fd_sc_hd__nand2_1 U19544 ( .A(j202_soc_core_memory0_ram_dout0[268]), 
        .B(n21605), .Y(n12817) );
  sky130_fd_sc_hd__nand2_1 U19545 ( .A(j202_soc_core_memory0_ram_dout0[460]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12818) );
  sky130_fd_sc_hd__nand4_1 U19546 ( .A(n12824), .B(n12823), .C(n12822), .D(
        n12821), .Y(n12820) );
  sky130_fd_sc_hd__nand2_1 U19547 ( .A(j202_soc_core_memory0_ram_dout0[138]), 
        .B(n21592), .Y(n12821) );
  sky130_fd_sc_hd__nand2_1 U19548 ( .A(j202_soc_core_memory0_ram_dout0[330]), 
        .B(n21593), .Y(n12822) );
  sky130_fd_sc_hd__nand2_1 U19549 ( .A(j202_soc_core_memory0_ram_dout0[170]), 
        .B(n21590), .Y(n12823) );
  sky130_fd_sc_hd__nand2_1 U19550 ( .A(j202_soc_core_memory0_ram_dout0[106]), 
        .B(n21591), .Y(n12824) );
  sky130_fd_sc_hd__nand4_1 U19551 ( .A(n12828), .B(n12829), .C(n12827), .D(
        n12826), .Y(n12825) );
  sky130_fd_sc_hd__nand2_1 U19552 ( .A(j202_soc_core_memory0_ram_dout0[458]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12826) );
  sky130_fd_sc_hd__nand2_1 U19553 ( .A(j202_soc_core_memory0_ram_dout0[426]), 
        .B(n21598), .Y(n12827) );
  sky130_fd_sc_hd__nand2_1 U19554 ( .A(j202_soc_core_memory0_ram_dout0[362]), 
        .B(n21596), .Y(n12828) );
  sky130_fd_sc_hd__nand2_1 U19555 ( .A(j202_soc_core_memory0_ram_dout0[394]), 
        .B(n21597), .Y(n12829) );
  sky130_fd_sc_hd__nand4_1 U19556 ( .A(n12835), .B(n12834), .C(n12833), .D(
        n12832), .Y(n12831) );
  sky130_fd_sc_hd__nand2_1 U19557 ( .A(j202_soc_core_memory0_ram_dout0[10]), 
        .B(n21733), .Y(n12832) );
  sky130_fd_sc_hd__nand2_1 U19558 ( .A(j202_soc_core_memory0_ram_dout0[202]), 
        .B(n21732), .Y(n12833) );
  sky130_fd_sc_hd__nand2_1 U19559 ( .A(j202_soc_core_memory0_ram_dout0[298]), 
        .B(n21603), .Y(n12834) );
  sky130_fd_sc_hd__nand2_1 U19560 ( .A(j202_soc_core_memory0_ram_dout0[42]), 
        .B(n21604), .Y(n12835) );
  sky130_fd_sc_hd__nand4_1 U19561 ( .A(n12839), .B(n12838), .C(n12837), .D(
        n19144), .Y(n12836) );
  sky130_fd_sc_hd__nand2_1 U19562 ( .A(j202_soc_core_memory0_ram_dout0[234]), 
        .B(n21735), .Y(n12837) );
  sky130_fd_sc_hd__nand2_1 U19563 ( .A(j202_soc_core_memory0_ram_dout0[74]), 
        .B(n21734), .Y(n12838) );
  sky130_fd_sc_hd__nand2_1 U19564 ( .A(j202_soc_core_memory0_ram_dout0[266]), 
        .B(n21605), .Y(n12839) );
  sky130_fd_sc_hd__nand2_1 U19565 ( .A(n12840), .B(n19172), .Y(n19196) );
  sky130_fd_sc_hd__nand2_1 U19566 ( .A(n11705), .B(n27452), .Y(n27437) );
  sky130_fd_sc_hd__nand2_1 U19567 ( .A(n11705), .B(n11157), .Y(n25240) );
  sky130_fd_sc_hd__a22oi_1 U19568 ( .A1(n25244), .A2(n26948), .B1(n11705), 
        .B2(n24650), .Y(n25245) );
  sky130_fd_sc_hd__and3_1 U19569 ( .A(n22311), .B(n19211), .C(n22310), .X(
        n12841) );
  sky130_fd_sc_hd__nand2_1 U19570 ( .A(n12850), .B(n12843), .Y(n21752) );
  sky130_fd_sc_hd__nand4_1 U19571 ( .A(n12845), .B(n12846), .C(n12847), .D(
        n12848), .Y(n12844) );
  sky130_fd_sc_hd__nand2_1 U19572 ( .A(j202_soc_core_memory0_ram_dout0[405]), 
        .B(n21597), .Y(n12845) );
  sky130_fd_sc_hd__nand2_1 U19573 ( .A(j202_soc_core_memory0_ram_dout0[373]), 
        .B(n21596), .Y(n12846) );
  sky130_fd_sc_hd__nand2_1 U19574 ( .A(j202_soc_core_memory0_ram_dout0[437]), 
        .B(n21598), .Y(n12847) );
  sky130_fd_sc_hd__nand2_1 U19575 ( .A(j202_soc_core_memory0_ram_dout0[469]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12848) );
  sky130_fd_sc_hd__nand4_1 U19576 ( .A(n15526), .B(n15527), .C(n15528), .D(
        n15529), .Y(n12851) );
  sky130_fd_sc_hd__nand4_1 U19577 ( .A(n15641), .B(n15640), .C(n15639), .D(
        n15638), .Y(n12852) );
  sky130_fd_sc_hd__nand2_1 U19578 ( .A(j202_soc_core_memory0_ram_dout0[377]), 
        .B(n21596), .Y(n12856) );
  sky130_fd_sc_hd__nand2_1 U19579 ( .A(j202_soc_core_memory0_ram_dout0[473]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12857) );
  sky130_fd_sc_hd__nand2_1 U19580 ( .A(j202_soc_core_memory0_ram_dout0[441]), 
        .B(n21598), .Y(n12858) );
  sky130_fd_sc_hd__nand2_1 U19581 ( .A(j202_soc_core_memory0_ram_dout0[57]), 
        .B(n21604), .Y(n12860) );
  sky130_fd_sc_hd__nand2_1 U19582 ( .A(j202_soc_core_memory0_ram_dout0[185]), 
        .B(n21590), .Y(n12861) );
  sky130_fd_sc_hd__nand2_1 U19583 ( .A(j202_soc_core_memory0_ram_dout0[313]), 
        .B(n21603), .Y(n12862) );
  sky130_fd_sc_hd__nand4_1 U19584 ( .A(n12868), .B(n12867), .C(n12866), .D(
        n12865), .Y(n12864) );
  sky130_fd_sc_hd__nand2_1 U19585 ( .A(j202_soc_core_memory0_ram_dout0[217]), 
        .B(n21732), .Y(n12865) );
  sky130_fd_sc_hd__nand2_1 U19586 ( .A(j202_soc_core_memory0_ram_dout0[121]), 
        .B(n21591), .Y(n12866) );
  sky130_fd_sc_hd__nand2_1 U19587 ( .A(j202_soc_core_memory0_ram_dout0[153]), 
        .B(n21592), .Y(n12867) );
  sky130_fd_sc_hd__nand2_1 U19588 ( .A(j202_soc_core_memory0_ram_dout0[89]), 
        .B(n21734), .Y(n12868) );
  sky130_fd_sc_hd__inv_1 U19589 ( .A(n12870), .Y(n12869) );
  sky130_fd_sc_hd__nand4_1 U19590 ( .A(n12874), .B(n12873), .C(n12872), .D(
        n12871), .Y(n12870) );
  sky130_fd_sc_hd__nand2_1 U19591 ( .A(j202_soc_core_memory0_ram_dout0[345]), 
        .B(n21593), .Y(n12871) );
  sky130_fd_sc_hd__nand2_1 U19592 ( .A(j202_soc_core_memory0_ram_dout0[281]), 
        .B(n21605), .Y(n12872) );
  sky130_fd_sc_hd__nand2_1 U19593 ( .A(j202_soc_core_memory0_ram_dout0[409]), 
        .B(n21597), .Y(n12873) );
  sky130_fd_sc_hd__nand2_1 U19594 ( .A(j202_soc_core_memory0_ram_dout0[249]), 
        .B(n21735), .Y(n12874) );
  sky130_fd_sc_hd__nand3_1 U19595 ( .A(n12911), .B(n15898), .C(n21776), .Y(
        n20962) );
  sky130_fd_sc_hd__nand3_1 U19596 ( .A(n12878), .B(n19158), .C(n21750), .Y(
        n20960) );
  sky130_fd_sc_hd__inv_1 U19597 ( .A(n29014), .Y(n25048) );
  sky130_fd_sc_hd__nand2_1 U19598 ( .A(n12882), .B(n27980), .Y(n12881) );
  sky130_fd_sc_hd__nand2_1 U19599 ( .A(n27169), .B(n12655), .Y(n12882) );
  sky130_fd_sc_hd__inv_2 U19600 ( .A(n13194), .Y(n24310) );
  sky130_fd_sc_hd__nand2_1 U19601 ( .A(j202_soc_core_memory0_ram_dout0[307]), 
        .B(n21603), .Y(n12885) );
  sky130_fd_sc_hd__nand2_1 U19602 ( .A(j202_soc_core_memory0_ram_dout0[51]), 
        .B(n21604), .Y(n12886) );
  sky130_fd_sc_hd__nand2_1 U19603 ( .A(j202_soc_core_memory0_ram_dout0[243]), 
        .B(n21735), .Y(n12887) );
  sky130_fd_sc_hd__nand2_1 U19604 ( .A(j202_soc_core_memory0_ram_dout0[19]), 
        .B(n21733), .Y(n12888) );
  sky130_fd_sc_hd__nand4_1 U19605 ( .A(n12890), .B(n12892), .C(n12893), .D(
        n12891), .Y(n12889) );
  sky130_fd_sc_hd__nand2_1 U19606 ( .A(j202_soc_core_memory0_ram_dout0[339]), 
        .B(n21593), .Y(n12890) );
  sky130_fd_sc_hd__nand2_1 U19607 ( .A(j202_soc_core_memory0_ram_dout0[179]), 
        .B(n21590), .Y(n12891) );
  sky130_fd_sc_hd__nand2_1 U19608 ( .A(j202_soc_core_memory0_ram_dout0[275]), 
        .B(n21605), .Y(n12892) );
  sky130_fd_sc_hd__nand2_1 U19609 ( .A(j202_soc_core_memory0_ram_dout0[403]), 
        .B(n21597), .Y(n12893) );
  sky130_fd_sc_hd__nand2_1 U19610 ( .A(j202_soc_core_memory0_ram_dout0[499]), 
        .B(n21771), .Y(n12894) );
  sky130_fd_sc_hd__nand2_1 U19611 ( .A(n12897), .B(n12896), .Y(n12895) );
  sky130_fd_sc_hd__nand2_1 U19612 ( .A(j202_soc_core_memory0_ram_dout0[371]), 
        .B(n21596), .Y(n12896) );
  sky130_fd_sc_hd__nand2_1 U19613 ( .A(j202_soc_core_memory0_ram_dout0[467]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n12897) );
  sky130_fd_sc_hd__inv_2 U19616 ( .A(n27619), .Y(n12902) );
  sky130_fd_sc_hd__nor2_1 U19632 ( .A(n20715), .B(n20716), .Y(n12913) );
  sky130_fd_sc_hd__inv_2 U19633 ( .A(n23256), .Y(n27274) );
  sky130_fd_sc_hd__inv_2 U19634 ( .A(n12917), .Y(n12999) );
  sky130_fd_sc_hd__nand2_1 U19635 ( .A(n12920), .B(n12919), .Y(n18821) );
  sky130_fd_sc_hd__nand2_1 U19636 ( .A(n18550), .B(n18551), .Y(n12919) );
  sky130_fd_sc_hd__xnor2_1 U19638 ( .A(n18551), .B(n18550), .Y(n12921) );
  sky130_fd_sc_hd__nand2_1 U19639 ( .A(n12923), .B(n12922), .Y(n18508) );
  sky130_fd_sc_hd__nand2_1 U19640 ( .A(n18475), .B(n18476), .Y(n12922) );
  sky130_fd_sc_hd__xor2_1 U19642 ( .A(n18474), .B(n12924), .X(n18438) );
  sky130_fd_sc_hd__xnor2_1 U19643 ( .A(n12925), .B(n18475), .Y(n12924) );
  sky130_fd_sc_hd__nand2_1 U19644 ( .A(n12931), .B(n12930), .Y(n18833) );
  sky130_fd_sc_hd__nand2_1 U19645 ( .A(n18745), .B(n18746), .Y(n12930) );
  sky130_fd_sc_hd__o21ai_1 U19646 ( .A1(n18746), .A2(n18745), .B1(n18744), .Y(
        n12931) );
  sky130_fd_sc_hd__nand2_1 U19647 ( .A(n12933), .B(n12932), .Y(n18743) );
  sky130_fd_sc_hd__nand2_1 U19648 ( .A(n18740), .B(n18739), .Y(n12932) );
  sky130_fd_sc_hd__o21ai_1 U19649 ( .A1(n18739), .A2(n18740), .B1(n18738), .Y(
        n12933) );
  sky130_fd_sc_hd__xnor2_1 U19650 ( .A(n18740), .B(n12934), .Y(n18797) );
  sky130_fd_sc_hd__xnor2_1 U19651 ( .A(n18739), .B(n18738), .Y(n12934) );
  sky130_fd_sc_hd__nand2_1 U19652 ( .A(n12940), .B(n13214), .Y(n24161) );
  sky130_fd_sc_hd__o21ai_1 U19653 ( .A1(n12940), .A2(n12939), .B1(n12936), .Y(
        n12935) );
  sky130_fd_sc_hd__nor2b_1 U19654 ( .B_N(n11153), .A(n24162), .Y(n12937) );
  sky130_fd_sc_hd__o21ai_1 U19655 ( .A1(n12351), .A2(n12939), .B1(n26726), .Y(
        n12938) );
  sky130_fd_sc_hd__or2_0 U19656 ( .A(n26443), .B(n24162), .X(n12939) );
  sky130_fd_sc_hd__nand3_1 U19657 ( .A(n21755), .B(n21750), .C(n21754), .Y(
        n13198) );
  sky130_fd_sc_hd__xnor2_1 U19658 ( .A(n12941), .B(n12944), .Y(n18125) );
  sky130_fd_sc_hd__xor2_1 U19659 ( .A(n18135), .B(n18134), .X(n12941) );
  sky130_fd_sc_hd__nand2_1 U19660 ( .A(n12943), .B(n12942), .Y(n18243) );
  sky130_fd_sc_hd__nand2_1 U19661 ( .A(n18134), .B(n18135), .Y(n12942) );
  sky130_fd_sc_hd__o21ai_1 U19662 ( .A1(n18135), .A2(n18134), .B1(n12945), .Y(
        n12943) );
  sky130_fd_sc_hd__inv_2 U19663 ( .A(n12945), .Y(n12944) );
  sky130_fd_sc_hd__o22ai_1 U19664 ( .A1(n18514), .A2(n18138), .B1(n18110), 
        .B2(n18424), .Y(n12945) );
  sky130_fd_sc_hd__nand2_1 U19665 ( .A(n18563), .B(n18564), .Y(n12946) );
  sky130_fd_sc_hd__nand2_1 U19666 ( .A(n12952), .B(n12948), .Y(n12947) );
  sky130_fd_sc_hd__nand2_1 U19667 ( .A(n12950), .B(n12949), .Y(n12948) );
  sky130_fd_sc_hd__xnor2_1 U19668 ( .A(n12952), .B(n12951), .Y(n18590) );
  sky130_fd_sc_hd__xnor2_1 U19669 ( .A(n18564), .B(n18563), .Y(n12951) );
  sky130_fd_sc_hd__nand2_1 U19670 ( .A(n18248), .B(n12953), .Y(n12952) );
  sky130_fd_sc_hd__o21ai_1 U19671 ( .A1(n18250), .A2(n18252), .B1(n18249), .Y(
        n12953) );
  sky130_fd_sc_hd__nand2_1 U19672 ( .A(n28996), .B(n24225), .Y(n12954) );
  sky130_fd_sc_hd__nand4_1 U19673 ( .A(n19255), .B(n19254), .C(n19256), .D(
        n12957), .Y(n12956) );
  sky130_fd_sc_hd__nand2_1 U19674 ( .A(j202_soc_core_memory0_ram_dout0[428]), 
        .B(n21598), .Y(n12957) );
  sky130_fd_sc_hd__nand2_1 U19675 ( .A(j202_soc_core_memory0_ram_dout0[413]), 
        .B(n21597), .Y(n12961) );
  sky130_fd_sc_hd__nand2_1 U19676 ( .A(j202_soc_core_memory0_ram_dout0[61]), 
        .B(n21604), .Y(n12962) );
  sky130_fd_sc_hd__nand2_1 U19677 ( .A(j202_soc_core_memory0_ram_dout0[317]), 
        .B(n21603), .Y(n12963) );
  sky130_fd_sc_hd__nand4_1 U19678 ( .A(n12968), .B(n12967), .C(n12965), .D(
        n12966), .Y(n12964) );
  sky130_fd_sc_hd__nand2_1 U19679 ( .A(j202_soc_core_memory0_ram_dout0[445]), 
        .B(n21598), .Y(n12965) );
  sky130_fd_sc_hd__nand2_1 U19680 ( .A(j202_soc_core_memory0_ram_dout0[221]), 
        .B(n21732), .Y(n12967) );
  sky130_fd_sc_hd__nand2_1 U19681 ( .A(j202_soc_core_memory0_ram_dout0[285]), 
        .B(n21605), .Y(n12968) );
  sky130_fd_sc_hd__nand2_1 U19682 ( .A(j202_soc_core_memory0_ram_dout0[253]), 
        .B(n21735), .Y(n12971) );
  sky130_fd_sc_hd__nand4_1 U19683 ( .A(n20566), .B(n20567), .C(n20696), .D(
        n20697), .Y(n12975) );
  sky130_fd_sc_hd__and2_0 U19685 ( .A(n20704), .B(n20695), .X(n12977) );
  sky130_fd_sc_hd__nand2_1 U19686 ( .A(n12980), .B(n26422), .Y(n12986) );
  sky130_fd_sc_hd__nand2_1 U19687 ( .A(n11669), .B(n12981), .Y(n12980) );
  sky130_fd_sc_hd__nand4_1 U19688 ( .A(n12982), .B(n12989), .C(n22716), .D(
        n22717), .Y(n12987) );
  sky130_fd_sc_hd__nor2_2 U19689 ( .A(n22713), .B(n26524), .Y(n12983) );
  sky130_fd_sc_hd__nor2_2 U19690 ( .A(n18276), .B(n18275), .Y(n22828) );
  sky130_fd_sc_hd__nand2_1 U19691 ( .A(n12991), .B(n18660), .Y(n13200) );
  sky130_fd_sc_hd__o22ai_1 U19692 ( .A1(n18660), .A2(n18351), .B1(n18299), 
        .B2(n12991), .Y(n18362) );
  sky130_fd_sc_hd__o22ai_1 U19693 ( .A1(n12991), .A2(n18200), .B1(n18660), 
        .B2(n18232), .Y(n18216) );
  sky130_fd_sc_hd__o22ai_1 U19694 ( .A1(n18660), .A2(n18299), .B1(n18306), 
        .B2(n12991), .Y(n18345) );
  sky130_fd_sc_hd__o22ai_1 U19695 ( .A1(n18660), .A2(n18200), .B1(n18137), 
        .B2(n12991), .Y(n18186) );
  sky130_fd_sc_hd__o22ai_1 U19696 ( .A1(n18660), .A2(n18109), .B1(n18059), 
        .B2(n12991), .Y(n18096) );
  sky130_fd_sc_hd__o22ai_1 U19697 ( .A1(n18660), .A2(n18305), .B1(n18232), 
        .B2(n12991), .Y(n18333) );
  sky130_fd_sc_hd__o22ai_1 U19698 ( .A1(n12991), .A2(n18019), .B1(n18660), 
        .B2(n18059), .Y(n18053) );
  sky130_fd_sc_hd__o22ai_1 U19699 ( .A1(n18660), .A2(n18473), .B1(n18402), 
        .B2(n12991), .Y(n18465) );
  sky130_fd_sc_hd__o22ai_1 U19700 ( .A1(n18660), .A2(n18402), .B1(n18351), 
        .B2(n12991), .Y(n18432) );
  sky130_fd_sc_hd__o22ai_1 U19701 ( .A1(n18660), .A2(n18306), .B1(n18305), 
        .B2(n12991), .Y(n18557) );
  sky130_fd_sc_hd__nand2_4 U19702 ( .A(n18660), .B(n17969), .Y(n12991) );
  sky130_fd_sc_hd__nand2_1 U19703 ( .A(n12993), .B(n12992), .Y(n18174) );
  sky130_fd_sc_hd__nand2_1 U19704 ( .A(n18073), .B(n18074), .Y(n12992) );
  sky130_fd_sc_hd__o21ai_1 U19705 ( .A1(n18074), .A2(n18073), .B1(n18072), .Y(
        n12993) );
  sky130_fd_sc_hd__nor2_2 U19706 ( .A(n18271), .B(n18272), .Y(n18908) );
  sky130_fd_sc_hd__nand2b_1 U19707 ( .A_N(n24060), .B(n22450), .Y(n12995) );
  sky130_fd_sc_hd__nand2b_1 U19708 ( .A_N(n25337), .B(n25336), .Y(n12996) );
  sky130_fd_sc_hd__nand2_1 U19709 ( .A(n12916), .B(n24637), .Y(n24136) );
  sky130_fd_sc_hd__nand2_1 U19710 ( .A(n12916), .B(n23271), .Y(n23272) );
  sky130_fd_sc_hd__nand2_1 U19711 ( .A(n25822), .B(n12997), .Y(
        j202_soc_core_j22_cpu_ml_maclj[18]) );
  sky130_fd_sc_hd__nand3_1 U19712 ( .A(n12916), .B(n25875), .C(n25254), .Y(
        n12997) );
  sky130_fd_sc_hd__a21oi_1 U19713 ( .A1(n12999), .A2(n24511), .B1(n26976), .Y(
        n24512) );
  sky130_fd_sc_hd__a21oi_1 U19714 ( .A1(n12999), .A2(n24551), .B1(n26976), .Y(
        n24552) );
  sky130_fd_sc_hd__a21oi_1 U19715 ( .A1(n12999), .A2(n26978), .B1(n26976), .Y(
        n26979) );
  sky130_fd_sc_hd__nand2_1 U19716 ( .A(n13002), .B(n13001), .Y(n18076) );
  sky130_fd_sc_hd__nand2_1 U19717 ( .A(n18089), .B(n18088), .Y(n13001) );
  sky130_fd_sc_hd__xnor2_1 U19719 ( .A(n18087), .B(n13003), .Y(n18092) );
  sky130_fd_sc_hd__xnor2_1 U19720 ( .A(n18088), .B(n18089), .Y(n13003) );
  sky130_fd_sc_hd__nand2_1 U19721 ( .A(n13006), .B(n13005), .Y(n13004) );
  sky130_fd_sc_hd__nand2_1 U19722 ( .A(j202_soc_core_memory0_ram_dout0[388]), 
        .B(n21597), .Y(n13005) );
  sky130_fd_sc_hd__nand2_1 U19723 ( .A(j202_soc_core_memory0_ram_dout0[292]), 
        .B(n21603), .Y(n13006) );
  sky130_fd_sc_hd__nor2_1 U19724 ( .A(n27688), .B(n27561), .Y(n13009) );
  sky130_fd_sc_hd__nand2_1 U19725 ( .A(j202_soc_core_memory0_ram_dout0[290]), 
        .B(n21603), .Y(n13010) );
  sky130_fd_sc_hd__nand3_1 U19727 ( .A(n19826), .B(n13022), .C(n19827), .Y(
        n13013) );
  sky130_fd_sc_hd__nand2_1 U19728 ( .A(n13013), .B(n13012), .Y(n26851) );
  sky130_fd_sc_hd__nand2_1 U19729 ( .A(n19825), .B(n13022), .Y(n13012) );
  sky130_fd_sc_hd__nand3_2 U19730 ( .A(n13018), .B(n13020), .C(n13015), .Y(
        n26904) );
  sky130_fd_sc_hd__nor2_1 U19731 ( .A(n13017), .B(n12125), .Y(n13016) );
  sky130_fd_sc_hd__nand2_1 U19732 ( .A(n13019), .B(n13023), .Y(n13018) );
  sky130_fd_sc_hd__inv_1 U19733 ( .A(n19827), .Y(n13019) );
  sky130_fd_sc_hd__inv_1 U19734 ( .A(n19826), .Y(n13021) );
  sky130_fd_sc_hd__nand2_1 U19735 ( .A(n13026), .B(n13025), .Y(n13024) );
  sky130_fd_sc_hd__nand2_1 U19736 ( .A(n13028), .B(n19769), .Y(n13025) );
  sky130_fd_sc_hd__nand2_1 U19737 ( .A(n19651), .B(n19664), .Y(n13026) );
  sky130_fd_sc_hd__nand2_1 U19738 ( .A(n19775), .B(n19776), .Y(n13028) );
  sky130_fd_sc_hd__nand4_1 U19740 ( .A(n13035), .B(n13037), .C(n13217), .D(
        n13222), .Y(n13030) );
  sky130_fd_sc_hd__nand4_1 U19741 ( .A(n13036), .B(n13220), .C(n13039), .D(
        n13221), .Y(n13031) );
  sky130_fd_sc_hd__nand2_1 U19744 ( .A(n24497), .B(n26379), .Y(n13032) );
  sky130_fd_sc_hd__nand2_1 U19745 ( .A(j202_soc_core_memory0_ram_dout0[175]), 
        .B(n21590), .Y(n13033) );
  sky130_fd_sc_hd__nand2_1 U19746 ( .A(j202_soc_core_memory0_ram_dout0[335]), 
        .B(n21593), .Y(n13034) );
  sky130_fd_sc_hd__nand2_1 U19747 ( .A(j202_soc_core_memory0_ram_dout0[271]), 
        .B(n21605), .Y(n13035) );
  sky130_fd_sc_hd__nand2_1 U19748 ( .A(j202_soc_core_memory0_ram_dout0[15]), 
        .B(n21733), .Y(n13036) );
  sky130_fd_sc_hd__nand2_1 U19749 ( .A(j202_soc_core_memory0_ram_dout0[47]), 
        .B(n21604), .Y(n13037) );
  sky130_fd_sc_hd__nand2_1 U19750 ( .A(j202_soc_core_memory0_ram_dout0[399]), 
        .B(n21597), .Y(n13038) );
  sky130_fd_sc_hd__nand2_1 U19751 ( .A(j202_soc_core_memory0_ram_dout0[431]), 
        .B(n21598), .Y(n13039) );
  sky130_fd_sc_hd__nand2_1 U19752 ( .A(j202_soc_core_memory0_ram_dout0[82]), 
        .B(n21734), .Y(n13040) );
  sky130_fd_sc_hd__nand2_1 U19753 ( .A(j202_soc_core_memory0_ram_dout0[146]), 
        .B(n21592), .Y(n13041) );
  sky130_fd_sc_hd__nand2_1 U19754 ( .A(j202_soc_core_memory0_ram_dout0[306]), 
        .B(n21603), .Y(n13042) );
  sky130_fd_sc_hd__nand2_1 U19756 ( .A(n27965), .B(n13049), .Y(n13047) );
  sky130_fd_sc_hd__nor2_1 U19757 ( .A(n11793), .B(n13051), .Y(n24351) );
  sky130_fd_sc_hd__and2_0 U19758 ( .A(n21316), .B(n20975), .X(n13052) );
  sky130_fd_sc_hd__nand2_1 U19760 ( .A(j202_soc_core_memory0_ram_dout0[94]), 
        .B(n21734), .Y(n13057) );
  sky130_fd_sc_hd__nand2_1 U19761 ( .A(j202_soc_core_memory0_ram_dout0[158]), 
        .B(n21592), .Y(n13058) );
  sky130_fd_sc_hd__nand2_1 U19762 ( .A(j202_soc_core_memory0_ram_dout0[190]), 
        .B(n21590), .Y(n13059) );
  sky130_fd_sc_hd__nand2_1 U19763 ( .A(j202_soc_core_memory0_ram_dout0[446]), 
        .B(n21598), .Y(n13060) );
  sky130_fd_sc_hd__nand2_1 U19764 ( .A(j202_soc_core_memory0_ram_dout0[478]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n13061) );
  sky130_fd_sc_hd__nand2_1 U19765 ( .A(j202_soc_core_memory0_ram_dout0[222]), 
        .B(n21732), .Y(n13062) );
  sky130_fd_sc_hd__nand2_1 U19766 ( .A(j202_soc_core_memory0_ram_dout0[126]), 
        .B(n21591), .Y(n13063) );
  sky130_fd_sc_hd__nand2_1 U19767 ( .A(n12642), .B(n24094), .Y(n27256) );
  sky130_fd_sc_hd__nand2_1 U19768 ( .A(n13065), .B(n29535), .Y(n24464) );
  sky130_fd_sc_hd__nand2_1 U19769 ( .A(n21914), .B(n22715), .Y(n13069) );
  sky130_fd_sc_hd__inv_2 U19770 ( .A(n29053), .Y(n22273) );
  sky130_fd_sc_hd__nand2_1 U19771 ( .A(j202_soc_core_memory0_ram_dout0[197]), 
        .B(n21732), .Y(n13073) );
  sky130_fd_sc_hd__nand3_1 U19772 ( .A(n13075), .B(n13271), .C(n13074), .Y(
        n13080) );
  sky130_fd_sc_hd__nand2_1 U19773 ( .A(n13077), .B(n23163), .Y(n13074) );
  sky130_fd_sc_hd__nand2_1 U19774 ( .A(n23154), .B(n23163), .Y(n13075) );
  sky130_fd_sc_hd__nand2b_1 U19775 ( .A_N(n23154), .B(n12677), .Y(n13078) );
  sky130_fd_sc_hd__nand2_1 U19776 ( .A(n27877), .B(n13083), .Y(n27568) );
  sky130_fd_sc_hd__nand2_1 U19777 ( .A(n11073), .B(n12278), .Y(n27694) );
  sky130_fd_sc_hd__inv_1 U19778 ( .A(n12438), .Y(n13082) );
  sky130_fd_sc_hd__nand4_1 U19779 ( .A(n13092), .B(n13097), .C(n13087), .D(
        n13085), .Y(n13084) );
  sky130_fd_sc_hd__nand2_1 U19780 ( .A(j202_soc_core_memory0_ram_dout0[148]), 
        .B(n21592), .Y(n13088) );
  sky130_fd_sc_hd__nand2_1 U19781 ( .A(j202_soc_core_memory0_ram_dout0[468]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n13089) );
  sky130_fd_sc_hd__nand2_1 U19782 ( .A(j202_soc_core_memory0_ram_dout0[180]), 
        .B(n21590), .Y(n13090) );
  sky130_fd_sc_hd__nand2_1 U19783 ( .A(j202_soc_core_memory0_ram_dout0[116]), 
        .B(n21591), .Y(n13091) );
  sky130_fd_sc_hd__nand2_1 U19784 ( .A(j202_soc_core_memory0_ram_dout0[372]), 
        .B(n21596), .Y(n13094) );
  sky130_fd_sc_hd__nand2_1 U19785 ( .A(j202_soc_core_memory0_ram_dout0[436]), 
        .B(n21598), .Y(n13095) );
  sky130_fd_sc_hd__nand2_1 U19786 ( .A(j202_soc_core_memory0_ram_dout0[340]), 
        .B(n21593), .Y(n13096) );
  sky130_fd_sc_hd__nand2_1 U19789 ( .A(j202_soc_core_memory0_ram_dout0[212]), 
        .B(n21732), .Y(n13100) );
  sky130_fd_sc_hd__nand2_1 U19790 ( .A(j202_soc_core_memory0_ram_dout0[244]), 
        .B(n21735), .Y(n13101) );
  sky130_fd_sc_hd__nand3_2 U19792 ( .A(n13104), .B(n13105), .C(n23000), .Y(
        n23001) );
  sky130_fd_sc_hd__nand2_1 U19793 ( .A(n26531), .B(n22999), .Y(n13104) );
  sky130_fd_sc_hd__nand2_1 U19794 ( .A(j202_soc_core_memory0_ram_dout0[440]), 
        .B(n21598), .Y(n13106) );
  sky130_fd_sc_hd__nand2_1 U19795 ( .A(j202_soc_core_memory0_ram_dout0[376]), 
        .B(n21596), .Y(n13107) );
  sky130_fd_sc_hd__nand2_1 U19796 ( .A(j202_soc_core_memory0_ram_dout0[408]), 
        .B(n21597), .Y(n13108) );
  sky130_fd_sc_hd__nand2_1 U19797 ( .A(j202_soc_core_memory0_ram_dout0[56]), 
        .B(n21604), .Y(n13109) );
  sky130_fd_sc_hd__nand2_1 U19798 ( .A(j202_soc_core_memory0_ram_dout0[280]), 
        .B(n21605), .Y(n13110) );
  sky130_fd_sc_hd__nand2_1 U19799 ( .A(j202_soc_core_memory0_ram_dout0[248]), 
        .B(n21735), .Y(n13111) );
  sky130_fd_sc_hd__nand2_1 U19800 ( .A(j202_soc_core_memory0_ram_dout0[88]), 
        .B(n21734), .Y(n13112) );
  sky130_fd_sc_hd__nand2_1 U19801 ( .A(j202_soc_core_memory0_ram_dout0[24]), 
        .B(n21733), .Y(n13113) );
  sky130_fd_sc_hd__nand2_1 U19802 ( .A(j202_soc_core_memory0_ram_dout0[216]), 
        .B(n21732), .Y(n13114) );
  sky130_fd_sc_hd__nand4_1 U19803 ( .A(n13116), .B(n12436), .C(n29015), .D(
        n11873), .Y(n23950) );
  sky130_fd_sc_hd__nand2_1 U19804 ( .A(j202_soc_core_memory0_ram_dout0[448]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n13117) );
  sky130_fd_sc_hd__nand2_1 U19805 ( .A(j202_soc_core_memory0_ram_dout0[416]), 
        .B(n21598), .Y(n13118) );
  sky130_fd_sc_hd__nand2_1 U19806 ( .A(j202_soc_core_memory0_ram_dout0[160]), 
        .B(n21590), .Y(n13119) );
  sky130_fd_sc_hd__nand2_1 U19807 ( .A(n21435), .B(n21436), .Y(n22704) );
  sky130_fd_sc_hd__nand3_2 U19808 ( .A(n13129), .B(n13126), .C(n13120), .Y(
        n17107) );
  sky130_fd_sc_hd__nand4_1 U19809 ( .A(n13125), .B(n13124), .C(n13123), .D(
        n13122), .Y(n13121) );
  sky130_fd_sc_hd__nand2_1 U19810 ( .A(j202_soc_core_memory0_ram_dout0[59]), 
        .B(n21604), .Y(n13122) );
  sky130_fd_sc_hd__nand2_1 U19811 ( .A(j202_soc_core_memory0_ram_dout0[251]), 
        .B(n21735), .Y(n13123) );
  sky130_fd_sc_hd__nand2_1 U19812 ( .A(j202_soc_core_memory0_ram_dout0[187]), 
        .B(n21590), .Y(n13124) );
  sky130_fd_sc_hd__nand2_1 U19813 ( .A(j202_soc_core_memory0_ram_dout0[219]), 
        .B(n21732), .Y(n13125) );
  sky130_fd_sc_hd__nand2_1 U19814 ( .A(j202_soc_core_memory0_ram_dout0[315]), 
        .B(n21603), .Y(n13127) );
  sky130_fd_sc_hd__nand2_1 U19815 ( .A(j202_soc_core_memory0_ram_dout0[155]), 
        .B(n21592), .Y(n13128) );
  sky130_fd_sc_hd__nand4_1 U19816 ( .A(n13134), .B(n13133), .C(n13132), .D(
        n13131), .Y(n13130) );
  sky130_fd_sc_hd__nand2_1 U19817 ( .A(j202_soc_core_memory0_ram_dout0[91]), 
        .B(n21734), .Y(n13131) );
  sky130_fd_sc_hd__nand2_1 U19818 ( .A(j202_soc_core_memory0_ram_dout0[123]), 
        .B(n21591), .Y(n13132) );
  sky130_fd_sc_hd__nand2_1 U19819 ( .A(j202_soc_core_memory0_ram_dout0[475]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n13133) );
  sky130_fd_sc_hd__nand2_1 U19820 ( .A(j202_soc_core_memory0_ram_dout0[283]), 
        .B(n21605), .Y(n13134) );
  sky130_fd_sc_hd__nand4_1 U19821 ( .A(n13139), .B(n13138), .C(n13137), .D(
        n13136), .Y(n13135) );
  sky130_fd_sc_hd__nand2_1 U19822 ( .A(j202_soc_core_memory0_ram_dout0[379]), 
        .B(n21596), .Y(n13136) );
  sky130_fd_sc_hd__nand2_1 U19823 ( .A(j202_soc_core_memory0_ram_dout0[347]), 
        .B(n21593), .Y(n13137) );
  sky130_fd_sc_hd__nand2_1 U19824 ( .A(j202_soc_core_memory0_ram_dout0[411]), 
        .B(n21597), .Y(n13138) );
  sky130_fd_sc_hd__nand2_1 U19825 ( .A(j202_soc_core_memory0_ram_dout0[27]), 
        .B(n21733), .Y(n13139) );
  sky130_fd_sc_hd__nand2_1 U19828 ( .A(j202_soc_core_memory0_ram_dout0[338]), 
        .B(n21593), .Y(n13154) );
  sky130_fd_sc_hd__nor2_1 U19830 ( .A(n21778), .B(n20562), .Y(n13156) );
  sky130_fd_sc_hd__inv_2 U19832 ( .A(n24354), .Y(n24257) );
  sky130_fd_sc_hd__nand4_1 U19833 ( .A(n24454), .B(n24456), .C(n24455), .D(
        n13159), .Y(n24457) );
  sky130_fd_sc_hd__nand2_1 U19834 ( .A(n13163), .B(n12234), .Y(n13235) );
  sky130_fd_sc_hd__nand4_1 U19835 ( .A(n12257), .B(n11059), .C(n12148), .D(
        n12155), .Y(n13163) );
  sky130_fd_sc_hd__nand2_1 U19836 ( .A(j202_soc_core_memory0_ram_dout0[267]), 
        .B(n21605), .Y(n13164) );
  sky130_fd_sc_hd__nand2_1 U19837 ( .A(j202_soc_core_memory0_ram_dout0[235]), 
        .B(n21735), .Y(n13165) );
  sky130_fd_sc_hd__nand2_1 U19838 ( .A(j202_soc_core_memory0_ram_dout0[363]), 
        .B(n21596), .Y(n13166) );
  sky130_fd_sc_hd__nand2_1 U19839 ( .A(j202_soc_core_memory0_ram_dout0[75]), 
        .B(n21734), .Y(n13167) );
  sky130_fd_sc_hd__nand2_1 U19840 ( .A(j202_soc_core_memory0_ram_dout0[299]), 
        .B(n21603), .Y(n13168) );
  sky130_fd_sc_hd__nand2_1 U19841 ( .A(j202_soc_core_memory0_ram_dout0[11]), 
        .B(n21733), .Y(n13169) );
  sky130_fd_sc_hd__nand2_1 U19842 ( .A(j202_soc_core_memory0_ram_dout0[43]), 
        .B(n21604), .Y(n13170) );
  sky130_fd_sc_hd__nand2_1 U19843 ( .A(j202_soc_core_memory0_ram_dout0[171]), 
        .B(n21590), .Y(n13171) );
  sky130_fd_sc_hd__nand2_1 U19844 ( .A(j202_soc_core_memory0_ram_dout0[203]), 
        .B(n21732), .Y(n13172) );
  sky130_fd_sc_hd__nand2_1 U19845 ( .A(j202_soc_core_memory0_ram_dout0[107]), 
        .B(n21591), .Y(n13173) );
  sky130_fd_sc_hd__nand2_1 U19846 ( .A(j202_soc_core_memory0_ram_dout0[139]), 
        .B(n21592), .Y(n13174) );
  sky130_fd_sc_hd__nand2_1 U19847 ( .A(j202_soc_core_memory0_ram_dout0[395]), 
        .B(n21597), .Y(n13175) );
  sky130_fd_sc_hd__nand2_1 U19848 ( .A(j202_soc_core_memory0_ram_dout0[331]), 
        .B(n21593), .Y(n13176) );
  sky130_fd_sc_hd__nand2_1 U19849 ( .A(j202_soc_core_memory0_ram_dout0[427]), 
        .B(n21598), .Y(n13177) );
  sky130_fd_sc_hd__nand2_1 U19850 ( .A(n24435), .B(n13179), .Y(n24418) );
  sky130_fd_sc_hd__o21a_1 U19851 ( .A1(n29075), .A2(n13179), .B1(n27772), .X(
        n24425) );
  sky130_fd_sc_hd__nand4_1 U19852 ( .A(n27895), .B(n27894), .C(n27893), .D(
        n13179), .Y(n27896) );
  sky130_fd_sc_hd__nand2_1 U19856 ( .A(j202_soc_core_memory0_ram_dout0[354]), 
        .B(n21596), .Y(n13183) );
  sky130_fd_sc_hd__nand2_1 U19857 ( .A(j202_soc_core_memory0_ram_dout0[450]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n13184) );
  sky130_fd_sc_hd__nand2_1 U19858 ( .A(j202_soc_core_memory0_ram_dout0[418]), 
        .B(n21598), .Y(n13185) );
  sky130_fd_sc_hd__nand2_1 U19859 ( .A(n27522), .B(n12291), .Y(n10493) );
  sky130_fd_sc_hd__nand2_1 U19860 ( .A(n12439), .B(n27980), .Y(n13186) );
  sky130_fd_sc_hd__inv_2 U19861 ( .A(n13229), .Y(n13190) );
  sky130_fd_sc_hd__nand2_1 U19862 ( .A(n11767), .B(n27980), .Y(n23959) );
  sky130_fd_sc_hd__nand2_1 U19863 ( .A(n11767), .B(n11793), .Y(n23158) );
  sky130_fd_sc_hd__inv_2 U19864 ( .A(n29070), .Y(n27298) );
  sky130_fd_sc_hd__nand3_1 U19865 ( .A(n27557), .B(n27565), .C(n13194), .Y(
        n27559) );
  sky130_fd_sc_hd__nand4_1 U19866 ( .A(n13208), .B(n13207), .C(n17338), .D(
        n13195), .Y(n13206) );
  sky130_fd_sc_hd__nand2_1 U19867 ( .A(j202_soc_core_memory0_ram_dout0[327]), 
        .B(n21593), .Y(n13195) );
  sky130_fd_sc_hd__nand2_1 U19868 ( .A(n24089), .B(n26443), .Y(n13197) );
  sky130_fd_sc_hd__nand2_1 U19869 ( .A(n13201), .B(n13200), .Y(n18698) );
  sky130_fd_sc_hd__nand2_1 U19870 ( .A(n13203), .B(n13202), .Y(n18572) );
  sky130_fd_sc_hd__nand2_1 U19871 ( .A(n18247), .B(n18246), .Y(n13202) );
  sky130_fd_sc_hd__nand2_1 U19873 ( .A(n18594), .B(n18595), .Y(n13204) );
  sky130_fd_sc_hd__nand2_1 U19875 ( .A(j202_soc_core_memory0_ram_dout0[295]), 
        .B(n21603), .Y(n13207) );
  sky130_fd_sc_hd__nand2_1 U19876 ( .A(j202_soc_core_memory0_ram_dout0[7]), 
        .B(n21733), .Y(n13208) );
  sky130_fd_sc_hd__nand4_1 U19877 ( .A(n13213), .B(n13212), .C(n13210), .D(
        n13211), .Y(n13209) );
  sky130_fd_sc_hd__nand2_1 U19878 ( .A(j202_soc_core_memory0_ram_dout0[167]), 
        .B(n21590), .Y(n13210) );
  sky130_fd_sc_hd__nand2_1 U19879 ( .A(j202_soc_core_memory0_ram_dout0[39]), 
        .B(n21604), .Y(n13211) );
  sky130_fd_sc_hd__nand2_1 U19880 ( .A(j202_soc_core_memory0_ram_dout0[231]), 
        .B(n21735), .Y(n13212) );
  sky130_fd_sc_hd__nand2_1 U19881 ( .A(j202_soc_core_memory0_ram_dout0[391]), 
        .B(n21597), .Y(n13213) );
  sky130_fd_sc_hd__nand2_1 U19882 ( .A(j202_soc_core_memory0_ram_dout0[239]), 
        .B(n21735), .Y(n13215) );
  sky130_fd_sc_hd__nand2_1 U19883 ( .A(j202_soc_core_memory0_ram_dout0[79]), 
        .B(n21734), .Y(n13216) );
  sky130_fd_sc_hd__nand2_1 U19884 ( .A(j202_soc_core_memory0_ram_dout0[303]), 
        .B(n21603), .Y(n13217) );
  sky130_fd_sc_hd__nand2_1 U19885 ( .A(j202_soc_core_memory0_ram_dout0[111]), 
        .B(n21591), .Y(n13218) );
  sky130_fd_sc_hd__nand2_1 U19886 ( .A(j202_soc_core_memory0_ram_dout0[367]), 
        .B(n21596), .Y(n13219) );
  sky130_fd_sc_hd__nand2_1 U19887 ( .A(j202_soc_core_memory0_ram_dout0[143]), 
        .B(n21592), .Y(n13220) );
  sky130_fd_sc_hd__nand2_1 U19888 ( .A(j202_soc_core_memory0_ram_dout0[463]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n13221) );
  sky130_fd_sc_hd__nand2_1 U19889 ( .A(j202_soc_core_memory0_ram_dout0[207]), 
        .B(n21732), .Y(n13222) );
  sky130_fd_sc_hd__and2_0 U19890 ( .A(n21677), .B(n18978), .X(n13223) );
  sky130_fd_sc_hd__nand2_1 U19891 ( .A(j202_soc_core_memory0_ram_dout0[13]), 
        .B(n21733), .Y(n13225) );
  sky130_fd_sc_hd__nand2_1 U19892 ( .A(n12475), .B(n11626), .Y(n13227) );
  sky130_fd_sc_hd__o21ai_1 U19893 ( .A1(n27977), .A2(n27976), .B1(n27975), .Y(
        n10568) );
  sky130_fd_sc_hd__nand2_1 U19894 ( .A(n13232), .B(n27949), .Y(n27976) );
  sky130_fd_sc_hd__nand3_1 U19895 ( .A(n11072), .B(n24110), .C(n12395), .Y(
        n13239) );
  sky130_fd_sc_hd__nand2b_1 U19896 ( .A_N(n27980), .B(n24093), .Y(n13240) );
  sky130_fd_sc_hd__nand2_1 U19897 ( .A(n16634), .B(n16631), .Y(n13241) );
  sky130_fd_sc_hd__nand3_1 U19898 ( .A(n16633), .B(n16632), .C(n16630), .Y(
        n13242) );
  sky130_fd_sc_hd__nand2_1 U19899 ( .A(n13258), .B(n13255), .Y(n13247) );
  sky130_fd_sc_hd__nand2_1 U19900 ( .A(n16634), .B(n16632), .Y(n13248) );
  sky130_fd_sc_hd__nand3_1 U19901 ( .A(n13252), .B(n16628), .C(n13253), .Y(
        n13250) );
  sky130_fd_sc_hd__nand2_1 U19902 ( .A(j202_soc_core_memory0_ram_dout0[444]), 
        .B(n21598), .Y(n13252) );
  sky130_fd_sc_hd__and2_0 U19903 ( .A(n16627), .B(n16646), .X(n13253) );
  sky130_fd_sc_hd__nand2_1 U19904 ( .A(j202_soc_core_memory0_ram_dout0[60]), 
        .B(n21604), .Y(n13255) );
  sky130_fd_sc_hd__nand2_1 U19905 ( .A(j202_soc_core_memory0_ram_dout0[316]), 
        .B(n21603), .Y(n13256) );
  sky130_fd_sc_hd__nand2_1 U19906 ( .A(j202_soc_core_memory0_ram_dout0[28]), 
        .B(n21733), .Y(n13257) );
  sky130_fd_sc_hd__nand2_1 U19907 ( .A(j202_soc_core_memory0_ram_dout0[252]), 
        .B(n21735), .Y(n13258) );
  sky130_fd_sc_hd__nand2_1 U19908 ( .A(n14979), .B(n12283), .Y(n13261) );
  sky130_fd_sc_hd__nand4_1 U19909 ( .A(n20402), .B(n20406), .C(n20403), .D(
        n20405), .Y(n13260) );
  sky130_fd_sc_hd__nand4_1 U19911 ( .A(n19332), .B(n19333), .C(n19331), .D(
        n19330), .Y(n13266) );
  sky130_fd_sc_hd__nand3b_1 U19912 ( .A_N(n13263), .B(n19326), .C(n19327), .Y(
        n13267) );
  sky130_fd_sc_hd__nand2_1 U19913 ( .A(n19329), .B(n19328), .Y(n13263) );
  sky130_fd_sc_hd__nand2_1 U19914 ( .A(n21781), .B(n13343), .Y(n21782) );
  sky130_fd_sc_hd__nand2_1 U19915 ( .A(n13265), .B(n13264), .Y(n21781) );
  sky130_fd_sc_hd__o2bb2ai_1 U19916 ( .B1(n27226), .B2(n27451), .A1_N(n12644), 
        .A2_N(n26379), .Y(j202_soc_core_j22_cpu_rf_N3140) );
  sky130_fd_sc_hd__nand2_1 U19917 ( .A(n12277), .B(n13269), .Y(n13268) );
  sky130_fd_sc_hd__inv_2 U19918 ( .A(n13272), .Y(n13271) );
  sky130_fd_sc_hd__a22oi_2 U19920 ( .A1(j202_soc_core_memory0_ram_dout0[449]), 
        .A2(j202_soc_core_memory0_ram_dout0_sel[14]), .B1(n21598), .B2(
        j202_soc_core_memory0_ram_dout0[417]), .Y(n19929) );
  sky130_fd_sc_hd__nand3_1 U19921 ( .A(n20827), .B(n20826), .C(n12248), .Y(
        n21519) );
  sky130_fd_sc_hd__clkinv_1 U19922 ( .A(n20804), .Y(n20807) );
  sky130_fd_sc_hd__clkinv_1 U19923 ( .A(n20201), .Y(n20204) );
  sky130_fd_sc_hd__nand2b_2 U19924 ( .A_N(n20201), .B(n17274), .Y(n20384) );
  sky130_fd_sc_hd__nand3_2 U19926 ( .A(n14741), .B(n14740), .C(n13339), .Y(
        n27354) );
  sky130_fd_sc_hd__o22a_1 U19927 ( .A1(n15326), .A2(n15557), .B1(n15325), .B2(
        n15708), .X(n15327) );
  sky130_fd_sc_hd__inv_2 U19928 ( .A(n16533), .Y(n17108) );
  sky130_fd_sc_hd__inv_2 U19929 ( .A(n12174), .Y(n16449) );
  sky130_fd_sc_hd__a2bb2oi_1 U19930 ( .B1(n26077), .B2(n26726), .A1_N(n26704), 
        .A2_N(n22729), .Y(n19029) );
  sky130_fd_sc_hd__and4_1 U19931 ( .A(n13773), .B(n13772), .C(n13771), .D(
        n13770), .X(n13785) );
  sky130_fd_sc_hd__nor2_1 U19932 ( .A(n13783), .B(n13782), .Y(n13784) );
  sky130_fd_sc_hd__a21oi_1 U19933 ( .A1(n22944), .A2(n22800), .B1(n22799), .Y(
        n22801) );
  sky130_fd_sc_hd__nor4_1 U19934 ( .A(n21611), .B(n21704), .C(n21131), .D(
        n21130), .Y(n21281) );
  sky130_fd_sc_hd__and3_1 U19935 ( .A(n12180), .B(n21648), .C(n20747), .X(
        n19295) );
  sky130_fd_sc_hd__buf_4 U19936 ( .A(n13794), .X(n23098) );
  sky130_fd_sc_hd__nand2_1 U19938 ( .A(n24500), .B(n22627), .Y(n26515) );
  sky130_fd_sc_hd__nand2_1 U19939 ( .A(n13387), .B(n20787), .Y(n17282) );
  sky130_fd_sc_hd__nand3_2 U19940 ( .A(n14005), .B(n14004), .C(n14003), .Y(
        n27443) );
  sky130_fd_sc_hd__nand3_2 U19941 ( .A(n13921), .B(n12215), .C(n13920), .Y(
        n26711) );
  sky130_fd_sc_hd__nand2_1 U19942 ( .A(n17193), .B(n17192), .Y(n20117) );
  sky130_fd_sc_hd__nor4_1 U19943 ( .A(n19830), .B(n20916), .C(n19900), .D(
        n20179), .Y(n19893) );
  sky130_fd_sc_hd__nand3_2 U19944 ( .A(n14085), .B(n14084), .C(n14083), .Y(
        n26603) );
  sky130_fd_sc_hd__a21oi_1 U19945 ( .A1(n21347), .A2(n21346), .B1(n21331), .Y(
        n21336) );
  sky130_fd_sc_hd__nand3_2 U19946 ( .A(n12210), .B(n14174), .C(n14173), .Y(
        n26725) );
  sky130_fd_sc_hd__inv_2 U19948 ( .A(n16436), .Y(n14755) );
  sky130_fd_sc_hd__nand3_2 U19949 ( .A(n15057), .B(n15056), .C(n15055), .Y(
        n26061) );
  sky130_fd_sc_hd__nor2_1 U19950 ( .A(n20363), .B(n20046), .Y(n20247) );
  sky130_fd_sc_hd__inv_2 U19951 ( .A(n17190), .Y(n20363) );
  sky130_fd_sc_hd__nand3_2 U19952 ( .A(n15135), .B(n13309), .C(n15134), .Y(
        n27183) );
  sky130_fd_sc_hd__a2bb2oi_1 U19953 ( .B1(n13752), .B2(
        j202_soc_core_intr_vec__3_), .A1_N(n10978), .A2_N(n14466), .Y(n13916)
         );
  sky130_fd_sc_hd__nor2_2 U19954 ( .A(n10921), .B(n14466), .Y(n16436) );
  sky130_fd_sc_hd__nor2_1 U19955 ( .A(n14031), .B(n14030), .Y(n14032) );
  sky130_fd_sc_hd__a21oi_1 U19956 ( .A1(j202_soc_core_j22_cpu_rf_gpr[0]), .A2(
        n16369), .B1(n14021), .Y(n14033) );
  sky130_fd_sc_hd__fah_1 U19957 ( .A(n18728), .B(n18727), .CI(n18726), .COUT(
        n18783), .SUM(n18744) );
  sky130_fd_sc_hd__nand2_1 U19958 ( .A(n28986), .B(n27824), .Y(n24189) );
  sky130_fd_sc_hd__nand3_2 U19959 ( .A(n15081), .B(n15080), .C(n15079), .Y(
        n26508) );
  sky130_fd_sc_hd__nor2_2 U19960 ( .A(n17289), .B(n17274), .Y(n16706) );
  sky130_fd_sc_hd__nor2_1 U19961 ( .A(n13623), .B(n13622), .Y(n13648) );
  sky130_fd_sc_hd__a21oi_2 U19962 ( .A1(n14835), .A2(n21012), .B1(n14834), .Y(
        n15413) );
  sky130_fd_sc_hd__o21ai_2 U19963 ( .A1(n22511), .A2(n20999), .B1(n21000), .Y(
        n21012) );
  sky130_fd_sc_hd__nand3_1 U19964 ( .A(n27822), .B(n24425), .C(n24424), .Y(
        n24438) );
  sky130_fd_sc_hd__nand3_1 U19966 ( .A(n22563), .B(n23824), .C(n23850), .Y(
        n24582) );
  sky130_fd_sc_hd__fah_1 U19967 ( .A(n18779), .B(n18778), .CI(n18777), .COUT(
        n18850), .SUM(n18839) );
  sky130_fd_sc_hd__a21oi_1 U19968 ( .A1(n22944), .A2(n22191), .B1(n22190), .Y(
        n22192) );
  sky130_fd_sc_hd__nand3_2 U19969 ( .A(n14614), .B(n12202), .C(n14613), .Y(
        n26728) );
  sky130_fd_sc_hd__inv_2 U19970 ( .A(n13680), .Y(n23126) );
  sky130_fd_sc_hd__nor2_1 U19971 ( .A(n19841), .B(n20218), .Y(n20329) );
  sky130_fd_sc_hd__nand2_1 U19972 ( .A(n19112), .B(n20117), .Y(n20218) );
  sky130_fd_sc_hd__inv_2 U19973 ( .A(n13667), .Y(n23076) );
  sky130_fd_sc_hd__nand2_1 U19974 ( .A(n17301), .B(n20623), .Y(n17211) );
  sky130_fd_sc_hd__nand3_2 U19975 ( .A(n14685), .B(n13308), .C(n14684), .Y(
        n27045) );
  sky130_fd_sc_hd__a21oi_1 U19976 ( .A1(n11774), .A2(n26863), .B1(n24654), .Y(
        n24691) );
  sky130_fd_sc_hd__nor2_2 U19977 ( .A(n12137), .B(
        j202_soc_core_bootrom_00_address_w[4]), .Y(n17273) );
  sky130_fd_sc_hd__nor2_2 U19978 ( .A(n17277), .B(
        j202_soc_core_bootrom_00_address_w[4]), .Y(n16616) );
  sky130_fd_sc_hd__o22ai_1 U19979 ( .A1(n18711), .A2(n18710), .B1(n18657), 
        .B2(n18712), .Y(n18755) );
  sky130_fd_sc_hd__nor2_1 U19980 ( .A(n29015), .B(n27523), .Y(n23584) );
  sky130_fd_sc_hd__nand2_1 U19982 ( .A(n17161), .B(n20787), .Y(n17168) );
  sky130_fd_sc_hd__nand2_1 U19983 ( .A(n28999), .B(n24225), .Y(n24208) );
  sky130_fd_sc_hd__fah_1 U19984 ( .A(n18788), .B(n18787), .CI(n18786), .COUT(
        n18837), .SUM(n18836) );
  sky130_fd_sc_hd__a21oi_1 U19986 ( .A1(n22944), .A2(n22943), .B1(n22942), .Y(
        n22945) );
  sky130_fd_sc_hd__o22a_1 U19987 ( .A1(n22318), .A2(n22317), .B1(n22978), .B2(
        n22316), .X(n22320) );
  sky130_fd_sc_hd__fah_1 U19988 ( .A(n18536), .B(n18535), .CI(n18534), .COUT(
        n18733), .SUM(n18528) );
  sky130_fd_sc_hd__nand2_1 U19989 ( .A(n21854), .B(n16513), .Y(n13975) );
  sky130_fd_sc_hd__o21ai_1 U19990 ( .A1(n22946), .A2(n22897), .B1(n22945), .Y(
        n22947) );
  sky130_fd_sc_hd__nand3_1 U19991 ( .A(n24135), .B(n24134), .C(n24133), .Y(
        n24637) );
  sky130_fd_sc_hd__fah_1 U19992 ( .A(n18743), .B(n18742), .CI(n18741), .COUT(
        n18745), .SUM(n18805) );
  sky130_fd_sc_hd__nand2_1 U19993 ( .A(n22174), .B(n22173), .Y(n26472) );
  sky130_fd_sc_hd__o2bb2ai_1 U19994 ( .B1(n27228), .B2(n27524), .A1_N(n27228), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N3168) );
  sky130_fd_sc_hd__o2bb2ai_1 U19995 ( .B1(n27225), .B2(n27524), .A1_N(n27225), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N2946) );
  sky130_fd_sc_hd__o2bb2ai_1 U19996 ( .B1(n27333), .B2(n27524), .A1_N(n26371), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N3057) );
  sky130_fd_sc_hd__o2bb2ai_1 U19997 ( .B1(n27226), .B2(n27524), .A1_N(n26379), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N3131) );
  sky130_fd_sc_hd__o2bb2ai_1 U19998 ( .B1(n27575), .B2(n27524), .A1_N(n11109), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N3094) );
  sky130_fd_sc_hd__o2bb2ai_1 U19999 ( .B1(n27219), .B2(n27524), .A1_N(n26369), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N2983) );
  sky130_fd_sc_hd__o2bb2ai_1 U20000 ( .B1(n27221), .B2(n27524), .A1_N(n26374), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N2872) );
  sky130_fd_sc_hd__fah_1 U20001 ( .A(n18386), .B(n18385), .CI(n18384), .COUT(
        n18582), .SUM(n18570) );
  sky130_fd_sc_hd__a21oi_2 U20002 ( .A1(n21516), .A2(n12173), .B1(n17841), .Y(
        n18997) );
  sky130_fd_sc_hd__nor3_1 U20003 ( .A(n27919), .B(n24409), .C(n24410), .Y(
        n24411) );
  sky130_fd_sc_hd__a21o_1 U20004 ( .A1(n17786), .A2(n17771), .B1(n17504), .X(
        n17932) );
  sky130_fd_sc_hd__fah_1 U20005 ( .A(n18347), .B(n18346), .CI(n18345), .COUT(
        n18394), .SUM(n18585) );
  sky130_fd_sc_hd__nand2_2 U20006 ( .A(n21843), .B(n29535), .Y(n24383) );
  sky130_fd_sc_hd__nand2_1 U20007 ( .A(n24382), .B(n24380), .Y(n24060) );
  sky130_fd_sc_hd__nand3_2 U20008 ( .A(n21841), .B(n21840), .C(n21839), .Y(
        n22458) );
  sky130_fd_sc_hd__nand3_2 U20009 ( .A(n13760), .B(n12203), .C(n13759), .Y(
        n22723) );
  sky130_fd_sc_hd__fah_1 U20010 ( .A(n18704), .B(n18703), .CI(n18702), .COUT(
        n18766), .SUM(n18723) );
  sky130_fd_sc_hd__nand2b_1 U20011 ( .A_N(n25547), .B(n26802), .Y(n25559) );
  sky130_fd_sc_hd__fah_1 U20012 ( .A(n18635), .B(n18634), .CI(n18633), .COUT(
        n18640), .SUM(n18772) );
  sky130_fd_sc_hd__fah_1 U20013 ( .A(n18684), .B(n18683), .CI(n18682), .COUT(
        n18735), .SUM(n18732) );
  sky130_fd_sc_hd__nand2_4 U20014 ( .A(n17395), .B(n17394), .Y(n17802) );
  sky130_fd_sc_hd__fah_1 U20016 ( .A(n18392), .B(n18391), .CI(n18390), .COUT(
        n18395), .SUM(n18581) );
  sky130_fd_sc_hd__nand2_1 U20017 ( .A(n21886), .B(n23042), .Y(n25289) );
  sky130_fd_sc_hd__o2bb2ai_1 U20018 ( .B1(n26378), .B2(n27524), .A1_N(n26378), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N3242) );
  sky130_fd_sc_hd__o2bb2ai_1 U20019 ( .B1(n27223), .B2(n27524), .A1_N(n27223), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N3020) );
  sky130_fd_sc_hd__nand2_1 U20020 ( .A(n15308), .B(n13294), .Y(n15545) );
  sky130_fd_sc_hd__fah_1 U20021 ( .A(n17881), .B(n17880), .CI(n17879), .COUT(
        n17886), .SUM(n17882) );
  sky130_fd_sc_hd__o22a_2 U20022 ( .A1(n22713), .A2(n26530), .B1(n21915), .B2(
        n26537), .X(n21817) );
  sky130_fd_sc_hd__nor2b_1 U20023 ( .B_N(n18353), .A(n17972), .Y(n17784) );
  sky130_fd_sc_hd__fah_1 U20024 ( .A(n18006), .B(n18005), .CI(n18004), .COUT(
        n18039), .SUM(n18014) );
  sky130_fd_sc_hd__fah_1 U20025 ( .A(n17935), .B(n17934), .CI(n17933), .COUT(
        n17993), .SUM(n17953) );
  sky130_fd_sc_hd__fah_1 U20026 ( .A(n18785), .B(n18784), .CI(n18783), .COUT(
        n18835), .SUM(n18834) );
  sky130_fd_sc_hd__nand2_1 U20027 ( .A(n19581), .B(n19580), .Y(n19585) );
  sky130_fd_sc_hd__fah_1 U20028 ( .A(n17777), .B(n17776), .CI(n17775), .COUT(
        n17852), .SUM(n17845) );
  sky130_fd_sc_hd__fah_1 U20029 ( .A(n17683), .B(n17682), .CI(n17681), .COUT(
        n17904), .SUM(n17673) );
  sky130_fd_sc_hd__nand2_2 U20030 ( .A(n17170), .B(n19355), .Y(n21206) );
  sky130_fd_sc_hd__o21ai_1 U20031 ( .A1(n11128), .A2(n23044), .B1(n23043), .Y(
        n23072) );
  sky130_fd_sc_hd__o21ai_2 U20032 ( .A1(n21821), .A2(n21824), .B1(n21822), .Y(
        n21516) );
  sky130_fd_sc_hd__o2bb2ai_1 U20033 ( .B1(n27215), .B2(n27524), .A1_N(n27215), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N2909) );
  sky130_fd_sc_hd__o2bb2ai_1 U20034 ( .B1(n11141), .B2(n27524), .A1_N(n11141), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N2687) );
  sky130_fd_sc_hd__o2bb2ai_1 U20035 ( .B1(n27211), .B2(n27524), .A1_N(n27211), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N3205) );
  sky130_fd_sc_hd__o2bb2ai_1 U20036 ( .B1(n27524), .B2(n26899), .A1_N(n26383), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N3318) );
  sky130_fd_sc_hd__o2bb2ai_1 U20037 ( .B1(n27209), .B2(n27524), .A1_N(n26360), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N2724) );
  sky130_fd_sc_hd__o2bb2ai_1 U20038 ( .B1(n27466), .B2(n27524), .A1_N(n25818), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N2761) );
  sky130_fd_sc_hd__o2bb2ai_1 U20039 ( .B1(n27213), .B2(n27524), .A1_N(n26362), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N2798) );
  sky130_fd_sc_hd__fah_1 U20040 ( .A(n17435), .B(n17434), .CI(n17433), .COUT(
        n17477), .SUM(n17571) );
  sky130_fd_sc_hd__fah_1 U20041 ( .A(n17780), .B(n17779), .CI(n17778), .COUT(
        n17844), .SUM(n17836) );
  sky130_fd_sc_hd__fah_1 U20042 ( .A(n17906), .B(n17904), .CI(n17905), .COUT(
        n17911), .SUM(n17898) );
  sky130_fd_sc_hd__nand2_1 U20043 ( .A(n17273), .B(n19381), .Y(n20804) );
  sky130_fd_sc_hd__fah_1 U20044 ( .A(n17967), .B(n17966), .CI(n17965), .COUT(
        n18000), .SUM(n17956) );
  sky130_fd_sc_hd__fah_1 U20045 ( .A(n17503), .B(n17502), .CI(n17501), .COUT(
        n17987), .SUM(n17483) );
  sky130_fd_sc_hd__o2bb2ai_1 U20046 ( .B1(n19719), .B2(n19735), .A1_N(n19718), 
        .A2_N(n19753), .Y(n19732) );
  sky130_fd_sc_hd__mux2_4 U20047 ( .A0(j202_soc_core_intc_core_00_rg_ipr[44]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[40]), .S(n26826), .X(n19746) );
  sky130_fd_sc_hd__fah_1 U20048 ( .A(n17665), .B(n17664), .CI(n17663), .COUT(
        n17681), .SUM(n17685) );
  sky130_fd_sc_hd__fah_1 U20049 ( .A(n18364), .B(n18363), .CI(n18362), .COUT(
        n18415), .SUM(n18357) );
  sky130_fd_sc_hd__o21ai_2 U20050 ( .A1(n26802), .A2(n24636), .B1(n22768), .Y(
        n22014) );
  sky130_fd_sc_hd__fah_1 U20051 ( .A(n18331), .B(n18330), .CI(n18329), .COUT(
        n18559), .SUM(n18567) );
  sky130_fd_sc_hd__xnor2_2 U20052 ( .A(n17396), .B(n21887), .Y(n17399) );
  sky130_fd_sc_hd__nor2b_1 U20053 ( .B_N(n18353), .A(n18151), .Y(n17725) );
  sky130_fd_sc_hd__a21o_1 U20054 ( .A1(n18148), .A2(n18151), .B1(n18150), .X(
        n18188) );
  sky130_fd_sc_hd__o21ai_1 U20056 ( .A1(n19744), .A2(n19746), .B1(n19687), .Y(
        n19688) );
  sky130_fd_sc_hd__nand2_2 U20057 ( .A(n19797), .B(n12205), .Y(n19799) );
  sky130_fd_sc_hd__o21ai_2 U20058 ( .A1(n17842), .A2(n18997), .B1(n18994), .Y(
        n21967) );
  sky130_fd_sc_hd__a21oi_2 U20059 ( .A1(n19608), .A2(n19607), .B1(n19606), .Y(
        n26837) );
  sky130_fd_sc_hd__nand2_1 U20060 ( .A(n19604), .B(n19603), .Y(n19608) );
  sky130_fd_sc_hd__o2bb2ai_1 U20061 ( .B1(n11141), .B2(n25157), .A1_N(n11141), 
        .A2_N(n12385), .Y(j202_soc_core_j22_cpu_rf_N2708) );
  sky130_fd_sc_hd__o2bb2ai_1 U20062 ( .B1(n27215), .B2(n25157), .A1_N(n27215), 
        .A2_N(n25158), .Y(j202_soc_core_j22_cpu_rf_N2930) );
  sky130_fd_sc_hd__o2bb2ai_1 U20063 ( .B1(n27211), .B2(n25157), .A1_N(n27211), 
        .A2_N(n12385), .Y(j202_soc_core_j22_cpu_rf_N3226) );
  sky130_fd_sc_hd__o2bb2ai_1 U20064 ( .B1(n27225), .B2(n25157), .A1_N(n27225), 
        .A2_N(n12385), .Y(j202_soc_core_j22_cpu_rf_N2967) );
  sky130_fd_sc_hd__o2bb2ai_1 U20065 ( .B1(n27228), .B2(n25157), .A1_N(n27228), 
        .A2_N(n25158), .Y(j202_soc_core_j22_cpu_rf_N3189) );
  sky130_fd_sc_hd__o2bb2ai_1 U20066 ( .B1(n26378), .B2(n25157), .A1_N(n26378), 
        .A2_N(n12385), .Y(j202_soc_core_j22_cpu_rf_N3263) );
  sky130_fd_sc_hd__o2bb2ai_1 U20067 ( .B1(n26899), .B2(n25157), .A1_N(n26383), 
        .A2_N(n12385), .Y(j202_soc_core_j22_cpu_rf_N3339) );
  sky130_fd_sc_hd__o2bb2ai_1 U20068 ( .B1(n27217), .B2(n25157), .A1_N(n25819), 
        .A2_N(n25158), .Y(j202_soc_core_j22_cpu_rf_N2856) );
  sky130_fd_sc_hd__o2bb2ai_1 U20069 ( .B1(n27226), .B2(n25157), .A1_N(n26379), 
        .A2_N(n12385), .Y(j202_soc_core_j22_cpu_rf_N3152) );
  sky130_fd_sc_hd__o2bb2ai_1 U20070 ( .B1(n27213), .B2(n25157), .A1_N(n26362), 
        .A2_N(n25158), .Y(j202_soc_core_j22_cpu_rf_N2819) );
  sky130_fd_sc_hd__o2bb2ai_1 U20071 ( .B1(n27221), .B2(n25157), .A1_N(n26374), 
        .A2_N(n25158), .Y(j202_soc_core_j22_cpu_rf_N2893) );
  sky130_fd_sc_hd__o2bb2ai_1 U20072 ( .B1(n27466), .B2(n25157), .A1_N(n25818), 
        .A2_N(n25158), .Y(j202_soc_core_j22_cpu_rf_N2782) );
  sky130_fd_sc_hd__o2bb2ai_1 U20073 ( .B1(n27219), .B2(n25157), .A1_N(n26369), 
        .A2_N(n25158), .Y(j202_soc_core_j22_cpu_rf_N3004) );
  sky130_fd_sc_hd__nand2_2 U20074 ( .A(n19764), .B(n19763), .Y(n25771) );
  sky130_fd_sc_hd__xnor2_2 U20075 ( .A(n19234), .B(n19233), .Y(n23241) );
  sky130_fd_sc_hd__fah_1 U20076 ( .A(n17548), .B(n17547), .CI(n17546), .COUT(
        n17577), .SUM(n17608) );
  sky130_fd_sc_hd__fah_1 U20077 ( .A(n18407), .B(n18406), .CI(n18405), .COUT(
        n18444), .SUM(n18414) );
  sky130_fd_sc_hd__fah_1 U20078 ( .A(n18071), .B(n18070), .CI(n18069), .COUT(
        n18120), .SUM(n18074) );
  sky130_fd_sc_hd__fah_1 U20079 ( .A(n17500), .B(n17499), .CI(n17498), .COUT(
        n17988), .SUM(n17482) );
  sky130_fd_sc_hd__fah_1 U20080 ( .A(n18410), .B(n18409), .CI(n18408), .COUT(
        n18443), .SUM(n18434) );
  sky130_fd_sc_hd__a21oi_1 U20081 ( .A1(n22661), .A2(n12178), .B1(n18904), .Y(
        n18905) );
  sky130_fd_sc_hd__xnor2_1 U20082 ( .A(j202_soc_core_j22_cpu_ml_bufa[16]), .B(
        j202_soc_core_j22_cpu_ml_bufa[15]), .Y(n17390) );
  sky130_fd_sc_hd__fah_1 U20083 ( .A(n17422), .B(n17421), .CI(n17420), .COUT(
        n17485), .SUM(n17479) );
  sky130_fd_sc_hd__fah_1 U20084 ( .A(n18679), .B(n18680), .CI(n18681), .COUT(
        n18736), .SUM(n18796) );
  sky130_fd_sc_hd__fah_1 U20085 ( .A(n17668), .B(n17667), .CI(n17666), .COUT(
        n17682), .SUM(n17684) );
  sky130_fd_sc_hd__nand3_1 U20086 ( .A(n23275), .B(n25336), .C(n23274), .Y(
        n23276) );
  sky130_fd_sc_hd__nand3_1 U20087 ( .A(n23275), .B(n25336), .C(n21518), .Y(
        n22613) );
  sky130_fd_sc_hd__nand2_4 U20088 ( .A(n25771), .B(n19766), .Y(n26831) );
  sky130_fd_sc_hd__a21oi_1 U20089 ( .A1(n23236), .A2(n26863), .B1(n24692), .Y(
        n25547) );
  sky130_fd_sc_hd__a22oi_2 U20090 ( .A1(j202_soc_core_memory0_ram_dout0[420]), 
        .A2(n21598), .B1(n21593), .B2(j202_soc_core_memory0_ram_dout0[324]), 
        .Y(n19328) );
  sky130_fd_sc_hd__a21oi_1 U20092 ( .A1(n23235), .A2(n26863), .B1(n25787), .Y(
        n25832) );
  sky130_fd_sc_hd__nand3_1 U20093 ( .A(n23244), .B(n26329), .C(n24478), .Y(
        n26514) );
  sky130_fd_sc_hd__a21boi_0 U20094 ( .A1(n24478), .A2(n23244), .B1_N(n26513), 
        .Y(n22635) );
  sky130_fd_sc_hd__clkinv_1 U20095 ( .A(n27222), .Y(n27223) );
  sky130_fd_sc_hd__a21o_2 U20096 ( .A1(n23450), .A2(n23449), .B1(n14849), .X(
        n26449) );
  sky130_fd_sc_hd__clkinv_1 U20097 ( .A(n26449), .Y(n26378) );
  sky130_fd_sc_hd__o21a_1 U20098 ( .A1(n24066), .A2(n26981), .B1(n25822), .X(
        n13281) );
  sky130_fd_sc_hd__o21a_1 U20099 ( .A1(n25182), .A2(n26981), .B1(n25822), .X(
        n13282) );
  sky130_fd_sc_hd__o21a_1 U20100 ( .A1(n24538), .A2(n26981), .B1(n25822), .X(
        n13283) );
  sky130_fd_sc_hd__o21a_1 U20101 ( .A1(n23262), .A2(n26981), .B1(n25822), .X(
        n13284) );
  sky130_fd_sc_hd__o21a_1 U20102 ( .A1(n25398), .A2(n26981), .B1(n25822), .X(
        n13285) );
  sky130_fd_sc_hd__o21a_1 U20103 ( .A1(n26101), .A2(n26981), .B1(n25822), .X(
        n13286) );
  sky130_fd_sc_hd__nor3_2 U20104 ( .A(n27660), .B(n27659), .C(n27658), .Y(
        n13289) );
  sky130_fd_sc_hd__and4_1 U20105 ( .A(n16339), .B(n16338), .C(n16337), .D(
        n16336), .X(n13290) );
  sky130_fd_sc_hd__and4_1 U20106 ( .A(n15974), .B(n15973), .C(n15972), .D(
        n15971), .X(n13291) );
  sky130_fd_sc_hd__and4_1 U20107 ( .A(n24124), .B(n17138), .C(n17155), .D(
        n27602), .X(n13292) );
  sky130_fd_sc_hd__a21o_2 U20108 ( .A1(n23522), .A2(n23521), .B1(n14849), .X(
        n27224) );
  sky130_fd_sc_hd__and4_1 U20109 ( .A(n14784), .B(n14783), .C(n14782), .D(
        n14781), .X(n13295) );
  sky130_fd_sc_hd__and4_1 U20110 ( .A(n14757), .B(n14756), .C(n14755), .D(
        n14754), .X(n13296) );
  sky130_fd_sc_hd__xor2_1 U20111 ( .A(j202_soc_core_qspi_wb_addr[11]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[11]), .X(n13297) );
  sky130_fd_sc_hd__xor2_1 U20112 ( .A(j202_soc_core_qspi_wb_addr[10]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[10]), .X(n13298) );
  sky130_fd_sc_hd__o21a_1 U20113 ( .A1(n23260), .A2(n26981), .B1(n25822), .X(
        n13299) );
  sky130_fd_sc_hd__nor2_1 U20114 ( .A(n23700), .B(n23705), .Y(n23794) );
  sky130_fd_sc_hd__xor2_1 U20115 ( .A(n26206), .B(n26205), .X(n13300) );
  sky130_fd_sc_hd__clkinv_1 U20116 ( .A(n18300), .Y(n22807) );
  sky130_fd_sc_hd__a21o_2 U20117 ( .A1(n23512), .A2(n23511), .B1(n14849), .X(
        n27227) );
  sky130_fd_sc_hd__nor2_2 U20118 ( .A(n15780), .B(n14849), .Y(n29356) );
  sky130_fd_sc_hd__clkinv_1 U20119 ( .A(n21095), .Y(n21650) );
  sky130_fd_sc_hd__clkinv_1 U20120 ( .A(n20908), .Y(n20794) );
  sky130_fd_sc_hd__inv_2 U20121 ( .A(j202_soc_core_j22_cpu_ml_bufa[12]), .Y(
        n17396) );
  sky130_fd_sc_hd__inv_2 U20122 ( .A(n13821), .Y(n14593) );
  sky130_fd_sc_hd__inv_2 U20123 ( .A(n14593), .Y(n16323) );
  sky130_fd_sc_hd__inv_2 U20124 ( .A(n14593), .Y(n16262) );
  sky130_fd_sc_hd__inv_2 U20125 ( .A(j202_soc_core_bootrom_00_address_w[11]), 
        .Y(n13393) );
  sky130_fd_sc_hd__inv_2 U20126 ( .A(n13393), .Y(n19354) );
  sky130_fd_sc_hd__and4_1 U20127 ( .A(n21274), .B(n21061), .C(n21270), .D(
        n21614), .X(n13304) );
  sky130_fd_sc_hd__and2_1 U20128 ( .A(n17067), .B(n14877), .X(n13306) );
  sky130_fd_sc_hd__and4_1 U20129 ( .A(n17007), .B(n15802), .C(n17049), .D(
        n16110), .X(n13307) );
  sky130_fd_sc_hd__and4_1 U20130 ( .A(n14678), .B(n14677), .C(n14676), .D(
        n14675), .X(n13308) );
  sky130_fd_sc_hd__and4_1 U20131 ( .A(n15127), .B(n15126), .C(n15125), .D(
        n15124), .X(n13309) );
  sky130_fd_sc_hd__o211ai_2 U20132 ( .A1(n23541), .A2(n23537), .B1(n23451), 
        .C1(n26449), .Y(n13310) );
  sky130_fd_sc_hd__inv_2 U20133 ( .A(n12169), .Y(n16443) );
  sky130_fd_sc_hd__inv_2 U20136 ( .A(n14770), .Y(n15982) );
  sky130_fd_sc_hd__inv_2 U20137 ( .A(n14770), .Y(n16493) );
  sky130_fd_sc_hd__inv_2 U20139 ( .A(n14496), .Y(n16470) );
  sky130_fd_sc_hd__inv_2 U20140 ( .A(n12163), .Y(n16324) );
  sky130_fd_sc_hd__inv_2 U20141 ( .A(n12163), .Y(n16431) );
  sky130_fd_sc_hd__inv_2 U20142 ( .A(n12174), .Y(n16279) );
  sky130_fd_sc_hd__clkinv_1 U20143 ( .A(j202_soc_core_j22_cpu_pc[3]), .Y(
        n20285) );
  sky130_fd_sc_hd__xor2_1 U20144 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]), .B(
        j202_soc_core_qspi_wb_addr[20]), .X(n13311) );
  sky130_fd_sc_hd__xor2_1 U20145 ( .A(j202_soc_core_qspi_wb_addr[13]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[13]), .X(n13312) );
  sky130_fd_sc_hd__xor2_1 U20146 ( .A(j202_soc_core_qspi_wb_addr[14]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]), .X(n13313) );
  sky130_fd_sc_hd__or2_1 U20147 ( .A(n17106), .B(n17105), .X(n13314) );
  sky130_fd_sc_hd__clkinv_1 U20148 ( .A(n24650), .Y(n25714) );
  sky130_fd_sc_hd__clkinv_1 U20149 ( .A(n27212), .Y(n26362) );
  sky130_fd_sc_hd__clkinv_1 U20150 ( .A(n27465), .Y(n25818) );
  sky130_fd_sc_hd__a21oi_1 U20151 ( .A1(n24637), .A2(n26802), .B1(n24636), .Y(
        n24638) );
  sky130_fd_sc_hd__o21a_1 U20152 ( .A1(n24660), .A2(n27892), .B1(n25813), .X(
        n13321) );
  sky130_fd_sc_hd__clkinv_1 U20154 ( .A(n22112), .Y(n22114) );
  sky130_fd_sc_hd__and4_1 U20155 ( .A(n14351), .B(n14350), .C(n14349), .D(
        n14348), .X(n13323) );
  sky130_fd_sc_hd__and4_1 U20156 ( .A(n13815), .B(n13814), .C(n13813), .D(
        n13812), .X(n13324) );
  sky130_fd_sc_hd__clkinv_1 U20157 ( .A(j202_soc_core_j22_cpu_pc[6]), .Y(
        n21555) );
  sky130_fd_sc_hd__clkinv_1 U20158 ( .A(j202_soc_core_j22_cpu_pc[5]), .Y(
        n21761) );
  sky130_fd_sc_hd__and4_1 U20159 ( .A(n15160), .B(n15159), .C(n15158), .D(
        n15157), .X(n13325) );
  sky130_fd_sc_hd__clkinv_1 U20160 ( .A(j202_soc_core_j22_cpu_pc[12]), .Y(
        n19496) );
  sky130_fd_sc_hd__clkinv_1 U20161 ( .A(j202_soc_core_j22_cpu_pc[11]), .Y(
        n21469) );
  sky130_fd_sc_hd__clkinv_1 U20162 ( .A(j202_soc_core_j22_cpu_pc[4]), .Y(
        n19453) );
  sky130_fd_sc_hd__clkinv_1 U20163 ( .A(j202_soc_core_j22_cpu_pc[8]), .Y(
        n21994) );
  sky130_fd_sc_hd__clkinv_1 U20164 ( .A(j202_soc_core_j22_cpu_pc[7]), .Y(
        n19078) );
  sky130_fd_sc_hd__and4_1 U20165 ( .A(n14628), .B(n14627), .C(n14626), .D(
        n14625), .X(n13326) );
  sky130_fd_sc_hd__and4_1 U20166 ( .A(n14638), .B(n14637), .C(n14636), .D(
        n14635), .X(n13327) );
  sky130_fd_sc_hd__clkinv_1 U20167 ( .A(j202_soc_core_j22_cpu_pc[9]), .Y(
        n22861) );
  sky130_fd_sc_hd__and2_1 U20168 ( .A(n24733), .B(n26450), .X(n13329) );
  sky130_fd_sc_hd__and4_1 U20169 ( .A(n14710), .B(n14709), .C(n14708), .D(
        n14707), .X(n13332) );
  sky130_fd_sc_hd__and4_1 U20170 ( .A(n14794), .B(n14793), .C(n14792), .D(
        n14791), .X(n13333) );
  sky130_fd_sc_hd__clkinv_1 U20171 ( .A(j202_soc_core_j22_cpu_pc[2]), .Y(
        n19203) );
  sky130_fd_sc_hd__and2_1 U20172 ( .A(n24497), .B(n26450), .X(n13336) );
  sky130_fd_sc_hd__clkinv_1 U20173 ( .A(j202_soc_core_j22_cpu_pc[13]), .Y(
        n21342) );
  sky130_fd_sc_hd__and4_1 U20174 ( .A(n15189), .B(n15188), .C(n15187), .D(
        n15186), .X(n13337) );
  sky130_fd_sc_hd__clkinv_1 U20175 ( .A(j202_soc_core_j22_cpu_pc[10]), .Y(
        n19213) );
  sky130_fd_sc_hd__clkinv_1 U20176 ( .A(j202_soc_core_j22_cpu_pc[14]), .Y(
        n21321) );
  sky130_fd_sc_hd__and4_1 U20177 ( .A(n14739), .B(n14738), .C(n14737), .D(
        n14736), .X(n13339) );
  sky130_fd_sc_hd__clkinv_1 U20178 ( .A(j202_soc_core_j22_cpu_pc[15]), .Y(
        n19063) );
  sky130_fd_sc_hd__and4_1 U20179 ( .A(n14822), .B(n14821), .C(n14820), .D(
        n14819), .X(n13340) );
  sky130_fd_sc_hd__and4_1 U20180 ( .A(n16361), .B(n16360), .C(n16359), .D(
        n16358), .X(n13341) );
  sky130_fd_sc_hd__and4_1 U20181 ( .A(n13710), .B(n13709), .C(n13708), .D(
        n13707), .X(n13345) );
  sky130_fd_sc_hd__nor2_1 U20182 ( .A(n20984), .B(n24575), .Y(n29056) );
  sky130_fd_sc_hd__clkinv_1 U20183 ( .A(n29056), .Y(n26211) );
  sky130_fd_sc_hd__nor2_2 U20184 ( .A(n24569), .B(n24807), .Y(n27983) );
  sky130_fd_sc_hd__inv_2 U20185 ( .A(n18619), .Y(n18140) );
  sky130_fd_sc_hd__nand2b_1 U20186 ( .A_N(n18353), .B(n22051), .Y(n18375) );
  sky130_fd_sc_hd__o21a_1 U20187 ( .A1(j202_soc_core_intc_core_00_rg_ipr[10]), 
        .A2(n25533), .B1(n19567), .X(n19569) );
  sky130_fd_sc_hd__clkbuf_1 U20188 ( .A(n17382), .X(n18617) );
  sky130_fd_sc_hd__inv_2 U20189 ( .A(n20669), .Y(n15705) );
  sky130_fd_sc_hd__clkinv_1 U20190 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[4]), .Y(n13384) );
  sky130_fd_sc_hd__a21oi_1 U20191 ( .A1(n22944), .A2(n19475), .B1(n19474), .Y(
        n19476) );
  sky130_fd_sc_hd__nor2_1 U20192 ( .A(n13386), .B(n13385), .Y(n21676) );
  sky130_fd_sc_hd__a2bb2oi_1 U20193 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[35]), .B2(n25485), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[38]), .A2_N(n24967), .Y(n19679) );
  sky130_fd_sc_hd__o22ai_1 U20194 ( .A1(n16492), .A2(n26567), .B1(n26565), 
        .B2(n13793), .Y(n14827) );
  sky130_fd_sc_hd__nor2_1 U20196 ( .A(n26398), .B(n25824), .Y(n22923) );
  sky130_fd_sc_hd__clkinv_1 U20197 ( .A(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n21677) );
  sky130_fd_sc_hd__nor2_1 U20198 ( .A(n24778), .B(n24783), .Y(n26085) );
  sky130_fd_sc_hd__nand2_1 U20199 ( .A(n11614), .B(n18892), .Y(n18893) );
  sky130_fd_sc_hd__clkinv_1 U20200 ( .A(n23922), .Y(n26409) );
  sky130_fd_sc_hd__inv_2 U20201 ( .A(n13676), .Y(n14496) );
  sky130_fd_sc_hd__nor2_1 U20202 ( .A(n23012), .B(n24778), .Y(n26443) );
  sky130_fd_sc_hd__nand2_1 U20203 ( .A(n17289), .B(n20623), .Y(n21722) );
  sky130_fd_sc_hd__nand2_1 U20204 ( .A(n25325), .B(n25323), .Y(n21502) );
  sky130_fd_sc_hd__clkinv_1 U20205 ( .A(j202_soc_core_memory0_ram_dout0_sel[7]), .Y(n13377) );
  sky130_fd_sc_hd__nand2_1 U20206 ( .A(n13503), .B(n13505), .Y(n13501) );
  sky130_fd_sc_hd__nor2_1 U20207 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .B(n13429), .Y(n21697) );
  sky130_fd_sc_hd__nor2_1 U20208 ( .A(n19054), .B(n19053), .Y(n22865) );
  sky130_fd_sc_hd__nand3_1 U20209 ( .A(n13655), .B(n13654), .C(n13653), .Y(
        n14846) );
  sky130_fd_sc_hd__nor2_1 U20210 ( .A(n24752), .B(n25094), .Y(n27863) );
  sky130_fd_sc_hd__nand2_1 U20211 ( .A(n11128), .B(n24499), .Y(n24051) );
  sky130_fd_sc_hd__nand2b_1 U20212 ( .A_N(n23260), .B(n11713), .Y(n22853) );
  sky130_fd_sc_hd__nor2_1 U20213 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__0_), 
        .B(j202_soc_core_j22_cpu_regop_M_Wm__3_), .Y(n24429) );
  sky130_fd_sc_hd__nand2_1 U20214 ( .A(n16048), .B(n20428), .Y(n20547) );
  sky130_fd_sc_hd__clkinv_1 U20216 ( .A(n28738), .Y(n28732) );
  sky130_fd_sc_hd__nor2_1 U20217 ( .A(n24750), .B(n25094), .Y(n27864) );
  sky130_fd_sc_hd__nand3_1 U20218 ( .A(n24760), .B(
        j202_soc_core_intc_core_00_bs_addr[8]), .C(n28886), .Y(n27306) );
  sky130_fd_sc_hd__nor2_1 U20219 ( .A(j202_soc_core_wbqspiflash_00_state[1]), 
        .B(n26042), .Y(n25954) );
  sky130_fd_sc_hd__nand2_1 U20220 ( .A(n24053), .B(n27450), .Y(n27438) );
  sky130_fd_sc_hd__nand2_1 U20221 ( .A(n27271), .B(n18871), .Y(n26863) );
  sky130_fd_sc_hd__nor2_1 U20222 ( .A(n13571), .B(n12763), .Y(n18879) );
  sky130_fd_sc_hd__clkinv_1 U20223 ( .A(n27226), .Y(n23082) );
  sky130_fd_sc_hd__nor2_1 U20224 ( .A(n24953), .B(n24952), .Y(n27835) );
  sky130_fd_sc_hd__nor2_1 U20225 ( .A(n28590), .B(n24975), .Y(n27861) );
  sky130_fd_sc_hd__nand2b_1 U20226 ( .A_N(n29056), .B(n26225), .Y(n28737) );
  sky130_fd_sc_hd__nor2_1 U20227 ( .A(n27924), .B(n23611), .Y(n27785) );
  sky130_fd_sc_hd__nor2_1 U20228 ( .A(n27721), .B(n16054), .Y(n27914) );
  sky130_fd_sc_hd__inv_1 U20229 ( .A(n16831), .Y(n17126) );
  sky130_fd_sc_hd__nand3_1 U20230 ( .A(start_n_reg[1]), .B(wbs_cyc_i), .C(
        wbs_stb_i), .Y(n13346) );
  sky130_fd_sc_hd__clkinv_1 U20231 ( .A(j202_soc_core_intc_core_00_rg_ie[14]), 
        .Y(n25498) );
  sky130_fd_sc_hd__nor2b_1 U20232 ( .B_N(n28776), .A(n24228), .Y(n28775) );
  sky130_fd_sc_hd__nand2_1 U20233 ( .A(n26042), .B(
        j202_soc_core_wbqspiflash_00_state[1]), .Y(n28243) );
  sky130_fd_sc_hd__nand2_1 U20234 ( .A(j202_soc_core_qspi_wb_wdat[25]), .B(
        n29594), .Y(n25203) );
  sky130_fd_sc_hd__clkinv_1 U20235 ( .A(n28519), .Y(n28539) );
  sky130_fd_sc_hd__clkinv_1 U20236 ( .A(n27751), .Y(n27988) );
  sky130_fd_sc_hd__nand2_1 U20237 ( .A(j202_soc_core_qspi_wb_wdat[27]), .B(
        n29594), .Y(n25649) );
  sky130_fd_sc_hd__nand2_1 U20238 ( .A(j202_soc_core_qspi_wb_wdat[21]), .B(
        n29594), .Y(n25427) );
  sky130_fd_sc_hd__a211oi_1 U20239 ( .A1(n25982), .A2(n27040), .B1(n25026), 
        .C1(n27719), .Y(n27874) );
  sky130_fd_sc_hd__clkinv_1 U20240 ( .A(n24575), .Y(n23907) );
  sky130_fd_sc_hd__nand2_1 U20241 ( .A(n23328), .B(n23327), .Y(n26861) );
  sky130_fd_sc_hd__clkinv_1 U20242 ( .A(n28967), .Y(n28281) );
  sky130_fd_sc_hd__nand2_1 U20243 ( .A(n24946), .B(n24955), .Y(n27833) );
  sky130_fd_sc_hd__clkinv_1 U20244 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[12]), .Y(n26307) );
  sky130_fd_sc_hd__nand2_1 U20245 ( .A(n25534), .B(n29594), .Y(n25532) );
  sky130_fd_sc_hd__nand2_1 U20246 ( .A(n25112), .B(j202_soc_core_aquc_SEL__2_), 
        .Y(n27593) );
  sky130_fd_sc_hd__clkinv_1 U20247 ( .A(n25350), .Y(n27193) );
  sky130_fd_sc_hd__inv_2 U20248 ( .A(n19040), .Y(n22234) );
  sky130_fd_sc_hd__nor3_1 U20249 ( .A(wb_rst_i), .B(wbs_ack_o), .C(n13346), 
        .Y(n23690) );
  sky130_fd_sc_hd__or3_1 U20250 ( .A(n26199), .B(n26200), .C(n28727), .X(
        n29244) );
  sky130_fd_sc_hd__nand3_1 U20251 ( .A(n21376), .B(n21375), .C(n21374), .Y(
        n29062) );
  sky130_fd_sc_hd__o31ai_1 U20252 ( .A1(n27659), .A2(n23454), .A3(n27658), 
        .B1(n29594), .Y(n10674) );
  sky130_fd_sc_hd__nand2b_1 U20253 ( .A_N(n29056), .B(n29593), .Y(n29237) );
  sky130_fd_sc_hd__and3_1 U20254 ( .A(n25024), .B(n23321), .C(n29594), .X(
        n29120) );
  sky130_fd_sc_hd__o2bb2ai_1 U20255 ( .B1(n27217), .B2(n27524), .A1_N(n25819), 
        .A2_N(n25810), .Y(j202_soc_core_j22_cpu_rf_N2835) );
  sky130_fd_sc_hd__o2bb2ai_1 U20256 ( .B1(n27223), .B2(n25157), .A1_N(n27223), 
        .A2_N(n25158), .Y(j202_soc_core_j22_cpu_rf_N3041) );
  sky130_fd_sc_hd__or3_1 U20257 ( .A(n28590), .B(n23943), .C(n26383), .X(
        n29112) );
  sky130_fd_sc_hd__nand2_1 U20258 ( .A(n28647), .B(n12142), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N311) );
  sky130_fd_sc_hd__clkbuf_1 U20259 ( .A(io_oeb[12]), .X(io_oeb[13]) );
  sky130_fd_sc_hd__clkbuf_1 U20260 ( .A(la_data_out[2]), .X(io_out[2]) );
  sky130_fd_sc_hd__clkbuf_1 U20261 ( .A(la_data_out[11]), .X(io_out[31]) );
  sky130_fd_sc_hd__nor2_1 U20262 ( .A(n28590), .B(n28298), .Y(n29083) );
  sky130_fd_sc_hd__nor2_1 U20263 ( .A(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[1]), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[0]), .Y(n13349) );
  sky130_fd_sc_hd__xnor2_1 U20264 ( .A(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[1]), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[1]), .Y(n13348) );
  sky130_fd_sc_hd__xnor2_1 U20265 ( .A(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[0]), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[0]), .Y(n13347) );
  sky130_fd_sc_hd__nand2_1 U20266 ( .A(n13348), .B(n13347), .Y(n13350) );
  sky130_fd_sc_hd__or4_1 U20267 ( .A(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[2]), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[2]), .C(n13349), 
        .D(n13350), .X(n24802) );
  sky130_fd_sc_hd__nand3_1 U20268 ( .A(n13351), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[2]), .C(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[2]), .Y(n24803) );
  sky130_fd_sc_hd__nand2_1 U20269 ( .A(n24802), .B(n24803), .Y(n29076) );
  sky130_fd_sc_hd__xnor2_1 U20270 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .B(
        j202_soc_core_bldc_core_00_pwm_period[10]), .Y(n13363) );
  sky130_fd_sc_hd__xnor2_1 U20271 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .B(
        j202_soc_core_bldc_core_00_pwm_period[0]), .Y(n13362) );
  sky130_fd_sc_hd__xor2_1 U20272 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[11]), .B(
        j202_soc_core_bldc_core_00_pwm_period[11]), .X(n13353) );
  sky130_fd_sc_hd__xor2_1 U20273 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]), .B(
        j202_soc_core_bldc_core_00_pwm_period[7]), .X(n13352) );
  sky130_fd_sc_hd__nor2_1 U20274 ( .A(n13353), .B(n13352), .Y(n13360) );
  sky130_fd_sc_hd__xnor2_1 U20275 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[3]), .B(n27846), .Y(
        n13355) );
  sky130_fd_sc_hd__xnor2_1 U20276 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[2]), .B(n24966), .Y(
        n13354) );
  sky130_fd_sc_hd__nor2_1 U20277 ( .A(n13355), .B(n13354), .Y(n13359) );
  sky130_fd_sc_hd__xnor2_1 U20278 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .B(n27150), .Y(
        n13357) );
  sky130_fd_sc_hd__xnor2_1 U20279 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]), .B(n25624), .Y(
        n13356) );
  sky130_fd_sc_hd__nor2_1 U20280 ( .A(n13357), .B(n13356), .Y(n13358) );
  sky130_fd_sc_hd__and3_1 U20281 ( .A(n13360), .B(n13359), .C(n13358), .X(
        n13361) );
  sky130_fd_sc_hd__and3_1 U20282 ( .A(n13363), .B(n13362), .C(n13361), .X(
        n13370) );
  sky130_fd_sc_hd__xnor2_1 U20283 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[4]), .B(
        j202_soc_core_bldc_core_00_pwm_period[4]), .Y(n13365) );
  sky130_fd_sc_hd__xnor2_1 U20284 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .B(
        j202_soc_core_bldc_core_00_pwm_period[1]), .Y(n13364) );
  sky130_fd_sc_hd__xnor2_1 U20285 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .B(
        j202_soc_core_bldc_core_00_pwm_period[6]), .Y(n13367) );
  sky130_fd_sc_hd__xnor2_1 U20286 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]), .B(
        j202_soc_core_bldc_core_00_pwm_period[5]), .Y(n13366) );
  sky130_fd_sc_hd__nand3_1 U20287 ( .A(n13370), .B(n13369), .C(n13368), .Y(
        n28581) );
  sky130_fd_sc_hd__nand2_1 U20288 ( .A(n28581), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .Y(n29008) );
  sky130_fd_sc_hd__nor2_1 U20289 ( .A(j202_soc_core_qspi_wb_ack), .B(n26131), 
        .Y(n25881) );
  sky130_fd_sc_hd__nor2_1 U20291 ( .A(j202_soc_core_memory0_ram_dout0_sel[14]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[13]), .Y(n13503) );
  sky130_fd_sc_hd__nor2_1 U20292 ( .A(j202_soc_core_memory0_ram_dout0_sel[7]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[6]), .Y(n13490) );
  sky130_fd_sc_hd__nand2_1 U20293 ( .A(n13490), .B(n13372), .Y(n13494) );
  sky130_fd_sc_hd__nor2_1 U20294 ( .A(j202_soc_core_memory0_ram_dout0_sel[4]), 
        .B(n13494), .Y(n13492) );
  sky130_fd_sc_hd__nand3_1 U20295 ( .A(n13492), .B(
        j202_soc_core_memory0_ram_dout0_sel[2]), .C(n13373), .Y(n13374) );
  sky130_fd_sc_hd__nor2_1 U20296 ( .A(j202_soc_core_memory0_ram_dout0_sel[3]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[2]), .Y(n13379) );
  sky130_fd_sc_hd__nand4_1 U20297 ( .A(n13492), .B(n13379), .C(
        j202_soc_core_memory0_ram_dout0_sel[0]), .D(n13375), .Y(n13376) );
  sky130_fd_sc_hd__nand2_1 U20298 ( .A(n13377), .B(
        j202_soc_core_memory0_ram_dout0_sel[6]), .Y(n13378) );
  sky130_fd_sc_hd__nand3_1 U20299 ( .A(n13492), .B(
        j202_soc_core_memory0_ram_dout0_sel[1]), .C(n13379), .Y(n13380) );
  sky130_fd_sc_hd__nand3_1 U20300 ( .A(n13381), .B(n11919), .C(
        j202_soc_core_j22_cpu_ma_M_area[1]), .Y(n13385) );
  sky130_fd_sc_hd__nor2_1 U20301 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[5]), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[3]), .Y(n13382) );
  sky130_fd_sc_hd__nand3_1 U20302 ( .A(n13451), .B(n13382), .C(n13384), .Y(
        n17184) );
  sky130_fd_sc_hd__nand2_1 U20303 ( .A(n17182), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[1]), .Y(n13383) );
  sky130_fd_sc_hd__a22oi_1 U20304 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[52]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[84]), .Y(n13508) );
  sky130_fd_sc_hd__and3_1 U20305 ( .A(n13384), .B(n13386), .C(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[3]), .X(n13450) );
  sky130_fd_sc_hd__nand3_1 U20306 ( .A(n13451), .B(n13450), .C(
        j202_soc_core_aquc_CE__1_), .Y(n20860) );
  sky130_fd_sc_hd__nand2_1 U20307 ( .A(n21675), .B(j202_soc_core_uart_div1[4]), 
        .Y(n13507) );
  sky130_fd_sc_hd__nand2_1 U20308 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[20]), .Y(n13506) );
  sky130_fd_sc_hd__nand4_1 U20309 ( .A(n13508), .B(n21677), .C(n13507), .D(
        n13506), .Y(n13461) );
  sky130_fd_sc_hd__nand2_1 U20310 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .B(n17277), .Y(n16170) );
  sky130_fd_sc_hd__nor2_1 U20311 ( .A(n19354), .B(n16170), .Y(n19085) );
  sky130_fd_sc_hd__inv_2 U20312 ( .A(j202_soc_core_bootrom_00_address_w[10]), 
        .Y(n17274) );
  sky130_fd_sc_hd__nand2_1 U20313 ( .A(n19085), .B(n16706), .Y(n16682) );
  sky130_fd_sc_hd__nor2_1 U20314 ( .A(n17175), .B(n16682), .Y(n15319) );
  sky130_fd_sc_hd__buf_2 U20315 ( .A(j202_soc_core_bootrom_00_address_w[10]), 
        .X(n19381) );
  sky130_fd_sc_hd__nand2_1 U20316 ( .A(n19381), .B(n17289), .Y(n14884) );
  sky130_fd_sc_hd__inv_2 U20317 ( .A(j202_soc_core_bootrom_00_address_w[11]), 
        .Y(n20787) );
  sky130_fd_sc_hd__nand2_1 U20318 ( .A(n16171), .B(n20787), .Y(n17165) );
  sky130_fd_sc_hd__nor2_1 U20319 ( .A(n14884), .B(n17165), .Y(n16840) );
  sky130_fd_sc_hd__nand2_1 U20320 ( .A(n16840), .B(n12137), .Y(n15350) );
  sky130_fd_sc_hd__nand2_1 U20321 ( .A(n15550), .B(n15350), .Y(n15383) );
  sky130_fd_sc_hd__nor2_1 U20322 ( .A(n17277), .B(n15423), .Y(n14863) );
  sky130_fd_sc_hd__nand2_1 U20323 ( .A(n14863), .B(n19354), .Y(n13391) );
  sky130_fd_sc_hd__nand2b_1 U20324 ( .A_N(n13391), .B(n13387), .Y(n15578) );
  sky130_fd_sc_hd__nand2_1 U20325 ( .A(n17273), .B(n19354), .Y(n17059) );
  sky130_fd_sc_hd__nor2_1 U20326 ( .A(n17314), .B(n15423), .Y(n13417) );
  sky130_fd_sc_hd__nand2b_1 U20327 ( .A_N(n17059), .B(n13417), .Y(n15538) );
  sky130_fd_sc_hd__nand2_1 U20328 ( .A(n15578), .B(n15538), .Y(n15596) );
  sky130_fd_sc_hd__nor2_1 U20329 ( .A(n17289), .B(n19381), .Y(n15838) );
  sky130_fd_sc_hd__nand2_1 U20330 ( .A(n15838), .B(n17314), .Y(n13394) );
  sky130_fd_sc_hd__nor2_1 U20331 ( .A(n13394), .B(n17059), .Y(n15321) );
  sky130_fd_sc_hd__nor2_1 U20332 ( .A(j202_soc_core_bootrom_00_address_w[11]), 
        .B(n14884), .Y(n16176) );
  sky130_fd_sc_hd__nand2_1 U20333 ( .A(n16176), .B(n13388), .Y(n15589) );
  sky130_fd_sc_hd__nand3_1 U20334 ( .A(n15364), .B(n15592), .C(n15589), .Y(
        n13392) );
  sky130_fd_sc_hd__nor2_1 U20335 ( .A(n17278), .B(n13389), .Y(n15365) );
  sky130_fd_sc_hd__nand2b_1 U20336 ( .A_N(n17059), .B(n14863), .Y(n15537) );
  sky130_fd_sc_hd__nor2_1 U20337 ( .A(n15365), .B(n13390), .Y(n13476) );
  sky130_fd_sc_hd__nand2b_1 U20338 ( .A_N(n13391), .B(n13388), .Y(n15595) );
  sky130_fd_sc_hd__nand2_1 U20339 ( .A(n13476), .B(n15595), .Y(n15608) );
  sky130_fd_sc_hd__nor3_1 U20340 ( .A(n15383), .B(n13392), .C(n15608), .Y(
        n13406) );
  sky130_fd_sc_hd__nor2_1 U20341 ( .A(n20788), .B(n20687), .Y(n16090) );
  sky130_fd_sc_hd__nand2b_1 U20342 ( .A_N(n16162), .B(n17273), .Y(n15610) );
  sky130_fd_sc_hd__nand2b_1 U20343 ( .A_N(n15610), .B(n17314), .Y(n15615) );
  sky130_fd_sc_hd__nand2_1 U20344 ( .A(n16706), .B(n17314), .Y(n13436) );
  sky130_fd_sc_hd__nand2b_1 U20345 ( .A_N(n17282), .B(n13431), .Y(n15593) );
  sky130_fd_sc_hd__nand2_1 U20346 ( .A(n16180), .B(n16171), .Y(n20633) );
  sky130_fd_sc_hd__nand2b_1 U20347 ( .A_N(n20633), .B(n17175), .Y(n15613) );
  sky130_fd_sc_hd__nand2_1 U20348 ( .A(n16616), .B(n20787), .Y(n19121) );
  sky130_fd_sc_hd__nand2b_1 U20349 ( .A_N(n19121), .B(n15425), .Y(n16722) );
  sky130_fd_sc_hd__nand2b_1 U20350 ( .A_N(n16722), .B(n12137), .Y(n15535) );
  sky130_fd_sc_hd__nand3_1 U20351 ( .A(n15344), .B(n15613), .C(n15535), .Y(
        n13412) );
  sky130_fd_sc_hd__inv_2 U20352 ( .A(n13398), .Y(n20623) );
  sky130_fd_sc_hd__inv_2 U20353 ( .A(j202_soc_core_bootrom_00_address_w[3]), 
        .Y(n20579) );
  sky130_fd_sc_hd__nor2_1 U20354 ( .A(n20623), .B(n20579), .Y(n15584) );
  sky130_fd_sc_hd__nand2b_1 U20355 ( .A_N(n17278), .B(n13395), .Y(n15359) );
  sky130_fd_sc_hd__nor2_1 U20356 ( .A(n14884), .B(n17282), .Y(n13471) );
  sky130_fd_sc_hd__nand2_1 U20357 ( .A(n13471), .B(n17277), .Y(n15341) );
  sky130_fd_sc_hd__nand2_1 U20358 ( .A(n15613), .B(n15341), .Y(n15243) );
  sky130_fd_sc_hd__nand2_1 U20359 ( .A(n16180), .B(n13388), .Y(n15594) );
  sky130_fd_sc_hd__nand2b_1 U20360 ( .A_N(n15594), .B(n17277), .Y(n15380) );
  sky130_fd_sc_hd__nand2b_1 U20361 ( .A_N(n17278), .B(n13294), .Y(n15614) );
  sky130_fd_sc_hd__nor2_1 U20362 ( .A(n19354), .B(n17314), .Y(n19380) );
  sky130_fd_sc_hd__nand3_1 U20363 ( .A(n19380), .B(n17273), .C(n15425), .Y(
        n15558) );
  sky130_fd_sc_hd__nand2_1 U20364 ( .A(n13419), .B(n15595), .Y(n15330) );
  sky130_fd_sc_hd__nor2_1 U20365 ( .A(n15423), .B(n17278), .Y(n15548) );
  sky130_fd_sc_hd__nor2_1 U20366 ( .A(n15330), .B(n15548), .Y(n13397) );
  sky130_fd_sc_hd__nand4_1 U20367 ( .A(n15380), .B(n13397), .C(n15537), .D(
        n15589), .Y(n13422) );
  sky130_fd_sc_hd__nand2_1 U20368 ( .A(n20788), .B(n20623), .Y(n15557) );
  sky130_fd_sc_hd__o31a_1 U20369 ( .A1(n15266), .A2(n15243), .A3(n13422), .B1(
        n15630), .X(n13399) );
  sky130_fd_sc_hd__a21oi_1 U20370 ( .A1(n13412), .A2(n15584), .B1(n13399), .Y(
        n13405) );
  sky130_fd_sc_hd__nand2_1 U20371 ( .A(n15595), .B(n15359), .Y(n15220) );
  sky130_fd_sc_hd__nand2b_1 U20372 ( .A_N(n17278), .B(n13417), .Y(n15564) );
  sky130_fd_sc_hd__nand2_1 U20373 ( .A(n15610), .B(n15564), .Y(n13400) );
  sky130_fd_sc_hd__nor2_1 U20374 ( .A(n15220), .B(n13400), .Y(n13402) );
  sky130_fd_sc_hd__nand2_1 U20375 ( .A(n13387), .B(n19354), .Y(n13430) );
  sky130_fd_sc_hd__nor2_1 U20376 ( .A(n13430), .B(n13401), .Y(n15366) );
  sky130_fd_sc_hd__nor2_1 U20377 ( .A(n15366), .B(n15596), .Y(n15251) );
  sky130_fd_sc_hd__nand2_1 U20378 ( .A(n16180), .B(n13387), .Y(n15256) );
  sky130_fd_sc_hd__nand3_1 U20379 ( .A(n13402), .B(n15251), .C(n15256), .Y(
        n13403) );
  sky130_fd_sc_hd__nand2_1 U20380 ( .A(n20579), .B(n20687), .Y(n15708) );
  sky130_fd_sc_hd__nand2_1 U20381 ( .A(n13403), .B(n17163), .Y(n13404) );
  sky130_fd_sc_hd__o211ai_1 U20382 ( .A1(n13406), .A2(n15384), .B1(n13405), 
        .C1(n13404), .Y(n13411) );
  sky130_fd_sc_hd__nor3_1 U20383 ( .A(j202_soc_core_bootrom_00_address_w[17]), 
        .B(j202_soc_core_bootrom_00_address_w[16]), .C(
        j202_soc_core_j22_cpu_ma_M_area[0]), .Y(n13410) );
  sky130_fd_sc_hd__nor2_1 U20384 ( .A(j202_soc_core_bootrom_00_address_w[14]), 
        .B(j202_soc_core_bootrom_00_address_w[13]), .Y(n13408) );
  sky130_fd_sc_hd__nor2_1 U20385 ( .A(j202_soc_core_bootrom_00_address_w[15]), 
        .B(j202_soc_core_bootrom_00_address_w[12]), .Y(n13407) );
  sky130_fd_sc_hd__nand4_1 U20386 ( .A(n13410), .B(n13409), .C(n13408), .D(
        n13407), .Y(n14965) );
  sky130_fd_sc_hd__nand2_1 U20387 ( .A(n17098), .B(
        j202_soc_core_bootrom_00_address_w[8]), .Y(n15493) );
  sky130_fd_sc_hd__nor2_2 U20388 ( .A(n15454), .B(n15493), .Y(n20908) );
  sky130_fd_sc_hd__nand2_1 U20389 ( .A(n13411), .B(n20908), .Y(n13511) );
  sky130_fd_sc_hd__nor2_1 U20390 ( .A(n19121), .B(n15432), .Y(n16182) );
  sky130_fd_sc_hd__nand2_1 U20391 ( .A(n16182), .B(n12137), .Y(n15533) );
  sky130_fd_sc_hd__nand2_1 U20392 ( .A(n16176), .B(n17302), .Y(n15242) );
  sky130_fd_sc_hd__nand2_1 U20393 ( .A(n15533), .B(n15242), .Y(n15310) );
  sky130_fd_sc_hd__nand3_1 U20394 ( .A(n16176), .B(n17273), .C(n17314), .Y(
        n15586) );
  sky130_fd_sc_hd__nand4_1 U20395 ( .A(n13414), .B(n13413), .C(n15586), .D(
        n15545), .Y(n13428) );
  sky130_fd_sc_hd__nand3b_1 U20396 ( .A_N(n16162), .B(n17302), .C(n17314), .Y(
        n15340) );
  sky130_fd_sc_hd__nor2_1 U20397 ( .A(n13438), .B(n15366), .Y(n13465) );
  sky130_fd_sc_hd__nand2b_1 U20398 ( .A_N(n15321), .B(n15614), .Y(n13415) );
  sky130_fd_sc_hd__nor2_1 U20399 ( .A(n17037), .B(n16162), .Y(n15347) );
  sky130_fd_sc_hd__nand2_1 U20400 ( .A(n15347), .B(n17277), .Y(n15560) );
  sky130_fd_sc_hd__nand2b_1 U20401 ( .A_N(n15256), .B(n17277), .Y(n15534) );
  sky130_fd_sc_hd__nand2_1 U20402 ( .A(n15341), .B(n15537), .Y(n13437) );
  sky130_fd_sc_hd__nand3_1 U20403 ( .A(n13464), .B(n13416), .C(n15538), .Y(
        n15569) );
  sky130_fd_sc_hd__and4b_1 U20404 ( .B(n13465), .C(n15381), .D(n15578), .A_N(
        n15569), .X(n13426) );
  sky130_fd_sc_hd__nor2_1 U20405 ( .A(n17314), .B(n15610), .Y(n15369) );
  sky130_fd_sc_hd__nand3_1 U20406 ( .A(n13417), .B(n13388), .C(n19354), .Y(
        n15612) );
  sky130_fd_sc_hd__nor2_1 U20407 ( .A(n15366), .B(n15321), .Y(n15331) );
  sky130_fd_sc_hd__nand2_1 U20408 ( .A(n15612), .B(n15331), .Y(n15226) );
  sky130_fd_sc_hd__a21oi_1 U20409 ( .A1(n16163), .A2(n13387), .B1(n15226), .Y(
        n13418) );
  sky130_fd_sc_hd__nand4_1 U20410 ( .A(n13479), .B(n13419), .C(n13418), .D(
        n15340), .Y(n13420) );
  sky130_fd_sc_hd__nand2_1 U20411 ( .A(n13420), .B(n15630), .Y(n13425) );
  sky130_fd_sc_hd__nand2b_1 U20412 ( .A_N(n15596), .B(n15359), .Y(n15254) );
  sky130_fd_sc_hd__nor2_1 U20413 ( .A(n17277), .B(n15594), .Y(n15258) );
  sky130_fd_sc_hd__nand2_1 U20414 ( .A(n15586), .B(n15530), .Y(n15323) );
  sky130_fd_sc_hd__nor4_1 U20415 ( .A(n13478), .B(n15254), .C(n15323), .D(
        n15383), .Y(n13421) );
  sky130_fd_sc_hd__nand3_1 U20416 ( .A(n15533), .B(n13421), .C(n15612), .Y(
        n13423) );
  sky130_fd_sc_hd__o211ai_1 U20418 ( .A1(n13426), .A2(n15708), .B1(n13425), 
        .C1(n13424), .Y(n13427) );
  sky130_fd_sc_hd__a21oi_1 U20419 ( .A1(n13428), .A2(n16090), .B1(n13427), .Y(
        n13449) );
  sky130_fd_sc_hd__nand2_1 U20420 ( .A(n13432), .B(n13431), .Y(n13433) );
  sky130_fd_sc_hd__nand3_1 U20421 ( .A(n15615), .B(n15589), .C(n13433), .Y(
        n15568) );
  sky130_fd_sc_hd__nor3_1 U20422 ( .A(n16840), .B(n15365), .C(n13438), .Y(
        n13434) );
  sky130_fd_sc_hd__nand4_1 U20423 ( .A(n15314), .B(n15551), .C(n13434), .D(
        n15534), .Y(n13447) );
  sky130_fd_sc_hd__nand2_1 U20424 ( .A(n15380), .B(n16722), .Y(n15351) );
  sky130_fd_sc_hd__nand2_1 U20425 ( .A(n15545), .B(n15340), .Y(n15580) );
  sky130_fd_sc_hd__nand2_1 U20426 ( .A(n15534), .B(n12192), .Y(n13435) );
  sky130_fd_sc_hd__nor2_1 U20427 ( .A(n13435), .B(n15254), .Y(n15324) );
  sky130_fd_sc_hd__nor4_1 U20429 ( .A(n15319), .B(n15351), .C(n15561), .D(
        n13437), .Y(n13442) );
  sky130_fd_sc_hd__nor2_1 U20430 ( .A(n15321), .B(n13438), .Y(n13440) );
  sky130_fd_sc_hd__nor2b_1 U20431 ( .B_N(n15564), .A(n15347), .Y(n13439) );
  sky130_fd_sc_hd__nand3_1 U20432 ( .A(n15344), .B(n13440), .C(n13439), .Y(
        n15316) );
  sky130_fd_sc_hd__nor3_1 U20433 ( .A(n16840), .B(n15316), .C(n15596), .Y(
        n13441) );
  sky130_fd_sc_hd__o22ai_1 U20434 ( .A1(n13442), .A2(n15708), .B1(n13441), 
        .B2(n15384), .Y(n13446) );
  sky130_fd_sc_hd__nand2_1 U20435 ( .A(n15593), .B(n15558), .Y(n13443) );
  sky130_fd_sc_hd__nand2_1 U20436 ( .A(n19085), .B(n15425), .Y(n20463) );
  sky130_fd_sc_hd__nand2b_1 U20437 ( .A_N(n20463), .B(n12137), .Y(n13466) );
  sky130_fd_sc_hd__nand2_1 U20438 ( .A(n13466), .B(n15537), .Y(n15581) );
  sky130_fd_sc_hd__nor2_1 U20439 ( .A(n13443), .B(n15581), .Y(n15373) );
  sky130_fd_sc_hd__nor2_1 U20440 ( .A(n15623), .B(n15319), .Y(n13444) );
  sky130_fd_sc_hd__a31oi_1 U20441 ( .A1(n15373), .A2(n13444), .A3(n15610), 
        .B1(n15557), .Y(n13445) );
  sky130_fd_sc_hd__a211oi_1 U20442 ( .A1(n13447), .A2(n15584), .B1(n13446), 
        .C1(n13445), .Y(n13448) );
  sky130_fd_sc_hd__o22a_1 U20443 ( .A1(n13449), .A2(n19856), .B1(n21124), .B2(
        n13448), .X(n13510) );
  sky130_fd_sc_hd__nor2_1 U20444 ( .A(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[0]), .B(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[1]), .Y(n23910) );
  sky130_fd_sc_hd__nand3_1 U20445 ( .A(n23910), .B(n23909), .C(n22296), .Y(
        n20149) );
  sky130_fd_sc_hd__nand2_1 U20446 ( .A(n13451), .B(n13450), .Y(n17203) );
  sky130_fd_sc_hd__nor3_1 U20447 ( .A(j202_soc_core_aquc_ADR__2_), .B(n20149), 
        .C(n17203), .Y(n13452) );
  sky130_fd_sc_hd__nand2_1 U20448 ( .A(n25677), .B(n13452), .Y(n13460) );
  sky130_fd_sc_hd__nor2_1 U20449 ( .A(j202_soc_core_aquc_ADR__6_), .B(
        j202_soc_core_aquc_ADR__5_), .Y(n13455) );
  sky130_fd_sc_hd__nor2_1 U20450 ( .A(j202_soc_core_aquc_ADR__7_), .B(n10960), 
        .Y(n13454) );
  sky130_fd_sc_hd__nand3_1 U20451 ( .A(n13455), .B(n13454), .C(n13453), .Y(
        n13459) );
  sky130_fd_sc_hd__nor2_1 U20452 ( .A(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[6]), .B(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[5]), .Y(n13457) );
  sky130_fd_sc_hd__nor2_1 U20453 ( .A(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[7]), .B(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[1]), .Y(n13456) );
  sky130_fd_sc_hd__nand3b_1 U20454 ( .A_N(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[0]), .B(n13457), 
        .C(n13456), .Y(n13458) );
  sky130_fd_sc_hd__mux2i_1 U20455 ( .A0(n13459), .A1(n13458), .S(n20149), .Y(
        n20147) );
  sky130_fd_sc_hd__mux2i_1 U20456 ( .A0(j202_soc_core_aquc_ADR__4_), .A1(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[4]), .S(n20149), 
        .Y(n20148) );
  sky130_fd_sc_hd__nand2_1 U20457 ( .A(n20147), .B(n20148), .Y(n19858) );
  sky130_fd_sc_hd__nor2_1 U20458 ( .A(n13460), .B(n19858), .Y(n15249) );
  sky130_fd_sc_hd__nand2_1 U20459 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_duty[8]), .Y(n13509) );
  sky130_fd_sc_hd__nand4b_1 U20460 ( .A_N(n13461), .B(n13511), .C(n13510), .D(
        n13509), .Y(n13484) );
  sky130_fd_sc_hd__nand2_1 U20461 ( .A(n13471), .B(n17314), .Y(n15577) );
  sky130_fd_sc_hd__nand2_1 U20462 ( .A(n15577), .B(n15595), .Y(n13463) );
  sky130_fd_sc_hd__nand4_1 U20463 ( .A(n15380), .B(n15564), .C(n15538), .D(
        n15589), .Y(n13462) );
  sky130_fd_sc_hd__nor2_1 U20464 ( .A(n13463), .B(n13462), .Y(n15532) );
  sky130_fd_sc_hd__a31oi_1 U20465 ( .A1(n13465), .A2(n15532), .A3(n13464), 
        .B1(n15708), .Y(n13475) );
  sky130_fd_sc_hd__nand2b_1 U20466 ( .A_N(n17282), .B(n15309), .Y(n15609) );
  sky130_fd_sc_hd__nand2_1 U20467 ( .A(n13466), .B(n15256), .Y(n15625) );
  sky130_fd_sc_hd__nor3_1 U20468 ( .A(n13467), .B(n15625), .C(n15608), .Y(
        n13470) );
  sky130_fd_sc_hd__nand2_1 U20469 ( .A(n15577), .B(n15589), .Y(n13469) );
  sky130_fd_sc_hd__nand2_1 U20470 ( .A(n13469), .B(n13468), .Y(n15221) );
  sky130_fd_sc_hd__a21oi_1 U20471 ( .A1(n13470), .A2(n15221), .B1(n15616), .Y(
        n13474) );
  sky130_fd_sc_hd__nand2_1 U20472 ( .A(n16180), .B(n15458), .Y(n16953) );
  sky130_fd_sc_hd__nand2b_1 U20473 ( .A_N(n13471), .B(n15564), .Y(n15332) );
  sky130_fd_sc_hd__nand2_1 U20474 ( .A(n15228), .B(n15593), .Y(n15318) );
  sky130_fd_sc_hd__nor4_1 U20475 ( .A(n20513), .B(n15570), .C(n15622), .D(
        n15318), .Y(n13472) );
  sky130_fd_sc_hd__a21oi_1 U20476 ( .A1(n15251), .A2(n13472), .B1(n15384), .Y(
        n13473) );
  sky130_fd_sc_hd__nor3_1 U20477 ( .A(n13475), .B(n13474), .C(n13473), .Y(
        n13483) );
  sky130_fd_sc_hd__nand4_1 U20478 ( .A(n13476), .B(n15578), .C(n15256), .D(
        n15340), .Y(n13477) );
  sky130_fd_sc_hd__nand2_1 U20480 ( .A(n15341), .B(n15564), .Y(n15539) );
  sky130_fd_sc_hd__nand4b_1 U20481 ( .A_N(n15539), .B(n13479), .C(n15380), .D(
        n15595), .Y(n13480) );
  sky130_fd_sc_hd__nand2_1 U20482 ( .A(n13480), .B(n15630), .Y(n15231) );
  sky130_fd_sc_hd__nor2_1 U20483 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .B(n15493), .Y(n13481) );
  sky130_fd_sc_hd__a31oi_1 U20484 ( .A1(n13483), .A2(n13482), .A3(n15231), 
        .B1(n21179), .Y(n13513) );
  sky130_fd_sc_hd__nor2_1 U20485 ( .A(n13484), .B(n13513), .Y(n13485) );
  sky130_fd_sc_hd__nand2_1 U20486 ( .A(n13486), .B(
        j202_soc_core_memory0_ram_dout0_sel[8]), .Y(n13488) );
  sky130_fd_sc_hd__nand2_1 U20487 ( .A(n13500), .B(
        j202_soc_core_memory0_ram_dout0_sel[9]), .Y(n13489) );
  sky130_fd_sc_hd__nand2_1 U20488 ( .A(n13490), .B(
        j202_soc_core_memory0_ram_dout0_sel[5]), .Y(n13491) );
  sky130_fd_sc_hd__nand2_1 U20489 ( .A(n13492), .B(
        j202_soc_core_memory0_ram_dout0_sel[3]), .Y(n13493) );
  sky130_fd_sc_hd__nand2_1 U20490 ( .A(n13495), .B(
        j202_soc_core_memory0_ram_dout0_sel[4]), .Y(n13497) );
  sky130_fd_sc_hd__nand2_1 U20491 ( .A(j202_soc_core_memory0_ram_dout0[500]), 
        .B(n21771), .Y(n13516) );
  sky130_fd_sc_hd__nand4_1 U20492 ( .A(n13508), .B(n21738), .C(n13507), .D(
        n13506), .Y(n13512) );
  sky130_fd_sc_hd__nand4b_1 U20493 ( .A_N(n13512), .B(n13511), .C(n13510), .D(
        n13509), .Y(n13514) );
  sky130_fd_sc_hd__nor2_1 U20494 ( .A(n13514), .B(n13513), .Y(n13515) );
  sky130_fd_sc_hd__nand2_1 U20495 ( .A(n13516), .B(n13515), .Y(n13517) );
  sky130_fd_sc_hd__nor2_1 U20497 ( .A(n13518), .B(n24815), .Y(n13519) );
  sky130_fd_sc_hd__nand2_1 U20498 ( .A(n24005), .B(n24320), .Y(n24321) );
  sky130_fd_sc_hd__mux2i_1 U20499 ( .A0(n13519), .A1(n24321), .S(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[1]), .Y(n13520) );
  sky130_fd_sc_hd__nor2_1 U20500 ( .A(j202_soc_core_ahb2apb_02_state[0]), .B(
        j202_soc_core_ahb2apb_02_state[1]), .Y(n24317) );
  sky130_fd_sc_hd__mux2i_1 U20501 ( .A0(n13520), .A1(n24317), .S(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[2]), .Y(n13522) );
  sky130_fd_sc_hd__nor2_1 U20502 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[4]), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[3]), .Y(n13521) );
  sky130_fd_sc_hd__nand2_1 U20503 ( .A(n13522), .B(n13521), .Y(n13523) );
  sky130_fd_sc_hd__mux2i_1 U20504 ( .A0(n13523), .A1(n10539), .S(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[5]), .Y(n13524) );
  sky130_fd_sc_hd__nor2_1 U20505 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[3]), .B(
        j202_soc_core_j22_cpu_ma_M_MEM[2]), .Y(n13527) );
  sky130_fd_sc_hd__nand2_1 U20506 ( .A(n26539), .B(n13527), .Y(n13525) );
  sky130_fd_sc_hd__nor2_1 U20507 ( .A(j202_soc_core_j22_cpu_memop_MEM__1_), 
        .B(j202_soc_core_j22_cpu_memop_MEM__3_), .Y(n18915) );
  sky130_fd_sc_hd__nor2_1 U20508 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[1]), .B(
        j202_soc_core_j22_cpu_ma_M_MEM[0]), .Y(n13526) );
  sky130_fd_sc_hd__nor2_1 U20509 ( .A(n12365), .B(
        j202_soc_core_j22_cpu_regop_We__1_), .Y(n13528) );
  sky130_fd_sc_hd__nand2_1 U20510 ( .A(n13528), .B(n23279), .Y(n13529) );
  sky130_fd_sc_hd__nand2_1 U20512 ( .A(n24113), .B(n23520), .Y(n13537) );
  sky130_fd_sc_hd__xnor2_1 U20514 ( .A(n12429), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__1_), .Y(n13534) );
  sky130_fd_sc_hd__xnor2_1 U20515 ( .A(n12427), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__3_), .Y(n13533) );
  sky130_fd_sc_hd__xnor2_1 U20516 ( .A(n12431), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__0_), .Y(n13532) );
  sky130_fd_sc_hd__xnor2_1 U20517 ( .A(n12425), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__2_), .Y(n13531) );
  sky130_fd_sc_hd__nand4_1 U20518 ( .A(n13534), .B(n13533), .C(n13532), .D(
        n13531), .Y(n13535) );
  sky130_fd_sc_hd__a21o_1 U20519 ( .A1(n13537), .A2(n13536), .B1(n13535), .X(
        n13544) );
  sky130_fd_sc_hd__nor2_1 U20520 ( .A(j202_soc_core_j22_cpu_regop_We__3_), .B(
        n23279), .Y(n23446) );
  sky130_fd_sc_hd__nand2_1 U20521 ( .A(n23446), .B(n12365), .Y(n13552) );
  sky130_fd_sc_hd__nand2_1 U20522 ( .A(n24113), .B(n23174), .Y(n13543) );
  sky130_fd_sc_hd__xnor2_1 U20523 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__0_), 
        .B(j202_soc_core_j22_cpu_regop_Rn__0_), .Y(n13541) );
  sky130_fd_sc_hd__xnor2_1 U20524 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__1_), 
        .B(j202_soc_core_j22_cpu_regop_Rn__1_), .Y(n13540) );
  sky130_fd_sc_hd__xnor2_1 U20525 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__3_), 
        .B(j202_soc_core_j22_cpu_regop_Rn__3_), .Y(n13539) );
  sky130_fd_sc_hd__xnor2_1 U20526 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__2_), 
        .B(j202_soc_core_j22_cpu_regop_Rn__2_), .Y(n13538) );
  sky130_fd_sc_hd__nand2_1 U20527 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__1_), 
        .B(j202_soc_core_j22_cpu_regop_M_Wm__2_), .Y(n23283) );
  sky130_fd_sc_hd__nand2_1 U20528 ( .A(n13545), .B(n24429), .Y(n13549) );
  sky130_fd_sc_hd__nor2_1 U20529 ( .A(j202_soc_core_j22_cpu_regop_We__1_), .B(
        n13552), .Y(n23525) );
  sky130_fd_sc_hd__nand2_1 U20530 ( .A(j202_soc_core_j22_cpu_regop_Ra__0_), 
        .B(j202_soc_core_j22_cpu_regop_Ra__1_), .Y(n14752) );
  sky130_fd_sc_hd__nand2_1 U20532 ( .A(n12506), .B(n12508), .Y(n13547) );
  sky130_fd_sc_hd__nand2_1 U20533 ( .A(n13706), .B(n13546), .Y(n16014) );
  sky130_fd_sc_hd__nand2_1 U20535 ( .A(n13548), .B(
        j202_soc_core_j22_cpu_regop_Rs__1_), .Y(n22034) );
  sky130_fd_sc_hd__nor2_1 U20536 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__3_), 
        .B(n13549), .Y(n23535) );
  sky130_fd_sc_hd__nor2_1 U20537 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__1_), 
        .B(j202_soc_core_j22_cpu_regop_M_Rn__0_), .Y(n23536) );
  sky130_fd_sc_hd__nand3_1 U20538 ( .A(n23535), .B(n23536), .C(n23534), .Y(
        n13550) );
  sky130_fd_sc_hd__nor2_1 U20539 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__1_), 
        .B(n13559), .Y(n23443) );
  sky130_fd_sc_hd__nand2_1 U20540 ( .A(n23443), .B(n24429), .Y(n13556) );
  sky130_fd_sc_hd__nand2_1 U20541 ( .A(n13550), .B(n13556), .Y(n23523) );
  sky130_fd_sc_hd__nand2_1 U20542 ( .A(n13551), .B(n23523), .Y(n13595) );
  sky130_fd_sc_hd__nor2_1 U20543 ( .A(j202_soc_core_j22_cpu_regop_Rn__2_), .B(
        j202_soc_core_j22_cpu_regop_Rn__3_), .Y(n13616) );
  sky130_fd_sc_hd__nor2_1 U20544 ( .A(j202_soc_core_j22_cpu_regop_Rn__0_), .B(
        j202_soc_core_j22_cpu_regop_Rn__1_), .Y(n13613) );
  sky130_fd_sc_hd__nand2_1 U20545 ( .A(n13616), .B(n13613), .Y(n14155) );
  sky130_fd_sc_hd__nor2_1 U20546 ( .A(n12429), .B(n12431), .Y(n13666) );
  sky130_fd_sc_hd__nor2_1 U20547 ( .A(n12427), .B(n12425), .Y(n13677) );
  sky130_fd_sc_hd__nand2_1 U20548 ( .A(n13666), .B(n13677), .Y(n14231) );
  sky130_fd_sc_hd__o22ai_1 U20549 ( .A1(n14155), .A2(n13552), .B1(n14231), 
        .B2(n23172), .Y(n23524) );
  sky130_fd_sc_hd__nand2_1 U20550 ( .A(n24113), .B(n23524), .Y(n13555) );
  sky130_fd_sc_hd__inv_2 U20551 ( .A(n14231), .Y(n16498) );
  sky130_fd_sc_hd__nor2_1 U20552 ( .A(n13750), .B(n14155), .Y(n13632) );
  sky130_fd_sc_hd__a21oi_1 U20553 ( .A1(n16498), .A2(n13553), .B1(n13632), .Y(
        n13554) );
  sky130_fd_sc_hd__nand2_1 U20554 ( .A(n13555), .B(n13554), .Y(n13558) );
  sky130_fd_sc_hd__nand2_1 U20555 ( .A(n13558), .B(n13557), .Y(n13594) );
  sky130_fd_sc_hd__nor2_1 U20556 ( .A(n12508), .B(n12507), .Y(n19044) );
  sky130_fd_sc_hd__nand2_1 U20557 ( .A(n13706), .B(n19044), .Y(n16008) );
  sky130_fd_sc_hd__nand2_1 U20558 ( .A(n13559), .B(
        j202_soc_core_j22_cpu_regop_M_Wm__1_), .Y(n13561) );
  sky130_fd_sc_hd__nand2b_1 U20559 ( .A_N(n16008), .B(n23485), .Y(n16035) );
  sky130_fd_sc_hd__nor2_1 U20560 ( .A(n12506), .B(n12509), .Y(n13697) );
  sky130_fd_sc_hd__nand2_1 U20561 ( .A(n13706), .B(n13697), .Y(n16010) );
  sky130_fd_sc_hd__nand2_1 U20562 ( .A(j202_soc_core_j22_cpu_regop_Rs__1_), 
        .B(j202_soc_core_j22_cpu_regop_Rs__0_), .Y(n19054) );
  sky130_fd_sc_hd__nor2_1 U20563 ( .A(n12505), .B(n19054), .Y(n19046) );
  sky130_fd_sc_hd__nand2_1 U20564 ( .A(n19046), .B(n13697), .Y(n22854) );
  sky130_fd_sc_hd__nand2_1 U20565 ( .A(n16010), .B(n22854), .Y(n13562) );
  sky130_fd_sc_hd__nand2_1 U20566 ( .A(n23507), .B(
        j202_soc_core_j22_cpu_regop_M_Wm__0_), .Y(n23281) );
  sky130_fd_sc_hd__nor2_1 U20567 ( .A(n13561), .B(n23281), .Y(n23554) );
  sky130_fd_sc_hd__nand2_1 U20568 ( .A(n13562), .B(n23554), .Y(n13567) );
  sky130_fd_sc_hd__nand2_1 U20569 ( .A(n12505), .B(n12506), .Y(n13698) );
  sky130_fd_sc_hd__nand3_1 U20570 ( .A(n13699), .B(n13563), .C(n12509), .Y(
        n14539) );
  sky130_fd_sc_hd__nand3_1 U20571 ( .A(n13563), .B(n19051), .C(n12509), .Y(
        n22856) );
  sky130_fd_sc_hd__nand2_1 U20572 ( .A(n14539), .B(n22856), .Y(n13565) );
  sky130_fd_sc_hd__nor2_1 U20573 ( .A(n23283), .B(n23281), .Y(n13564) );
  sky130_fd_sc_hd__nand2_1 U20574 ( .A(n13565), .B(n13564), .Y(n13566) );
  sky130_fd_sc_hd__nand3_1 U20575 ( .A(n16035), .B(n13567), .C(n13566), .Y(
        n13588) );
  sky130_fd_sc_hd__nand2_1 U20576 ( .A(j202_soc_core_j22_cpu_macop_MAC_[3]), 
        .B(j202_soc_core_j22_cpu_macop_MAC_[0]), .Y(n13568) );
  sky130_fd_sc_hd__nor2_1 U20577 ( .A(n24288), .B(n13568), .Y(n13569) );
  sky130_fd_sc_hd__nand2_1 U20578 ( .A(n13568), .B(n24288), .Y(n24018) );
  sky130_fd_sc_hd__nand3_1 U20579 ( .A(n24018), .B(
        j202_soc_core_j22_cpu_macop_MAC_[2]), .C(n24293), .Y(n23322) );
  sky130_fd_sc_hd__nand3_1 U20580 ( .A(n24019), .B(
        j202_soc_core_j22_cpu_macop_MAC_[4]), .C(n24288), .Y(n24272) );
  sky130_fd_sc_hd__o21a_1 U20581 ( .A1(n13569), .A2(n23322), .B1(n24272), .X(
        n24275) );
  sky130_fd_sc_hd__inv_2 U20582 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[0]), 
        .Y(n24282) );
  sky130_fd_sc_hd__nand2_1 U20583 ( .A(n17356), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .Y(n18868) );
  sky130_fd_sc_hd__nand3_1 U20584 ( .A(n18865), .B(n24282), .C(n22055), .Y(
        n24285) );
  sky130_fd_sc_hd__and3_1 U20585 ( .A(n13576), .B(n24116), .C(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[4]), .X(n23330) );
  sky130_fd_sc_hd__nand2_1 U20586 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]), .B(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .Y(n13573) );
  sky130_fd_sc_hd__nand2_1 U20587 ( .A(n23330), .B(n13573), .Y(n23323) );
  sky130_fd_sc_hd__nand2_1 U20588 ( .A(n13575), .B(n13574), .Y(n23329) );
  sky130_fd_sc_hd__nor2_1 U20589 ( .A(j202_soc_core_j22_cpu_ml_M_macop_MAC_[4]), .B(n13576), .Y(n13580) );
  sky130_fd_sc_hd__o211ai_1 U20590 ( .A1(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .A2(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[3]), .B1(n23329), .C1(n13580), 
        .Y(n23326) );
  sky130_fd_sc_hd__nand2_1 U20591 ( .A(n23323), .B(n23326), .Y(n24290) );
  sky130_fd_sc_hd__o22ai_1 U20592 ( .A1(n24275), .A2(n13578), .B1(n24290), 
        .B2(n27456), .Y(n13581) );
  sky130_fd_sc_hd__nand2_1 U20593 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .B(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[3]), .Y(n23327) );
  sky130_fd_sc_hd__nand2_1 U20594 ( .A(n13581), .B(n27450), .Y(n13583) );
  sky130_fd_sc_hd__nand4_1 U20595 ( .A(n24019), .B(n26398), .C(n24293), .D(
        n24288), .Y(n13582) );
  sky130_fd_sc_hd__nand2_1 U20596 ( .A(n13583), .B(n13582), .Y(n13587) );
  sky130_fd_sc_hd__a21oi_1 U20597 ( .A1(n13584), .A2(n22055), .B1(n11166), .Y(
        n13585) );
  sky130_fd_sc_hd__nor2_1 U20598 ( .A(j202_soc_core_j22_cpu_macop_MAC_[4]), 
        .B(n24288), .Y(n24276) );
  sky130_fd_sc_hd__nand4_1 U20599 ( .A(n13585), .B(n18867), .C(n24276), .D(
        n18868), .Y(n13586) );
  sky130_fd_sc_hd__nand2_1 U20600 ( .A(n13587), .B(n13586), .Y(n24274) );
  sky130_fd_sc_hd__nor2_1 U20601 ( .A(n13588), .B(n24274), .Y(n13593) );
  sky130_fd_sc_hd__nand2_1 U20602 ( .A(n27910), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[3]), .Y(n26781) );
  sky130_fd_sc_hd__inv_2 U20603 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[0]), .Y(
        n26727) );
  sky130_fd_sc_hd__nor2_1 U20604 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .B(n26727), .Y(n26750) );
  sky130_fd_sc_hd__nand2_1 U20605 ( .A(n26750), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n13728) );
  sky130_fd_sc_hd__nor2_1 U20607 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[2]), 
        .B(n12381), .Y(n26749) );
  sky130_fd_sc_hd__nand3_1 U20608 ( .A(n26691), .B(n26682), .C(n26749), .Y(
        n13589) );
  sky130_fd_sc_hd__o21a_1 U20609 ( .A1(n26781), .A2(n13728), .B1(n13589), .X(
        n13592) );
  sky130_fd_sc_hd__nand2_1 U20610 ( .A(n26679), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n13590) );
  sky130_fd_sc_hd__nand2_1 U20611 ( .A(n26744), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[5]), .Y(n26757) );
  sky130_fd_sc_hd__nor2_1 U20612 ( .A(n13590), .B(n26757), .Y(n26783) );
  sky130_fd_sc_hd__nand2_1 U20613 ( .A(n26783), .B(n26727), .Y(n13591) );
  sky130_fd_sc_hd__nand2_1 U20614 ( .A(n24280), .B(
        j202_soc_core_j22_cpu_memop_MEM__1_), .Y(n18898) );
  sky130_fd_sc_hd__nand2_1 U20615 ( .A(n24279), .B(n27721), .Y(n19071) );
  sky130_fd_sc_hd__xnor2_1 U20616 ( .A(j202_soc_core_j22_cpu_regop_We__1_), 
        .B(j202_soc_core_j22_cpu_regop_We__3_), .Y(n13597) );
  sky130_fd_sc_hd__nand2_1 U20617 ( .A(n12366), .B(
        j202_soc_core_j22_cpu_regop_We__2_), .Y(n13596) );
  sky130_fd_sc_hd__o22ai_1 U20618 ( .A1(n18898), .A2(n19071), .B1(n13597), 
        .B2(n13596), .Y(n13599) );
  sky130_fd_sc_hd__nand2_1 U20619 ( .A(n22024), .B(
        j202_soc_core_j22_cpu_opst[0]), .Y(n24260) );
  sky130_fd_sc_hd__nand3_1 U20620 ( .A(n23862), .B(n22275), .C(n23195), .Y(
        n23194) );
  sky130_fd_sc_hd__nor2_1 U20621 ( .A(n24260), .B(n23194), .Y(n13598) );
  sky130_fd_sc_hd__nor3_1 U20622 ( .A(j202_soc_core_j22_cpu_istall), .B(n27919), .C(n12200), .Y(n13600) );
  sky130_fd_sc_hd__nand2_1 U20623 ( .A(n24113), .B(
        j202_soc_core_j22_cpu_ifetchl), .Y(n23487) );
  sky130_fd_sc_hd__inv_1 U20624 ( .A(j202_soc_core_j22_cpu_regop_Rn__3_), .Y(
        n13604) );
  sky130_fd_sc_hd__nand2_1 U20625 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[148]), .Y(n13610) );
  sky130_fd_sc_hd__nand2_1 U20626 ( .A(j202_soc_core_j22_cpu_regop_Rn__3_), 
        .B(j202_soc_core_j22_cpu_regop_Rn__0_), .Y(n13624) );
  sky130_fd_sc_hd__nand3_1 U20627 ( .A(n13636), .B(
        j202_soc_core_j22_cpu_regop_Rn__1_), .C(n13625), .Y(n23121) );
  sky130_fd_sc_hd__nand2_1 U20628 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[372]), .Y(n13609) );
  sky130_fd_sc_hd__nand3_1 U20629 ( .A(n13616), .B(
        j202_soc_core_j22_cpu_regop_Rn__0_), .C(
        j202_soc_core_j22_cpu_regop_Rn__1_), .Y(n23104) );
  sky130_fd_sc_hd__nor2_1 U20630 ( .A(n13638), .B(n23104), .Y(n13605) );
  sky130_fd_sc_hd__inv_2 U20631 ( .A(n13605), .Y(n14476) );
  sky130_fd_sc_hd__nand2_1 U20632 ( .A(n11116), .B(
        j202_soc_core_j22_cpu_rf_gpr[116]), .Y(n13608) );
  sky130_fd_sc_hd__nand3_1 U20633 ( .A(n13613), .B(
        j202_soc_core_j22_cpu_regop_Rn__2_), .C(
        j202_soc_core_j22_cpu_regop_Rn__3_), .Y(n23080) );
  sky130_fd_sc_hd__nor2_1 U20634 ( .A(n13638), .B(n23080), .Y(n13606) );
  sky130_fd_sc_hd__inv_2 U20635 ( .A(n13606), .Y(n15062) );
  sky130_fd_sc_hd__nand2_1 U20636 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[404]), .Y(n13607) );
  sky130_fd_sc_hd__nand4_1 U20637 ( .A(n13610), .B(n13609), .C(n13608), .D(
        n13607), .Y(n13623) );
  sky130_fd_sc_hd__nand2_1 U20638 ( .A(n13751), .B(n25782), .Y(n13612) );
  sky130_fd_sc_hd__nand2_1 U20639 ( .A(n13611), .B(n13750), .Y(n14749) );
  sky130_fd_sc_hd__a21oi_1 U20640 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[20]), .B1(n16436), .Y(n13621) );
  sky130_fd_sc_hd__nand3_1 U20641 ( .A(n13613), .B(
        j202_soc_core_j22_cpu_regop_Rn__3_), .C(n13625), .Y(n23129) );
  sky130_fd_sc_hd__nand2_1 U20642 ( .A(n16431), .B(
        j202_soc_core_j22_cpu_rf_gpr[276]), .Y(n13620) );
  sky130_fd_sc_hd__nand3_1 U20643 ( .A(n13616), .B(
        j202_soc_core_j22_cpu_regop_Rn__0_), .C(n13614), .Y(n23036) );
  sky130_fd_sc_hd__nor2_1 U20644 ( .A(n13638), .B(n23036), .Y(n13615) );
  sky130_fd_sc_hd__inv_2 U20645 ( .A(n13615), .Y(n14642) );
  sky130_fd_sc_hd__nand2_1 U20646 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[52]), .Y(n13619) );
  sky130_fd_sc_hd__nand3_1 U20647 ( .A(n13616), .B(
        j202_soc_core_j22_cpu_regop_Rn__1_), .C(n10964), .Y(n23088) );
  sky130_fd_sc_hd__nor2_1 U20648 ( .A(n13638), .B(n23088), .Y(n13617) );
  sky130_fd_sc_hd__inv_2 U20649 ( .A(n13617), .Y(n14668) );
  sky130_fd_sc_hd__nand2_1 U20650 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[84]), .Y(n13618) );
  sky130_fd_sc_hd__nand4_1 U20651 ( .A(n13621), .B(n13620), .C(n13619), .D(
        n13618), .Y(n13622) );
  sky130_fd_sc_hd__nand2_1 U20652 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[436]), .Y(n13631) );
  sky130_fd_sc_hd__nand2_1 U20653 ( .A(j202_soc_core_j22_cpu_regop_Rn__1_), 
        .B(j202_soc_core_j22_cpu_regop_Rn__2_), .Y(n13635) );
  sky130_fd_sc_hd__nand2_1 U20654 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[244]), .Y(n13630) );
  sky130_fd_sc_hd__nand2_1 U20655 ( .A(n13626), .B(n13625), .Y(n23495) );
  sky130_fd_sc_hd__nand2_1 U20656 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[308]), .Y(n13629) );
  sky130_fd_sc_hd__nand2_1 U20657 ( .A(n13627), .B(n10964), .Y(n23513) );
  sky130_fd_sc_hd__nand2_1 U20658 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_rf_gpr[212]), .Y(n13628) );
  sky130_fd_sc_hd__nand2_1 U20659 ( .A(n13633), .B(n14752), .Y(n13634) );
  sky130_fd_sc_hd__inv_2 U20660 ( .A(n13634), .Y(n14465) );
  sky130_fd_sc_hd__nand2_1 U20662 ( .A(n13641), .B(n13636), .Y(n23445) );
  sky130_fd_sc_hd__nand2_1 U20663 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[500]), .Y(n13645) );
  sky130_fd_sc_hd__nor2_1 U20664 ( .A(j202_soc_core_j22_cpu_regop_Rn__0_), .B(
        j202_soc_core_j22_cpu_regop_Rn__2_), .Y(n13637) );
  sky130_fd_sc_hd__nand3_1 U20665 ( .A(n13637), .B(
        j202_soc_core_j22_cpu_regop_Rn__1_), .C(
        j202_soc_core_j22_cpu_regop_Rn__3_), .Y(n23171) );
  sky130_fd_sc_hd__nand2_1 U20666 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[340]), .Y(n13644) );
  sky130_fd_sc_hd__nor2_1 U20667 ( .A(j202_soc_core_j22_cpu_regop_Rn__3_), .B(
        j202_soc_core_j22_cpu_regop_Rn__1_), .Y(n13639) );
  sky130_fd_sc_hd__nand3_1 U20668 ( .A(n13639), .B(
        j202_soc_core_j22_cpu_regop_Rn__0_), .C(
        j202_soc_core_j22_cpu_regop_Rn__2_), .Y(n23097) );
  sky130_fd_sc_hd__nand2_1 U20669 ( .A(n15128), .B(
        j202_soc_core_j22_cpu_rf_gpr[180]), .Y(n13643) );
  sky130_fd_sc_hd__nand3_1 U20670 ( .A(n13641), .B(
        j202_soc_core_j22_cpu_regop_Rn__3_), .C(n10964), .Y(n23500) );
  sky130_fd_sc_hd__nor2_1 U20671 ( .A(n13638), .B(n23500), .Y(n13821) );
  sky130_fd_sc_hd__nand2_1 U20672 ( .A(n16323), .B(
        j202_soc_core_j22_cpu_rf_gpr[468]), .Y(n13642) );
  sky130_fd_sc_hd__nand4_1 U20673 ( .A(n13645), .B(n13644), .C(n13643), .D(
        n13642), .Y(n13646) );
  sky130_fd_sc_hd__a21oi_1 U20674 ( .A1(j202_soc_core_j22_cpu_rf_gpr[20]), 
        .A2(n16369), .B1(n13646), .Y(n13647) );
  sky130_fd_sc_hd__inv_2 U20675 ( .A(n26717), .Y(n26417) );
  sky130_fd_sc_hd__nand3_1 U20676 ( .A(n26744), .B(n26727), .C(
        j202_soc_core_j22_cpu_exuop_EXU_[4]), .Y(n27908) );
  sky130_fd_sc_hd__nand2_1 U20677 ( .A(j202_soc_core_j22_cpu_rfuo_sr__t_), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n13650) );
  sky130_fd_sc_hd__nand2_1 U20678 ( .A(n13650), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[4]), .Y(n13652) );
  sky130_fd_sc_hd__nor2_1 U20679 ( .A(n13652), .B(n13651), .Y(n13655) );
  sky130_fd_sc_hd__nand2_1 U20680 ( .A(n12381), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n27909) );
  sky130_fd_sc_hd__nor2_1 U20681 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[2]), 
        .B(n12382), .Y(n24774) );
  sky130_fd_sc_hd__nand2_1 U20682 ( .A(n24774), .B(n23928), .Y(n13653) );
  sky130_fd_sc_hd__nor2_1 U20683 ( .A(n27908), .B(n14846), .Y(n23698) );
  sky130_fd_sc_hd__nand2b_2 U20684 ( .A_N(n14847), .B(n23698), .Y(n22592) );
  sky130_fd_sc_hd__nand3_1 U20685 ( .A(n13603), .B(
        j202_soc_core_j22_cpu_memop_Ma__1_), .C(n13656), .Y(n22590) );
  sky130_fd_sc_hd__nand2_1 U20686 ( .A(n12430), .B(n12431), .Y(n13659) );
  sky130_fd_sc_hd__nand2_1 U20687 ( .A(n12428), .B(n12425), .Y(n13682) );
  sky130_fd_sc_hd__nand2_1 U20688 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[180]), .Y(n13663) );
  sky130_fd_sc_hd__nand2_1 U20689 ( .A(n12431), .B(n12429), .Y(n13658) );
  sky130_fd_sc_hd__nor2_1 U20690 ( .A(n13658), .B(n13682), .Y(n13657) );
  sky130_fd_sc_hd__inv_2 U20691 ( .A(n13657), .Y(n14770) );
  sky130_fd_sc_hd__nand2_1 U20692 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[244]), .Y(n13662) );
  sky130_fd_sc_hd__nand2_1 U20693 ( .A(n12425), .B(n12427), .Y(n13675) );
  sky130_fd_sc_hd__nand2_1 U20694 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[500]), .Y(n13661) );
  sky130_fd_sc_hd__nand2_1 U20695 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[436]), .Y(n13660) );
  sky130_fd_sc_hd__nand4_1 U20696 ( .A(n13663), .B(n13662), .C(n13661), .D(
        n13660), .Y(n13673) );
  sky130_fd_sc_hd__nand2_1 U20697 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[20]), .Y(n13671) );
  sky130_fd_sc_hd__nand2_1 U20698 ( .A(n12430), .B(n12428), .Y(n13664) );
  sky130_fd_sc_hd__nand2_1 U20699 ( .A(n12426), .B(n12431), .Y(n13684) );
  sky130_fd_sc_hd__nand2_1 U20700 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[52]), .Y(n13670) );
  sky130_fd_sc_hd__nand2_1 U20701 ( .A(n12428), .B(n12429), .Y(n13665) );
  sky130_fd_sc_hd__nand2_1 U20702 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[116]), .Y(n13669) );
  sky130_fd_sc_hd__nor2_1 U20703 ( .A(n13675), .B(n13681), .Y(n13667) );
  sky130_fd_sc_hd__nand2_1 U20704 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[404]), .Y(n13668) );
  sky130_fd_sc_hd__nand4_1 U20705 ( .A(n13671), .B(n13670), .C(n13669), .D(
        n13668), .Y(n13672) );
  sky130_fd_sc_hd__nor2_1 U20706 ( .A(n13673), .B(n13672), .Y(n13696) );
  sky130_fd_sc_hd__nand2_1 U20707 ( .A(n12430), .B(n12427), .Y(n13674) );
  sky130_fd_sc_hd__nor2_1 U20708 ( .A(n13674), .B(n13684), .Y(n14725) );
  sky130_fd_sc_hd__nor2_1 U20709 ( .A(n13675), .B(n13687), .Y(n14724) );
  sky130_fd_sc_hd__a22oi_1 U20710 ( .A1(n11160), .A2(
        j202_soc_core_j22_cpu_rf_gpr[308]), .B1(n23502), .B2(
        j202_soc_core_j22_cpu_rf_gpr[468]), .Y(n13695) );
  sky130_fd_sc_hd__nor2_1 U20711 ( .A(n13682), .B(n13687), .Y(n13676) );
  sky130_fd_sc_hd__a22oi_1 U20713 ( .A1(n16470), .A2(
        j202_soc_core_j22_cpu_rf_gpr[212]), .B1(n23089), .B2(
        j202_soc_core_j22_cpu_rf_gpr[84]), .Y(n13694) );
  sky130_fd_sc_hd__nand2_1 U20714 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[276]), .Y(n13692) );
  sky130_fd_sc_hd__nor2_1 U20715 ( .A(n13682), .B(n13681), .Y(n13683) );
  sky130_fd_sc_hd__nand2_1 U20716 ( .A(n16471), .B(
        j202_soc_core_j22_cpu_rf_gpr[148]), .Y(n13691) );
  sky130_fd_sc_hd__nand2_1 U20717 ( .A(n12429), .B(n12427), .Y(n13685) );
  sky130_fd_sc_hd__nor2_1 U20718 ( .A(n13685), .B(n13684), .Y(n13686) );
  sky130_fd_sc_hd__nand2_1 U20719 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[372]), .Y(n13690) );
  sky130_fd_sc_hd__nand2_1 U20720 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[340]), .Y(n13689) );
  sky130_fd_sc_hd__and4_1 U20721 ( .A(n13692), .B(n13691), .C(n13690), .D(
        n13689), .X(n13693) );
  sky130_fd_sc_hd__nand4_1 U20722 ( .A(n13696), .B(n13695), .C(n13694), .D(
        n13693), .Y(n22149) );
  sky130_fd_sc_hd__nand2_1 U20723 ( .A(n22149), .B(n16513), .Y(n13712) );
  sky130_fd_sc_hd__nand2_1 U20724 ( .A(n13697), .B(n12505), .Y(n19050) );
  sky130_fd_sc_hd__nand2_1 U20725 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[20]), .Y(n13705) );
  sky130_fd_sc_hd__nor2_1 U20726 ( .A(n12509), .B(n13698), .Y(n19052) );
  sky130_fd_sc_hd__nand2_1 U20727 ( .A(n19052), .B(n13699), .Y(n16007) );
  sky130_fd_sc_hd__inv_2 U20728 ( .A(n16007), .Y(n16514) );
  sky130_fd_sc_hd__nand2_1 U20729 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[20]), .Y(n13704) );
  sky130_fd_sc_hd__nor2_1 U20730 ( .A(n12350), .B(n13700), .Y(n13701) );
  sky130_fd_sc_hd__nand2_2 U20731 ( .A(n13701), .B(n10920), .Y(n16516) );
  sky130_fd_sc_hd__nor2_1 U20732 ( .A(n12508), .B(n12506), .Y(n19045) );
  sky130_fd_sc_hd__nand2_1 U20733 ( .A(n19045), .B(n12505), .Y(n19053) );
  sky130_fd_sc_hd__nand2_1 U20734 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[500]), .Y(n13703) );
  sky130_fd_sc_hd__and4_1 U20735 ( .A(n13705), .B(n13704), .C(n16516), .D(
        n13703), .X(n13711) );
  sky130_fd_sc_hd__inv_2 U20736 ( .A(n16008), .Y(n16519) );
  sky130_fd_sc_hd__nand2_1 U20737 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[20]), .Y(n13710) );
  sky130_fd_sc_hd__inv_2 U20738 ( .A(n16014), .Y(n16520) );
  sky130_fd_sc_hd__nand2_1 U20739 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[20]), .Y(n13709) );
  sky130_fd_sc_hd__inv_2 U20740 ( .A(n16010), .Y(n16521) );
  sky130_fd_sc_hd__nand2_1 U20741 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[20]), .Y(n13708) );
  sky130_fd_sc_hd__nand2_1 U20742 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[20]), .Y(n13707) );
  sky130_fd_sc_hd__nand3_1 U20743 ( .A(n13712), .B(n13711), .C(n13345), .Y(
        n27419) );
  sky130_fd_sc_hd__nand2_1 U20744 ( .A(n22515), .B(n27419), .Y(n13723) );
  sky130_fd_sc_hd__nor2_1 U20745 ( .A(n26727), .B(n14846), .Y(n23701) );
  sky130_fd_sc_hd__nand2_1 U20746 ( .A(j202_soc_core_j22_cpu_pc[17]), .B(
        j202_soc_core_j22_cpu_pc[18]), .Y(n15030) );
  sky130_fd_sc_hd__nand2_1 U20747 ( .A(j202_soc_core_j22_cpu_pc[7]), .B(
        j202_soc_core_j22_cpu_pc[8]), .Y(n13713) );
  sky130_fd_sc_hd__nand2_1 U20748 ( .A(j202_soc_core_j22_cpu_pc[5]), .B(
        j202_soc_core_j22_cpu_pc[6]), .Y(n19077) );
  sky130_fd_sc_hd__nor2_1 U20749 ( .A(n13713), .B(n19077), .Y(n13715) );
  sky130_fd_sc_hd__nand2_1 U20750 ( .A(j202_soc_core_j22_cpu_pc[3]), .B(
        j202_soc_core_j22_cpu_pc[4]), .Y(n13714) );
  sky130_fd_sc_hd__nand2_1 U20751 ( .A(j202_soc_core_j22_cpu_pc[1]), .B(
        j202_soc_core_j22_cpu_pc[2]), .Y(n20284) );
  sky130_fd_sc_hd__nor2_1 U20752 ( .A(n13714), .B(n20284), .Y(n19076) );
  sky130_fd_sc_hd__nand2_1 U20753 ( .A(n13715), .B(n19076), .Y(n20989) );
  sky130_fd_sc_hd__nand2_1 U20754 ( .A(j202_soc_core_j22_cpu_pc[11]), .B(
        j202_soc_core_j22_cpu_pc[12]), .Y(n13716) );
  sky130_fd_sc_hd__nand2_1 U20755 ( .A(j202_soc_core_j22_cpu_pc[9]), .B(
        j202_soc_core_j22_cpu_pc[10]), .Y(n21352) );
  sky130_fd_sc_hd__nor2_1 U20756 ( .A(n13716), .B(n21352), .Y(n20990) );
  sky130_fd_sc_hd__nand2_1 U20757 ( .A(j202_soc_core_j22_cpu_pc[15]), .B(
        j202_soc_core_j22_cpu_pc[16]), .Y(n13717) );
  sky130_fd_sc_hd__nand2_1 U20758 ( .A(j202_soc_core_j22_cpu_pc[13]), .B(
        j202_soc_core_j22_cpu_pc[14]), .Y(n20991) );
  sky130_fd_sc_hd__nor2_1 U20759 ( .A(n13717), .B(n20991), .Y(n13718) );
  sky130_fd_sc_hd__nand2_1 U20760 ( .A(n20990), .B(n13718), .Y(n13719) );
  sky130_fd_sc_hd__nor2_1 U20761 ( .A(n20989), .B(n13719), .Y(n16029) );
  sky130_fd_sc_hd__nor2_1 U20762 ( .A(n15030), .B(n21009), .Y(n15766) );
  sky130_fd_sc_hd__nand2_1 U20763 ( .A(n15766), .B(
        j202_soc_core_j22_cpu_pc[19]), .Y(n13721) );
  sky130_fd_sc_hd__xor2_1 U20764 ( .A(n13721), .B(n13720), .X(n24542) );
  sky130_fd_sc_hd__nand2_1 U20765 ( .A(n22596), .B(n24542), .Y(n13722) );
  sky130_fd_sc_hd__nand2_1 U20766 ( .A(n26727), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n19013) );
  sky130_fd_sc_hd__nand2_1 U20767 ( .A(n13725), .B(n12382), .Y(n13727) );
  sky130_fd_sc_hd__nand2_1 U20768 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n19003) );
  sky130_fd_sc_hd__nand2_1 U20769 ( .A(n26744), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[4]), .Y(n13726) );
  sky130_fd_sc_hd__nand3_1 U20770 ( .A(n13727), .B(n19003), .C(n13726), .Y(
        n14008) );
  sky130_fd_sc_hd__nor2_1 U20771 ( .A(n13724), .B(n14008), .Y(n14006) );
  sky130_fd_sc_hd__nor2_1 U20772 ( .A(n12381), .B(n26781), .Y(n26739) );
  sky130_fd_sc_hd__nand2_1 U20773 ( .A(n13728), .B(n27910), .Y(n13729) );
  sky130_fd_sc_hd__nor2_1 U20774 ( .A(n26739), .B(n13729), .Y(n13788) );
  sky130_fd_sc_hd__o21ai_1 U20775 ( .A1(j202_soc_core_j22_cpu_exuop_EXU_[0]), 
        .A2(j202_soc_core_j22_cpu_exuop_EXU_[4]), .B1(
        j202_soc_core_j22_cpu_exuop_EXU_[3]), .Y(n13730) );
  sky130_fd_sc_hd__nand2_1 U20776 ( .A(n13730), .B(n27909), .Y(n13789) );
  sky130_fd_sc_hd__nor2_1 U20777 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[2]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[4]), .Y(n26755) );
  sky130_fd_sc_hd__nand2_1 U20778 ( .A(n12381), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[0]), .Y(n26782) );
  sky130_fd_sc_hd__nand2_1 U20779 ( .A(n12381), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[3]), .Y(n13731) );
  sky130_fd_sc_hd__nand3_1 U20780 ( .A(n26755), .B(n26782), .C(n13731), .Y(
        n13791) );
  sky130_fd_sc_hd__nor2_1 U20781 ( .A(n13789), .B(n13732), .Y(n13733) );
  sky130_fd_sc_hd__nand3_1 U20782 ( .A(n14006), .B(n13788), .C(n13733), .Y(
        n16289) );
  sky130_fd_sc_hd__inv_2 U20783 ( .A(n16289), .Y(n16492) );
  sky130_fd_sc_hd__nand2_1 U20784 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[131]), .Y(n13737) );
  sky130_fd_sc_hd__nand2_1 U20785 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[355]), .Y(n13736) );
  sky130_fd_sc_hd__nand2_1 U20786 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[99]), .Y(n13735) );
  sky130_fd_sc_hd__nand2_1 U20787 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[67]), .Y(n13734) );
  sky130_fd_sc_hd__nand4_1 U20788 ( .A(n13737), .B(n13736), .C(n13735), .D(
        n13734), .Y(n13742) );
  sky130_fd_sc_hd__nand2_1 U20789 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[291]), .Y(n13740) );
  sky130_fd_sc_hd__nand2_1 U20790 ( .A(n11154), .B(
        j202_soc_core_j22_cpu_rf_gpr[259]), .Y(n13739) );
  sky130_fd_sc_hd__nand2_1 U20791 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[387]), .Y(n13738) );
  sky130_fd_sc_hd__nand3_1 U20792 ( .A(n13740), .B(n13739), .C(n13738), .Y(
        n13741) );
  sky130_fd_sc_hd__nor2_1 U20793 ( .A(n13742), .B(n13741), .Y(n13760) );
  sky130_fd_sc_hd__nand2_1 U20794 ( .A(n16369), .B(
        j202_soc_core_j22_cpu_rf_gpr[3]), .Y(n13746) );
  sky130_fd_sc_hd__nand2_1 U20795 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[419]), .Y(n13745) );
  sky130_fd_sc_hd__nand2_1 U20796 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[227]), .Y(n13744) );
  sky130_fd_sc_hd__nand2_1 U20797 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_rf_gpr[195]), .Y(n13743) );
  sky130_fd_sc_hd__nand2_1 U20798 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[35]), .Y(n13749) );
  sky130_fd_sc_hd__nand2_1 U20799 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[163]), .Y(n13748) );
  sky130_fd_sc_hd__nand2_1 U20800 ( .A(n14393), .B(n10931), .Y(n13747) );
  sky130_fd_sc_hd__nand3_1 U20801 ( .A(n13749), .B(n13748), .C(n13747), .Y(
        n13758) );
  sky130_fd_sc_hd__nand2_1 U20802 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[483]), .Y(n13756) );
  sky130_fd_sc_hd__a2bb2oi_1 U20803 ( .B1(n13752), .B2(
        j202_soc_core_intr_vec__1_), .A1_N(n21413), .A2_N(n14749), .Y(n13755)
         );
  sky130_fd_sc_hd__nand2_1 U20804 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[323]), .Y(n13754) );
  sky130_fd_sc_hd__nand2_1 U20805 ( .A(n16323), .B(
        j202_soc_core_j22_cpu_rf_gpr[451]), .Y(n13753) );
  sky130_fd_sc_hd__nand4_1 U20806 ( .A(n13756), .B(n13755), .C(n13754), .D(
        n13753), .Y(n13757) );
  sky130_fd_sc_hd__nor2_1 U20807 ( .A(n13758), .B(n13757), .Y(n13759) );
  sky130_fd_sc_hd__inv_2 U20808 ( .A(n22723), .Y(n26713) );
  sky130_fd_sc_hd__nand2_1 U20809 ( .A(n11154), .B(
        j202_soc_core_j22_cpu_rf_gpr[258]), .Y(n13764) );
  sky130_fd_sc_hd__nand2_1 U20810 ( .A(n13821), .B(
        j202_soc_core_j22_cpu_rf_gpr[450]), .Y(n13763) );
  sky130_fd_sc_hd__nand2_1 U20811 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[386]), .Y(n13762) );
  sky130_fd_sc_hd__nand2_1 U20812 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[130]), .Y(n13761) );
  sky130_fd_sc_hd__nand4_1 U20813 ( .A(n13764), .B(n13763), .C(n13762), .D(
        n13761), .Y(n13769) );
  sky130_fd_sc_hd__nand2_1 U20814 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[418]), .Y(n13767) );
  sky130_fd_sc_hd__nand2_1 U20815 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[98]), .Y(n13766) );
  sky130_fd_sc_hd__nand2_1 U20816 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[34]), .Y(n13765) );
  sky130_fd_sc_hd__nand3_1 U20817 ( .A(n13767), .B(n13766), .C(n13765), .Y(
        n13768) );
  sky130_fd_sc_hd__nor2_1 U20818 ( .A(n13769), .B(n13768), .Y(n13786) );
  sky130_fd_sc_hd__nand2_1 U20819 ( .A(n16369), .B(
        j202_soc_core_j22_cpu_rf_gpr[2]), .Y(n13773) );
  sky130_fd_sc_hd__nand2_1 U20820 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[226]), .Y(n13772) );
  sky130_fd_sc_hd__nand2_1 U20821 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[290]), .Y(n13771) );
  sky130_fd_sc_hd__nand2_1 U20822 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_rf_gpr[194]), .Y(n13770) );
  sky130_fd_sc_hd__nand2_1 U20823 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[66]), .Y(n13777) );
  sky130_fd_sc_hd__nand2_1 U20824 ( .A(n13774), .B(
        j202_soc_core_j22_cpu_rf_tmp[2]), .Y(n13776) );
  sky130_fd_sc_hd__nand2_1 U20825 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[162]), .Y(n13775) );
  sky130_fd_sc_hd__nand3_1 U20826 ( .A(n13777), .B(n13776), .C(n13775), .Y(
        n13783) );
  sky130_fd_sc_hd__nand2_1 U20827 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[482]), .Y(n13781) );
  sky130_fd_sc_hd__a2bb2oi_1 U20828 ( .B1(n13752), .B2(
        j202_soc_core_intr_vec__0_), .A1_N(n10930), .A2_N(n14466), .Y(n13780)
         );
  sky130_fd_sc_hd__nand2_1 U20829 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[322]), .Y(n13779) );
  sky130_fd_sc_hd__nand2_1 U20830 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[354]), .Y(n13778) );
  sky130_fd_sc_hd__nand4_1 U20831 ( .A(n13781), .B(n13780), .C(n13779), .D(
        n13778), .Y(n13782) );
  sky130_fd_sc_hd__inv_2 U20832 ( .A(n23920), .Y(n25229) );
  sky130_fd_sc_hd__nor2_1 U20833 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .B(n26744), .Y(n16261) );
  sky130_fd_sc_hd__o22ai_1 U20834 ( .A1(n16492), .A2(n26713), .B1(n25229), 
        .B2(n13793), .Y(n14121) );
  sky130_fd_sc_hd__xnor2_1 U20835 ( .A(j202_soc_core_j22_cpu_rfuo_sr__m_), .B(
        j202_soc_core_j22_cpu_rfuo_sr__q_), .Y(n13792) );
  sky130_fd_sc_hd__nand2_1 U20836 ( .A(n13792), .B(n16261), .Y(n13787) );
  sky130_fd_sc_hd__nand2_1 U20837 ( .A(n13788), .B(n13787), .Y(n14009) );
  sky130_fd_sc_hd__inv_2 U20838 ( .A(n16322), .Y(n14742) );
  sky130_fd_sc_hd__o21a_1 U20839 ( .A1(n13793), .A2(n13792), .B1(n13791), .X(
        n14059) );
  sky130_fd_sc_hd__nand2_2 U20840 ( .A(n14006), .B(n14059), .Y(n16529) );
  sky130_fd_sc_hd__inv_2 U20841 ( .A(n16529), .Y(n16320) );
  sky130_fd_sc_hd__nand2_1 U20842 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[163]), .Y(n13798) );
  sky130_fd_sc_hd__nand2_1 U20843 ( .A(n15982), .B(
        j202_soc_core_j22_cpu_rf_gpr[227]), .Y(n13797) );
  sky130_fd_sc_hd__nand2_1 U20844 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[483]), .Y(n13796) );
  sky130_fd_sc_hd__nand2_1 U20845 ( .A(n15983), .B(
        j202_soc_core_j22_cpu_rf_gpr[419]), .Y(n13795) );
  sky130_fd_sc_hd__nand4_1 U20846 ( .A(n13798), .B(n13797), .C(n13796), .D(
        n13795), .Y(n13804) );
  sky130_fd_sc_hd__nand2_1 U20847 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[3]), .Y(n13802) );
  sky130_fd_sc_hd__nand2_1 U20848 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[35]), .Y(n13801) );
  sky130_fd_sc_hd__nand2_1 U20849 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[99]), .Y(n13800) );
  sky130_fd_sc_hd__nand2_1 U20850 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[387]), .Y(n13799) );
  sky130_fd_sc_hd__nand4_1 U20851 ( .A(n13802), .B(n13801), .C(n13800), .D(
        n13799), .Y(n13803) );
  sky130_fd_sc_hd__nor2_1 U20852 ( .A(n13804), .B(n13803), .Y(n13811) );
  sky130_fd_sc_hd__a22oi_1 U20853 ( .A1(n11160), .A2(
        j202_soc_core_j22_cpu_rf_gpr[291]), .B1(n23502), .B2(
        j202_soc_core_j22_cpu_rf_gpr[451]), .Y(n13810) );
  sky130_fd_sc_hd__inv_2 U20854 ( .A(n14496), .Y(n23515) );
  sky130_fd_sc_hd__a22oi_1 U20855 ( .A1(n23515), .A2(
        j202_soc_core_j22_cpu_rf_gpr[195]), .B1(n23089), .B2(
        j202_soc_core_j22_cpu_rf_gpr[67]), .Y(n13809) );
  sky130_fd_sc_hd__nand2_1 U20856 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[259]), .Y(n13808) );
  sky130_fd_sc_hd__inv_2 U20857 ( .A(n23109), .Y(n23113) );
  sky130_fd_sc_hd__nand2_1 U20858 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[131]), .Y(n13807) );
  sky130_fd_sc_hd__nand2_1 U20859 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[355]), .Y(n13806) );
  sky130_fd_sc_hd__nand2_1 U20860 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[323]), .Y(n13805) );
  sky130_fd_sc_hd__nand4_1 U20861 ( .A(n13811), .B(n13810), .C(n13809), .D(
        n12221), .Y(n21410) );
  sky130_fd_sc_hd__nand2_1 U20862 ( .A(n21410), .B(n16513), .Y(n13820) );
  sky130_fd_sc_hd__nand2_1 U20863 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[3]), .Y(n13815) );
  sky130_fd_sc_hd__nand2_1 U20864 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[3]), .Y(n13814) );
  sky130_fd_sc_hd__nand2_1 U20865 ( .A(n13701), .B(n10931), .Y(n13813) );
  sky130_fd_sc_hd__nand2_1 U20866 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[483]), .Y(n13812) );
  sky130_fd_sc_hd__nand2_1 U20867 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[3]), .Y(n13819) );
  sky130_fd_sc_hd__nand2_1 U20868 ( .A(n16519), .B(j202_soc_core_j22_cpu_pc[3]), .Y(n13818) );
  sky130_fd_sc_hd__nand2_1 U20869 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[3]), .Y(n13817) );
  sky130_fd_sc_hd__nand2_1 U20870 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[3]), .Y(n13816) );
  sky130_fd_sc_hd__mux2i_1 U20872 ( .A0(n14742), .A1(n16320), .S(n27429), .Y(
        n14122) );
  sky130_fd_sc_hd__nor2_1 U20873 ( .A(n14121), .B(n14122), .Y(n19416) );
  sky130_fd_sc_hd__nand2_1 U20874 ( .A(n11114), .B(
        j202_soc_core_j22_cpu_rf_gpr[388]), .Y(n13825) );
  sky130_fd_sc_hd__nand2_1 U20875 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[452]), .Y(n13824) );
  sky130_fd_sc_hd__nand2_1 U20876 ( .A(n16431), .B(
        j202_soc_core_j22_cpu_rf_gpr[260]), .Y(n13823) );
  sky130_fd_sc_hd__nand2_1 U20877 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[132]), .Y(n13822) );
  sky130_fd_sc_hd__nand4_1 U20878 ( .A(n13825), .B(n13824), .C(n13823), .D(
        n13822), .Y(n13830) );
  sky130_fd_sc_hd__nand2_1 U20879 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[420]), .Y(n13828) );
  sky130_fd_sc_hd__nand2_1 U20880 ( .A(n11116), .B(
        j202_soc_core_j22_cpu_rf_gpr[100]), .Y(n13827) );
  sky130_fd_sc_hd__nand2_1 U20881 ( .A(n11152), .B(
        j202_soc_core_j22_cpu_rf_gpr[36]), .Y(n13826) );
  sky130_fd_sc_hd__nand3_1 U20882 ( .A(n13828), .B(n13827), .C(n13826), .Y(
        n13829) );
  sky130_fd_sc_hd__nor2_1 U20883 ( .A(n13830), .B(n13829), .Y(n13845) );
  sky130_fd_sc_hd__nand2_1 U20884 ( .A(n16369), .B(
        j202_soc_core_j22_cpu_rf_gpr[4]), .Y(n13834) );
  sky130_fd_sc_hd__nand2_1 U20885 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[228]), .Y(n13833) );
  sky130_fd_sc_hd__nand2_1 U20886 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[292]), .Y(n13832) );
  sky130_fd_sc_hd__nand2_1 U20887 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_rf_gpr[196]), .Y(n13831) );
  sky130_fd_sc_hd__nand2_1 U20888 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[68]), .Y(n13837) );
  sky130_fd_sc_hd__nand2_1 U20889 ( .A(n13774), .B(
        j202_soc_core_j22_cpu_rf_tmp[4]), .Y(n13836) );
  sky130_fd_sc_hd__nand2_1 U20890 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[164]), .Y(n13835) );
  sky130_fd_sc_hd__nand3_1 U20891 ( .A(n13837), .B(n13836), .C(n13835), .Y(
        n13843) );
  sky130_fd_sc_hd__nand2_1 U20892 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[484]), .Y(n13841) );
  sky130_fd_sc_hd__a2bb2oi_1 U20893 ( .B1(n13752), .B2(
        j202_soc_core_intr_vec__2_), .A1_N(n10982), .A2_N(n14466), .Y(n13840)
         );
  sky130_fd_sc_hd__nand2_1 U20894 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[324]), .Y(n13839) );
  sky130_fd_sc_hd__nand2_1 U20895 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[356]), .Y(n13838) );
  sky130_fd_sc_hd__nand4_1 U20896 ( .A(n13841), .B(n13840), .C(n13839), .D(
        n13838), .Y(n13842) );
  sky130_fd_sc_hd__nor2_1 U20897 ( .A(n13843), .B(n13842), .Y(n13844) );
  sky130_fd_sc_hd__o22ai_1 U20898 ( .A1(n16492), .A2(n27007), .B1(n26713), 
        .B2(n13793), .Y(n14123) );
  sky130_fd_sc_hd__nand2_1 U20899 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[164]), .Y(n13849) );
  sky130_fd_sc_hd__nand2_1 U20900 ( .A(n15982), .B(
        j202_soc_core_j22_cpu_rf_gpr[228]), .Y(n13848) );
  sky130_fd_sc_hd__nand2_1 U20901 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[484]), .Y(n13847) );
  sky130_fd_sc_hd__nand2_1 U20902 ( .A(n15983), .B(
        j202_soc_core_j22_cpu_rf_gpr[420]), .Y(n13846) );
  sky130_fd_sc_hd__nand4_1 U20903 ( .A(n13849), .B(n13848), .C(n13847), .D(
        n13846), .Y(n13855) );
  sky130_fd_sc_hd__nand2_1 U20904 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[4]), .Y(n13853) );
  sky130_fd_sc_hd__nand2_1 U20905 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[36]), .Y(n13852) );
  sky130_fd_sc_hd__nand2_1 U20906 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[100]), .Y(n13851) );
  sky130_fd_sc_hd__nand2_1 U20907 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[388]), .Y(n13850) );
  sky130_fd_sc_hd__nand4_1 U20908 ( .A(n13853), .B(n13852), .C(n13851), .D(
        n13850), .Y(n13854) );
  sky130_fd_sc_hd__nor2_1 U20909 ( .A(n13855), .B(n13854), .Y(n13867) );
  sky130_fd_sc_hd__nand2_1 U20910 ( .A(n16469), .B(
        j202_soc_core_j22_cpu_rf_gpr[68]), .Y(n13859) );
  sky130_fd_sc_hd__nand2_1 U20911 ( .A(n16470), .B(
        j202_soc_core_j22_cpu_rf_gpr[196]), .Y(n13858) );
  sky130_fd_sc_hd__nand2_1 U20912 ( .A(n11160), .B(
        j202_soc_core_j22_cpu_rf_gpr[292]), .Y(n13857) );
  sky130_fd_sc_hd__nand2_1 U20913 ( .A(n14414), .B(
        j202_soc_core_j22_cpu_rf_gpr[452]), .Y(n13856) );
  sky130_fd_sc_hd__and4_1 U20914 ( .A(n13859), .B(n13858), .C(n13857), .D(
        n13856), .X(n13866) );
  sky130_fd_sc_hd__nand2_1 U20915 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[260]), .Y(n13864) );
  sky130_fd_sc_hd__nand2_1 U20916 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[132]), .Y(n13863) );
  sky130_fd_sc_hd__nand2_1 U20917 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[356]), .Y(n13862) );
  sky130_fd_sc_hd__nand2_1 U20918 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[324]), .Y(n13861) );
  sky130_fd_sc_hd__and4_1 U20919 ( .A(n13864), .B(n13863), .C(n13862), .D(
        n13861), .X(n13865) );
  sky130_fd_sc_hd__nand3_1 U20920 ( .A(n13867), .B(n13866), .C(n13865), .Y(
        n19449) );
  sky130_fd_sc_hd__a22oi_1 U20921 ( .A1(n29563), .A2(
        j202_soc_core_j22_cpu_rf_gpr[484]), .B1(n29567), .B2(
        j202_soc_core_j22_cpu_rf_vbr[4]), .Y(n13872) );
  sky130_fd_sc_hd__o2bb2ai_1 U20922 ( .B1(n19451), .B2(n14539), .A1_N(n13701), 
        .A2_N(n10981), .Y(n13868) );
  sky130_fd_sc_hd__a21oi_1 U20923 ( .A1(n16012), .A2(
        j202_soc_core_j22_cpu_rf_gbr[4]), .B1(n13868), .Y(n13871) );
  sky130_fd_sc_hd__o22a_1 U20924 ( .A1(n19450), .A2(n16010), .B1(n16007), .B2(
        n19456), .X(n13870) );
  sky130_fd_sc_hd__o22a_1 U20925 ( .A1(n19457), .A2(n16014), .B1(n19453), .B2(
        n16008), .X(n13869) );
  sky130_fd_sc_hd__nand4_1 U20926 ( .A(n13872), .B(n13871), .C(n13870), .D(
        n13869), .Y(n13873) );
  sky130_fd_sc_hd__a21oi_2 U20927 ( .A1(n19449), .A2(n16513), .B1(n13873), .Y(
        n26791) );
  sky130_fd_sc_hd__mux2i_1 U20928 ( .A0(n16320), .A1(n14742), .S(n26791), .Y(
        n14124) );
  sky130_fd_sc_hd__nor2_1 U20929 ( .A(n14123), .B(n14124), .Y(n19418) );
  sky130_fd_sc_hd__nor2_1 U20930 ( .A(n19416), .B(n19418), .Y(n21530) );
  sky130_fd_sc_hd__nand2_1 U20931 ( .A(n16324), .B(
        j202_soc_core_j22_cpu_rf_gpr[262]), .Y(n13877) );
  sky130_fd_sc_hd__nand2_1 U20932 ( .A(n16323), .B(
        j202_soc_core_j22_cpu_rf_gpr[454]), .Y(n13876) );
  sky130_fd_sc_hd__nand2_1 U20933 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[134]), .Y(n13875) );
  sky130_fd_sc_hd__nand2_1 U20934 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[102]), .Y(n13874) );
  sky130_fd_sc_hd__nand4_1 U20935 ( .A(n13877), .B(n13876), .C(n13875), .D(
        n13874), .Y(n13882) );
  sky130_fd_sc_hd__nand2_1 U20936 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[230]), .Y(n13880) );
  sky130_fd_sc_hd__nand2_1 U20937 ( .A(n11152), .B(
        j202_soc_core_j22_cpu_rf_gpr[38]), .Y(n13879) );
  sky130_fd_sc_hd__nand2_1 U20938 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[390]), .Y(n13878) );
  sky130_fd_sc_hd__nand3_1 U20939 ( .A(n13880), .B(n13879), .C(n13878), .Y(
        n13881) );
  sky130_fd_sc_hd__nor2_1 U20940 ( .A(n13882), .B(n13881), .Y(n13897) );
  sky130_fd_sc_hd__nand2_1 U20941 ( .A(n16369), .B(
        j202_soc_core_j22_cpu_rf_gpr[6]), .Y(n13886) );
  sky130_fd_sc_hd__nand2_1 U20942 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[198]), .Y(n13885) );
  sky130_fd_sc_hd__nand2_1 U20943 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[422]), .Y(n13884) );
  sky130_fd_sc_hd__nand2_1 U20944 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[294]), .Y(n13883) );
  sky130_fd_sc_hd__nand2_1 U20945 ( .A(n11155), .B(
        j202_soc_core_j22_cpu_rf_gpr[70]), .Y(n13889) );
  sky130_fd_sc_hd__nand2_1 U20946 ( .A(n14393), .B(n10983), .Y(n13888) );
  sky130_fd_sc_hd__nand2_1 U20947 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[166]), .Y(n13887) );
  sky130_fd_sc_hd__nand3_1 U20948 ( .A(n13889), .B(n13888), .C(n13887), .Y(
        n13895) );
  sky130_fd_sc_hd__nand2_1 U20949 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[486]), .Y(n13893) );
  sky130_fd_sc_hd__a2bb2oi_1 U20950 ( .B1(n13752), .B2(
        j202_soc_core_intr_vec__4_), .A1_N(n13940), .A2_N(n14749), .Y(n13892)
         );
  sky130_fd_sc_hd__nand2_1 U20951 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[326]), .Y(n13891) );
  sky130_fd_sc_hd__nand2_1 U20952 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[358]), .Y(n13890) );
  sky130_fd_sc_hd__nand4_1 U20953 ( .A(n13893), .B(n13892), .C(n13891), .D(
        n13890), .Y(n13894) );
  sky130_fd_sc_hd__nor2_1 U20954 ( .A(n13895), .B(n13894), .Y(n13896) );
  sky130_fd_sc_hd__nand2_1 U20955 ( .A(n16324), .B(
        j202_soc_core_j22_cpu_rf_gpr[261]), .Y(n13901) );
  sky130_fd_sc_hd__nand2_1 U20956 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[453]), .Y(n13900) );
  sky130_fd_sc_hd__nand2_1 U20957 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[389]), .Y(n13899) );
  sky130_fd_sc_hd__nand2_1 U20958 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[133]), .Y(n13898) );
  sky130_fd_sc_hd__nand4_1 U20959 ( .A(n13901), .B(n13900), .C(n13899), .D(
        n13898), .Y(n13906) );
  sky130_fd_sc_hd__nand2_1 U20960 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[421]), .Y(n13904) );
  sky130_fd_sc_hd__nand2_1 U20961 ( .A(n11116), .B(
        j202_soc_core_j22_cpu_rf_gpr[101]), .Y(n13903) );
  sky130_fd_sc_hd__nand2_1 U20962 ( .A(n11152), .B(
        j202_soc_core_j22_cpu_rf_gpr[37]), .Y(n13902) );
  sky130_fd_sc_hd__nand3_1 U20963 ( .A(n13904), .B(n13903), .C(n13902), .Y(
        n13905) );
  sky130_fd_sc_hd__nor2_1 U20964 ( .A(n13906), .B(n13905), .Y(n13921) );
  sky130_fd_sc_hd__nand2_1 U20965 ( .A(n16369), .B(
        j202_soc_core_j22_cpu_rf_gpr[5]), .Y(n13910) );
  sky130_fd_sc_hd__nand2_1 U20966 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[229]), .Y(n13909) );
  sky130_fd_sc_hd__nand2_1 U20967 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[293]), .Y(n13908) );
  sky130_fd_sc_hd__nand2_1 U20968 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[197]), .Y(n13907) );
  sky130_fd_sc_hd__nand2_1 U20969 ( .A(n11155), .B(
        j202_soc_core_j22_cpu_rf_gpr[69]), .Y(n13913) );
  sky130_fd_sc_hd__nand2_1 U20970 ( .A(n13774), .B(
        j202_soc_core_j22_cpu_rf_tmp[5]), .Y(n13912) );
  sky130_fd_sc_hd__nand2_1 U20971 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[165]), .Y(n13911) );
  sky130_fd_sc_hd__nand3_1 U20972 ( .A(n13913), .B(n13912), .C(n13911), .Y(
        n13919) );
  sky130_fd_sc_hd__nand2_1 U20973 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[485]), .Y(n13917) );
  sky130_fd_sc_hd__nand2_1 U20974 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[325]), .Y(n13915) );
  sky130_fd_sc_hd__nand2_1 U20975 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[357]), .Y(n13914) );
  sky130_fd_sc_hd__nand4_1 U20976 ( .A(n13917), .B(n13916), .C(n13915), .D(
        n13914), .Y(n13918) );
  sky130_fd_sc_hd__nor2_1 U20977 ( .A(n13919), .B(n13918), .Y(n13920) );
  sky130_fd_sc_hd__inv_2 U20978 ( .A(n26711), .Y(n26577) );
  sky130_fd_sc_hd__nand2_1 U20979 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[166]), .Y(n13925) );
  sky130_fd_sc_hd__nand2_1 U20980 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[230]), .Y(n13924) );
  sky130_fd_sc_hd__nand2_1 U20981 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[486]), .Y(n13923) );
  sky130_fd_sc_hd__nand2_1 U20982 ( .A(n15983), .B(
        j202_soc_core_j22_cpu_rf_gpr[422]), .Y(n13922) );
  sky130_fd_sc_hd__nand4_1 U20983 ( .A(n13925), .B(n13924), .C(n13923), .D(
        n13922), .Y(n13931) );
  sky130_fd_sc_hd__nand2_1 U20984 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[6]), .Y(n13929) );
  sky130_fd_sc_hd__nand2_1 U20985 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[38]), .Y(n13928) );
  sky130_fd_sc_hd__nand2_1 U20986 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[102]), .Y(n13927) );
  sky130_fd_sc_hd__nand2_1 U20987 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[390]), .Y(n13926) );
  sky130_fd_sc_hd__nand4_1 U20988 ( .A(n13929), .B(n13928), .C(n13927), .D(
        n13926), .Y(n13930) );
  sky130_fd_sc_hd__nor2_1 U20989 ( .A(n13931), .B(n13930), .Y(n13939) );
  sky130_fd_sc_hd__a22oi_1 U20990 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[294]), .B1(n23502), .B2(
        j202_soc_core_j22_cpu_rf_gpr[454]), .Y(n13938) );
  sky130_fd_sc_hd__inv_2 U20991 ( .A(n29568), .Y(n16469) );
  sky130_fd_sc_hd__a22oi_1 U20992 ( .A1(n16470), .A2(
        j202_soc_core_j22_cpu_rf_gpr[198]), .B1(n16469), .B2(
        j202_soc_core_j22_cpu_rf_gpr[70]), .Y(n13937) );
  sky130_fd_sc_hd__nand2_1 U20993 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[262]), .Y(n13935) );
  sky130_fd_sc_hd__nand2_1 U20994 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[134]), .Y(n13934) );
  sky130_fd_sc_hd__nand2_1 U20995 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[358]), .Y(n13933) );
  sky130_fd_sc_hd__nand2_1 U20996 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[326]), .Y(n13932) );
  sky130_fd_sc_hd__and4_1 U20997 ( .A(n13935), .B(n13934), .C(n13933), .D(
        n13932), .X(n13936) );
  sky130_fd_sc_hd__nand4_1 U20998 ( .A(n13939), .B(n13938), .C(n13937), .D(
        n13936), .Y(n21563) );
  sky130_fd_sc_hd__nand2_1 U20999 ( .A(n21563), .B(n16513), .Y(n13949) );
  sky130_fd_sc_hd__o22ai_1 U21000 ( .A1(n13940), .A2(n16007), .B1(n16008), 
        .B2(n21555), .Y(n13942) );
  sky130_fd_sc_hd__a22o_1 U21001 ( .A1(n29563), .A2(
        j202_soc_core_j22_cpu_rf_gpr[486]), .B1(n29567), .B2(
        j202_soc_core_j22_cpu_rf_vbr[6]), .X(n13941) );
  sky130_fd_sc_hd__nor2_1 U21002 ( .A(n13942), .B(n13941), .Y(n13948) );
  sky130_fd_sc_hd__a2bb2oi_1 U21003 ( .B1(n13701), .B2(n10983), .A1_N(n21553), 
        .A2_N(n14539), .Y(n13943) );
  sky130_fd_sc_hd__o21ai_1 U21004 ( .A1(n21554), .A2(n11095), .B1(n13943), .Y(
        n13946) );
  sky130_fd_sc_hd__o22ai_1 U21005 ( .A1(n13944), .A2(n16014), .B1(n16010), 
        .B2(n21552), .Y(n13945) );
  sky130_fd_sc_hd__nor2_1 U21006 ( .A(n13946), .B(n13945), .Y(n13947) );
  sky130_fd_sc_hd__o22ai_1 U21007 ( .A1(n16492), .A2(n26577), .B1(n27007), 
        .B2(n13793), .Y(n14125) );
  sky130_fd_sc_hd__nand2_1 U21008 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[165]), .Y(n13953) );
  sky130_fd_sc_hd__nand2_1 U21009 ( .A(n15982), .B(
        j202_soc_core_j22_cpu_rf_gpr[229]), .Y(n13952) );
  sky130_fd_sc_hd__nand2_1 U21010 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[485]), .Y(n13951) );
  sky130_fd_sc_hd__nand2_1 U21011 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[421]), .Y(n13950) );
  sky130_fd_sc_hd__nand4_1 U21012 ( .A(n13953), .B(n13952), .C(n13951), .D(
        n13950), .Y(n13959) );
  sky130_fd_sc_hd__nand2_1 U21013 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[5]), .Y(n13957) );
  sky130_fd_sc_hd__nand2_1 U21014 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[37]), .Y(n13956) );
  sky130_fd_sc_hd__nand2_1 U21015 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[101]), .Y(n13955) );
  sky130_fd_sc_hd__nand2_1 U21016 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[389]), .Y(n13954) );
  sky130_fd_sc_hd__nand4_1 U21017 ( .A(n13957), .B(n13956), .C(n13955), .D(
        n13954), .Y(n13958) );
  sky130_fd_sc_hd__nor2_1 U21018 ( .A(n13959), .B(n13958), .Y(n13966) );
  sky130_fd_sc_hd__a22oi_1 U21019 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[293]), .B1(n23502), .B2(
        j202_soc_core_j22_cpu_rf_gpr[453]), .Y(n13965) );
  sky130_fd_sc_hd__a22oi_1 U21020 ( .A1(n16470), .A2(
        j202_soc_core_j22_cpu_rf_gpr[197]), .B1(n23089), .B2(
        j202_soc_core_j22_cpu_rf_gpr[69]), .Y(n13964) );
  sky130_fd_sc_hd__nand2_1 U21021 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[261]), .Y(n13963) );
  sky130_fd_sc_hd__nand2_1 U21022 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[133]), .Y(n13962) );
  sky130_fd_sc_hd__nand2_1 U21023 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[357]), .Y(n13961) );
  sky130_fd_sc_hd__nand2_1 U21024 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[325]), .Y(n13960) );
  sky130_fd_sc_hd__nand4_1 U21025 ( .A(n13966), .B(n13965), .C(n13964), .D(
        n12222), .Y(n21854) );
  sky130_fd_sc_hd__nand2_1 U21026 ( .A(n16519), .B(j202_soc_core_j22_cpu_pc[5]), .Y(n13970) );
  sky130_fd_sc_hd__nand2_1 U21027 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[5]), .Y(n13969) );
  sky130_fd_sc_hd__nand2_1 U21028 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[485]), .Y(n13968) );
  sky130_fd_sc_hd__nand2_1 U21029 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[5]), .Y(n13967) );
  sky130_fd_sc_hd__a2bb2oi_1 U21030 ( .B1(n13701), .B2(n10977), .A1_N(n21856), 
        .A2_N(n14539), .Y(n13971) );
  sky130_fd_sc_hd__o21ai_1 U21031 ( .A1(n21857), .A2(n11095), .B1(n13971), .Y(
        n13973) );
  sky130_fd_sc_hd__o22ai_1 U21032 ( .A1(n21861), .A2(n16014), .B1(n16010), 
        .B2(n21855), .Y(n13972) );
  sky130_fd_sc_hd__nor2_1 U21033 ( .A(n13973), .B(n13972), .Y(n13974) );
  sky130_fd_sc_hd__mux2i_1 U21034 ( .A0(n14742), .A1(n16320), .S(n27415), .Y(
        n14126) );
  sky130_fd_sc_hd__nor2_1 U21035 ( .A(n14125), .B(n14126), .Y(n21756) );
  sky130_fd_sc_hd__nor2_1 U21036 ( .A(n21526), .B(n21756), .Y(n14130) );
  sky130_fd_sc_hd__nand2_1 U21037 ( .A(n21530), .B(n14130), .Y(n14132) );
  sky130_fd_sc_hd__nand2_1 U21038 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[161]), .Y(n13979) );
  sky130_fd_sc_hd__nand2_1 U21039 ( .A(n15982), .B(
        j202_soc_core_j22_cpu_rf_gpr[225]), .Y(n13978) );
  sky130_fd_sc_hd__nand2_1 U21040 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[481]), .Y(n13977) );
  sky130_fd_sc_hd__nand2_1 U21041 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[417]), .Y(n13976) );
  sky130_fd_sc_hd__nand4_1 U21042 ( .A(n13979), .B(n13978), .C(n13977), .D(
        n13976), .Y(n13985) );
  sky130_fd_sc_hd__nand2_1 U21043 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[1]), .Y(n13983) );
  sky130_fd_sc_hd__nand2_1 U21044 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[33]), .Y(n13982) );
  sky130_fd_sc_hd__nand2_1 U21045 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[97]), .Y(n13981) );
  sky130_fd_sc_hd__nand2_1 U21046 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[385]), .Y(n13980) );
  sky130_fd_sc_hd__nand4_1 U21047 ( .A(n13983), .B(n13982), .C(n13981), .D(
        n13980), .Y(n13984) );
  sky130_fd_sc_hd__nor2_1 U21048 ( .A(n13985), .B(n13984), .Y(n13994) );
  sky130_fd_sc_hd__a22oi_1 U21049 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[289]), .B1(n14414), .B2(
        j202_soc_core_j22_cpu_rf_gpr[449]), .Y(n13993) );
  sky130_fd_sc_hd__a22oi_1 U21050 ( .A1(n16470), .A2(
        j202_soc_core_j22_cpu_rf_gpr[193]), .B1(n23089), .B2(
        j202_soc_core_j22_cpu_rf_gpr[65]), .Y(n13992) );
  sky130_fd_sc_hd__nand2_1 U21051 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[257]), .Y(n13990) );
  sky130_fd_sc_hd__nand2_1 U21052 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[129]), .Y(n13989) );
  sky130_fd_sc_hd__nand2_1 U21053 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[353]), .Y(n13988) );
  sky130_fd_sc_hd__nand2_1 U21054 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[321]), .Y(n13987) );
  sky130_fd_sc_hd__and4_1 U21055 ( .A(n13990), .B(n13989), .C(n13988), .D(
        n13987), .X(n13991) );
  sky130_fd_sc_hd__nand4_1 U21056 ( .A(n13994), .B(n13993), .C(n13992), .D(
        n13991), .Y(n22779) );
  sky130_fd_sc_hd__nand2_1 U21057 ( .A(n22779), .B(n16513), .Y(n14005) );
  sky130_fd_sc_hd__nand2_1 U21058 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[1]), .Y(n13998) );
  sky130_fd_sc_hd__nand2_1 U21059 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[1]), .Y(n13997) );
  sky130_fd_sc_hd__nand2_1 U21060 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[481]), .Y(n13996) );
  sky130_fd_sc_hd__nand2_1 U21061 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[1]), .Y(n13995) );
  sky130_fd_sc_hd__and4_1 U21062 ( .A(n13998), .B(n13997), .C(n13996), .D(
        n13995), .X(n14004) );
  sky130_fd_sc_hd__a2bb2oi_1 U21063 ( .B1(n13701), .B2(n10922), .A1_N(n24273), 
        .A2_N(n14539), .Y(n13999) );
  sky130_fd_sc_hd__o21ai_1 U21064 ( .A1(n22781), .A2(n11095), .B1(n13999), .Y(
        n14002) );
  sky130_fd_sc_hd__o22ai_1 U21065 ( .A1(n14000), .A2(n16014), .B1(n16008), 
        .B2(n22782), .Y(n14001) );
  sky130_fd_sc_hd__nor2_1 U21066 ( .A(n14002), .B(n14001), .Y(n14003) );
  sky130_fd_sc_hd__o21ai_1 U21067 ( .A1(n14008), .A2(n27443), .B1(n14007), .Y(
        n14060) );
  sky130_fd_sc_hd__nand2_1 U21068 ( .A(n26750), .B(n12382), .Y(n19413) );
  sky130_fd_sc_hd__nor2_1 U21069 ( .A(n23928), .B(n19413), .Y(n14010) );
  sky130_fd_sc_hd__a211oi_1 U21070 ( .A1(n14011), .A2(n23928), .B1(n14010), 
        .C1(n14009), .Y(n14012) );
  sky130_fd_sc_hd__nand2_1 U21071 ( .A(n14060), .B(n14012), .Y(n21923) );
  sky130_fd_sc_hd__nand2_1 U21072 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[416]), .Y(n14016) );
  sky130_fd_sc_hd__nand2_1 U21073 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[224]), .Y(n14015) );
  sky130_fd_sc_hd__nand2_1 U21074 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[288]), .Y(n14014) );
  sky130_fd_sc_hd__nand2_1 U21075 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_rf_gpr[192]), .Y(n14013) );
  sky130_fd_sc_hd__and4_1 U21076 ( .A(n14016), .B(n14015), .C(n14014), .D(
        n14013), .X(n14034) );
  sky130_fd_sc_hd__nand2_1 U21077 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[480]), .Y(n14020) );
  sky130_fd_sc_hd__a2bb2oi_1 U21078 ( .B1(j202_soc_core_j22_cpu_rf_tmp[0]), 
        .B2(n13774), .A1_N(n14466), .A2_N(n10980), .Y(n14019) );
  sky130_fd_sc_hd__nand2_1 U21079 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[160]), .Y(n14018) );
  sky130_fd_sc_hd__nand2_1 U21080 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[320]), .Y(n14017) );
  sky130_fd_sc_hd__nand4_1 U21081 ( .A(n14020), .B(n14019), .C(n14018), .D(
        n14017), .Y(n14021) );
  sky130_fd_sc_hd__nand2_1 U21082 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[352]), .Y(n14025) );
  sky130_fd_sc_hd__nand2_1 U21083 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[448]), .Y(n14024) );
  sky130_fd_sc_hd__nand2_1 U21084 ( .A(n11154), .B(
        j202_soc_core_j22_cpu_rf_gpr[256]), .Y(n14023) );
  sky130_fd_sc_hd__nand2_1 U21085 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[384]), .Y(n14022) );
  sky130_fd_sc_hd__nand4_1 U21086 ( .A(n14025), .B(n14024), .C(n14023), .D(
        n14022), .Y(n14031) );
  sky130_fd_sc_hd__nand2_1 U21087 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[128]), .Y(n14029) );
  sky130_fd_sc_hd__nand2_1 U21088 ( .A(n11116), .B(
        j202_soc_core_j22_cpu_rf_gpr[96]), .Y(n14028) );
  sky130_fd_sc_hd__nand2_1 U21089 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[32]), .Y(n14027) );
  sky130_fd_sc_hd__nand2_1 U21090 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[64]), .Y(n14026) );
  sky130_fd_sc_hd__nand4_1 U21091 ( .A(n14029), .B(n14028), .C(n14027), .D(
        n14026), .Y(n14030) );
  sky130_fd_sc_hd__inv_2 U21092 ( .A(n26723), .Y(n25789) );
  sky130_fd_sc_hd__o22ai_1 U21093 ( .A1(n13793), .A2(n23928), .B1(n16492), 
        .B2(n25789), .Y(n14061) );
  sky130_fd_sc_hd__nand2_1 U21094 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[160]), .Y(n14038) );
  sky130_fd_sc_hd__nand2_1 U21095 ( .A(n15982), .B(
        j202_soc_core_j22_cpu_rf_gpr[224]), .Y(n14037) );
  sky130_fd_sc_hd__nand2_1 U21096 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[480]), .Y(n14036) );
  sky130_fd_sc_hd__nand2_1 U21097 ( .A(n15983), .B(
        j202_soc_core_j22_cpu_rf_gpr[416]), .Y(n14035) );
  sky130_fd_sc_hd__nand4_1 U21098 ( .A(n14038), .B(n14037), .C(n14036), .D(
        n14035), .Y(n14044) );
  sky130_fd_sc_hd__nand2_1 U21099 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[0]), .Y(n14042) );
  sky130_fd_sc_hd__nand2_1 U21100 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[32]), .Y(n14041) );
  sky130_fd_sc_hd__nand2_1 U21101 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[96]), .Y(n14040) );
  sky130_fd_sc_hd__nand2_1 U21102 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[384]), .Y(n14039) );
  sky130_fd_sc_hd__nand4_1 U21103 ( .A(n14042), .B(n14041), .C(n14040), .D(
        n14039), .Y(n14043) );
  sky130_fd_sc_hd__nor2_1 U21104 ( .A(n14044), .B(n14043), .Y(n14051) );
  sky130_fd_sc_hd__a22oi_1 U21105 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[288]), .B1(n14414), .B2(
        j202_soc_core_j22_cpu_rf_gpr[448]), .Y(n14050) );
  sky130_fd_sc_hd__a22oi_1 U21106 ( .A1(n16470), .A2(
        j202_soc_core_j22_cpu_rf_gpr[192]), .B1(n23089), .B2(
        j202_soc_core_j22_cpu_rf_gpr[64]), .Y(n14049) );
  sky130_fd_sc_hd__nand2_1 U21107 ( .A(n23130), .B(
        j202_soc_core_j22_cpu_rf_gpr[256]), .Y(n14048) );
  sky130_fd_sc_hd__nand2_1 U21108 ( .A(n16471), .B(
        j202_soc_core_j22_cpu_rf_gpr[128]), .Y(n14047) );
  sky130_fd_sc_hd__nand2_1 U21109 ( .A(n13686), .B(
        j202_soc_core_j22_cpu_rf_gpr[352]), .Y(n14046) );
  sky130_fd_sc_hd__nand2_1 U21110 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[320]), .Y(n14045) );
  sky130_fd_sc_hd__nand4_1 U21111 ( .A(n14051), .B(n14050), .C(n14049), .D(
        n12223), .Y(n21960) );
  sky130_fd_sc_hd__o22ai_1 U21112 ( .A1(n21954), .A2(n16007), .B1(n16008), 
        .B2(n23720), .Y(n14053) );
  sky130_fd_sc_hd__a22o_1 U21113 ( .A1(n29563), .A2(
        j202_soc_core_j22_cpu_rf_gpr[480]), .B1(n29567), .B2(
        j202_soc_core_j22_cpu_rf_vbr[0]), .X(n14052) );
  sky130_fd_sc_hd__nor2_1 U21114 ( .A(n14053), .B(n14052), .Y(n14058) );
  sky130_fd_sc_hd__a2bb2oi_1 U21115 ( .B1(n13701), .B2(n10979), .A1_N(n23928), 
        .A2_N(n14539), .Y(n14054) );
  sky130_fd_sc_hd__o22ai_1 U21117 ( .A1(n21955), .A2(n16014), .B1(n16010), 
        .B2(n21950), .Y(n14055) );
  sky130_fd_sc_hd__nor2_1 U21118 ( .A(n14056), .B(n14055), .Y(n14057) );
  sky130_fd_sc_hd__nor2_1 U21119 ( .A(n14061), .B(n14062), .Y(n21919) );
  sky130_fd_sc_hd__nand2_1 U21120 ( .A(n14062), .B(n14061), .Y(n21920) );
  sky130_fd_sc_hd__nand2_1 U21121 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[225]), .Y(n14067) );
  sky130_fd_sc_hd__nand2_1 U21122 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[193]), .Y(n14066) );
  sky130_fd_sc_hd__nand2_1 U21123 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[417]), .Y(n14065) );
  sky130_fd_sc_hd__nand2_1 U21124 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[289]), .Y(n14064) );
  sky130_fd_sc_hd__and4_1 U21125 ( .A(n14067), .B(n14066), .C(n14065), .D(
        n14064), .X(n14085) );
  sky130_fd_sc_hd__nand2_1 U21126 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[481]), .Y(n14071) );
  sky130_fd_sc_hd__a2bb2oi_1 U21127 ( .B1(j202_soc_core_j22_cpu_rf_tmp[1]), 
        .B2(n13774), .A1_N(n14466), .A2_N(n10923), .Y(n14070) );
  sky130_fd_sc_hd__nand2_1 U21128 ( .A(n15128), .B(
        j202_soc_core_j22_cpu_rf_gpr[161]), .Y(n14069) );
  sky130_fd_sc_hd__nand2_1 U21129 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[321]), .Y(n14068) );
  sky130_fd_sc_hd__nand4_1 U21130 ( .A(n14071), .B(n14070), .C(n14069), .D(
        n14068), .Y(n14072) );
  sky130_fd_sc_hd__a21oi_1 U21131 ( .A1(j202_soc_core_j22_cpu_rf_gpr[1]), .A2(
        n16285), .B1(n14072), .Y(n14084) );
  sky130_fd_sc_hd__nand2_1 U21132 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[449]), .Y(n14076) );
  sky130_fd_sc_hd__nand2_1 U21133 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[353]), .Y(n14075) );
  sky130_fd_sc_hd__nand2_1 U21134 ( .A(n11154), .B(
        j202_soc_core_j22_cpu_rf_gpr[257]), .Y(n14074) );
  sky130_fd_sc_hd__nand2_1 U21135 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[385]), .Y(n14073) );
  sky130_fd_sc_hd__nand4_1 U21136 ( .A(n14076), .B(n14075), .C(n14074), .D(
        n14073), .Y(n14082) );
  sky130_fd_sc_hd__nand2_1 U21137 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[129]), .Y(n14080) );
  sky130_fd_sc_hd__nand2_1 U21138 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[97]), .Y(n14079) );
  sky130_fd_sc_hd__nand2_1 U21139 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[33]), .Y(n14078) );
  sky130_fd_sc_hd__nand2_1 U21140 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[65]), .Y(n14077) );
  sky130_fd_sc_hd__nand4_1 U21141 ( .A(n14080), .B(n14079), .C(n14078), .D(
        n14077), .Y(n14081) );
  sky130_fd_sc_hd__nor2_1 U21142 ( .A(n14082), .B(n14081), .Y(n14083) );
  sky130_fd_sc_hd__inv_2 U21143 ( .A(n26603), .Y(n25743) );
  sky130_fd_sc_hd__o22ai_1 U21144 ( .A1(n16492), .A2(n25743), .B1(n25789), 
        .B2(n13793), .Y(n14115) );
  sky130_fd_sc_hd__mux2i_1 U21145 ( .A0(n14742), .A1(n16320), .S(n27443), .Y(
        n14116) );
  sky130_fd_sc_hd__nor2_1 U21146 ( .A(n14115), .B(n14116), .Y(n20275) );
  sky130_fd_sc_hd__o22ai_1 U21147 ( .A1(n13793), .A2(n25743), .B1(n25229), 
        .B2(n16492), .Y(n14117) );
  sky130_fd_sc_hd__nand2_1 U21148 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[162]), .Y(n14089) );
  sky130_fd_sc_hd__nand2_1 U21149 ( .A(n15982), .B(
        j202_soc_core_j22_cpu_rf_gpr[226]), .Y(n14088) );
  sky130_fd_sc_hd__nand2_1 U21150 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[482]), .Y(n14087) );
  sky130_fd_sc_hd__nand2_1 U21151 ( .A(n15983), .B(
        j202_soc_core_j22_cpu_rf_gpr[418]), .Y(n14086) );
  sky130_fd_sc_hd__nand4_1 U21152 ( .A(n14089), .B(n14088), .C(n14087), .D(
        n14086), .Y(n14095) );
  sky130_fd_sc_hd__nand2_1 U21153 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[2]), .Y(n14093) );
  sky130_fd_sc_hd__nand2_1 U21154 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[34]), .Y(n14092) );
  sky130_fd_sc_hd__nand2_1 U21155 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[98]), .Y(n14091) );
  sky130_fd_sc_hd__nand2_1 U21156 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[386]), .Y(n14090) );
  sky130_fd_sc_hd__nand4_1 U21157 ( .A(n14093), .B(n14092), .C(n14091), .D(
        n14090), .Y(n14094) );
  sky130_fd_sc_hd__nor2_1 U21158 ( .A(n14095), .B(n14094), .Y(n14106) );
  sky130_fd_sc_hd__nand2_1 U21159 ( .A(n16469), .B(
        j202_soc_core_j22_cpu_rf_gpr[66]), .Y(n14099) );
  sky130_fd_sc_hd__nand2_1 U21160 ( .A(n16470), .B(
        j202_soc_core_j22_cpu_rf_gpr[194]), .Y(n14098) );
  sky130_fd_sc_hd__nand2_1 U21161 ( .A(n11160), .B(
        j202_soc_core_j22_cpu_rf_gpr[290]), .Y(n14097) );
  sky130_fd_sc_hd__nand2_1 U21162 ( .A(n14414), .B(
        j202_soc_core_j22_cpu_rf_gpr[450]), .Y(n14096) );
  sky130_fd_sc_hd__and4_1 U21163 ( .A(n14099), .B(n14098), .C(n14097), .D(
        n14096), .X(n14105) );
  sky130_fd_sc_hd__nand2_1 U21164 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[258]), .Y(n14103) );
  sky130_fd_sc_hd__nand2_1 U21165 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[130]), .Y(n14102) );
  sky130_fd_sc_hd__nand2_1 U21166 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[354]), .Y(n14101) );
  sky130_fd_sc_hd__nand2_1 U21167 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[322]), .Y(n14100) );
  sky130_fd_sc_hd__and4_1 U21168 ( .A(n14103), .B(n14102), .C(n14101), .D(
        n14100), .X(n14104) );
  sky130_fd_sc_hd__nand3_1 U21169 ( .A(n14106), .B(n14105), .C(n14104), .Y(
        n19210) );
  sky130_fd_sc_hd__a22oi_1 U21170 ( .A1(n16514), .A2(
        j202_soc_core_j22_cpu_rf_tmp[2]), .B1(n29567), .B2(
        j202_soc_core_j22_cpu_rf_vbr[2]), .Y(n14112) );
  sky130_fd_sc_hd__a22oi_1 U21171 ( .A1(n10929), .A2(n13701), .B1(n29563), 
        .B2(j202_soc_core_j22_cpu_rf_gpr[482]), .Y(n14111) );
  sky130_fd_sc_hd__o22a_1 U21172 ( .A1(n14107), .A2(n16014), .B1(n19203), .B2(
        n16008), .X(n14110) );
  sky130_fd_sc_hd__o22a_1 U21173 ( .A1(n19202), .A2(n16010), .B1(n14108), .B2(
        n11095), .X(n14109) );
  sky130_fd_sc_hd__nand4_1 U21174 ( .A(n14112), .B(n14111), .C(n14110), .D(
        n14109), .Y(n14113) );
  sky130_fd_sc_hd__a21oi_1 U21175 ( .A1(n19210), .A2(n16513), .B1(n14113), .Y(
        n25237) );
  sky130_fd_sc_hd__nand2_1 U21176 ( .A(n25237), .B(n16322), .Y(n14114) );
  sky130_fd_sc_hd__o21ai_1 U21177 ( .A1(n16320), .A2(n25237), .B1(n14114), .Y(
        n14118) );
  sky130_fd_sc_hd__nor2_1 U21178 ( .A(n14117), .B(n14118), .Y(n17259) );
  sky130_fd_sc_hd__nor2_1 U21179 ( .A(n20275), .B(n17259), .Y(n14120) );
  sky130_fd_sc_hd__nand2_1 U21180 ( .A(n14116), .B(n14115), .Y(n20276) );
  sky130_fd_sc_hd__nand2_1 U21181 ( .A(n14118), .B(n14117), .Y(n17260) );
  sky130_fd_sc_hd__o21ai_1 U21182 ( .A1(n20276), .A2(n17259), .B1(n17260), .Y(
        n14119) );
  sky130_fd_sc_hd__nand2_1 U21183 ( .A(n14122), .B(n14121), .Y(n20286) );
  sky130_fd_sc_hd__nand2_1 U21184 ( .A(n14124), .B(n14123), .Y(n19419) );
  sky130_fd_sc_hd__o21ai_1 U21185 ( .A1(n20286), .A2(n19418), .B1(n19419), .Y(
        n21529) );
  sky130_fd_sc_hd__nand2_1 U21186 ( .A(n14126), .B(n14125), .Y(n21757) );
  sky130_fd_sc_hd__nand2_1 U21187 ( .A(n14128), .B(n14127), .Y(n21527) );
  sky130_fd_sc_hd__o21ai_1 U21188 ( .A1(n21757), .A2(n21526), .B1(n21527), .Y(
        n14129) );
  sky130_fd_sc_hd__a21oi_1 U21189 ( .A1(n14130), .A2(n21529), .B1(n14129), .Y(
        n14131) );
  sky130_fd_sc_hd__nand2_1 U21190 ( .A(n11114), .B(
        j202_soc_core_j22_cpu_rf_gpr[397]), .Y(n14136) );
  sky130_fd_sc_hd__nand2_1 U21191 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[461]), .Y(n14135) );
  sky130_fd_sc_hd__nand2_1 U21192 ( .A(n16324), .B(
        j202_soc_core_j22_cpu_rf_gpr[269]), .Y(n14134) );
  sky130_fd_sc_hd__nand2_1 U21193 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[141]), .Y(n14133) );
  sky130_fd_sc_hd__nand4_1 U21194 ( .A(n14136), .B(n14135), .C(n14134), .D(
        n14133), .Y(n14142) );
  sky130_fd_sc_hd__a21oi_1 U21195 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[13]), .B1(n16436), .Y(n14140) );
  sky130_fd_sc_hd__nand2_1 U21196 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[109]), .Y(n14139) );
  sky130_fd_sc_hd__nand2_1 U21197 ( .A(n11152), .B(
        j202_soc_core_j22_cpu_rf_gpr[45]), .Y(n14138) );
  sky130_fd_sc_hd__nand2_1 U21198 ( .A(n11155), .B(
        j202_soc_core_j22_cpu_rf_gpr[77]), .Y(n14137) );
  sky130_fd_sc_hd__nand4_1 U21199 ( .A(n14140), .B(n14139), .C(n14138), .D(
        n14137), .Y(n14141) );
  sky130_fd_sc_hd__nor2_1 U21200 ( .A(n14142), .B(n14141), .Y(n14154) );
  sky130_fd_sc_hd__nand2_1 U21201 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[429]), .Y(n14147) );
  sky130_fd_sc_hd__nand2_1 U21202 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[237]), .Y(n14146) );
  sky130_fd_sc_hd__nand2_1 U21203 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[205]), .Y(n14145) );
  sky130_fd_sc_hd__nand2_1 U21204 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[301]), .Y(n14144) );
  sky130_fd_sc_hd__nand2_1 U21205 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[493]), .Y(n14151) );
  sky130_fd_sc_hd__nand2_1 U21206 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[173]), .Y(n14150) );
  sky130_fd_sc_hd__nand2_1 U21207 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[333]), .Y(n14149) );
  sky130_fd_sc_hd__nand2_1 U21208 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[365]), .Y(n14148) );
  sky130_fd_sc_hd__nand4_1 U21209 ( .A(n14151), .B(n14150), .C(n14149), .D(
        n14148), .Y(n14152) );
  sky130_fd_sc_hd__a21oi_1 U21210 ( .A1(j202_soc_core_j22_cpu_rf_gpr[13]), 
        .A2(n16285), .B1(n14152), .Y(n14153) );
  sky130_fd_sc_hd__a22oi_1 U21211 ( .A1(n11114), .A2(
        j202_soc_core_j22_cpu_rf_gpr[398]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_rf_gpr[462]), .Y(n14160) );
  sky130_fd_sc_hd__a22oi_1 U21212 ( .A1(n11154), .A2(
        j202_soc_core_j22_cpu_rf_gpr[270]), .B1(n11113), .B2(
        j202_soc_core_j22_cpu_rf_gpr[142]), .Y(n14159) );
  sky130_fd_sc_hd__nor2_1 U21213 ( .A(n13638), .B(n14155), .Y(n14758) );
  sky130_fd_sc_hd__o21ai_1 U21214 ( .A1(n14156), .A2(n14758), .B1(
        j202_soc_core_j22_cpu_rf_gpr[14]), .Y(n14158) );
  sky130_fd_sc_hd__a22oi_1 U21215 ( .A1(n11155), .A2(
        j202_soc_core_j22_cpu_rf_gpr[78]), .B1(n11116), .B2(
        j202_soc_core_j22_cpu_rf_gpr[110]), .Y(n14157) );
  sky130_fd_sc_hd__nand2_1 U21216 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[238]), .Y(n14163) );
  sky130_fd_sc_hd__nand2_1 U21217 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[302]), .Y(n14162) );
  sky130_fd_sc_hd__nand2_1 U21218 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[430]), .Y(n14161) );
  sky130_fd_sc_hd__nand3_1 U21219 ( .A(n14163), .B(n14162), .C(n14161), .Y(
        n14167) );
  sky130_fd_sc_hd__nand2_1 U21220 ( .A(n11152), .B(
        j202_soc_core_j22_cpu_rf_gpr[46]), .Y(n14165) );
  sky130_fd_sc_hd__nand2_1 U21221 ( .A(n13774), .B(
        j202_soc_core_j22_cpu_rf_tmp[14]), .Y(n14164) );
  sky130_fd_sc_hd__nand3_1 U21222 ( .A(n14755), .B(n14165), .C(n14164), .Y(
        n14166) );
  sky130_fd_sc_hd__nor2_1 U21223 ( .A(n14167), .B(n14166), .Y(n14174) );
  sky130_fd_sc_hd__nand2_1 U21224 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[494]), .Y(n14171) );
  sky130_fd_sc_hd__nand2_1 U21225 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[174]), .Y(n14170) );
  sky130_fd_sc_hd__nand2_1 U21226 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[334]), .Y(n14169) );
  sky130_fd_sc_hd__nand2_1 U21227 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[366]), .Y(n14168) );
  sky130_fd_sc_hd__nand4_1 U21228 ( .A(n14171), .B(n14170), .C(n14169), .D(
        n14168), .Y(n14172) );
  sky130_fd_sc_hd__a21oi_1 U21229 ( .A1(n16248), .A2(
        j202_soc_core_j22_cpu_rf_gpr[206]), .B1(n14172), .Y(n14173) );
  sky130_fd_sc_hd__inv_2 U21230 ( .A(n26725), .Y(n26565) );
  sky130_fd_sc_hd__o22ai_1 U21231 ( .A1(n13793), .A2(n26708), .B1(n26565), 
        .B2(n16492), .Y(n14564) );
  sky130_fd_sc_hd__nand2_1 U21232 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[174]), .Y(n14178) );
  sky130_fd_sc_hd__nand2_1 U21233 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[238]), .Y(n14177) );
  sky130_fd_sc_hd__nand2_1 U21234 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[494]), .Y(n14176) );
  sky130_fd_sc_hd__nand2_1 U21235 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[430]), .Y(n14175) );
  sky130_fd_sc_hd__nand4_1 U21236 ( .A(n14178), .B(n14177), .C(n14176), .D(
        n14175), .Y(n14184) );
  sky130_fd_sc_hd__nand2_1 U21237 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[14]), .Y(n14182) );
  sky130_fd_sc_hd__nand2_1 U21238 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[46]), .Y(n14181) );
  sky130_fd_sc_hd__nand2_1 U21239 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[110]), .Y(n14180) );
  sky130_fd_sc_hd__nand2_1 U21240 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[398]), .Y(n14179) );
  sky130_fd_sc_hd__nand4_1 U21241 ( .A(n14182), .B(n14181), .C(n14180), .D(
        n14179), .Y(n14183) );
  sky130_fd_sc_hd__nor2_1 U21242 ( .A(n14184), .B(n14183), .Y(n14192) );
  sky130_fd_sc_hd__a22oi_1 U21243 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[302]), .B1(n23502), .B2(
        j202_soc_core_j22_cpu_rf_gpr[462]), .Y(n14191) );
  sky130_fd_sc_hd__a22oi_1 U21244 ( .A1(n23515), .A2(
        j202_soc_core_j22_cpu_rf_gpr[206]), .B1(n23089), .B2(
        j202_soc_core_j22_cpu_rf_gpr[78]), .Y(n14190) );
  sky130_fd_sc_hd__nand2_1 U21245 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[270]), .Y(n14188) );
  sky130_fd_sc_hd__nand2_1 U21246 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[142]), .Y(n14187) );
  sky130_fd_sc_hd__nand2_1 U21247 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[366]), .Y(n14186) );
  sky130_fd_sc_hd__nand2_1 U21248 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[334]), .Y(n14185) );
  sky130_fd_sc_hd__and4_1 U21249 ( .A(n14188), .B(n14187), .C(n14186), .D(
        n14185), .X(n14189) );
  sky130_fd_sc_hd__nand4_1 U21250 ( .A(n14192), .B(n14191), .C(n14190), .D(
        n14189), .Y(n21573) );
  sky130_fd_sc_hd__nand2_1 U21251 ( .A(n21573), .B(n16513), .Y(n14202) );
  sky130_fd_sc_hd__nand2_1 U21252 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[14]), .Y(n14195) );
  sky130_fd_sc_hd__nand2_1 U21253 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[14]), .Y(n14194) );
  sky130_fd_sc_hd__nand2_1 U21254 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[494]), .Y(n14193) );
  sky130_fd_sc_hd__and4_1 U21255 ( .A(n14195), .B(n14194), .C(n16516), .D(
        n14193), .X(n14201) );
  sky130_fd_sc_hd__nand2_1 U21256 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[14]), .Y(n14199) );
  sky130_fd_sc_hd__nand2_1 U21257 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[14]), .Y(n14198) );
  sky130_fd_sc_hd__nand2_1 U21258 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[14]), .Y(n14197) );
  sky130_fd_sc_hd__nand2_1 U21259 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[14]), .Y(n14196) );
  sky130_fd_sc_hd__and4_1 U21260 ( .A(n14199), .B(n14198), .C(n14197), .D(
        n14196), .X(n14200) );
  sky130_fd_sc_hd__nand3_1 U21261 ( .A(n14202), .B(n14201), .C(n14200), .Y(
        n27361) );
  sky130_fd_sc_hd__nand2_1 U21262 ( .A(n27361), .B(n16529), .Y(n14203) );
  sky130_fd_sc_hd__nor2_1 U21264 ( .A(n14564), .B(n14565), .Y(n21332) );
  sky130_fd_sc_hd__nand2_1 U21265 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[396]), .Y(n14208) );
  sky130_fd_sc_hd__nand2_1 U21266 ( .A(n16323), .B(
        j202_soc_core_j22_cpu_rf_gpr[460]), .Y(n14207) );
  sky130_fd_sc_hd__nand2_1 U21267 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[76]), .Y(n14206) );
  sky130_fd_sc_hd__nand2_1 U21268 ( .A(n11154), .B(
        j202_soc_core_j22_cpu_rf_gpr[268]), .Y(n14205) );
  sky130_fd_sc_hd__nand4_1 U21269 ( .A(n14208), .B(n14207), .C(n14206), .D(
        n14205), .Y(n14214) );
  sky130_fd_sc_hd__a21oi_1 U21270 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[12]), .B1(n16436), .Y(n14212) );
  sky130_fd_sc_hd__nand2_1 U21271 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[140]), .Y(n14211) );
  sky130_fd_sc_hd__nand2_1 U21272 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[108]), .Y(n14210) );
  sky130_fd_sc_hd__nand2_1 U21273 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[44]), .Y(n14209) );
  sky130_fd_sc_hd__nand4_1 U21274 ( .A(n14212), .B(n14211), .C(n14210), .D(
        n14209), .Y(n14213) );
  sky130_fd_sc_hd__nor2_1 U21275 ( .A(n14214), .B(n14213), .Y(n14226) );
  sky130_fd_sc_hd__nand2_1 U21276 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[428]), .Y(n14218) );
  sky130_fd_sc_hd__nand2_1 U21277 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[236]), .Y(n14217) );
  sky130_fd_sc_hd__nand2_1 U21278 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[204]), .Y(n14216) );
  sky130_fd_sc_hd__nand2_1 U21279 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[300]), .Y(n14215) );
  sky130_fd_sc_hd__and4_1 U21280 ( .A(n14218), .B(n14217), .C(n14216), .D(
        n14215), .X(n14225) );
  sky130_fd_sc_hd__nand2_1 U21281 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[492]), .Y(n14222) );
  sky130_fd_sc_hd__nand2_1 U21282 ( .A(n15128), .B(
        j202_soc_core_j22_cpu_rf_gpr[172]), .Y(n14221) );
  sky130_fd_sc_hd__nand2_1 U21283 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[332]), .Y(n14220) );
  sky130_fd_sc_hd__nand2_1 U21284 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[364]), .Y(n14219) );
  sky130_fd_sc_hd__nand4_1 U21285 ( .A(n14222), .B(n14221), .C(n14220), .D(
        n14219), .Y(n14223) );
  sky130_fd_sc_hd__a21oi_1 U21286 ( .A1(j202_soc_core_j22_cpu_rf_gpr[12]), 
        .A2(n16285), .B1(n14223), .Y(n14224) );
  sky130_fd_sc_hd__nand3_1 U21287 ( .A(n14226), .B(n14225), .C(n14224), .Y(
        n26709) );
  sky130_fd_sc_hd__o22ai_1 U21288 ( .A1(n16492), .A2(n26708), .B1(n26426), 
        .B2(n13793), .Y(n14562) );
  sky130_fd_sc_hd__nand2_1 U21289 ( .A(n13794), .B(
        j202_soc_core_j22_cpu_rf_gpr[173]), .Y(n14230) );
  sky130_fd_sc_hd__nand2_1 U21290 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[237]), .Y(n14229) );
  sky130_fd_sc_hd__nand2_1 U21291 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[493]), .Y(n14228) );
  sky130_fd_sc_hd__nand2_1 U21292 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[429]), .Y(n14227) );
  sky130_fd_sc_hd__nand4_1 U21293 ( .A(n14230), .B(n14229), .C(n14228), .D(
        n14227), .Y(n14237) );
  sky130_fd_sc_hd__nand2_1 U21294 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[13]), .Y(n14235) );
  sky130_fd_sc_hd__nand2_1 U21295 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[45]), .Y(n14234) );
  sky130_fd_sc_hd__nand2_1 U21296 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[109]), .Y(n14233) );
  sky130_fd_sc_hd__nand2_1 U21297 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[397]), .Y(n14232) );
  sky130_fd_sc_hd__nand4_1 U21298 ( .A(n14235), .B(n14234), .C(n14233), .D(
        n14232), .Y(n14236) );
  sky130_fd_sc_hd__nor2_1 U21299 ( .A(n14237), .B(n14236), .Y(n14245) );
  sky130_fd_sc_hd__a22oi_1 U21300 ( .A1(n11160), .A2(
        j202_soc_core_j22_cpu_rf_gpr[301]), .B1(n14414), .B2(
        j202_soc_core_j22_cpu_rf_gpr[461]), .Y(n14244) );
  sky130_fd_sc_hd__a22oi_1 U21301 ( .A1(n23515), .A2(
        j202_soc_core_j22_cpu_rf_gpr[205]), .B1(n16469), .B2(
        j202_soc_core_j22_cpu_rf_gpr[77]), .Y(n14243) );
  sky130_fd_sc_hd__nand2_1 U21302 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[269]), .Y(n14241) );
  sky130_fd_sc_hd__nand2_1 U21303 ( .A(n16471), .B(
        j202_soc_core_j22_cpu_rf_gpr[141]), .Y(n14240) );
  sky130_fd_sc_hd__nand2_1 U21304 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[365]), .Y(n14239) );
  sky130_fd_sc_hd__nand2_1 U21305 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[333]), .Y(n14238) );
  sky130_fd_sc_hd__and4_1 U21306 ( .A(n14241), .B(n14240), .C(n14239), .D(
        n14238), .X(n14242) );
  sky130_fd_sc_hd__nand4_1 U21307 ( .A(n14245), .B(n14244), .C(n14243), .D(
        n14242), .Y(n21853) );
  sky130_fd_sc_hd__nand2_1 U21308 ( .A(n21853), .B(n16513), .Y(n14255) );
  sky130_fd_sc_hd__nand2_1 U21309 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[13]), .Y(n14248) );
  sky130_fd_sc_hd__nand2_1 U21310 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[13]), .Y(n14247) );
  sky130_fd_sc_hd__nand2_1 U21311 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[493]), .Y(n14246) );
  sky130_fd_sc_hd__and4_1 U21312 ( .A(n14248), .B(n14247), .C(n16516), .D(
        n14246), .X(n14254) );
  sky130_fd_sc_hd__nand2_1 U21313 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[13]), .Y(n14252) );
  sky130_fd_sc_hd__nand2_1 U21314 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[13]), .Y(n14251) );
  sky130_fd_sc_hd__nand2_1 U21315 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[13]), .Y(n14250) );
  sky130_fd_sc_hd__nand2_1 U21316 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[13]), .Y(n14249) );
  sky130_fd_sc_hd__and4_1 U21317 ( .A(n14252), .B(n14251), .C(n14250), .D(
        n14249), .X(n14253) );
  sky130_fd_sc_hd__nand3_1 U21318 ( .A(n14255), .B(n14254), .C(n14253), .Y(
        n27365) );
  sky130_fd_sc_hd__nand2_1 U21319 ( .A(n27365), .B(n16529), .Y(n14256) );
  sky130_fd_sc_hd__o21ai_1 U21320 ( .A1(n14742), .A2(n27365), .B1(n14256), .Y(
        n14563) );
  sky130_fd_sc_hd__nor2_1 U21321 ( .A(n14562), .B(n14563), .Y(n21330) );
  sky130_fd_sc_hd__nor2_1 U21322 ( .A(n21332), .B(n21330), .Y(n14567) );
  sky130_fd_sc_hd__nand2_1 U21323 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[427]), .Y(n14260) );
  sky130_fd_sc_hd__nand2_1 U21324 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[235]), .Y(n14259) );
  sky130_fd_sc_hd__nand2_1 U21325 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[299]), .Y(n14258) );
  sky130_fd_sc_hd__nand2_1 U21326 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[203]), .Y(n14257) );
  sky130_fd_sc_hd__nand2_1 U21327 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[491]), .Y(n14264) );
  sky130_fd_sc_hd__a2bb2oi_1 U21328 ( .B1(j202_soc_core_j22_cpu_rf_tmp[11]), 
        .B2(n13774), .A1_N(n14466), .A2_N(n10990), .Y(n14263) );
  sky130_fd_sc_hd__nand2_1 U21329 ( .A(n15128), .B(
        j202_soc_core_j22_cpu_rf_gpr[171]), .Y(n14262) );
  sky130_fd_sc_hd__nand2_1 U21330 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[331]), .Y(n14261) );
  sky130_fd_sc_hd__nand4_1 U21331 ( .A(n14264), .B(n14263), .C(n14262), .D(
        n14261), .Y(n14265) );
  sky130_fd_sc_hd__a21oi_1 U21332 ( .A1(j202_soc_core_j22_cpu_rf_gpr[11]), 
        .A2(n16285), .B1(n14265), .Y(n14277) );
  sky130_fd_sc_hd__nand2_1 U21333 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[363]), .Y(n14269) );
  sky130_fd_sc_hd__nand2_1 U21334 ( .A(n16323), .B(
        j202_soc_core_j22_cpu_rf_gpr[459]), .Y(n14268) );
  sky130_fd_sc_hd__nand2_1 U21335 ( .A(n16324), .B(
        j202_soc_core_j22_cpu_rf_gpr[267]), .Y(n14267) );
  sky130_fd_sc_hd__nand2_1 U21336 ( .A(n11114), .B(
        j202_soc_core_j22_cpu_rf_gpr[395]), .Y(n14266) );
  sky130_fd_sc_hd__nand4_1 U21337 ( .A(n14269), .B(n14268), .C(n14267), .D(
        n14266), .Y(n14275) );
  sky130_fd_sc_hd__nand2_1 U21338 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[139]), .Y(n14273) );
  sky130_fd_sc_hd__nand2_1 U21339 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[107]), .Y(n14272) );
  sky130_fd_sc_hd__nand2_1 U21340 ( .A(n11155), .B(
        j202_soc_core_j22_cpu_rf_gpr[75]), .Y(n14271) );
  sky130_fd_sc_hd__nand2_1 U21341 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[43]), .Y(n14270) );
  sky130_fd_sc_hd__nand4_1 U21342 ( .A(n14273), .B(n14272), .C(n14271), .D(
        n14270), .Y(n14274) );
  sky130_fd_sc_hd__nor2_1 U21343 ( .A(n14275), .B(n14274), .Y(n14276) );
  sky130_fd_sc_hd__nand3_1 U21344 ( .A(n12259), .B(n14277), .C(n14276), .Y(
        n26720) );
  sky130_fd_sc_hd__nand2_1 U21345 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[172]), .Y(n14281) );
  sky130_fd_sc_hd__nand2_1 U21346 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[236]), .Y(n14280) );
  sky130_fd_sc_hd__nand2_1 U21347 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[492]), .Y(n14279) );
  sky130_fd_sc_hd__nand2_1 U21348 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[428]), .Y(n14278) );
  sky130_fd_sc_hd__nand4_1 U21349 ( .A(n14281), .B(n14280), .C(n14279), .D(
        n14278), .Y(n14287) );
  sky130_fd_sc_hd__nand2_1 U21350 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[12]), .Y(n14285) );
  sky130_fd_sc_hd__nand2_1 U21351 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[44]), .Y(n14284) );
  sky130_fd_sc_hd__nand2_1 U21352 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[108]), .Y(n14283) );
  sky130_fd_sc_hd__nand2_1 U21353 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[396]), .Y(n14282) );
  sky130_fd_sc_hd__nand4_1 U21354 ( .A(n14285), .B(n14284), .C(n14283), .D(
        n14282), .Y(n14286) );
  sky130_fd_sc_hd__nor2_1 U21355 ( .A(n14287), .B(n14286), .Y(n14296) );
  sky130_fd_sc_hd__a22oi_1 U21356 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[300]), .B1(n14414), .B2(
        j202_soc_core_j22_cpu_rf_gpr[460]), .Y(n14295) );
  sky130_fd_sc_hd__a22oi_1 U21357 ( .A1(n16470), .A2(
        j202_soc_core_j22_cpu_rf_gpr[204]), .B1(n16469), .B2(
        j202_soc_core_j22_cpu_rf_gpr[76]), .Y(n14294) );
  sky130_fd_sc_hd__nand2_1 U21358 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[268]), .Y(n14292) );
  sky130_fd_sc_hd__nand2_1 U21359 ( .A(n16471), .B(
        j202_soc_core_j22_cpu_rf_gpr[140]), .Y(n14291) );
  sky130_fd_sc_hd__nand2_1 U21360 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[364]), .Y(n14290) );
  sky130_fd_sc_hd__nand2_1 U21361 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[332]), .Y(n14289) );
  sky130_fd_sc_hd__and4_1 U21362 ( .A(n14292), .B(n14291), .C(n14290), .D(
        n14289), .X(n14293) );
  sky130_fd_sc_hd__nand4_1 U21363 ( .A(n14296), .B(n14295), .C(n14294), .D(
        n14293), .Y(n19494) );
  sky130_fd_sc_hd__nand2_1 U21364 ( .A(n19494), .B(n16513), .Y(n14306) );
  sky130_fd_sc_hd__nand2_1 U21365 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[12]), .Y(n14299) );
  sky130_fd_sc_hd__nand2_1 U21366 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[12]), .Y(n14298) );
  sky130_fd_sc_hd__nand2_1 U21367 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[492]), .Y(n14297) );
  sky130_fd_sc_hd__and4_1 U21368 ( .A(n14299), .B(n14298), .C(n16516), .D(
        n14297), .X(n14305) );
  sky130_fd_sc_hd__nand2_1 U21369 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[12]), .Y(n14303) );
  sky130_fd_sc_hd__nand2_1 U21370 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[12]), .Y(n14302) );
  sky130_fd_sc_hd__nand2_1 U21371 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[12]), .Y(n14301) );
  sky130_fd_sc_hd__nand2_1 U21372 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[12]), .Y(n14300) );
  sky130_fd_sc_hd__and4_1 U21373 ( .A(n14303), .B(n14302), .C(n14301), .D(
        n14300), .X(n14304) );
  sky130_fd_sc_hd__nand3_1 U21374 ( .A(n14306), .B(n14305), .C(n14304), .Y(
        n27372) );
  sky130_fd_sc_hd__nand2_1 U21375 ( .A(n27372), .B(n16529), .Y(n14307) );
  sky130_fd_sc_hd__nand2_1 U21377 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[234]), .Y(n14311) );
  sky130_fd_sc_hd__nand2_1 U21378 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[426]), .Y(n14310) );
  sky130_fd_sc_hd__nand2_1 U21379 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[202]), .Y(n14309) );
  sky130_fd_sc_hd__nand2_1 U21380 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[298]), .Y(n14308) );
  sky130_fd_sc_hd__and4_1 U21381 ( .A(n14311), .B(n14310), .C(n14309), .D(
        n14308), .X(n14329) );
  sky130_fd_sc_hd__nand2_1 U21382 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[490]), .Y(n14315) );
  sky130_fd_sc_hd__a2bb2oi_1 U21383 ( .B1(j202_soc_core_j22_cpu_rf_tmp[10]), 
        .B2(n13774), .A1_N(n14466), .A2_N(n10988), .Y(n14314) );
  sky130_fd_sc_hd__nand2_1 U21384 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[170]), .Y(n14313) );
  sky130_fd_sc_hd__nand2_1 U21385 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[330]), .Y(n14312) );
  sky130_fd_sc_hd__nand4_1 U21386 ( .A(n14315), .B(n14314), .C(n14313), .D(
        n14312), .Y(n14316) );
  sky130_fd_sc_hd__a21oi_1 U21387 ( .A1(j202_soc_core_j22_cpu_rf_gpr[10]), 
        .A2(n16369), .B1(n14316), .Y(n14328) );
  sky130_fd_sc_hd__nand2_1 U21388 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[362]), .Y(n14320) );
  sky130_fd_sc_hd__nand2_1 U21389 ( .A(n16323), .B(
        j202_soc_core_j22_cpu_rf_gpr[458]), .Y(n14319) );
  sky130_fd_sc_hd__nand2_1 U21390 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[138]), .Y(n14318) );
  sky130_fd_sc_hd__nand2_1 U21391 ( .A(n16431), .B(
        j202_soc_core_j22_cpu_rf_gpr[266]), .Y(n14317) );
  sky130_fd_sc_hd__nand4_1 U21392 ( .A(n14320), .B(n14319), .C(n14318), .D(
        n14317), .Y(n14326) );
  sky130_fd_sc_hd__nand2_1 U21393 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[394]), .Y(n14324) );
  sky130_fd_sc_hd__nand2_1 U21394 ( .A(n11116), .B(
        j202_soc_core_j22_cpu_rf_gpr[106]), .Y(n14323) );
  sky130_fd_sc_hd__nand2_1 U21395 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[74]), .Y(n14322) );
  sky130_fd_sc_hd__nand2_1 U21396 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[42]), .Y(n14321) );
  sky130_fd_sc_hd__nand4_1 U21397 ( .A(n14324), .B(n14323), .C(n14322), .D(
        n14321), .Y(n14325) );
  sky130_fd_sc_hd__nor2_1 U21398 ( .A(n14326), .B(n14325), .Y(n14327) );
  sky130_fd_sc_hd__nand3_1 U21399 ( .A(n14329), .B(n14328), .C(n14327), .Y(
        n26722) );
  sky130_fd_sc_hd__inv_2 U21400 ( .A(n26722), .Y(n26325) );
  sky130_fd_sc_hd__nand2_1 U21401 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[171]), .Y(n14333) );
  sky130_fd_sc_hd__nand2_1 U21402 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[235]), .Y(n14332) );
  sky130_fd_sc_hd__nand2_1 U21403 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[491]), .Y(n14331) );
  sky130_fd_sc_hd__nand2_1 U21404 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[427]), .Y(n14330) );
  sky130_fd_sc_hd__nand4_1 U21405 ( .A(n14333), .B(n14332), .C(n14331), .D(
        n14330), .Y(n14339) );
  sky130_fd_sc_hd__nand2_1 U21406 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[11]), .Y(n14337) );
  sky130_fd_sc_hd__nand2_1 U21407 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[43]), .Y(n14336) );
  sky130_fd_sc_hd__nand2_1 U21408 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[107]), .Y(n14335) );
  sky130_fd_sc_hd__nand2_1 U21409 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[395]), .Y(n14334) );
  sky130_fd_sc_hd__nand4_1 U21410 ( .A(n14337), .B(n14336), .C(n14335), .D(
        n14334), .Y(n14338) );
  sky130_fd_sc_hd__nor2_1 U21411 ( .A(n14339), .B(n14338), .Y(n14347) );
  sky130_fd_sc_hd__a22oi_1 U21412 ( .A1(n11160), .A2(
        j202_soc_core_j22_cpu_rf_gpr[299]), .B1(n23502), .B2(
        j202_soc_core_j22_cpu_rf_gpr[459]), .Y(n14346) );
  sky130_fd_sc_hd__a22oi_1 U21413 ( .A1(n16470), .A2(
        j202_soc_core_j22_cpu_rf_gpr[203]), .B1(n16469), .B2(
        j202_soc_core_j22_cpu_rf_gpr[75]), .Y(n14345) );
  sky130_fd_sc_hd__nand2_1 U21414 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[267]), .Y(n14343) );
  sky130_fd_sc_hd__nand2_1 U21415 ( .A(n16471), .B(
        j202_soc_core_j22_cpu_rf_gpr[139]), .Y(n14342) );
  sky130_fd_sc_hd__nand2_1 U21416 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[363]), .Y(n14341) );
  sky130_fd_sc_hd__nand2_1 U21417 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[331]), .Y(n14340) );
  sky130_fd_sc_hd__and4_1 U21418 ( .A(n14343), .B(n14342), .C(n14341), .D(
        n14340), .X(n14344) );
  sky130_fd_sc_hd__nand4_1 U21419 ( .A(n14347), .B(n14346), .C(n14345), .D(
        n14344), .Y(n21467) );
  sky130_fd_sc_hd__nand2_1 U21420 ( .A(n21467), .B(n16513), .Y(n14357) );
  sky130_fd_sc_hd__nand2_1 U21421 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[11]), .Y(n14351) );
  sky130_fd_sc_hd__nand2_1 U21422 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[11]), .Y(n14350) );
  sky130_fd_sc_hd__nand2_1 U21423 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[491]), .Y(n14349) );
  sky130_fd_sc_hd__nand2_1 U21424 ( .A(n13701), .B(n10989), .Y(n14348) );
  sky130_fd_sc_hd__nand2_1 U21425 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[11]), .Y(n14355) );
  sky130_fd_sc_hd__nand2_1 U21426 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[11]), .Y(n14354) );
  sky130_fd_sc_hd__nand2_1 U21427 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[11]), .Y(n14353) );
  sky130_fd_sc_hd__nand2_1 U21428 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[11]), .Y(n14352) );
  sky130_fd_sc_hd__and4_1 U21429 ( .A(n14355), .B(n14354), .C(n14353), .D(
        n14352), .X(n14356) );
  sky130_fd_sc_hd__nand3_1 U21430 ( .A(n14357), .B(n13323), .C(n14356), .Y(
        n27377) );
  sky130_fd_sc_hd__nand2_1 U21431 ( .A(n27377), .B(n16529), .Y(n14358) );
  sky130_fd_sc_hd__o21ai_1 U21432 ( .A1(n14742), .A2(n27377), .B1(n14358), .Y(
        n14559) );
  sky130_fd_sc_hd__nand2_1 U21433 ( .A(n14567), .B(n21324), .Y(n14569) );
  sky130_fd_sc_hd__nand2_1 U21434 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[231]), .Y(n14362) );
  sky130_fd_sc_hd__nand2_1 U21435 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[423]), .Y(n14361) );
  sky130_fd_sc_hd__nand2_1 U21436 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_rf_gpr[199]), .Y(n14360) );
  sky130_fd_sc_hd__nand2_1 U21437 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[295]), .Y(n14359) );
  sky130_fd_sc_hd__nand2_1 U21438 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[487]), .Y(n14367) );
  sky130_fd_sc_hd__a2bb2oi_1 U21439 ( .B1(j202_soc_core_j22_cpu_rf_tmp[7]), 
        .B2(n13774), .A1_N(n14466), .A2_N(n14363), .Y(n14366) );
  sky130_fd_sc_hd__nand2_1 U21440 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[327]), .Y(n14365) );
  sky130_fd_sc_hd__nand2_1 U21441 ( .A(n15128), .B(
        j202_soc_core_j22_cpu_rf_gpr[167]), .Y(n14364) );
  sky130_fd_sc_hd__nand4_1 U21442 ( .A(n14367), .B(n14366), .C(n14365), .D(
        n14364), .Y(n14368) );
  sky130_fd_sc_hd__a21oi_1 U21443 ( .A1(j202_soc_core_j22_cpu_rf_gpr[7]), .A2(
        n16285), .B1(n14368), .Y(n14380) );
  sky130_fd_sc_hd__nand2_1 U21444 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[359]), .Y(n14372) );
  sky130_fd_sc_hd__nand2_1 U21445 ( .A(n16323), .B(
        j202_soc_core_j22_cpu_rf_gpr[455]), .Y(n14371) );
  sky130_fd_sc_hd__nand2_1 U21446 ( .A(n16324), .B(
        j202_soc_core_j22_cpu_rf_gpr[263]), .Y(n14370) );
  sky130_fd_sc_hd__nand2_1 U21447 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[103]), .Y(n14369) );
  sky130_fd_sc_hd__nand4_1 U21448 ( .A(n14372), .B(n14371), .C(n14370), .D(
        n14369), .Y(n14378) );
  sky130_fd_sc_hd__nand2_1 U21449 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[135]), .Y(n14376) );
  sky130_fd_sc_hd__nand2_1 U21450 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[391]), .Y(n14375) );
  sky130_fd_sc_hd__nand2_1 U21451 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[71]), .Y(n14374) );
  sky130_fd_sc_hd__nand2_1 U21452 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[39]), .Y(n14373) );
  sky130_fd_sc_hd__nand4_1 U21453 ( .A(n14376), .B(n14375), .C(n14374), .D(
        n14373), .Y(n14377) );
  sky130_fd_sc_hd__nor2_1 U21454 ( .A(n14378), .B(n14377), .Y(n14379) );
  sky130_fd_sc_hd__inv_2 U21455 ( .A(n26729), .Y(n25798) );
  sky130_fd_sc_hd__nand2_1 U21456 ( .A(n16324), .B(
        j202_soc_core_j22_cpu_rf_gpr[264]), .Y(n14384) );
  sky130_fd_sc_hd__nand2_1 U21457 ( .A(n16323), .B(
        j202_soc_core_j22_cpu_rf_gpr[456]), .Y(n14383) );
  sky130_fd_sc_hd__nand2_1 U21458 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[136]), .Y(n14382) );
  sky130_fd_sc_hd__nand2_1 U21459 ( .A(n11155), .B(
        j202_soc_core_j22_cpu_rf_gpr[72]), .Y(n14381) );
  sky130_fd_sc_hd__nand2_1 U21460 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[424]), .Y(n14387) );
  sky130_fd_sc_hd__nand2_1 U21461 ( .A(n11114), .B(
        j202_soc_core_j22_cpu_rf_gpr[392]), .Y(n14386) );
  sky130_fd_sc_hd__nand2_1 U21462 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[104]), .Y(n14385) );
  sky130_fd_sc_hd__nand3_1 U21463 ( .A(n14387), .B(n14386), .C(n14385), .Y(
        n14388) );
  sky130_fd_sc_hd__nand2_1 U21464 ( .A(n16285), .B(
        j202_soc_core_j22_cpu_rf_gpr[8]), .Y(n14392) );
  sky130_fd_sc_hd__nand2_1 U21465 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_rf_gpr[200]), .Y(n14391) );
  sky130_fd_sc_hd__nand2_1 U21466 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[296]), .Y(n14390) );
  sky130_fd_sc_hd__nand2_1 U21467 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[232]), .Y(n14389) );
  sky130_fd_sc_hd__nand2_1 U21468 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[40]), .Y(n14396) );
  sky130_fd_sc_hd__nand2_1 U21469 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[168]), .Y(n14395) );
  sky130_fd_sc_hd__nand2_1 U21470 ( .A(n14393), .B(n10984), .Y(n14394) );
  sky130_fd_sc_hd__nand3_1 U21471 ( .A(n14396), .B(n14395), .C(n14394), .Y(
        n14402) );
  sky130_fd_sc_hd__nand2_1 U21472 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[488]), .Y(n14400) );
  sky130_fd_sc_hd__a2bb2oi_1 U21473 ( .B1(n13752), .B2(
        j202_soc_core_intr_vec__6_), .A1_N(n21997), .A2_N(n14749), .Y(n14399)
         );
  sky130_fd_sc_hd__nand2_1 U21474 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[328]), .Y(n14398) );
  sky130_fd_sc_hd__nand2_1 U21475 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[360]), .Y(n14397) );
  sky130_fd_sc_hd__nand4_1 U21476 ( .A(n14400), .B(n14399), .C(n14398), .D(
        n14397), .Y(n14401) );
  sky130_fd_sc_hd__nor2_1 U21477 ( .A(n14402), .B(n14401), .Y(n14403) );
  sky130_fd_sc_hd__o22ai_1 U21478 ( .A1(n13793), .A2(n25798), .B1(n25821), 
        .B2(n16492), .Y(n14550) );
  sky130_fd_sc_hd__nand2_1 U21479 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[168]), .Y(n14407) );
  sky130_fd_sc_hd__nand2_1 U21480 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[232]), .Y(n14406) );
  sky130_fd_sc_hd__nand2_1 U21481 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[488]), .Y(n14405) );
  sky130_fd_sc_hd__nand2_1 U21482 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[424]), .Y(n14404) );
  sky130_fd_sc_hd__nand4_1 U21483 ( .A(n14407), .B(n14406), .C(n14405), .D(
        n14404), .Y(n14413) );
  sky130_fd_sc_hd__nand2_1 U21484 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[8]), .Y(n14411) );
  sky130_fd_sc_hd__nand2_1 U21485 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[40]), .Y(n14410) );
  sky130_fd_sc_hd__nand2_1 U21486 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[104]), .Y(n14409) );
  sky130_fd_sc_hd__nand2_1 U21487 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[392]), .Y(n14408) );
  sky130_fd_sc_hd__nand4_1 U21488 ( .A(n14411), .B(n14410), .C(n14409), .D(
        n14408), .Y(n14412) );
  sky130_fd_sc_hd__nor2_1 U21489 ( .A(n14413), .B(n14412), .Y(n14422) );
  sky130_fd_sc_hd__a22oi_1 U21490 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[296]), .B1(n14414), .B2(
        j202_soc_core_j22_cpu_rf_gpr[456]), .Y(n14421) );
  sky130_fd_sc_hd__a22oi_1 U21491 ( .A1(n13676), .A2(
        j202_soc_core_j22_cpu_rf_gpr[200]), .B1(n23089), .B2(
        j202_soc_core_j22_cpu_rf_gpr[72]), .Y(n14420) );
  sky130_fd_sc_hd__nand2_1 U21492 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[264]), .Y(n14418) );
  sky130_fd_sc_hd__nand2_1 U21493 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[136]), .Y(n14417) );
  sky130_fd_sc_hd__nand2_1 U21494 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[360]), .Y(n14416) );
  sky130_fd_sc_hd__nand2_1 U21495 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[328]), .Y(n14415) );
  sky130_fd_sc_hd__and4_1 U21496 ( .A(n14418), .B(n14417), .C(n14416), .D(
        n14415), .X(n14419) );
  sky130_fd_sc_hd__nand4_1 U21497 ( .A(n14422), .B(n14421), .C(n14420), .D(
        n14419), .Y(n21990) );
  sky130_fd_sc_hd__nand2_1 U21498 ( .A(n21990), .B(n16513), .Y(n14430) );
  sky130_fd_sc_hd__o22ai_1 U21499 ( .A1(n21997), .A2(n16007), .B1(n16010), 
        .B2(n21991), .Y(n14424) );
  sky130_fd_sc_hd__a22o_1 U21500 ( .A1(n29563), .A2(
        j202_soc_core_j22_cpu_rf_gpr[488]), .B1(n29567), .B2(
        j202_soc_core_j22_cpu_rf_vbr[8]), .X(n14423) );
  sky130_fd_sc_hd__nor2_1 U21501 ( .A(n14424), .B(n14423), .Y(n14429) );
  sky130_fd_sc_hd__a2bb2oi_1 U21502 ( .B1(n13701), .B2(n10984), .A1_N(n21992), 
        .A2_N(n14539), .Y(n14425) );
  sky130_fd_sc_hd__o21ai_1 U21503 ( .A1(n21993), .A2(n11095), .B1(n14425), .Y(
        n14427) );
  sky130_fd_sc_hd__o22ai_1 U21504 ( .A1(n21998), .A2(n16014), .B1(n16008), 
        .B2(n21994), .Y(n14426) );
  sky130_fd_sc_hd__nor2_1 U21505 ( .A(n14427), .B(n14426), .Y(n14428) );
  sky130_fd_sc_hd__nand3_2 U21506 ( .A(n14430), .B(n14429), .C(n14428), .Y(
        n27396) );
  sky130_fd_sc_hd__mux2i_1 U21507 ( .A0(n14742), .A1(n16320), .S(n27396), .Y(
        n14551) );
  sky130_fd_sc_hd__nor2_1 U21508 ( .A(n14550), .B(n14551), .Y(n22582) );
  sky130_fd_sc_hd__o22ai_1 U21509 ( .A1(n16492), .A2(n25798), .B1(n11145), 
        .B2(n13793), .Y(n14548) );
  sky130_fd_sc_hd__nand2_1 U21510 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[167]), .Y(n14434) );
  sky130_fd_sc_hd__nand2_1 U21511 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[231]), .Y(n14433) );
  sky130_fd_sc_hd__nand2_1 U21512 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[487]), .Y(n14432) );
  sky130_fd_sc_hd__nand2_1 U21513 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[423]), .Y(n14431) );
  sky130_fd_sc_hd__nand4_1 U21514 ( .A(n14434), .B(n14433), .C(n14432), .D(
        n14431), .Y(n14440) );
  sky130_fd_sc_hd__nand2_1 U21515 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[7]), .Y(n14438) );
  sky130_fd_sc_hd__nand2_1 U21516 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[39]), .Y(n14437) );
  sky130_fd_sc_hd__nand2_1 U21517 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[103]), .Y(n14436) );
  sky130_fd_sc_hd__nand2_1 U21518 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[391]), .Y(n14435) );
  sky130_fd_sc_hd__nand4_1 U21519 ( .A(n14438), .B(n14437), .C(n14436), .D(
        n14435), .Y(n14439) );
  sky130_fd_sc_hd__nor2_1 U21520 ( .A(n14440), .B(n14439), .Y(n14451) );
  sky130_fd_sc_hd__nand2_1 U21521 ( .A(n16469), .B(
        j202_soc_core_j22_cpu_rf_gpr[71]), .Y(n14444) );
  sky130_fd_sc_hd__nand2_1 U21522 ( .A(n16470), .B(
        j202_soc_core_j22_cpu_rf_gpr[199]), .Y(n14443) );
  sky130_fd_sc_hd__nand2_1 U21523 ( .A(n11160), .B(
        j202_soc_core_j22_cpu_rf_gpr[295]), .Y(n14442) );
  sky130_fd_sc_hd__nand2_1 U21524 ( .A(n14414), .B(
        j202_soc_core_j22_cpu_rf_gpr[455]), .Y(n14441) );
  sky130_fd_sc_hd__and4_1 U21525 ( .A(n14444), .B(n14443), .C(n14442), .D(
        n14441), .X(n14450) );
  sky130_fd_sc_hd__nand2_1 U21526 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[263]), .Y(n14448) );
  sky130_fd_sc_hd__nand2_1 U21527 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[135]), .Y(n14447) );
  sky130_fd_sc_hd__nand2_1 U21528 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[359]), .Y(n14446) );
  sky130_fd_sc_hd__nand2_1 U21529 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[327]), .Y(n14445) );
  sky130_fd_sc_hd__and4_1 U21530 ( .A(n14448), .B(n14447), .C(n14446), .D(
        n14445), .X(n14449) );
  sky130_fd_sc_hd__nand3_1 U21531 ( .A(n14451), .B(n14450), .C(n14449), .Y(
        n19041) );
  sky130_fd_sc_hd__a22oi_1 U21532 ( .A1(n29563), .A2(
        j202_soc_core_j22_cpu_rf_gpr[487]), .B1(n29567), .B2(
        j202_soc_core_j22_cpu_rf_vbr[7]), .Y(n14458) );
  sky130_fd_sc_hd__o2bb2ai_1 U21533 ( .B1(n19043), .B2(n14539), .A1_N(n13701), 
        .A2_N(j202_soc_core_j22_cpu_regop_imm__7_), .Y(n14452) );
  sky130_fd_sc_hd__a21oi_1 U21534 ( .A1(n16012), .A2(
        j202_soc_core_j22_cpu_rf_gbr[7]), .B1(n14452), .Y(n14457) );
  sky130_fd_sc_hd__o22a_1 U21535 ( .A1(n19078), .A2(n16008), .B1(n16007), .B2(
        n14453), .X(n14456) );
  sky130_fd_sc_hd__o22a_1 U21536 ( .A1(n14454), .A2(n16014), .B1(n19042), .B2(
        n16010), .X(n14455) );
  sky130_fd_sc_hd__nand4_1 U21537 ( .A(n14458), .B(n14457), .C(n14456), .D(
        n14455), .Y(n14459) );
  sky130_fd_sc_hd__nand2_1 U21538 ( .A(n26790), .B(n16322), .Y(n14460) );
  sky130_fd_sc_hd__o21ai_1 U21539 ( .A1(n16320), .A2(n26790), .B1(n14460), .Y(
        n14549) );
  sky130_fd_sc_hd__nor2_1 U21540 ( .A(n14548), .B(n14549), .Y(n22587) );
  sky130_fd_sc_hd__nor2_1 U21541 ( .A(n22582), .B(n22587), .Y(n21479) );
  sky130_fd_sc_hd__nand2_1 U21542 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[425]), .Y(n14464) );
  sky130_fd_sc_hd__nand2_1 U21543 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[233]), .Y(n14463) );
  sky130_fd_sc_hd__nand2_1 U21544 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[201]), .Y(n14462) );
  sky130_fd_sc_hd__nand2_1 U21545 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[297]), .Y(n14461) );
  sky130_fd_sc_hd__and4_1 U21546 ( .A(n14464), .B(n14463), .C(n14462), .D(
        n14461), .X(n14485) );
  sky130_fd_sc_hd__nand2_1 U21547 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[489]), .Y(n14470) );
  sky130_fd_sc_hd__a2bb2oi_1 U21548 ( .B1(j202_soc_core_j22_cpu_rf_tmp[9]), 
        .B2(n13774), .A1_N(n14466), .A2_N(n10986), .Y(n14469) );
  sky130_fd_sc_hd__nand2_1 U21549 ( .A(n15128), .B(
        j202_soc_core_j22_cpu_rf_gpr[169]), .Y(n14468) );
  sky130_fd_sc_hd__nand2_1 U21550 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[329]), .Y(n14467) );
  sky130_fd_sc_hd__nand4_1 U21551 ( .A(n14470), .B(n14469), .C(n14468), .D(
        n14467), .Y(n14471) );
  sky130_fd_sc_hd__a21oi_1 U21552 ( .A1(j202_soc_core_j22_cpu_rf_gpr[9]), .A2(
        n16285), .B1(n14471), .Y(n14484) );
  sky130_fd_sc_hd__nand2_1 U21553 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[361]), .Y(n14475) );
  sky130_fd_sc_hd__nand2_1 U21554 ( .A(n16323), .B(
        j202_soc_core_j22_cpu_rf_gpr[457]), .Y(n14474) );
  sky130_fd_sc_hd__nand2_1 U21555 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[137]), .Y(n14473) );
  sky130_fd_sc_hd__nand2_1 U21556 ( .A(n16431), .B(
        j202_soc_core_j22_cpu_rf_gpr[265]), .Y(n14472) );
  sky130_fd_sc_hd__nand4_1 U21557 ( .A(n14475), .B(n14474), .C(n14473), .D(
        n14472), .Y(n14482) );
  sky130_fd_sc_hd__nand2_1 U21558 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[393]), .Y(n14480) );
  sky130_fd_sc_hd__nand2_1 U21559 ( .A(n11116), .B(
        j202_soc_core_j22_cpu_rf_gpr[105]), .Y(n14479) );
  sky130_fd_sc_hd__nand2_1 U21560 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[41]), .Y(n14478) );
  sky130_fd_sc_hd__nand2_1 U21561 ( .A(n11155), .B(
        j202_soc_core_j22_cpu_rf_gpr[73]), .Y(n14477) );
  sky130_fd_sc_hd__nand4_1 U21562 ( .A(n14480), .B(n14479), .C(n14478), .D(
        n14477), .Y(n14481) );
  sky130_fd_sc_hd__nor2_1 U21563 ( .A(n14482), .B(n14481), .Y(n14483) );
  sky130_fd_sc_hd__inv_2 U21564 ( .A(n26721), .Y(n25788) );
  sky130_fd_sc_hd__o22ai_1 U21565 ( .A1(n16492), .A2(n26325), .B1(n25788), 
        .B2(n13793), .Y(n14554) );
  sky130_fd_sc_hd__nand2_1 U21566 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[170]), .Y(n14489) );
  sky130_fd_sc_hd__nand2_1 U21567 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[234]), .Y(n14488) );
  sky130_fd_sc_hd__nand2_1 U21568 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[490]), .Y(n14487) );
  sky130_fd_sc_hd__nand2_1 U21569 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[426]), .Y(n14486) );
  sky130_fd_sc_hd__nand4_1 U21570 ( .A(n14489), .B(n14488), .C(n14487), .D(
        n14486), .Y(n14495) );
  sky130_fd_sc_hd__nand2_1 U21571 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[10]), .Y(n14493) );
  sky130_fd_sc_hd__nand2_1 U21572 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[42]), .Y(n14492) );
  sky130_fd_sc_hd__nand2_1 U21573 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[106]), .Y(n14491) );
  sky130_fd_sc_hd__nand2_1 U21574 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[394]), .Y(n14490) );
  sky130_fd_sc_hd__nand4_1 U21575 ( .A(n14493), .B(n14492), .C(n14491), .D(
        n14490), .Y(n14494) );
  sky130_fd_sc_hd__nor2_1 U21576 ( .A(n14495), .B(n14494), .Y(n14504) );
  sky130_fd_sc_hd__a22oi_1 U21577 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[298]), .B1(n14414), .B2(
        j202_soc_core_j22_cpu_rf_gpr[458]), .Y(n14503) );
  sky130_fd_sc_hd__a22oi_1 U21578 ( .A1(n23515), .A2(
        j202_soc_core_j22_cpu_rf_gpr[202]), .B1(n16469), .B2(
        j202_soc_core_j22_cpu_rf_gpr[74]), .Y(n14502) );
  sky130_fd_sc_hd__nand2_1 U21579 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[266]), .Y(n14500) );
  sky130_fd_sc_hd__nand2_1 U21580 ( .A(n16471), .B(
        j202_soc_core_j22_cpu_rf_gpr[138]), .Y(n14499) );
  sky130_fd_sc_hd__nand2_1 U21581 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[362]), .Y(n14498) );
  sky130_fd_sc_hd__nand2_1 U21582 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[330]), .Y(n14497) );
  sky130_fd_sc_hd__and4_1 U21583 ( .A(n14500), .B(n14499), .C(n14498), .D(
        n14497), .X(n14501) );
  sky130_fd_sc_hd__nand4_1 U21584 ( .A(n14504), .B(n14503), .C(n14502), .D(
        n14501), .Y(n19212) );
  sky130_fd_sc_hd__nand2_1 U21585 ( .A(n19212), .B(n16513), .Y(n14515) );
  sky130_fd_sc_hd__nand2_1 U21586 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[10]), .Y(n14508) );
  sky130_fd_sc_hd__nand2_1 U21587 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[10]), .Y(n14507) );
  sky130_fd_sc_hd__nand2_1 U21588 ( .A(n13701), .B(n10987), .Y(n14506) );
  sky130_fd_sc_hd__nand2_1 U21589 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[490]), .Y(n14505) );
  sky130_fd_sc_hd__and4_1 U21590 ( .A(n14508), .B(n14507), .C(n14506), .D(
        n14505), .X(n14514) );
  sky130_fd_sc_hd__nand2_1 U21591 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[10]), .Y(n14512) );
  sky130_fd_sc_hd__nand2_1 U21592 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[10]), .Y(n14511) );
  sky130_fd_sc_hd__nand2_1 U21593 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[10]), .Y(n14510) );
  sky130_fd_sc_hd__nand2_1 U21594 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[10]), .Y(n14509) );
  sky130_fd_sc_hd__and4_1 U21595 ( .A(n14512), .B(n14511), .C(n14510), .D(
        n14509), .X(n14513) );
  sky130_fd_sc_hd__nand3_1 U21596 ( .A(n14515), .B(n14514), .C(n14513), .Y(
        n27383) );
  sky130_fd_sc_hd__nand2_1 U21597 ( .A(n27383), .B(n16529), .Y(n14516) );
  sky130_fd_sc_hd__nor2_1 U21599 ( .A(n14554), .B(n14555), .Y(n22329) );
  sky130_fd_sc_hd__o22ai_1 U21600 ( .A1(n16492), .A2(n25788), .B1(n25821), 
        .B2(n13793), .Y(n14552) );
  sky130_fd_sc_hd__nand2_1 U21601 ( .A(n13794), .B(
        j202_soc_core_j22_cpu_rf_gpr[169]), .Y(n14520) );
  sky130_fd_sc_hd__nand2_1 U21602 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[233]), .Y(n14519) );
  sky130_fd_sc_hd__nand2_1 U21603 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[489]), .Y(n14518) );
  sky130_fd_sc_hd__nand2_1 U21604 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[425]), .Y(n14517) );
  sky130_fd_sc_hd__nand4_1 U21605 ( .A(n14520), .B(n14519), .C(n14518), .D(
        n14517), .Y(n14526) );
  sky130_fd_sc_hd__nand2_1 U21606 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[9]), .Y(n14524) );
  sky130_fd_sc_hd__nand2_1 U21607 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[41]), .Y(n14523) );
  sky130_fd_sc_hd__nand2_1 U21608 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[105]), .Y(n14522) );
  sky130_fd_sc_hd__nand2_1 U21609 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[393]), .Y(n14521) );
  sky130_fd_sc_hd__nand4_1 U21610 ( .A(n14524), .B(n14523), .C(n14522), .D(
        n14521), .Y(n14525) );
  sky130_fd_sc_hd__nor2_1 U21611 ( .A(n14526), .B(n14525), .Y(n14534) );
  sky130_fd_sc_hd__a22oi_1 U21612 ( .A1(n11160), .A2(
        j202_soc_core_j22_cpu_rf_gpr[297]), .B1(n23502), .B2(
        j202_soc_core_j22_cpu_rf_gpr[457]), .Y(n14533) );
  sky130_fd_sc_hd__a22oi_1 U21613 ( .A1(n23515), .A2(
        j202_soc_core_j22_cpu_rf_gpr[201]), .B1(n16469), .B2(
        j202_soc_core_j22_cpu_rf_gpr[73]), .Y(n14532) );
  sky130_fd_sc_hd__nand2_1 U21614 ( .A(n13680), .B(
        j202_soc_core_j22_cpu_rf_gpr[265]), .Y(n14530) );
  sky130_fd_sc_hd__nand2_1 U21615 ( .A(n16471), .B(
        j202_soc_core_j22_cpu_rf_gpr[137]), .Y(n14529) );
  sky130_fd_sc_hd__nand2_1 U21616 ( .A(n13686), .B(
        j202_soc_core_j22_cpu_rf_gpr[361]), .Y(n14528) );
  sky130_fd_sc_hd__nand2_1 U21617 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[329]), .Y(n14527) );
  sky130_fd_sc_hd__and4_1 U21618 ( .A(n14530), .B(n14529), .C(n14528), .D(
        n14527), .X(n14531) );
  sky130_fd_sc_hd__nand4_1 U21619 ( .A(n14534), .B(n14533), .C(n14532), .D(
        n14531), .Y(n22874) );
  sky130_fd_sc_hd__nand2_1 U21620 ( .A(n22874), .B(n16513), .Y(n14546) );
  sky130_fd_sc_hd__nand2_1 U21621 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[9]), .Y(n14538) );
  sky130_fd_sc_hd__nand2_1 U21622 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[9]), .Y(n14537) );
  sky130_fd_sc_hd__nand2_1 U21623 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[489]), .Y(n14536) );
  sky130_fd_sc_hd__nand2_1 U21624 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[9]), .Y(n14535) );
  sky130_fd_sc_hd__and4_1 U21625 ( .A(n14538), .B(n14537), .C(n14536), .D(
        n14535), .X(n14545) );
  sky130_fd_sc_hd__a2bb2oi_1 U21626 ( .B1(n13701), .B2(n10985), .A1_N(n22857), 
        .A2_N(n14539), .Y(n14540) );
  sky130_fd_sc_hd__o22ai_1 U21628 ( .A1(n14541), .A2(n16014), .B1(n16008), 
        .B2(n22861), .Y(n14542) );
  sky130_fd_sc_hd__nor2_1 U21629 ( .A(n14543), .B(n14542), .Y(n14544) );
  sky130_fd_sc_hd__nand3_1 U21630 ( .A(n14546), .B(n14545), .C(n14544), .Y(
        n27389) );
  sky130_fd_sc_hd__nand2_1 U21631 ( .A(n27389), .B(n16529), .Y(n14547) );
  sky130_fd_sc_hd__o21ai_1 U21632 ( .A1(n14742), .A2(n27389), .B1(n14547), .Y(
        n14553) );
  sky130_fd_sc_hd__nor2_1 U21633 ( .A(n14552), .B(n14553), .Y(n21478) );
  sky130_fd_sc_hd__nor2_1 U21634 ( .A(n22329), .B(n21478), .Y(n14557) );
  sky130_fd_sc_hd__nand2_1 U21635 ( .A(n21479), .B(n14557), .Y(n21326) );
  sky130_fd_sc_hd__nor2_1 U21636 ( .A(n14569), .B(n21326), .Y(n14571) );
  sky130_fd_sc_hd__nand2_1 U21637 ( .A(n14549), .B(n14548), .Y(n22585) );
  sky130_fd_sc_hd__nand2_1 U21638 ( .A(n14551), .B(n14550), .Y(n22583) );
  sky130_fd_sc_hd__o21ai_1 U21639 ( .A1(n22585), .A2(n22582), .B1(n22583), .Y(
        n21480) );
  sky130_fd_sc_hd__nand2_1 U21640 ( .A(n14553), .B(n14552), .Y(n22325) );
  sky130_fd_sc_hd__nand2_1 U21641 ( .A(n14555), .B(n14554), .Y(n22330) );
  sky130_fd_sc_hd__o21ai_1 U21642 ( .A1(n22325), .A2(n22329), .B1(n22330), .Y(
        n14556) );
  sky130_fd_sc_hd__a21oi_1 U21643 ( .A1(n14557), .A2(n21480), .B1(n14556), .Y(
        n21325) );
  sky130_fd_sc_hd__nand2_1 U21644 ( .A(n14559), .B(n14558), .Y(n21370) );
  sky130_fd_sc_hd__nand2_1 U21645 ( .A(n14561), .B(n14560), .Y(n21360) );
  sky130_fd_sc_hd__o21ai_1 U21646 ( .A1(n21370), .A2(n21359), .B1(n21360), .Y(
        n21327) );
  sky130_fd_sc_hd__nand2_1 U21647 ( .A(n14563), .B(n14562), .Y(n21345) );
  sky130_fd_sc_hd__nand2_1 U21648 ( .A(n14565), .B(n14564), .Y(n21333) );
  sky130_fd_sc_hd__a21oi_1 U21650 ( .A1(n14567), .A2(n21327), .B1(n14566), .Y(
        n14568) );
  sky130_fd_sc_hd__o21ai_1 U21651 ( .A1(n14569), .A2(n21325), .B1(n14568), .Y(
        n14570) );
  sky130_fd_sc_hd__a21o_4 U21652 ( .A1(n18998), .A2(n14571), .B1(n14570), .X(
        n22513) );
  sky130_fd_sc_hd__nand2_1 U21653 ( .A(n11114), .B(
        j202_soc_core_j22_cpu_rf_gpr[403]), .Y(n14575) );
  sky130_fd_sc_hd__nand2_1 U21654 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[371]), .Y(n14574) );
  sky130_fd_sc_hd__nand2_1 U21655 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[115]), .Y(n14573) );
  sky130_fd_sc_hd__nand2_1 U21656 ( .A(n11152), .B(
        j202_soc_core_j22_cpu_rf_gpr[51]), .Y(n14572) );
  sky130_fd_sc_hd__nand4_1 U21657 ( .A(n14575), .B(n14574), .C(n14573), .D(
        n14572), .Y(n14581) );
  sky130_fd_sc_hd__a21oi_1 U21658 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[19]), .B1(n16436), .Y(n14579) );
  sky130_fd_sc_hd__nand2_1 U21659 ( .A(n11155), .B(
        j202_soc_core_j22_cpu_rf_gpr[83]), .Y(n14578) );
  sky130_fd_sc_hd__nand2_1 U21660 ( .A(n16431), .B(
        j202_soc_core_j22_cpu_rf_gpr[275]), .Y(n14577) );
  sky130_fd_sc_hd__nand2_1 U21661 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[147]), .Y(n14576) );
  sky130_fd_sc_hd__nand4_1 U21662 ( .A(n14579), .B(n14578), .C(n14577), .D(
        n14576), .Y(n14580) );
  sky130_fd_sc_hd__nor2_1 U21663 ( .A(n14581), .B(n14580), .Y(n14592) );
  sky130_fd_sc_hd__nand2_1 U21664 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[435]), .Y(n14585) );
  sky130_fd_sc_hd__nand2_1 U21665 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[307]), .Y(n14584) );
  sky130_fd_sc_hd__nand2_1 U21666 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[211]), .Y(n14583) );
  sky130_fd_sc_hd__nand2_1 U21667 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[243]), .Y(n14582) );
  sky130_fd_sc_hd__nand2_1 U21668 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[499]), .Y(n14589) );
  sky130_fd_sc_hd__nand2_1 U21669 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[339]), .Y(n14588) );
  sky130_fd_sc_hd__nand2_1 U21670 ( .A(n15128), .B(
        j202_soc_core_j22_cpu_rf_gpr[179]), .Y(n14587) );
  sky130_fd_sc_hd__nand2_1 U21671 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[467]), .Y(n14586) );
  sky130_fd_sc_hd__nand4_1 U21672 ( .A(n14589), .B(n14588), .C(n14587), .D(
        n14586), .Y(n14590) );
  sky130_fd_sc_hd__a21oi_1 U21673 ( .A1(j202_soc_core_j22_cpu_rf_gpr[19]), 
        .A2(n16285), .B1(n14590), .Y(n14591) );
  sky130_fd_sc_hd__inv_2 U21674 ( .A(n26719), .Y(n25403) );
  sky130_fd_sc_hd__nand2_1 U21675 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[402]), .Y(n14597) );
  sky130_fd_sc_hd__nand2_1 U21676 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[466]), .Y(n14596) );
  sky130_fd_sc_hd__nand2_1 U21677 ( .A(n11154), .B(
        j202_soc_core_j22_cpu_rf_gpr[274]), .Y(n14595) );
  sky130_fd_sc_hd__nand2_1 U21678 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[146]), .Y(n14594) );
  sky130_fd_sc_hd__nand4_1 U21679 ( .A(n14597), .B(n14596), .C(n14595), .D(
        n14594), .Y(n14603) );
  sky130_fd_sc_hd__a21oi_1 U21680 ( .A1(j202_soc_core_j22_cpu_rf_tmp[18]), 
        .A2(n13774), .B1(n16436), .Y(n14601) );
  sky130_fd_sc_hd__nand2_1 U21681 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[114]), .Y(n14600) );
  sky130_fd_sc_hd__nand2_1 U21682 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[50]), .Y(n14599) );
  sky130_fd_sc_hd__nand2_1 U21683 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[82]), .Y(n14598) );
  sky130_fd_sc_hd__nand4_1 U21684 ( .A(n14601), .B(n14600), .C(n14599), .D(
        n14598), .Y(n14602) );
  sky130_fd_sc_hd__nor2_1 U21685 ( .A(n14603), .B(n14602), .Y(n14614) );
  sky130_fd_sc_hd__nand2_1 U21686 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[434]), .Y(n14607) );
  sky130_fd_sc_hd__nand2_1 U21687 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[242]), .Y(n14606) );
  sky130_fd_sc_hd__nand2_1 U21688 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[210]), .Y(n14605) );
  sky130_fd_sc_hd__nand2_1 U21689 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[306]), .Y(n14604) );
  sky130_fd_sc_hd__nand2_1 U21690 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[498]), .Y(n14611) );
  sky130_fd_sc_hd__nand2_1 U21691 ( .A(n15128), .B(
        j202_soc_core_j22_cpu_rf_gpr[178]), .Y(n14610) );
  sky130_fd_sc_hd__nand2_1 U21692 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[338]), .Y(n14609) );
  sky130_fd_sc_hd__nand2_1 U21693 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[370]), .Y(n14608) );
  sky130_fd_sc_hd__nand4_1 U21694 ( .A(n14611), .B(n14610), .C(n14609), .D(
        n14608), .Y(n14612) );
  sky130_fd_sc_hd__a21oi_1 U21695 ( .A1(j202_soc_core_j22_cpu_rf_gpr[18]), 
        .A2(n16285), .B1(n14612), .Y(n14613) );
  sky130_fd_sc_hd__o22ai_1 U21696 ( .A1(n16492), .A2(n25403), .B1(n26571), 
        .B2(n13793), .Y(n14836) );
  sky130_fd_sc_hd__nand2_1 U21697 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[179]), .Y(n14618) );
  sky130_fd_sc_hd__nand2_1 U21698 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[243]), .Y(n14617) );
  sky130_fd_sc_hd__nand2_1 U21699 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[499]), .Y(n14616) );
  sky130_fd_sc_hd__nand2_1 U21700 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[435]), .Y(n14615) );
  sky130_fd_sc_hd__nand4_1 U21701 ( .A(n14618), .B(n14617), .C(n14616), .D(
        n14615), .Y(n14624) );
  sky130_fd_sc_hd__nand2_1 U21702 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[19]), .Y(n14622) );
  sky130_fd_sc_hd__nand2_1 U21703 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[51]), .Y(n14621) );
  sky130_fd_sc_hd__nand2_1 U21704 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[115]), .Y(n14620) );
  sky130_fd_sc_hd__nand2_1 U21705 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[403]), .Y(n14619) );
  sky130_fd_sc_hd__nand4_1 U21706 ( .A(n14622), .B(n14621), .C(n14620), .D(
        n14619), .Y(n14623) );
  sky130_fd_sc_hd__nor2_1 U21707 ( .A(n14624), .B(n14623), .Y(n14631) );
  sky130_fd_sc_hd__a22oi_1 U21708 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[307]), .B1(n14414), .B2(
        j202_soc_core_j22_cpu_rf_gpr[467]), .Y(n14630) );
  sky130_fd_sc_hd__a22oi_1 U21709 ( .A1(n23515), .A2(
        j202_soc_core_j22_cpu_rf_gpr[211]), .B1(n16469), .B2(
        j202_soc_core_j22_cpu_rf_gpr[83]), .Y(n14629) );
  sky130_fd_sc_hd__nand2_1 U21710 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[275]), .Y(n14628) );
  sky130_fd_sc_hd__nand2_1 U21711 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[147]), .Y(n14627) );
  sky130_fd_sc_hd__nand2_1 U21712 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[371]), .Y(n14626) );
  sky130_fd_sc_hd__nand2_1 U21713 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[339]), .Y(n14625) );
  sky130_fd_sc_hd__nand4_1 U21714 ( .A(n14631), .B(n14630), .C(n14629), .D(
        n13326), .Y(n22970) );
  sky130_fd_sc_hd__nand2_1 U21715 ( .A(n22970), .B(n16513), .Y(n14640) );
  sky130_fd_sc_hd__nand2_1 U21716 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[19]), .Y(n14634) );
  sky130_fd_sc_hd__nand2_1 U21717 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[19]), .Y(n14633) );
  sky130_fd_sc_hd__nand2_1 U21718 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[499]), .Y(n14632) );
  sky130_fd_sc_hd__and4_1 U21719 ( .A(n14634), .B(n14633), .C(n16516), .D(
        n14632), .X(n14639) );
  sky130_fd_sc_hd__nand2_1 U21720 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[19]), .Y(n14638) );
  sky130_fd_sc_hd__nand2_1 U21721 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[19]), .Y(n14637) );
  sky130_fd_sc_hd__nand2_1 U21722 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[19]), .Y(n14636) );
  sky130_fd_sc_hd__nand2_1 U21723 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[19]), .Y(n14635) );
  sky130_fd_sc_hd__nand3_1 U21724 ( .A(n14640), .B(n14639), .C(n13327), .Y(
        n27425) );
  sky130_fd_sc_hd__nand2_1 U21725 ( .A(n27425), .B(n16529), .Y(n14641) );
  sky130_fd_sc_hd__o21ai_1 U21726 ( .A1(n14742), .A2(n27425), .B1(n14641), .Y(
        n14837) );
  sky130_fd_sc_hd__nor2_1 U21727 ( .A(n14836), .B(n14837), .Y(n15772) );
  sky130_fd_sc_hd__a22oi_1 U21728 ( .A1(n11116), .A2(
        j202_soc_core_j22_cpu_rf_gpr[111]), .B1(n11152), .B2(
        j202_soc_core_j22_cpu_rf_gpr[47]), .Y(n14646) );
  sky130_fd_sc_hd__nand2_1 U21729 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[207]), .Y(n14645) );
  sky130_fd_sc_hd__nand2_1 U21730 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[303]), .Y(n14644) );
  sky130_fd_sc_hd__nand2_1 U21731 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[431]), .Y(n14643) );
  sky130_fd_sc_hd__nand2_1 U21732 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[239]), .Y(n14651) );
  sky130_fd_sc_hd__o22ai_1 U21733 ( .A1(n14752), .A2(n14647), .B1(n19066), 
        .B2(n14749), .Y(n14648) );
  sky130_fd_sc_hd__a21oi_1 U21734 ( .A1(n16363), .A2(
        j202_soc_core_j22_cpu_rf_gpr[335]), .B1(n14648), .Y(n14650) );
  sky130_fd_sc_hd__nand2_1 U21735 ( .A(n15128), .B(
        j202_soc_core_j22_cpu_rf_gpr[175]), .Y(n14649) );
  sky130_fd_sc_hd__and4_1 U21736 ( .A(n14651), .B(n14650), .C(n14755), .D(
        n14649), .X(n14663) );
  sky130_fd_sc_hd__nand2_1 U21737 ( .A(n14758), .B(
        j202_soc_core_j22_cpu_rf_gpr[15]), .Y(n14655) );
  sky130_fd_sc_hd__nand2_1 U21738 ( .A(n11154), .B(
        j202_soc_core_j22_cpu_rf_gpr[271]), .Y(n14654) );
  sky130_fd_sc_hd__nand2_1 U21739 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[143]), .Y(n14653) );
  sky130_fd_sc_hd__nand2_1 U21740 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[79]), .Y(n14652) );
  sky130_fd_sc_hd__nand4_1 U21741 ( .A(n14655), .B(n14654), .C(n14653), .D(
        n14652), .Y(n14661) );
  sky130_fd_sc_hd__nand2_1 U21742 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[495]), .Y(n14659) );
  sky130_fd_sc_hd__nand2_1 U21743 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[367]), .Y(n14658) );
  sky130_fd_sc_hd__nand2_1 U21744 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[399]), .Y(n14657) );
  sky130_fd_sc_hd__nand2_1 U21745 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[463]), .Y(n14656) );
  sky130_fd_sc_hd__nand4_1 U21746 ( .A(n14659), .B(n14658), .C(n14657), .D(
        n14656), .Y(n14660) );
  sky130_fd_sc_hd__nor2_1 U21747 ( .A(n14661), .B(n14660), .Y(n14662) );
  sky130_fd_sc_hd__nand3_2 U21748 ( .A(n12195), .B(n14663), .C(n14662), .Y(
        n26726) );
  sky130_fd_sc_hd__inv_2 U21749 ( .A(n26726), .Y(n26567) );
  sky130_fd_sc_hd__nand2_1 U21750 ( .A(n16431), .B(
        j202_soc_core_j22_cpu_rf_gpr[272]), .Y(n14667) );
  sky130_fd_sc_hd__nand2_1 U21751 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[368]), .Y(n14666) );
  sky130_fd_sc_hd__nand2_1 U21752 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[144]), .Y(n14665) );
  sky130_fd_sc_hd__nand2_1 U21753 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[400]), .Y(n14664) );
  sky130_fd_sc_hd__nand4_1 U21754 ( .A(n14667), .B(n14666), .C(n14665), .D(
        n14664), .Y(n14674) );
  sky130_fd_sc_hd__a21oi_1 U21755 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[16]), .B1(n16436), .Y(n14672) );
  sky130_fd_sc_hd__nand2_1 U21756 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[112]), .Y(n14671) );
  sky130_fd_sc_hd__nand2_1 U21757 ( .A(n11152), .B(
        j202_soc_core_j22_cpu_rf_gpr[48]), .Y(n14670) );
  sky130_fd_sc_hd__nand2_1 U21758 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[80]), .Y(n14669) );
  sky130_fd_sc_hd__nand4_1 U21759 ( .A(n14672), .B(n14671), .C(n14670), .D(
        n14669), .Y(n14673) );
  sky130_fd_sc_hd__nor2_1 U21760 ( .A(n14674), .B(n14673), .Y(n14685) );
  sky130_fd_sc_hd__nand2_1 U21761 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[432]), .Y(n14678) );
  sky130_fd_sc_hd__nand2_1 U21762 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[240]), .Y(n14677) );
  sky130_fd_sc_hd__nand2_1 U21763 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_rf_gpr[208]), .Y(n14676) );
  sky130_fd_sc_hd__nand2_1 U21764 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[304]), .Y(n14675) );
  sky130_fd_sc_hd__nand2_1 U21765 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[496]), .Y(n14682) );
  sky130_fd_sc_hd__nand2_1 U21766 ( .A(n15128), .B(
        j202_soc_core_j22_cpu_rf_gpr[176]), .Y(n14681) );
  sky130_fd_sc_hd__nand2_1 U21767 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[336]), .Y(n14680) );
  sky130_fd_sc_hd__nand2_1 U21768 ( .A(n13821), .B(
        j202_soc_core_j22_cpu_rf_gpr[464]), .Y(n14679) );
  sky130_fd_sc_hd__nand4_1 U21769 ( .A(n14682), .B(n14681), .C(n14680), .D(
        n14679), .Y(n14683) );
  sky130_fd_sc_hd__a21oi_1 U21770 ( .A1(j202_soc_core_j22_cpu_rf_gpr[16]), 
        .A2(n16285), .B1(n14683), .Y(n14684) );
  sky130_fd_sc_hd__o22ai_1 U21771 ( .A1(n13793), .A2(n26567), .B1(n26581), 
        .B2(n16492), .Y(n14828) );
  sky130_fd_sc_hd__nand2_1 U21772 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[176]), .Y(n14689) );
  sky130_fd_sc_hd__nand2_1 U21773 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[240]), .Y(n14688) );
  sky130_fd_sc_hd__nand2_1 U21774 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[496]), .Y(n14687) );
  sky130_fd_sc_hd__nand2_1 U21775 ( .A(n15983), .B(
        j202_soc_core_j22_cpu_rf_gpr[432]), .Y(n14686) );
  sky130_fd_sc_hd__nand4_1 U21776 ( .A(n14689), .B(n14688), .C(n14687), .D(
        n14686), .Y(n14695) );
  sky130_fd_sc_hd__nand2_1 U21777 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[16]), .Y(n14693) );
  sky130_fd_sc_hd__nand2_1 U21778 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[48]), .Y(n14692) );
  sky130_fd_sc_hd__nand2_1 U21779 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[112]), .Y(n14691) );
  sky130_fd_sc_hd__nand2_1 U21780 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[400]), .Y(n14690) );
  sky130_fd_sc_hd__nand4_1 U21781 ( .A(n14693), .B(n14692), .C(n14691), .D(
        n14690), .Y(n14694) );
  sky130_fd_sc_hd__nor2_1 U21782 ( .A(n14695), .B(n14694), .Y(n14703) );
  sky130_fd_sc_hd__a22oi_1 U21783 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[304]), .B1(n14414), .B2(
        j202_soc_core_j22_cpu_rf_gpr[464]), .Y(n14702) );
  sky130_fd_sc_hd__a22oi_1 U21784 ( .A1(n23515), .A2(
        j202_soc_core_j22_cpu_rf_gpr[208]), .B1(n23089), .B2(
        j202_soc_core_j22_cpu_rf_gpr[80]), .Y(n14701) );
  sky130_fd_sc_hd__nand2_1 U21785 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[272]), .Y(n14699) );
  sky130_fd_sc_hd__nand2_1 U21786 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[144]), .Y(n14698) );
  sky130_fd_sc_hd__nand2_1 U21787 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[368]), .Y(n14697) );
  sky130_fd_sc_hd__nand2_1 U21788 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[336]), .Y(n14696) );
  sky130_fd_sc_hd__and4_1 U21789 ( .A(n14699), .B(n14698), .C(n14697), .D(
        n14696), .X(n14700) );
  sky130_fd_sc_hd__nand4_1 U21790 ( .A(n14703), .B(n14702), .C(n14701), .D(
        n14700), .Y(n22538) );
  sky130_fd_sc_hd__nand2_1 U21791 ( .A(n22538), .B(n16513), .Y(n14712) );
  sky130_fd_sc_hd__nand2_1 U21792 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[16]), .Y(n14706) );
  sky130_fd_sc_hd__nand2_1 U21793 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[16]), .Y(n14705) );
  sky130_fd_sc_hd__nand2_1 U21794 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[496]), .Y(n14704) );
  sky130_fd_sc_hd__and4_1 U21795 ( .A(n14706), .B(n14705), .C(n16516), .D(
        n14704), .X(n14711) );
  sky130_fd_sc_hd__nand2_1 U21796 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[16]), .Y(n14710) );
  sky130_fd_sc_hd__nand2_1 U21797 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[16]), .Y(n14709) );
  sky130_fd_sc_hd__nand2_1 U21798 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[16]), .Y(n14708) );
  sky130_fd_sc_hd__nand2_1 U21799 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[16]), .Y(n14707) );
  sky130_fd_sc_hd__nand3_1 U21800 ( .A(n14712), .B(n14711), .C(n13332), .Y(
        n27447) );
  sky130_fd_sc_hd__nand2_1 U21801 ( .A(n27447), .B(n16529), .Y(n14713) );
  sky130_fd_sc_hd__o21ai_1 U21802 ( .A1(n14742), .A2(n27447), .B1(n14713), .Y(
        n14829) );
  sky130_fd_sc_hd__nand2_1 U21803 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[175]), .Y(n14717) );
  sky130_fd_sc_hd__nand2_1 U21804 ( .A(n15982), .B(
        j202_soc_core_j22_cpu_rf_gpr[239]), .Y(n14716) );
  sky130_fd_sc_hd__nand2_1 U21805 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[495]), .Y(n14715) );
  sky130_fd_sc_hd__nand2_1 U21806 ( .A(n15983), .B(
        j202_soc_core_j22_cpu_rf_gpr[431]), .Y(n14714) );
  sky130_fd_sc_hd__nand4_1 U21807 ( .A(n14717), .B(n14716), .C(n14715), .D(
        n14714), .Y(n14723) );
  sky130_fd_sc_hd__nand2_1 U21808 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[15]), .Y(n14721) );
  sky130_fd_sc_hd__nand2_1 U21809 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[47]), .Y(n14720) );
  sky130_fd_sc_hd__nand2_1 U21810 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[111]), .Y(n14719) );
  sky130_fd_sc_hd__nand2_1 U21811 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[399]), .Y(n14718) );
  sky130_fd_sc_hd__nand4_1 U21812 ( .A(n14721), .B(n14720), .C(n14719), .D(
        n14718), .Y(n14722) );
  sky130_fd_sc_hd__nor2_1 U21813 ( .A(n14723), .B(n14722), .Y(n14732) );
  sky130_fd_sc_hd__a22oi_1 U21814 ( .A1(n14725), .A2(
        j202_soc_core_j22_cpu_rf_gpr[303]), .B1(n14724), .B2(
        j202_soc_core_j22_cpu_rf_gpr[463]), .Y(n14731) );
  sky130_fd_sc_hd__a22oi_1 U21815 ( .A1(n23515), .A2(
        j202_soc_core_j22_cpu_rf_gpr[207]), .B1(n23089), .B2(
        j202_soc_core_j22_cpu_rf_gpr[79]), .Y(n14730) );
  sky130_fd_sc_hd__nand2_1 U21816 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[271]), .Y(n14729) );
  sky130_fd_sc_hd__nand2_1 U21817 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[143]), .Y(n14728) );
  sky130_fd_sc_hd__nand2_1 U21818 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[367]), .Y(n14727) );
  sky130_fd_sc_hd__nand2_1 U21819 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[335]), .Y(n14726) );
  sky130_fd_sc_hd__nand4_1 U21820 ( .A(n14732), .B(n14731), .C(n14730), .D(
        n12224), .Y(n19062) );
  sky130_fd_sc_hd__nand2_1 U21821 ( .A(n19062), .B(n16513), .Y(n14741) );
  sky130_fd_sc_hd__nand2_1 U21822 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[15]), .Y(n14735) );
  sky130_fd_sc_hd__nand2_1 U21823 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[15]), .Y(n14734) );
  sky130_fd_sc_hd__nand2_1 U21824 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[495]), .Y(n14733) );
  sky130_fd_sc_hd__and4_1 U21825 ( .A(n14735), .B(n14734), .C(n16516), .D(
        n14733), .X(n14740) );
  sky130_fd_sc_hd__nand2_1 U21826 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[15]), .Y(n14739) );
  sky130_fd_sc_hd__nand2_1 U21827 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[15]), .Y(n14738) );
  sky130_fd_sc_hd__nand2_1 U21828 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[15]), .Y(n14737) );
  sky130_fd_sc_hd__nand2_1 U21829 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[15]), .Y(n14736) );
  sky130_fd_sc_hd__nand2_1 U21830 ( .A(n27354), .B(n16320), .Y(n14743) );
  sky130_fd_sc_hd__o21a_1 U21831 ( .A1(n27354), .A2(n16322), .B1(n14743), .X(
        n14826) );
  sky130_fd_sc_hd__nor2_1 U21832 ( .A(n14827), .B(n14826), .Y(n20997) );
  sky130_fd_sc_hd__nor2_1 U21833 ( .A(n20999), .B(n20997), .Y(n21013) );
  sky130_fd_sc_hd__a22oi_1 U21834 ( .A1(n11116), .A2(
        j202_soc_core_j22_cpu_rf_gpr[113]), .B1(n11152), .B2(
        j202_soc_core_j22_cpu_rf_gpr[49]), .Y(n14748) );
  sky130_fd_sc_hd__nand2_1 U21835 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[305]), .Y(n14747) );
  sky130_fd_sc_hd__nand2_1 U21836 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[433]), .Y(n14746) );
  sky130_fd_sc_hd__nand2_1 U21837 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[241]), .Y(n14745) );
  sky130_fd_sc_hd__nand2_1 U21838 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_rf_gpr[209]), .Y(n14757) );
  sky130_fd_sc_hd__o22ai_1 U21839 ( .A1(n14752), .A2(n14751), .B1(n14750), 
        .B2(n14749), .Y(n14753) );
  sky130_fd_sc_hd__a21oi_1 U21840 ( .A1(n16278), .A2(
        j202_soc_core_j22_cpu_rf_gpr[177]), .B1(n14753), .Y(n14756) );
  sky130_fd_sc_hd__nand2_1 U21841 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[337]), .Y(n14754) );
  sky130_fd_sc_hd__nand2_1 U21842 ( .A(n14758), .B(
        j202_soc_core_j22_cpu_rf_gpr[17]), .Y(n14762) );
  sky130_fd_sc_hd__nand2_1 U21843 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[145]), .Y(n14761) );
  sky130_fd_sc_hd__nand2_1 U21844 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[81]), .Y(n14760) );
  sky130_fd_sc_hd__nand2_1 U21845 ( .A(n11154), .B(
        j202_soc_core_j22_cpu_rf_gpr[273]), .Y(n14759) );
  sky130_fd_sc_hd__nand4_1 U21846 ( .A(n14762), .B(n14761), .C(n14760), .D(
        n14759), .Y(n14768) );
  sky130_fd_sc_hd__nand2_1 U21847 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[497]), .Y(n14766) );
  sky130_fd_sc_hd__nand2_1 U21848 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[369]), .Y(n14765) );
  sky130_fd_sc_hd__nand2_1 U21849 ( .A(n11114), .B(
        j202_soc_core_j22_cpu_rf_gpr[401]), .Y(n14764) );
  sky130_fd_sc_hd__nand2_1 U21850 ( .A(n16323), .B(
        j202_soc_core_j22_cpu_rf_gpr[465]), .Y(n14763) );
  sky130_fd_sc_hd__nand4_1 U21851 ( .A(n14766), .B(n14765), .C(n14764), .D(
        n14763), .Y(n14767) );
  sky130_fd_sc_hd__nor2_1 U21852 ( .A(n14768), .B(n14767), .Y(n14769) );
  sky130_fd_sc_hd__o22ai_1 U21853 ( .A1(n16492), .A2(n25128), .B1(n26581), 
        .B2(n13793), .Y(n14830) );
  sky130_fd_sc_hd__nand2_1 U21854 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[177]), .Y(n14774) );
  sky130_fd_sc_hd__nand2_1 U21855 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[241]), .Y(n14773) );
  sky130_fd_sc_hd__nand2_1 U21856 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[497]), .Y(n14772) );
  sky130_fd_sc_hd__nand2_1 U21857 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[433]), .Y(n14771) );
  sky130_fd_sc_hd__nand4_1 U21858 ( .A(n14774), .B(n14773), .C(n14772), .D(
        n14771), .Y(n14780) );
  sky130_fd_sc_hd__nand2_1 U21859 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[17]), .Y(n14778) );
  sky130_fd_sc_hd__nand2_1 U21860 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[49]), .Y(n14777) );
  sky130_fd_sc_hd__nand2_1 U21861 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[113]), .Y(n14776) );
  sky130_fd_sc_hd__nand2_1 U21862 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[401]), .Y(n14775) );
  sky130_fd_sc_hd__nand4_1 U21863 ( .A(n14778), .B(n14777), .C(n14776), .D(
        n14775), .Y(n14779) );
  sky130_fd_sc_hd__nor2_1 U21864 ( .A(n14780), .B(n14779), .Y(n14787) );
  sky130_fd_sc_hd__a22oi_1 U21865 ( .A1(n11160), .A2(
        j202_soc_core_j22_cpu_rf_gpr[305]), .B1(n14414), .B2(
        j202_soc_core_j22_cpu_rf_gpr[465]), .Y(n14786) );
  sky130_fd_sc_hd__a22oi_1 U21866 ( .A1(n23515), .A2(
        j202_soc_core_j22_cpu_rf_gpr[209]), .B1(n23089), .B2(
        j202_soc_core_j22_cpu_rf_gpr[81]), .Y(n14785) );
  sky130_fd_sc_hd__nand2_1 U21867 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[273]), .Y(n14784) );
  sky130_fd_sc_hd__nand2_1 U21868 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[145]), .Y(n14783) );
  sky130_fd_sc_hd__nand2_1 U21869 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[369]), .Y(n14782) );
  sky130_fd_sc_hd__nand2_1 U21870 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[337]), .Y(n14781) );
  sky130_fd_sc_hd__nand4_1 U21871 ( .A(n14787), .B(n14786), .C(n14785), .D(
        n13295), .Y(n22814) );
  sky130_fd_sc_hd__nand2_1 U21872 ( .A(n22814), .B(n16513), .Y(n14796) );
  sky130_fd_sc_hd__nand2_1 U21873 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[17]), .Y(n14790) );
  sky130_fd_sc_hd__nand2_1 U21874 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[17]), .Y(n14789) );
  sky130_fd_sc_hd__nand2_1 U21875 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[497]), .Y(n14788) );
  sky130_fd_sc_hd__and4_1 U21876 ( .A(n14790), .B(n14789), .C(n16516), .D(
        n14788), .X(n14795) );
  sky130_fd_sc_hd__nand2_1 U21877 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[17]), .Y(n14794) );
  sky130_fd_sc_hd__nand2_1 U21878 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[17]), .Y(n14793) );
  sky130_fd_sc_hd__nand2_1 U21879 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[17]), .Y(n14792) );
  sky130_fd_sc_hd__nand2_1 U21880 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[17]), .Y(n14791) );
  sky130_fd_sc_hd__nand3_1 U21881 ( .A(n14796), .B(n14795), .C(n13333), .Y(
        n24613) );
  sky130_fd_sc_hd__nand2_1 U21882 ( .A(n24613), .B(n16529), .Y(n14797) );
  sky130_fd_sc_hd__o22ai_1 U21884 ( .A1(n13793), .A2(n25128), .B1(n26571), 
        .B2(n16492), .Y(n14832) );
  sky130_fd_sc_hd__nand2_1 U21885 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[178]), .Y(n14801) );
  sky130_fd_sc_hd__nand2_1 U21886 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[242]), .Y(n14800) );
  sky130_fd_sc_hd__nand2_1 U21887 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[498]), .Y(n14799) );
  sky130_fd_sc_hd__nand2_1 U21888 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[434]), .Y(n14798) );
  sky130_fd_sc_hd__nand4_1 U21889 ( .A(n14801), .B(n14800), .C(n14799), .D(
        n14798), .Y(n14807) );
  sky130_fd_sc_hd__nand2_1 U21890 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[18]), .Y(n14805) );
  sky130_fd_sc_hd__nand2_1 U21891 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[50]), .Y(n14804) );
  sky130_fd_sc_hd__nand2_1 U21892 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[114]), .Y(n14803) );
  sky130_fd_sc_hd__nand2_1 U21893 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[402]), .Y(n14802) );
  sky130_fd_sc_hd__nand4_1 U21894 ( .A(n14805), .B(n14804), .C(n14803), .D(
        n14802), .Y(n14806) );
  sky130_fd_sc_hd__nor2_1 U21895 ( .A(n14807), .B(n14806), .Y(n14815) );
  sky130_fd_sc_hd__a22oi_1 U21896 ( .A1(n11160), .A2(
        j202_soc_core_j22_cpu_rf_gpr[306]), .B1(n14414), .B2(
        j202_soc_core_j22_cpu_rf_gpr[466]), .Y(n14814) );
  sky130_fd_sc_hd__a22oi_1 U21897 ( .A1(n16470), .A2(
        j202_soc_core_j22_cpu_rf_gpr[210]), .B1(n16469), .B2(
        j202_soc_core_j22_cpu_rf_gpr[82]), .Y(n14813) );
  sky130_fd_sc_hd__nand2_1 U21898 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[274]), .Y(n14811) );
  sky130_fd_sc_hd__nand2_1 U21899 ( .A(n16471), .B(
        j202_soc_core_j22_cpu_rf_gpr[146]), .Y(n14810) );
  sky130_fd_sc_hd__nand2_1 U21900 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[370]), .Y(n14809) );
  sky130_fd_sc_hd__nand2_1 U21901 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[338]), .Y(n14808) );
  sky130_fd_sc_hd__and4_1 U21902 ( .A(n14811), .B(n14810), .C(n14809), .D(
        n14808), .X(n14812) );
  sky130_fd_sc_hd__nand4_1 U21903 ( .A(n14815), .B(n14814), .C(n14813), .D(
        n14812), .Y(n22213) );
  sky130_fd_sc_hd__nand2_1 U21904 ( .A(n22213), .B(n16513), .Y(n14824) );
  sky130_fd_sc_hd__nand2_1 U21905 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[18]), .Y(n14818) );
  sky130_fd_sc_hd__nand2_1 U21906 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[18]), .Y(n14817) );
  sky130_fd_sc_hd__nand2_1 U21907 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[498]), .Y(n14816) );
  sky130_fd_sc_hd__and4_1 U21908 ( .A(n14818), .B(n14817), .C(n16516), .D(
        n14816), .X(n14823) );
  sky130_fd_sc_hd__nand2_1 U21909 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[18]), .Y(n14822) );
  sky130_fd_sc_hd__nand2_1 U21910 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[18]), .Y(n14821) );
  sky130_fd_sc_hd__nand2_1 U21911 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[18]), .Y(n14820) );
  sky130_fd_sc_hd__nand2_1 U21912 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[18]), .Y(n14819) );
  sky130_fd_sc_hd__nand3_1 U21913 ( .A(n14824), .B(n14823), .C(n13340), .Y(
        n27432) );
  sky130_fd_sc_hd__nand2_1 U21914 ( .A(n27432), .B(n16529), .Y(n14825) );
  sky130_fd_sc_hd__o21ai_1 U21915 ( .A1(n14742), .A2(n27432), .B1(n14825), .Y(
        n14833) );
  sky130_fd_sc_hd__nor2_1 U21916 ( .A(n14832), .B(n14833), .Y(n15512) );
  sky130_fd_sc_hd__nor2_1 U21917 ( .A(n21014), .B(n15512), .Y(n14835) );
  sky130_fd_sc_hd__nand2_1 U21918 ( .A(n21013), .B(n14835), .Y(n15412) );
  sky130_fd_sc_hd__nor2_1 U21919 ( .A(n15772), .B(n15412), .Y(n14839) );
  sky130_fd_sc_hd__nand2_1 U21920 ( .A(n14827), .B(n14826), .Y(n22511) );
  sky130_fd_sc_hd__nand2_1 U21921 ( .A(n14829), .B(n14828), .Y(n21000) );
  sky130_fd_sc_hd__nand2_1 U21922 ( .A(n14831), .B(n14830), .Y(n21015) );
  sky130_fd_sc_hd__nand2_1 U21923 ( .A(n14833), .B(n14832), .Y(n15513) );
  sky130_fd_sc_hd__nand2_1 U21925 ( .A(n14837), .B(n14836), .Y(n15773) );
  sky130_fd_sc_hd__a21oi_1 U21927 ( .A1(n22513), .A2(n14839), .B1(n14838), .Y(
        n14845) );
  sky130_fd_sc_hd__o22ai_1 U21928 ( .A1(n16492), .A2(n26417), .B1(n25403), 
        .B2(n13793), .Y(n14841) );
  sky130_fd_sc_hd__nand2_1 U21929 ( .A(n27419), .B(n16529), .Y(n14840) );
  sky130_fd_sc_hd__nor2_1 U21931 ( .A(n14841), .B(n14842), .Y(n15194) );
  sky130_fd_sc_hd__nand2_1 U21932 ( .A(n14842), .B(n14841), .Y(n15193) );
  sky130_fd_sc_hd__nand2_1 U21933 ( .A(n14843), .B(n15193), .Y(n14844) );
  sky130_fd_sc_hd__xor2_1 U21934 ( .A(n14845), .B(n14844), .X(n24531) );
  sky130_fd_sc_hd__nand2_1 U21935 ( .A(n24531), .B(n12158), .Y(n14848) );
  sky130_fd_sc_hd__nor2_1 U21936 ( .A(n23861), .B(n14849), .Y(n23490) );
  sky130_fd_sc_hd__nor2_1 U21937 ( .A(j202_soc_core_j22_cpu_opst[4]), .B(
        n23862), .Y(n23196) );
  sky130_fd_sc_hd__nor2_1 U21938 ( .A(n22024), .B(n14850), .Y(n23860) );
  sky130_fd_sc_hd__nand2_1 U21939 ( .A(n23196), .B(
        j202_soc_core_j22_cpu_opst[1]), .Y(n23197) );
  sky130_fd_sc_hd__nor2_1 U21940 ( .A(n24260), .B(n23197), .Y(n23564) );
  sky130_fd_sc_hd__nor3_1 U21941 ( .A(n23860), .B(n27914), .C(n23564), .Y(
        n14851) );
  sky130_fd_sc_hd__nand2_1 U21942 ( .A(n23860), .B(n27978), .Y(n27817) );
  sky130_fd_sc_hd__nor2_1 U21943 ( .A(j202_soc_core_j22_cpu_opst[3]), .B(
        n22275), .Y(n22025) );
  sky130_fd_sc_hd__nor2_1 U21944 ( .A(j202_soc_core_j22_cpu_opst[0]), .B(
        j202_soc_core_j22_cpu_opst[2]), .Y(n27904) );
  sky130_fd_sc_hd__nand2_1 U21945 ( .A(n22025), .B(n27904), .Y(n24470) );
  sky130_fd_sc_hd__nand2_1 U21946 ( .A(n27817), .B(n24470), .Y(n27931) );
  sky130_fd_sc_hd__nand2_1 U21947 ( .A(n27931), .B(
        j202_soc_core_j22_cpu_opst[1]), .Y(n27166) );
  sky130_fd_sc_hd__nand3_1 U21948 ( .A(n23490), .B(n14851), .C(n27166), .Y(
        n14855) );
  sky130_fd_sc_hd__nor2_1 U21949 ( .A(j202_soc_core_j22_cpu_istall), .B(n14852), .Y(n23488) );
  sky130_fd_sc_hd__o21ai_1 U21950 ( .A1(n24474), .A2(n12200), .B1(n20428), .Y(
        n14853) );
  sky130_fd_sc_hd__nand2_1 U21951 ( .A(n23488), .B(n14853), .Y(n14854) );
  sky130_fd_sc_hd__nand2_1 U21952 ( .A(n14855), .B(n14854), .Y(n28965) );
  sky130_fd_sc_hd__a22oi_1 U21953 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[56]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[88]), .Y(n14973) );
  sky130_fd_sc_hd__nand2_1 U21954 ( .A(n21675), .B(j202_soc_core_uart_div0[0]), 
        .Y(n14972) );
  sky130_fd_sc_hd__nand2_1 U21955 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[24]), .Y(n14971) );
  sky130_fd_sc_hd__nand4_1 U21956 ( .A(n14973), .B(n21677), .C(n14972), .D(
        n14971), .Y(n14969) );
  sky130_fd_sc_hd__nor2_1 U21957 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(n15454), .Y(n16126) );
  sky130_fd_sc_hd__nand2_1 U21958 ( .A(n16126), .B(n17277), .Y(n14936) );
  sky130_fd_sc_hd__nand2_1 U21959 ( .A(n17274), .B(n20788), .Y(n17279) );
  sky130_fd_sc_hd__nor2_1 U21960 ( .A(n17289), .B(n17279), .Y(n17067) );
  sky130_fd_sc_hd__nand2b_1 U21961 ( .A_N(n14936), .B(n17067), .Y(n16057) );
  sky130_fd_sc_hd__nor2_1 U21962 ( .A(n17293), .B(n17279), .Y(n14951) );
  sky130_fd_sc_hd__nor2_1 U21963 ( .A(n14936), .B(n14856), .Y(n17083) );
  sky130_fd_sc_hd__nand2_1 U21964 ( .A(n15454), .B(n20687), .Y(n14899) );
  sky130_fd_sc_hd__nor2_1 U21965 ( .A(n17277), .B(n14899), .Y(n14894) );
  sky130_fd_sc_hd__nand2_1 U21966 ( .A(n14894), .B(n15838), .Y(n15863) );
  sky130_fd_sc_hd__nand2b_1 U21967 ( .A_N(n15863), .B(n20579), .Y(n16098) );
  sky130_fd_sc_hd__nand2b_1 U21968 ( .A_N(n17083), .B(n16098), .Y(n17031) );
  sky130_fd_sc_hd__nand2_1 U21969 ( .A(n17274), .B(n20579), .Y(n17290) );
  sky130_fd_sc_hd__nand2_1 U21970 ( .A(n17271), .B(n17293), .Y(n14950) );
  sky130_fd_sc_hd__nor2_1 U21971 ( .A(n14936), .B(n14950), .Y(n15864) );
  sky130_fd_sc_hd__nor2_1 U21972 ( .A(n17314), .B(n14899), .Y(n14877) );
  sky130_fd_sc_hd__nor2_1 U21973 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .B(n13398), .Y(n17066) );
  sky130_fd_sc_hd__nand2_1 U21974 ( .A(n17066), .B(n17314), .Y(n14928) );
  sky130_fd_sc_hd__nor2_1 U21975 ( .A(n14857), .B(n14928), .Y(n15881) );
  sky130_fd_sc_hd__nor2_1 U21976 ( .A(n13306), .B(n15881), .Y(n14905) );
  sky130_fd_sc_hd__nand2_1 U21977 ( .A(n17066), .B(n17277), .Y(n15855) );
  sky130_fd_sc_hd__nand2_1 U21978 ( .A(n14858), .B(n14951), .Y(n14961) );
  sky130_fd_sc_hd__nand2_1 U21979 ( .A(n16126), .B(n17314), .Y(n14898) );
  sky130_fd_sc_hd__nand2b_1 U21980 ( .A_N(n14898), .B(n17067), .Y(n14859) );
  sky130_fd_sc_hd__nor2_1 U21981 ( .A(n17293), .B(n17290), .Y(n16564) );
  sky130_fd_sc_hd__nand2b_1 U21982 ( .A_N(n14936), .B(n16564), .Y(n14939) );
  sky130_fd_sc_hd__nand2b_1 U21983 ( .A_N(n14950), .B(n17066), .Y(n17073) );
  sky130_fd_sc_hd__nand2_1 U21984 ( .A(n14877), .B(n14951), .Y(n14862) );
  sky130_fd_sc_hd__nor2_1 U21985 ( .A(n14898), .B(n14950), .Y(n14946) );
  sky130_fd_sc_hd__nor3b_1 U21986 ( .C_N(n17073), .A(n14895), .B(n14946), .Y(
        n15821) );
  sky130_fd_sc_hd__nand2_1 U21987 ( .A(n16564), .B(n15871), .Y(n16099) );
  sky130_fd_sc_hd__nand2_1 U21988 ( .A(n14877), .B(n17271), .Y(n16091) );
  sky130_fd_sc_hd__nor2_1 U21989 ( .A(n17293), .B(n16091), .Y(n17071) );
  sky130_fd_sc_hd__nor2b_1 U21990 ( .B_N(n16099), .A(n17071), .Y(n15811) );
  sky130_fd_sc_hd__nor2_1 U21991 ( .A(n15786), .B(n14860), .Y(n15880) );
  sky130_fd_sc_hd__nand3_1 U21992 ( .A(n15821), .B(n15811), .C(n14900), .Y(
        n15865) );
  sky130_fd_sc_hd__nand2b_1 U21993 ( .A_N(n15855), .B(n16564), .Y(n14896) );
  sky130_fd_sc_hd__nand4b_1 U21994 ( .A_N(n15864), .B(n14905), .C(n16105), .D(
        n14896), .Y(n17029) );
  sky130_fd_sc_hd__nand2b_1 U21995 ( .A_N(n14898), .B(n16564), .Y(n14943) );
  sky130_fd_sc_hd__nand2_1 U21996 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .B(n20623), .Y(n14918) );
  sky130_fd_sc_hd__nor2_1 U21997 ( .A(n17277), .B(n14918), .Y(n14902) );
  sky130_fd_sc_hd__nand2_1 U21998 ( .A(n17067), .B(n14902), .Y(n16063) );
  sky130_fd_sc_hd__nand2_1 U21999 ( .A(n14943), .B(n16063), .Y(n17069) );
  sky130_fd_sc_hd__nor4b_1 U22000 ( .D_N(n16057), .A(n17031), .B(n17029), .C(
        n17069), .Y(n14869) );
  sky130_fd_sc_hd__nand2_1 U22001 ( .A(n14861), .B(n17314), .Y(n17088) );
  sky130_fd_sc_hd__nand2_1 U22002 ( .A(n16063), .B(n14862), .Y(n14904) );
  sky130_fd_sc_hd__nand2_1 U22003 ( .A(n19381), .B(n20788), .Y(n17169) );
  sky130_fd_sc_hd__nor2_1 U22004 ( .A(n17289), .B(n17169), .Y(n15870) );
  sky130_fd_sc_hd__nand2_1 U22005 ( .A(n14877), .B(n15870), .Y(n17010) );
  sky130_fd_sc_hd__nand2b_1 U22006 ( .A_N(n15855), .B(n17067), .Y(n17082) );
  sky130_fd_sc_hd__nand2_1 U22007 ( .A(n14863), .B(n16126), .Y(n14941) );
  sky130_fd_sc_hd__nand3_1 U22008 ( .A(n17082), .B(n16057), .C(n14941), .Y(
        n17030) );
  sky130_fd_sc_hd__and4_1 U22009 ( .A(n17088), .B(n14865), .C(n17010), .D(
        n14864), .X(n17028) );
  sky130_fd_sc_hd__nand2_1 U22010 ( .A(n16564), .B(n14902), .Y(n14897) );
  sky130_fd_sc_hd__nor2_1 U22011 ( .A(n17314), .B(n14918), .Y(n15818) );
  sky130_fd_sc_hd__nand2_1 U22012 ( .A(n14951), .B(n15818), .Y(n14954) );
  sky130_fd_sc_hd__nand2_1 U22013 ( .A(n14897), .B(n14954), .Y(n14944) );
  sky130_fd_sc_hd__nand2_1 U22014 ( .A(n19125), .B(n17293), .Y(n15854) );
  sky130_fd_sc_hd__nand2b_1 U22015 ( .A_N(n15854), .B(n14877), .Y(n17014) );
  sky130_fd_sc_hd__nand2_1 U22016 ( .A(n14951), .B(n14894), .Y(n15814) );
  sky130_fd_sc_hd__nand2_1 U22017 ( .A(n16091), .B(n15814), .Y(n17085) );
  sky130_fd_sc_hd__nor4b_1 U22018 ( .D_N(n14866), .A(n13306), .B(n16102), .C(
        n17085), .Y(n14867) );
  sky130_fd_sc_hd__a21oi_1 U22019 ( .A1(n17028), .A2(n14867), .B1(n17059), .Y(
        n14868) );
  sky130_fd_sc_hd__o21bai_1 U22020 ( .A1(n17278), .A2(n14869), .B1_N(n14868), 
        .Y(n14913) );
  sky130_fd_sc_hd__nand2_1 U22021 ( .A(n19125), .B(n17289), .Y(n15845) );
  sky130_fd_sc_hd__nor2_1 U22022 ( .A(n14918), .B(n15845), .Y(n17046) );
  sky130_fd_sc_hd__nand2_1 U22023 ( .A(n17046), .B(n17314), .Y(n15796) );
  sky130_fd_sc_hd__nand2_1 U22024 ( .A(n14894), .B(n16706), .Y(n15844) );
  sky130_fd_sc_hd__nand2_1 U22025 ( .A(n15796), .B(n15844), .Y(n17009) );
  sky130_fd_sc_hd__nor2_1 U22026 ( .A(n16119), .B(n17009), .Y(n16114) );
  sky130_fd_sc_hd__nand2_1 U22027 ( .A(n15870), .B(n14902), .Y(n17013) );
  sky130_fd_sc_hd__nor2_1 U22028 ( .A(n15845), .B(n15855), .Y(n17047) );
  sky130_fd_sc_hd__nor2_1 U22029 ( .A(n15854), .B(n14928), .Y(n15803) );
  sky130_fd_sc_hd__nor2_1 U22030 ( .A(n17047), .B(n15803), .Y(n17007) );
  sky130_fd_sc_hd__nor2_1 U22031 ( .A(n17169), .B(n15855), .Y(n15869) );
  sky130_fd_sc_hd__nand2b_1 U22032 ( .A_N(n15854), .B(n15818), .Y(n17049) );
  sky130_fd_sc_hd__nor2_1 U22033 ( .A(n17293), .B(n17169), .Y(n16197) );
  sky130_fd_sc_hd__nand2_1 U22034 ( .A(n14877), .B(n16197), .Y(n14917) );
  sky130_fd_sc_hd__nand2_1 U22035 ( .A(n17014), .B(n14917), .Y(n15853) );
  sky130_fd_sc_hd__nand2b_1 U22036 ( .A_N(n14898), .B(n15870), .Y(n16078) );
  sky130_fd_sc_hd__a211o_1 U22037 ( .A1(n15869), .A2(n17289), .B1(n15874), 
        .C1(n16118), .X(n15856) );
  sky130_fd_sc_hd__a22oi_1 U22038 ( .A1(n17273), .A2(n14872), .B1(n13388), 
        .B2(n14871), .Y(n17054) );
  sky130_fd_sc_hd__nand2_1 U22039 ( .A(n16197), .B(n14902), .Y(n15801) );
  sky130_fd_sc_hd__nor2_1 U22040 ( .A(n14936), .B(n14873), .Y(n15795) );
  sky130_fd_sc_hd__nand2b_1 U22041 ( .A_N(n14898), .B(n16197), .Y(n14929) );
  sky130_fd_sc_hd__nand2_1 U22042 ( .A(n17044), .B(n14874), .Y(n15849) );
  sky130_fd_sc_hd__nand2_1 U22043 ( .A(n14929), .B(n15849), .Y(n14916) );
  sky130_fd_sc_hd__nor3_1 U22044 ( .A(n14875), .B(n15795), .C(n14916), .Y(
        n17006) );
  sky130_fd_sc_hd__nand2b_1 U22045 ( .A_N(n19125), .B(n14884), .Y(n14876) );
  sky130_fd_sc_hd__nand2_1 U22046 ( .A(n14894), .B(n14876), .Y(n17048) );
  sky130_fd_sc_hd__nor2_1 U22047 ( .A(n15845), .B(n14885), .Y(n14882) );
  sky130_fd_sc_hd__nor2_1 U22048 ( .A(n14878), .B(n14882), .Y(n17042) );
  sky130_fd_sc_hd__nand2_1 U22049 ( .A(n17044), .B(n14879), .Y(n15802) );
  sky130_fd_sc_hd__nand2_1 U22050 ( .A(n16197), .B(n15818), .Y(n16110) );
  sky130_fd_sc_hd__a31oi_1 U22051 ( .A1(n17006), .A2(n17042), .A3(n13307), 
        .B1(n17055), .Y(n14892) );
  sky130_fd_sc_hd__nor2_1 U22052 ( .A(n14880), .B(n15854), .Y(n16111) );
  sky130_fd_sc_hd__nor2_1 U22053 ( .A(n14884), .B(n14928), .Y(n17045) );
  sky130_fd_sc_hd__nand2_1 U22054 ( .A(n15869), .B(n17293), .Y(n16113) );
  sky130_fd_sc_hd__nand2b_1 U22055 ( .A_N(n14936), .B(n16197), .Y(n15789) );
  sky130_fd_sc_hd__nor2_1 U22056 ( .A(n14881), .B(n15854), .Y(n16073) );
  sky130_fd_sc_hd__nand2_1 U22057 ( .A(n16073), .B(n17277), .Y(n16077) );
  sky130_fd_sc_hd__nand3_1 U22058 ( .A(n16113), .B(n15789), .C(n16077), .Y(
        n15800) );
  sky130_fd_sc_hd__nor4_1 U22059 ( .A(n14882), .B(n16111), .C(n17045), .D(
        n15800), .Y(n14883) );
  sky130_fd_sc_hd__nand2_1 U22060 ( .A(n14894), .B(n16197), .Y(n14919) );
  sky130_fd_sc_hd__a21oi_1 U22061 ( .A1(n14883), .A2(n14919), .B1(n17037), .Y(
        n14891) );
  sky130_fd_sc_hd__o21a_1 U22062 ( .A1(n14885), .A2(n14884), .B1(n17049), .X(
        n14925) );
  sky130_fd_sc_hd__o21a_1 U22063 ( .A1(n14886), .A2(n15854), .B1(n14925), .X(
        n14887) );
  sky130_fd_sc_hd__a31oi_1 U22064 ( .A1(n14887), .A2(n14919), .A3(n15789), 
        .B1(n17078), .Y(n14890) );
  sky130_fd_sc_hd__nor2_1 U22065 ( .A(n17277), .B(
        j202_soc_core_bootrom_00_address_w[9]), .Y(n14952) );
  sky130_fd_sc_hd__nand2b_1 U22066 ( .A_N(n15845), .B(n14952), .Y(n14927) );
  sky130_fd_sc_hd__nor2_1 U22067 ( .A(n20687), .B(n14927), .Y(n15858) );
  sky130_fd_sc_hd__nand2b_1 U22068 ( .A_N(n17046), .B(n17013), .Y(n16116) );
  sky130_fd_sc_hd__nor4b_1 U22069 ( .D_N(n13307), .A(n16111), .B(n15858), .C(
        n16116), .Y(n14888) );
  sky130_fd_sc_hd__inv_1 U22070 ( .A(n13387), .Y(n17039) );
  sky130_fd_sc_hd__a31oi_1 U22071 ( .A1(n14888), .A2(n14917), .A3(n17048), 
        .B1(n17039), .Y(n14889) );
  sky130_fd_sc_hd__or4_1 U22072 ( .A(n14892), .B(n14891), .C(n14890), .D(
        n14889), .X(n14893) );
  sky130_fd_sc_hd__nor2b_1 U22073 ( .B_N(n17054), .A(n14893), .Y(n14911) );
  sky130_fd_sc_hd__nand2_1 U22074 ( .A(n15818), .B(n15838), .Y(n17081) );
  sky130_fd_sc_hd__nand2b_1 U22075 ( .A_N(n17081), .B(n20788), .Y(n14942) );
  sky130_fd_sc_hd__nand2_1 U22076 ( .A(n14894), .B(n15870), .Y(n14920) );
  sky130_fd_sc_hd__nand2_1 U22077 ( .A(n14942), .B(n14920), .Y(n15836) );
  sky130_fd_sc_hd__nor3_1 U22078 ( .A(n14895), .B(n16055), .C(n15836), .Y(
        n16096) );
  sky130_fd_sc_hd__nand2_1 U22079 ( .A(n16096), .B(n14900), .Y(n17032) );
  sky130_fd_sc_hd__nand2b_1 U22080 ( .A_N(n14928), .B(n14951), .Y(n14934) );
  sky130_fd_sc_hd__nand2_1 U22081 ( .A(n14934), .B(n14896), .Y(n17070) );
  sky130_fd_sc_hd__nor2_1 U22082 ( .A(n14937), .B(n14898), .Y(n17075) );
  sky130_fd_sc_hd__nand2b_1 U22083 ( .A_N(n15863), .B(n20788), .Y(n14940) );
  sky130_fd_sc_hd__nand2b_1 U22084 ( .A_N(n13306), .B(n14940), .Y(n14960) );
  sky130_fd_sc_hd__o21ai_1 U22085 ( .A1(n14899), .A2(n14950), .B1(n15840), .Y(
        n16056) );
  sky130_fd_sc_hd__nor4_1 U22086 ( .A(n14903), .B(n17032), .C(n17070), .D(
        n16056), .Y(n14909) );
  sky130_fd_sc_hd__nand2_1 U22087 ( .A(n14951), .B(n14902), .Y(n17025) );
  sky130_fd_sc_hd__nand2_1 U22088 ( .A(n17025), .B(n14900), .Y(n15810) );
  sky130_fd_sc_hd__or4_1 U22089 ( .A(n16055), .B(n15817), .C(n17083), .D(
        n15810), .X(n14907) );
  sky130_fd_sc_hd__nor2_1 U22090 ( .A(n20788), .B(n17081), .Y(n14962) );
  sky130_fd_sc_hd__nor2_1 U22091 ( .A(n14901), .B(n14962), .Y(n16058) );
  sky130_fd_sc_hd__nand2_1 U22093 ( .A(n16172), .B(n14902), .Y(n15813) );
  sky130_fd_sc_hd__nor4b_2 U22094 ( .D_N(n15813), .A(n14904), .B(n14903), .C(
        n16095), .Y(n16093) );
  sky130_fd_sc_hd__nand3b_1 U22095 ( .A_N(n14906), .B(n16093), .C(n14905), .Y(
        n17034) );
  sky130_fd_sc_hd__o21a_1 U22097 ( .A1(n17039), .A2(n14909), .B1(n14908), .X(
        n14910) );
  sky130_fd_sc_hd__mux2i_1 U22098 ( .A0(n14911), .A1(n14910), .S(
        j202_soc_core_bootrom_00_address_w[11]), .Y(n14912) );
  sky130_fd_sc_hd__o21ai_1 U22099 ( .A1(n14913), .A2(n14912), .B1(n17061), .Y(
        n14968) );
  sky130_fd_sc_hd__nand2b_1 U22100 ( .A_N(n15869), .B(n14927), .Y(n14914) );
  sky130_fd_sc_hd__nand2_1 U22101 ( .A(n17013), .B(n14919), .Y(n15847) );
  sky130_fd_sc_hd__nor2_1 U22102 ( .A(n14914), .B(n15847), .Y(n17005) );
  sky130_fd_sc_hd__a21oi_1 U22103 ( .A1(n15870), .A2(n16126), .B1(n15857), .Y(
        n16121) );
  sky130_fd_sc_hd__a31oi_1 U22104 ( .A1(n17005), .A2(n14915), .A3(n16121), 
        .B1(n17039), .Y(n14933) );
  sky130_fd_sc_hd__nor2b_1 U22105 ( .B_N(n14917), .A(n14916), .Y(n14924) );
  sky130_fd_sc_hd__nand2b_1 U22106 ( .A_N(n16119), .B(n14924), .Y(n16075) );
  sky130_fd_sc_hd__nor2b_1 U22107 ( .B_N(n14920), .A(n16075), .Y(n15797) );
  sky130_fd_sc_hd__nand2_1 U22108 ( .A(n16197), .B(n15837), .Y(n17012) );
  sky130_fd_sc_hd__a31oi_1 U22109 ( .A1(n15797), .A2(n17012), .A3(n14919), 
        .B1(n17078), .Y(n14932) );
  sky130_fd_sc_hd__nand2_1 U22110 ( .A(n14920), .B(n16110), .Y(n16081) );
  sky130_fd_sc_hd__nand2_1 U22111 ( .A(n16073), .B(n17314), .Y(n14926) );
  sky130_fd_sc_hd__nor4_1 U22112 ( .A(n14922), .B(n14921), .C(n16081), .D(
        n16117), .Y(n14923) );
  sky130_fd_sc_hd__a21oi_1 U22113 ( .A1(n14924), .A2(n14923), .B1(n17055), .Y(
        n16085) );
  sky130_fd_sc_hd__o211ai_1 U22114 ( .A1(n20623), .A2(n14927), .B1(n14926), 
        .C1(n14925), .Y(n16080) );
  sky130_fd_sc_hd__a31oi_1 U22115 ( .A1(n15870), .A2(n15454), .A3(n14928), 
        .B1(n16080), .Y(n14930) );
  sky130_fd_sc_hd__a21oi_1 U22116 ( .A1(n14930), .A2(n14929), .B1(n17037), .Y(
        n14931) );
  sky130_fd_sc_hd__or3_1 U22117 ( .A(n14932), .B(n16085), .C(n14931), .X(
        n17022) );
  sky130_fd_sc_hd__nor2_1 U22118 ( .A(j202_soc_core_bootrom_00_address_w[11]), 
        .B(n17061), .Y(n17021) );
  sky130_fd_sc_hd__o21ai_1 U22119 ( .A1(n14933), .A2(n17022), .B1(n17021), .Y(
        n14967) );
  sky130_fd_sc_hd__nor2_1 U22120 ( .A(n14935), .B(n17076), .Y(n16064) );
  sky130_fd_sc_hd__o21ai_1 U22121 ( .A1(n15855), .A2(n17290), .B1(n16064), .Y(
        n17033) );
  sky130_fd_sc_hd__nand3_1 U22122 ( .A(n16063), .B(n15814), .C(n16099), .Y(
        n17065) );
  sky130_fd_sc_hd__nor4_1 U22124 ( .A(n16056), .B(n17033), .C(n17065), .D(
        n14938), .Y(n14959) );
  sky130_fd_sc_hd__nor2_1 U22125 ( .A(n15881), .B(n15864), .Y(n16065) );
  sky130_fd_sc_hd__nand4_1 U22126 ( .A(n17088), .B(n16093), .C(n14940), .D(
        n14939), .Y(n14948) );
  sky130_fd_sc_hd__nor2_1 U22127 ( .A(n20579), .B(n14941), .Y(n15867) );
  sky130_fd_sc_hd__nand2b_1 U22128 ( .A_N(n15867), .B(n14942), .Y(n16067) );
  sky130_fd_sc_hd__nor2_1 U22129 ( .A(n14945), .B(n14944), .Y(n16059) );
  sky130_fd_sc_hd__nand2_1 U22130 ( .A(n16059), .B(n14947), .Y(n15833) );
  sky130_fd_sc_hd__nor3_1 U22131 ( .A(n14948), .B(n16067), .C(n15833), .Y(
        n14949) );
  sky130_fd_sc_hd__nand2_1 U22132 ( .A(n16065), .B(n14949), .Y(n14957) );
  sky130_fd_sc_hd__nand2b_1 U22133 ( .A_N(n14951), .B(n14950), .Y(n14953) );
  sky130_fd_sc_hd__nand2_1 U22134 ( .A(n14953), .B(n14952), .Y(n14955) );
  sky130_fd_sc_hd__nor2_1 U22135 ( .A(n15882), .B(n15867), .Y(n15822) );
  sky130_fd_sc_hd__a21oi_1 U22136 ( .A1(n14955), .A2(n15822), .B1(n17037), .Y(
        n14956) );
  sky130_fd_sc_hd__a21oi_1 U22137 ( .A1(n14957), .A2(n13387), .B1(n14956), .Y(
        n14958) );
  sky130_fd_sc_hd__nand2b_1 U22139 ( .A_N(n14960), .B(n17073), .Y(n15816) );
  sky130_fd_sc_hd__nand2_1 U22140 ( .A(n15813), .B(n14961), .Y(n15819) );
  sky130_fd_sc_hd__a31oi_1 U22142 ( .A1(n17077), .A2(n16091), .A3(n17025), 
        .B1(n17078), .Y(n14963) );
  sky130_fd_sc_hd__nand2_1 U22143 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .B(n19354), .Y(n15830) );
  sky130_fd_sc_hd__o21ai_1 U22144 ( .A1(n14964), .A2(n14963), .B1(n17094), .Y(
        n14966) );
  sky130_fd_sc_hd__a31oi_1 U22145 ( .A1(n14968), .A2(n14967), .A3(n14966), 
        .B1(n14965), .Y(n14974) );
  sky130_fd_sc_hd__nor2_1 U22146 ( .A(n14969), .B(n14974), .Y(n14970) );
  sky130_fd_sc_hd__nand2_1 U22147 ( .A(j202_soc_core_memory0_ram_dout0[504]), 
        .B(n21771), .Y(n14977) );
  sky130_fd_sc_hd__nand4_1 U22148 ( .A(n14973), .B(n21738), .C(n14972), .D(
        n14971), .Y(n14975) );
  sky130_fd_sc_hd__nor2_1 U22149 ( .A(n14975), .B(n14974), .Y(n14976) );
  sky130_fd_sc_hd__nand2_1 U22150 ( .A(n14977), .B(n14976), .Y(n14978) );
  sky130_fd_sc_hd__nand2_1 U22151 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[152]), .Y(n14983) );
  sky130_fd_sc_hd__nand2_1 U22152 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[376]), .Y(n14982) );
  sky130_fd_sc_hd__nand2_1 U22153 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[120]), .Y(n14981) );
  sky130_fd_sc_hd__nand2_1 U22154 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[88]), .Y(n14980) );
  sky130_fd_sc_hd__nand4_1 U22155 ( .A(n14983), .B(n14982), .C(n14981), .D(
        n14980), .Y(n14989) );
  sky130_fd_sc_hd__a21oi_1 U22156 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[24]), .B1(n16436), .Y(n14987) );
  sky130_fd_sc_hd__nand2_1 U22157 ( .A(n11114), .B(
        j202_soc_core_j22_cpu_rf_gpr[408]), .Y(n14986) );
  sky130_fd_sc_hd__nand2_1 U22158 ( .A(n16324), .B(
        j202_soc_core_j22_cpu_rf_gpr[280]), .Y(n14985) );
  sky130_fd_sc_hd__nand2_1 U22159 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[56]), .Y(n14984) );
  sky130_fd_sc_hd__nand4_1 U22160 ( .A(n14987), .B(n14986), .C(n14985), .D(
        n14984), .Y(n14988) );
  sky130_fd_sc_hd__nor2_1 U22161 ( .A(n14989), .B(n14988), .Y(n15001) );
  sky130_fd_sc_hd__nand2_1 U22162 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[440]), .Y(n14993) );
  sky130_fd_sc_hd__nand2_1 U22163 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_rf_gpr[216]), .Y(n14992) );
  sky130_fd_sc_hd__nand2_1 U22164 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[312]), .Y(n14991) );
  sky130_fd_sc_hd__nand2_1 U22165 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[248]), .Y(n14990) );
  sky130_fd_sc_hd__and4_1 U22166 ( .A(n14993), .B(n14992), .C(n14991), .D(
        n14990), .X(n15000) );
  sky130_fd_sc_hd__nand2_1 U22167 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[504]), .Y(n14997) );
  sky130_fd_sc_hd__nand2_1 U22168 ( .A(n15128), .B(
        j202_soc_core_j22_cpu_rf_gpr[184]), .Y(n14996) );
  sky130_fd_sc_hd__nand2_1 U22169 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[344]), .Y(n14995) );
  sky130_fd_sc_hd__nand2_1 U22170 ( .A(n16323), .B(
        j202_soc_core_j22_cpu_rf_gpr[472]), .Y(n14994) );
  sky130_fd_sc_hd__nand4_1 U22171 ( .A(n14997), .B(n14996), .C(n14995), .D(
        n14994), .Y(n14998) );
  sky130_fd_sc_hd__a21oi_1 U22172 ( .A1(j202_soc_core_j22_cpu_rf_gpr[24]), 
        .A2(n16285), .B1(n14998), .Y(n14999) );
  sky130_fd_sc_hd__nand3_1 U22173 ( .A(n15001), .B(n15000), .C(n14999), .Y(
        n25871) );
  sky130_fd_sc_hd__inv_2 U22174 ( .A(n25871), .Y(n26701) );
  sky130_fd_sc_hd__nand2_1 U22175 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[184]), .Y(n15005) );
  sky130_fd_sc_hd__nand2_1 U22176 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[248]), .Y(n15004) );
  sky130_fd_sc_hd__nand2_1 U22177 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[504]), .Y(n15003) );
  sky130_fd_sc_hd__nand2_1 U22178 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[440]), .Y(n15002) );
  sky130_fd_sc_hd__nand4_1 U22179 ( .A(n15005), .B(n15004), .C(n15003), .D(
        n15002), .Y(n15011) );
  sky130_fd_sc_hd__nand2_1 U22180 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[24]), .Y(n15009) );
  sky130_fd_sc_hd__nand2_1 U22181 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[56]), .Y(n15008) );
  sky130_fd_sc_hd__nand2_1 U22182 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[120]), .Y(n15007) );
  sky130_fd_sc_hd__nand2_1 U22183 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[408]), .Y(n15006) );
  sky130_fd_sc_hd__nand4_1 U22184 ( .A(n15009), .B(n15008), .C(n15007), .D(
        n15006), .Y(n15010) );
  sky130_fd_sc_hd__nor2_1 U22185 ( .A(n15011), .B(n15010), .Y(n15019) );
  sky130_fd_sc_hd__a22oi_1 U22186 ( .A1(n11160), .A2(
        j202_soc_core_j22_cpu_rf_gpr[312]), .B1(n23502), .B2(
        j202_soc_core_j22_cpu_rf_gpr[472]), .Y(n15018) );
  sky130_fd_sc_hd__a22oi_1 U22187 ( .A1(n23515), .A2(
        j202_soc_core_j22_cpu_rf_gpr[216]), .B1(n16469), .B2(
        j202_soc_core_j22_cpu_rf_gpr[88]), .Y(n15017) );
  sky130_fd_sc_hd__nand2_1 U22188 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[280]), .Y(n15015) );
  sky130_fd_sc_hd__nand2_1 U22189 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[152]), .Y(n15014) );
  sky130_fd_sc_hd__nand2_1 U22190 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[376]), .Y(n15013) );
  sky130_fd_sc_hd__nand2_1 U22191 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[344]), .Y(n15012) );
  sky130_fd_sc_hd__and4_1 U22192 ( .A(n15015), .B(n15014), .C(n15013), .D(
        n15012), .X(n15016) );
  sky130_fd_sc_hd__nand4_1 U22193 ( .A(n15019), .B(n15018), .C(n15017), .D(
        n15016), .Y(n22568) );
  sky130_fd_sc_hd__nand2_1 U22194 ( .A(n22568), .B(n16513), .Y(n15029) );
  sky130_fd_sc_hd__nand2_1 U22195 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[24]), .Y(n15022) );
  sky130_fd_sc_hd__nand2_1 U22196 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[24]), .Y(n15021) );
  sky130_fd_sc_hd__nand2_1 U22197 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[504]), .Y(n15020) );
  sky130_fd_sc_hd__and4_1 U22198 ( .A(n15022), .B(n15021), .C(n16516), .D(
        n15020), .X(n15028) );
  sky130_fd_sc_hd__nand2_1 U22199 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[24]), .Y(n15026) );
  sky130_fd_sc_hd__nand2_1 U22200 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[24]), .Y(n15025) );
  sky130_fd_sc_hd__nand2_1 U22201 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[24]), .Y(n15024) );
  sky130_fd_sc_hd__nand2_1 U22202 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[24]), .Y(n15023) );
  sky130_fd_sc_hd__and4_1 U22203 ( .A(n15026), .B(n15025), .C(n15024), .D(
        n15023), .X(n15027) );
  sky130_fd_sc_hd__nand3_1 U22204 ( .A(n15029), .B(n15028), .C(n15027), .Y(
        n27392) );
  sky130_fd_sc_hd__nand2_1 U22205 ( .A(n22515), .B(n27392), .Y(n15035) );
  sky130_fd_sc_hd__nand2_1 U22206 ( .A(j202_soc_core_j22_cpu_pc[19]), .B(
        j202_soc_core_j22_cpu_pc[20]), .Y(n15031) );
  sky130_fd_sc_hd__nor2_1 U22207 ( .A(n15031), .B(n15030), .Y(n15297) );
  sky130_fd_sc_hd__nand2_1 U22208 ( .A(j202_soc_core_j22_cpu_pc[21]), .B(
        j202_soc_core_j22_cpu_pc[22]), .Y(n15299) );
  sky130_fd_sc_hd__nor2_1 U22209 ( .A(n15301), .B(n15299), .Y(n15032) );
  sky130_fd_sc_hd__nand2_1 U22210 ( .A(n15297), .B(n15032), .Y(n16027) );
  sky130_fd_sc_hd__nor2_1 U22211 ( .A(n16027), .B(n21009), .Y(n15033) );
  sky130_fd_sc_hd__xnor2_1 U22212 ( .A(n16028), .B(n15033), .Y(n25851) );
  sky130_fd_sc_hd__nand2_1 U22213 ( .A(n22596), .B(n25851), .Y(n15034) );
  sky130_fd_sc_hd__o211a_2 U22214 ( .A1(n26701), .A2(n11143), .B1(n15035), 
        .C1(n15034), .X(n15214) );
  sky130_fd_sc_hd__nand2_1 U22215 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[151]), .Y(n15039) );
  sky130_fd_sc_hd__nand2_1 U22216 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[375]), .Y(n15038) );
  sky130_fd_sc_hd__nand2_1 U22217 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[55]), .Y(n15037) );
  sky130_fd_sc_hd__nand2_1 U22218 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[87]), .Y(n15036) );
  sky130_fd_sc_hd__nand4_1 U22219 ( .A(n15039), .B(n15038), .C(n15037), .D(
        n15036), .Y(n15045) );
  sky130_fd_sc_hd__a21oi_1 U22220 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[23]), .B1(n16436), .Y(n15043) );
  sky130_fd_sc_hd__nand2_1 U22221 ( .A(n11114), .B(
        j202_soc_core_j22_cpu_rf_gpr[407]), .Y(n15042) );
  sky130_fd_sc_hd__nand2_1 U22222 ( .A(n16324), .B(
        j202_soc_core_j22_cpu_rf_gpr[279]), .Y(n15041) );
  sky130_fd_sc_hd__nand2_1 U22223 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[119]), .Y(n15040) );
  sky130_fd_sc_hd__nand4_1 U22224 ( .A(n15043), .B(n15042), .C(n15041), .D(
        n15040), .Y(n15044) );
  sky130_fd_sc_hd__nor2_1 U22225 ( .A(n15045), .B(n15044), .Y(n15057) );
  sky130_fd_sc_hd__nand2_1 U22226 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[439]), .Y(n15049) );
  sky130_fd_sc_hd__nand2_1 U22227 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[215]), .Y(n15048) );
  sky130_fd_sc_hd__nand2_1 U22228 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[311]), .Y(n15047) );
  sky130_fd_sc_hd__nand2_1 U22229 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[247]), .Y(n15046) );
  sky130_fd_sc_hd__and4_1 U22230 ( .A(n15049), .B(n15048), .C(n15047), .D(
        n15046), .X(n15056) );
  sky130_fd_sc_hd__nand2_1 U22231 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[503]), .Y(n15053) );
  sky130_fd_sc_hd__nand2_1 U22232 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[183]), .Y(n15052) );
  sky130_fd_sc_hd__nand2_1 U22233 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[343]), .Y(n15051) );
  sky130_fd_sc_hd__nand2_1 U22234 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[471]), .Y(n15050) );
  sky130_fd_sc_hd__nand4_1 U22235 ( .A(n15053), .B(n15052), .C(n15051), .D(
        n15050), .Y(n15054) );
  sky130_fd_sc_hd__a21oi_1 U22236 ( .A1(j202_soc_core_j22_cpu_rf_gpr[23]), 
        .A2(n16285), .B1(n15054), .Y(n15055) );
  sky130_fd_sc_hd__inv_2 U22237 ( .A(n26061), .Y(n26704) );
  sky130_fd_sc_hd__nand2_1 U22238 ( .A(n16431), .B(
        j202_soc_core_j22_cpu_rf_gpr[278]), .Y(n15061) );
  sky130_fd_sc_hd__nand2_1 U22239 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[374]), .Y(n15060) );
  sky130_fd_sc_hd__nand2_1 U22240 ( .A(n11116), .B(
        j202_soc_core_j22_cpu_rf_gpr[118]), .Y(n15059) );
  sky130_fd_sc_hd__nand2_1 U22241 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[54]), .Y(n15058) );
  sky130_fd_sc_hd__nand4_1 U22242 ( .A(n15061), .B(n15060), .C(n15059), .D(
        n15058), .Y(n15069) );
  sky130_fd_sc_hd__a21oi_1 U22243 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[22]), .B1(n16436), .Y(n15067) );
  sky130_fd_sc_hd__nand2_1 U22244 ( .A(n11114), .B(
        j202_soc_core_j22_cpu_rf_gpr[406]), .Y(n15066) );
  sky130_fd_sc_hd__nand2_1 U22245 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[150]), .Y(n15065) );
  sky130_fd_sc_hd__nand2_1 U22246 ( .A(n11155), .B(
        j202_soc_core_j22_cpu_rf_gpr[86]), .Y(n15064) );
  sky130_fd_sc_hd__nand4_1 U22247 ( .A(n15067), .B(n15066), .C(n15065), .D(
        n15064), .Y(n15068) );
  sky130_fd_sc_hd__nor2_1 U22248 ( .A(n15069), .B(n15068), .Y(n15081) );
  sky130_fd_sc_hd__nand2_1 U22249 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[310]), .Y(n15073) );
  sky130_fd_sc_hd__nand2_1 U22250 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[214]), .Y(n15072) );
  sky130_fd_sc_hd__nand2_1 U22251 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[438]), .Y(n15071) );
  sky130_fd_sc_hd__nand2_1 U22252 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[246]), .Y(n15070) );
  sky130_fd_sc_hd__and4_1 U22253 ( .A(n15073), .B(n15072), .C(n15071), .D(
        n15070), .X(n15080) );
  sky130_fd_sc_hd__nand2_1 U22254 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[502]), .Y(n15077) );
  sky130_fd_sc_hd__nand2_1 U22255 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[182]), .Y(n15076) );
  sky130_fd_sc_hd__nand2_1 U22256 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[342]), .Y(n15075) );
  sky130_fd_sc_hd__nand2_1 U22257 ( .A(n16323), .B(
        j202_soc_core_j22_cpu_rf_gpr[470]), .Y(n15074) );
  sky130_fd_sc_hd__nand4_1 U22258 ( .A(n15077), .B(n15076), .C(n15075), .D(
        n15074), .Y(n15078) );
  sky130_fd_sc_hd__a21oi_1 U22259 ( .A1(j202_soc_core_j22_cpu_rf_gpr[22]), 
        .A2(n16369), .B1(n15078), .Y(n15079) );
  sky130_fd_sc_hd__inv_2 U22260 ( .A(n26508), .Y(n26703) );
  sky130_fd_sc_hd__o22ai_1 U22261 ( .A1(n16492), .A2(n26704), .B1(n26703), 
        .B2(n13793), .Y(n15203) );
  sky130_fd_sc_hd__nand2_1 U22262 ( .A(n16469), .B(
        j202_soc_core_j22_cpu_rf_gpr[87]), .Y(n15085) );
  sky130_fd_sc_hd__nand2_1 U22263 ( .A(n23515), .B(
        j202_soc_core_j22_cpu_rf_gpr[215]), .Y(n15084) );
  sky130_fd_sc_hd__nand2_1 U22264 ( .A(n11160), .B(
        j202_soc_core_j22_cpu_rf_gpr[311]), .Y(n15083) );
  sky130_fd_sc_hd__nand2_1 U22265 ( .A(n23502), .B(
        j202_soc_core_j22_cpu_rf_gpr[471]), .Y(n15082) );
  sky130_fd_sc_hd__nand4_1 U22266 ( .A(n15085), .B(n15084), .C(n15083), .D(
        n15082), .Y(n15091) );
  sky130_fd_sc_hd__nand2_1 U22267 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[279]), .Y(n15089) );
  sky130_fd_sc_hd__nand2_1 U22268 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[343]), .Y(n15088) );
  sky130_fd_sc_hd__nand2_1 U22269 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[375]), .Y(n15087) );
  sky130_fd_sc_hd__nand2_1 U22270 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[151]), .Y(n15086) );
  sky130_fd_sc_hd__nand4_1 U22271 ( .A(n15089), .B(n15088), .C(n15087), .D(
        n15086), .Y(n15090) );
  sky130_fd_sc_hd__nor2_1 U22272 ( .A(n15091), .B(n15090), .Y(n15103) );
  sky130_fd_sc_hd__nand2_1 U22273 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[183]), .Y(n15095) );
  sky130_fd_sc_hd__nand2_1 U22274 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[247]), .Y(n15094) );
  sky130_fd_sc_hd__nand2_1 U22275 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[503]), .Y(n15093) );
  sky130_fd_sc_hd__nand2_1 U22276 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[439]), .Y(n15092) );
  sky130_fd_sc_hd__nand4_1 U22277 ( .A(n15095), .B(n15094), .C(n15093), .D(
        n15092), .Y(n15101) );
  sky130_fd_sc_hd__nand2_1 U22278 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[23]), .Y(n15099) );
  sky130_fd_sc_hd__nand2_1 U22279 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[55]), .Y(n15098) );
  sky130_fd_sc_hd__nand2_1 U22280 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[119]), .Y(n15097) );
  sky130_fd_sc_hd__nand2_1 U22281 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[407]), .Y(n15096) );
  sky130_fd_sc_hd__nand4_1 U22282 ( .A(n15099), .B(n15098), .C(n15097), .D(
        n15096), .Y(n15100) );
  sky130_fd_sc_hd__nor2_1 U22283 ( .A(n15101), .B(n15100), .Y(n15102) );
  sky130_fd_sc_hd__nand2_1 U22284 ( .A(n15103), .B(n15102), .Y(n22040) );
  sky130_fd_sc_hd__nand2_1 U22285 ( .A(n22040), .B(n16513), .Y(n15112) );
  sky130_fd_sc_hd__nand2_1 U22286 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[23]), .Y(n15106) );
  sky130_fd_sc_hd__nand2_1 U22287 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[23]), .Y(n15105) );
  sky130_fd_sc_hd__nand2_1 U22288 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[503]), .Y(n15104) );
  sky130_fd_sc_hd__and4_1 U22289 ( .A(n15106), .B(n15105), .C(n16516), .D(
        n15104), .X(n15111) );
  sky130_fd_sc_hd__nand2_1 U22290 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[23]), .Y(n15110) );
  sky130_fd_sc_hd__nand2_1 U22291 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[23]), .Y(n15109) );
  sky130_fd_sc_hd__nand2_1 U22292 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[23]), .Y(n15108) );
  sky130_fd_sc_hd__nand2_1 U22293 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[23]), .Y(n15107) );
  sky130_fd_sc_hd__nand3_1 U22294 ( .A(n15112), .B(n15111), .C(n12219), .Y(
        n27399) );
  sky130_fd_sc_hd__nand2_1 U22295 ( .A(n27399), .B(n16529), .Y(n15113) );
  sky130_fd_sc_hd__o21ai_1 U22296 ( .A1(n14742), .A2(n27399), .B1(n15113), .Y(
        n15204) );
  sky130_fd_sc_hd__nor2_1 U22297 ( .A(n15203), .B(n15204), .Y(n15899) );
  sky130_fd_sc_hd__nor2_1 U22298 ( .A(n15194), .B(n15772), .Y(n15415) );
  sky130_fd_sc_hd__nand2_1 U22299 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[405]), .Y(n15117) );
  sky130_fd_sc_hd__nand2_1 U22300 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[469]), .Y(n15116) );
  sky130_fd_sc_hd__nand2_1 U22301 ( .A(n11154), .B(
        j202_soc_core_j22_cpu_rf_gpr[277]), .Y(n15115) );
  sky130_fd_sc_hd__nand2_1 U22302 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[149]), .Y(n15114) );
  sky130_fd_sc_hd__nand4_1 U22303 ( .A(n15117), .B(n15116), .C(n15115), .D(
        n15114), .Y(n15123) );
  sky130_fd_sc_hd__a21oi_1 U22304 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[21]), .B1(n16436), .Y(n15121) );
  sky130_fd_sc_hd__nand2_1 U22305 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[117]), .Y(n15120) );
  sky130_fd_sc_hd__nand2_1 U22306 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[53]), .Y(n15119) );
  sky130_fd_sc_hd__nand2_1 U22307 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[85]), .Y(n15118) );
  sky130_fd_sc_hd__nand4_1 U22308 ( .A(n15121), .B(n15120), .C(n15119), .D(
        n15118), .Y(n15122) );
  sky130_fd_sc_hd__nor2_1 U22309 ( .A(n15123), .B(n15122), .Y(n15135) );
  sky130_fd_sc_hd__nand2_1 U22310 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[437]), .Y(n15127) );
  sky130_fd_sc_hd__nand2_1 U22311 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[245]), .Y(n15126) );
  sky130_fd_sc_hd__nand2_1 U22312 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_rf_gpr[213]), .Y(n15125) );
  sky130_fd_sc_hd__nand2_1 U22313 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[309]), .Y(n15124) );
  sky130_fd_sc_hd__nand2_1 U22314 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[501]), .Y(n15132) );
  sky130_fd_sc_hd__nand2_1 U22315 ( .A(n15128), .B(
        j202_soc_core_j22_cpu_rf_gpr[181]), .Y(n15131) );
  sky130_fd_sc_hd__nand2_1 U22316 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[341]), .Y(n15130) );
  sky130_fd_sc_hd__nand2_1 U22317 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[373]), .Y(n15129) );
  sky130_fd_sc_hd__nand4_1 U22318 ( .A(n15132), .B(n15131), .C(n15130), .D(
        n15129), .Y(n15133) );
  sky130_fd_sc_hd__a21oi_1 U22319 ( .A1(j202_soc_core_j22_cpu_rf_gpr[21]), 
        .A2(n16285), .B1(n15133), .Y(n15134) );
  sky130_fd_sc_hd__inv_2 U22320 ( .A(n27183), .Y(n26570) );
  sky130_fd_sc_hd__o22ai_1 U22321 ( .A1(n16492), .A2(n26703), .B1(n26570), 
        .B2(n13793), .Y(n15197) );
  sky130_fd_sc_hd__nand2_1 U22322 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[182]), .Y(n15139) );
  sky130_fd_sc_hd__nand2_1 U22323 ( .A(n15982), .B(
        j202_soc_core_j22_cpu_rf_gpr[246]), .Y(n15138) );
  sky130_fd_sc_hd__nand2_1 U22324 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[502]), .Y(n15137) );
  sky130_fd_sc_hd__nand2_1 U22325 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[438]), .Y(n15136) );
  sky130_fd_sc_hd__nand4_1 U22326 ( .A(n15139), .B(n15138), .C(n15137), .D(
        n15136), .Y(n15145) );
  sky130_fd_sc_hd__nand2_1 U22327 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[22]), .Y(n15143) );
  sky130_fd_sc_hd__nand2_1 U22328 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[54]), .Y(n15142) );
  sky130_fd_sc_hd__nand2_1 U22329 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[118]), .Y(n15141) );
  sky130_fd_sc_hd__nand2_1 U22330 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[406]), .Y(n15140) );
  sky130_fd_sc_hd__nand4_1 U22331 ( .A(n15143), .B(n15142), .C(n15141), .D(
        n15140), .Y(n15144) );
  sky130_fd_sc_hd__nor2_1 U22332 ( .A(n15145), .B(n15144), .Y(n15153) );
  sky130_fd_sc_hd__a22oi_1 U22333 ( .A1(n11160), .A2(
        j202_soc_core_j22_cpu_rf_gpr[310]), .B1(n23502), .B2(
        j202_soc_core_j22_cpu_rf_gpr[470]), .Y(n15152) );
  sky130_fd_sc_hd__a22oi_1 U22334 ( .A1(n16470), .A2(
        j202_soc_core_j22_cpu_rf_gpr[214]), .B1(n16469), .B2(
        j202_soc_core_j22_cpu_rf_gpr[86]), .Y(n15151) );
  sky130_fd_sc_hd__nand2_1 U22335 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[278]), .Y(n15149) );
  sky130_fd_sc_hd__nand2_1 U22336 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[150]), .Y(n15148) );
  sky130_fd_sc_hd__nand2_1 U22337 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[374]), .Y(n15147) );
  sky130_fd_sc_hd__nand2_1 U22338 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[342]), .Y(n15146) );
  sky130_fd_sc_hd__and4_1 U22339 ( .A(n15149), .B(n15148), .C(n15147), .D(
        n15146), .X(n15150) );
  sky130_fd_sc_hd__nand4_1 U22340 ( .A(n15153), .B(n15152), .C(n15151), .D(
        n15150), .Y(n22345) );
  sky130_fd_sc_hd__nand2_1 U22341 ( .A(n22345), .B(n16513), .Y(n15162) );
  sky130_fd_sc_hd__nand2_1 U22342 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[22]), .Y(n15156) );
  sky130_fd_sc_hd__nand2_1 U22343 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[22]), .Y(n15155) );
  sky130_fd_sc_hd__nand2_1 U22344 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[502]), .Y(n15154) );
  sky130_fd_sc_hd__and4_1 U22345 ( .A(n15156), .B(n15155), .C(n16516), .D(
        n15154), .X(n15161) );
  sky130_fd_sc_hd__nand2_1 U22346 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[22]), .Y(n15160) );
  sky130_fd_sc_hd__nand2_1 U22347 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[22]), .Y(n15159) );
  sky130_fd_sc_hd__nand2_1 U22348 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[22]), .Y(n15158) );
  sky130_fd_sc_hd__nand2_1 U22349 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[22]), .Y(n15157) );
  sky130_fd_sc_hd__nand3_1 U22350 ( .A(n15162), .B(n15161), .C(n13325), .Y(
        n27405) );
  sky130_fd_sc_hd__nand2_1 U22351 ( .A(n27405), .B(n16529), .Y(n15163) );
  sky130_fd_sc_hd__nor2_1 U22353 ( .A(n15197), .B(n15198), .Y(n15418) );
  sky130_fd_sc_hd__o22ai_1 U22354 ( .A1(n16492), .A2(n26570), .B1(n26417), 
        .B2(n13793), .Y(n15195) );
  sky130_fd_sc_hd__nand2_1 U22355 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[181]), .Y(n15168) );
  sky130_fd_sc_hd__nand2_1 U22356 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[245]), .Y(n15167) );
  sky130_fd_sc_hd__nand2_1 U22357 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[501]), .Y(n15166) );
  sky130_fd_sc_hd__nand2_1 U22358 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[437]), .Y(n15165) );
  sky130_fd_sc_hd__nand4_1 U22359 ( .A(n15168), .B(n15167), .C(n15166), .D(
        n15165), .Y(n15174) );
  sky130_fd_sc_hd__nand2_1 U22360 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[21]), .Y(n15172) );
  sky130_fd_sc_hd__nand2_1 U22361 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[53]), .Y(n15171) );
  sky130_fd_sc_hd__nand2_1 U22362 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[117]), .Y(n15170) );
  sky130_fd_sc_hd__nand2_1 U22363 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[405]), .Y(n15169) );
  sky130_fd_sc_hd__nand4_1 U22364 ( .A(n15172), .B(n15171), .C(n15170), .D(
        n15169), .Y(n15173) );
  sky130_fd_sc_hd__nor2_1 U22365 ( .A(n15174), .B(n15173), .Y(n15182) );
  sky130_fd_sc_hd__a22oi_1 U22366 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[309]), .B1(n14414), .B2(
        j202_soc_core_j22_cpu_rf_gpr[469]), .Y(n15181) );
  sky130_fd_sc_hd__a22oi_1 U22367 ( .A1(n16470), .A2(
        j202_soc_core_j22_cpu_rf_gpr[213]), .B1(n23089), .B2(
        j202_soc_core_j22_cpu_rf_gpr[85]), .Y(n15180) );
  sky130_fd_sc_hd__nand2_1 U22368 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[277]), .Y(n15178) );
  sky130_fd_sc_hd__nand2_1 U22369 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[149]), .Y(n15177) );
  sky130_fd_sc_hd__nand2_1 U22370 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[373]), .Y(n15176) );
  sky130_fd_sc_hd__nand2_1 U22371 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[341]), .Y(n15175) );
  sky130_fd_sc_hd__and4_1 U22372 ( .A(n15178), .B(n15177), .C(n15176), .D(
        n15175), .X(n15179) );
  sky130_fd_sc_hd__nand4_1 U22373 ( .A(n15182), .B(n15181), .C(n15180), .D(
        n15179), .Y(n22121) );
  sky130_fd_sc_hd__nand2_1 U22374 ( .A(n22121), .B(n16513), .Y(n15191) );
  sky130_fd_sc_hd__nand2_1 U22375 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[21]), .Y(n15185) );
  sky130_fd_sc_hd__nand2_1 U22376 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[21]), .Y(n15184) );
  sky130_fd_sc_hd__nand2_1 U22377 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[501]), .Y(n15183) );
  sky130_fd_sc_hd__and4_1 U22378 ( .A(n15185), .B(n15184), .C(n16516), .D(
        n15183), .X(n15190) );
  sky130_fd_sc_hd__nand2_1 U22379 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[21]), .Y(n15189) );
  sky130_fd_sc_hd__nand2_1 U22380 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[21]), .Y(n15188) );
  sky130_fd_sc_hd__nand2_1 U22381 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[21]), .Y(n15187) );
  sky130_fd_sc_hd__nand2_1 U22382 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[21]), .Y(n15186) );
  sky130_fd_sc_hd__nand3_1 U22383 ( .A(n15191), .B(n15190), .C(n13337), .Y(
        n27412) );
  sky130_fd_sc_hd__nand2_1 U22384 ( .A(n27412), .B(n16529), .Y(n15192) );
  sky130_fd_sc_hd__nor2_1 U22386 ( .A(n15195), .B(n15196), .Y(n15663) );
  sky130_fd_sc_hd__nor2_1 U22387 ( .A(n15418), .B(n15663), .Y(n15200) );
  sky130_fd_sc_hd__nand2_1 U22388 ( .A(n15415), .B(n15200), .Y(n15202) );
  sky130_fd_sc_hd__nor2_1 U22389 ( .A(n15202), .B(n15412), .Y(n16533) );
  sky130_fd_sc_hd__nor2_1 U22390 ( .A(n15899), .B(n17108), .Y(n15206) );
  sky130_fd_sc_hd__nand2_1 U22392 ( .A(n15196), .B(n15195), .Y(n15664) );
  sky130_fd_sc_hd__nand2_1 U22393 ( .A(n15198), .B(n15197), .Y(n15419) );
  sky130_fd_sc_hd__a21oi_1 U22395 ( .A1(n15200), .A2(n15414), .B1(n15199), .Y(
        n15201) );
  sky130_fd_sc_hd__o21ai_2 U22396 ( .A1(n15202), .A2(n15413), .B1(n15201), .Y(
        n16554) );
  sky130_fd_sc_hd__inv_2 U22397 ( .A(n16554), .Y(n17110) );
  sky130_fd_sc_hd__nand2_1 U22398 ( .A(n15204), .B(n15203), .Y(n15953) );
  sky130_fd_sc_hd__a21oi_1 U22400 ( .A1(n22513), .A2(n15206), .B1(n15205), .Y(
        n15212) );
  sky130_fd_sc_hd__o22ai_1 U22401 ( .A1(n16492), .A2(n26701), .B1(n26704), 
        .B2(n13793), .Y(n15208) );
  sky130_fd_sc_hd__nand2_1 U22402 ( .A(n27392), .B(n16529), .Y(n15207) );
  sky130_fd_sc_hd__o21ai_1 U22403 ( .A1(n14742), .A2(n27392), .B1(n15207), .Y(
        n15209) );
  sky130_fd_sc_hd__nor2_1 U22404 ( .A(n15208), .B(n15209), .Y(n15952) );
  sky130_fd_sc_hd__nand2_1 U22405 ( .A(n15209), .B(n15208), .Y(n15951) );
  sky130_fd_sc_hd__nand2_1 U22406 ( .A(n15210), .B(n15951), .Y(n15211) );
  sky130_fd_sc_hd__xor2_1 U22407 ( .A(n15212), .B(n15211), .X(n23831) );
  sky130_fd_sc_hd__nand2_1 U22408 ( .A(n23831), .B(n12158), .Y(n15213) );
  sky130_fd_sc_hd__nand2_1 U22409 ( .A(j202_soc_core_memory0_ram_dout0[55]), 
        .B(n21604), .Y(n15218) );
  sky130_fd_sc_hd__nand2_1 U22410 ( .A(j202_soc_core_memory0_ram_dout0[375]), 
        .B(n21596), .Y(n15217) );
  sky130_fd_sc_hd__nand2_1 U22411 ( .A(j202_soc_core_memory0_ram_dout0[439]), 
        .B(n21598), .Y(n15216) );
  sky130_fd_sc_hd__nand2_1 U22412 ( .A(j202_soc_core_memory0_ram_dout0[407]), 
        .B(n21597), .Y(n15215) );
  sky130_fd_sc_hd__nand4_1 U22413 ( .A(n15218), .B(n15217), .C(n15216), .D(
        n15215), .Y(n15219) );
  sky130_fd_sc_hd__nand2_1 U22414 ( .A(j202_soc_core_memory0_ram_dout0[215]), 
        .B(n21732), .Y(n15275) );
  sky130_fd_sc_hd__nand3_1 U22415 ( .A(n15363), .B(n15381), .C(n15615), .Y(
        n15224) );
  sky130_fd_sc_hd__nor2_1 U22416 ( .A(n15581), .B(n15369), .Y(n15223) );
  sky130_fd_sc_hd__nand3_1 U22417 ( .A(n15223), .B(n15222), .C(n15221), .Y(
        n15547) );
  sky130_fd_sc_hd__nand4_1 U22419 ( .A(n15532), .B(n15359), .C(n15545), .D(
        n15560), .Y(n15225) );
  sky130_fd_sc_hd__nand2_1 U22420 ( .A(n15225), .B(n17163), .Y(n15337) );
  sky130_fd_sc_hd__nand3_1 U22421 ( .A(n15228), .B(n15227), .C(n15313), .Y(
        n15230) );
  sky130_fd_sc_hd__a21oi_1 U22422 ( .A1(n15609), .A2(n16953), .B1(n15708), .Y(
        n15229) );
  sky130_fd_sc_hd__a21oi_1 U22423 ( .A1(n15230), .A2(n16090), .B1(n15229), .Y(
        n15232) );
  sky130_fd_sc_hd__nand4_1 U22424 ( .A(n15233), .B(n15337), .C(n15232), .D(
        n15231), .Y(n15234) );
  sky130_fd_sc_hd__nand2_1 U22425 ( .A(n15234), .B(n13481), .Y(n15291) );
  sky130_fd_sc_hd__nand2_1 U22426 ( .A(n21675), .B(j202_soc_core_uart_div1[7]), 
        .Y(n15285) );
  sky130_fd_sc_hd__nand2_1 U22427 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[23]), .Y(n15284) );
  sky130_fd_sc_hd__nand3_1 U22428 ( .A(n15285), .B(n21677), .C(n15284), .Y(
        n15237) );
  sky130_fd_sc_hd__nand2_1 U22429 ( .A(n21699), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[55]), .Y(n15236) );
  sky130_fd_sc_hd__nand2_1 U22430 ( .A(n21666), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[87]), .Y(n15235) );
  sky130_fd_sc_hd__nand2_1 U22431 ( .A(n15236), .B(n15235), .Y(n15286) );
  sky130_fd_sc_hd__nor2_1 U22432 ( .A(n15237), .B(n15286), .Y(n15250) );
  sky130_fd_sc_hd__nand2_1 U22433 ( .A(n15340), .B(n15589), .Y(n15238) );
  sky130_fd_sc_hd__o21ai_1 U22434 ( .A1(n15238), .A2(n15383), .B1(n16090), .Y(
        n15247) );
  sky130_fd_sc_hd__nand2_1 U22435 ( .A(n17302), .B(n16163), .Y(n15239) );
  sky130_fd_sc_hd__nand2b_1 U22436 ( .A_N(n20804), .B(n19380), .Y(n18952) );
  sky130_fd_sc_hd__nand3_1 U22437 ( .A(n15533), .B(n15239), .C(n18952), .Y(
        n15240) );
  sky130_fd_sc_hd__o21ai_1 U22438 ( .A1(n15625), .A2(n15240), .B1(n17163), .Y(
        n15246) );
  sky130_fd_sc_hd__nand3_1 U22439 ( .A(n15593), .B(n15586), .C(n15589), .Y(
        n15241) );
  sky130_fd_sc_hd__nand2_1 U22440 ( .A(n15341), .B(n15558), .Y(n15320) );
  sky130_fd_sc_hd__o21ai_1 U22441 ( .A1(n15241), .A2(n15320), .B1(n15630), .Y(
        n15245) );
  sky130_fd_sc_hd__nand2_1 U22442 ( .A(n15535), .B(n15242), .Y(n15556) );
  sky130_fd_sc_hd__nand4_1 U22444 ( .A(n15247), .B(n15246), .C(n15245), .D(
        n15244), .Y(n15248) );
  sky130_fd_sc_hd__nand2_1 U22445 ( .A(n15248), .B(n20908), .Y(n15289) );
  sky130_fd_sc_hd__nand2_1 U22446 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_duty[11]), .Y(n15288) );
  sky130_fd_sc_hd__nand4_1 U22447 ( .A(n15291), .B(n15250), .C(n15289), .D(
        n15288), .Y(n15265) );
  sky130_fd_sc_hd__nand2_1 U22448 ( .A(n15251), .B(n15545), .Y(n15379) );
  sky130_fd_sc_hd__nand3_1 U22449 ( .A(n15594), .B(n15537), .C(n16722), .Y(
        n15252) );
  sky130_fd_sc_hd__nor3_1 U22450 ( .A(n15253), .B(n15379), .C(n15252), .Y(
        n15263) );
  sky130_fd_sc_hd__nand4_1 U22451 ( .A(n15255), .B(n15592), .C(n15534), .D(
        n15593), .Y(n15261) );
  sky130_fd_sc_hd__nand2_1 U22452 ( .A(n15256), .B(n15614), .Y(n15361) );
  sky130_fd_sc_hd__nand3_1 U22453 ( .A(n15533), .B(n15586), .C(n15614), .Y(
        n15257) );
  sky130_fd_sc_hd__nand2_1 U22454 ( .A(n15380), .B(n15359), .Y(n15317) );
  sky130_fd_sc_hd__nor2_1 U22455 ( .A(n15257), .B(n15317), .Y(n15583) );
  sky130_fd_sc_hd__nor2_1 U22456 ( .A(n15570), .B(n15258), .Y(n15590) );
  sky130_fd_sc_hd__nand3_1 U22457 ( .A(n15583), .B(n15590), .C(n15564), .Y(
        n15259) );
  sky130_fd_sc_hd__a21oi_1 U22458 ( .A1(n15261), .A2(n15630), .B1(n15260), .Y(
        n15262) );
  sky130_fd_sc_hd__o21a_1 U22459 ( .A1(n15384), .A2(n15263), .B1(n15262), .X(
        n15264) );
  sky130_fd_sc_hd__nor2_1 U22460 ( .A(n19856), .B(n15264), .Y(n15292) );
  sky130_fd_sc_hd__nor2_1 U22461 ( .A(n15265), .B(n15292), .Y(n15274) );
  sky130_fd_sc_hd__nand2_1 U22462 ( .A(n15381), .B(n15564), .Y(n15571) );
  sky130_fd_sc_hd__nor2_1 U22463 ( .A(n15266), .B(n15571), .Y(n15629) );
  sky130_fd_sc_hd__nor2_1 U22464 ( .A(n15347), .B(n15365), .Y(n15267) );
  sky130_fd_sc_hd__nand4_1 U22465 ( .A(n15324), .B(n15267), .C(n15564), .D(
        n15537), .Y(n15269) );
  sky130_fd_sc_hd__a31oi_1 U22466 ( .A1(n15380), .A2(n15564), .A3(n15558), 
        .B1(n15557), .Y(n15268) );
  sky130_fd_sc_hd__a21oi_1 U22467 ( .A1(n15269), .A2(n17163), .B1(n15268), .Y(
        n15272) );
  sky130_fd_sc_hd__nand2_1 U22468 ( .A(n15612), .B(n15537), .Y(n15360) );
  sky130_fd_sc_hd__nand2b_1 U22469 ( .A_N(n15366), .B(n15350), .Y(n15587) );
  sky130_fd_sc_hd__nor4_1 U22470 ( .A(n15347), .B(n15568), .C(n15360), .D(
        n15587), .Y(n15270) );
  sky130_fd_sc_hd__nand2b_1 U22471 ( .A_N(n15270), .B(n15584), .Y(n15271) );
  sky130_fd_sc_hd__o211ai_1 U22472 ( .A1(n15629), .A2(n15384), .B1(n15272), 
        .C1(n15271), .Y(n15273) );
  sky130_fd_sc_hd__nand2_1 U22473 ( .A(n15273), .B(n21697), .Y(n15294) );
  sky130_fd_sc_hd__nand2_1 U22474 ( .A(j202_soc_core_memory0_ram_dout0[343]), 
        .B(n21593), .Y(n15277) );
  sky130_fd_sc_hd__nand2_1 U22475 ( .A(j202_soc_core_memory0_ram_dout0[183]), 
        .B(n21590), .Y(n15276) );
  sky130_fd_sc_hd__nand2_1 U22476 ( .A(n15277), .B(n15276), .Y(n15278) );
  sky130_fd_sc_hd__nand2_1 U22477 ( .A(j202_soc_core_memory0_ram_dout0[87]), 
        .B(n21734), .Y(n15283) );
  sky130_fd_sc_hd__nand2_1 U22478 ( .A(j202_soc_core_memory0_ram_dout0[151]), 
        .B(n21592), .Y(n15282) );
  sky130_fd_sc_hd__nand2_1 U22479 ( .A(j202_soc_core_memory0_ram_dout0[119]), 
        .B(n21591), .Y(n15281) );
  sky130_fd_sc_hd__nand2_1 U22480 ( .A(j202_soc_core_memory0_ram_dout0[23]), 
        .B(n21733), .Y(n15280) );
  sky130_fd_sc_hd__nand2_1 U22481 ( .A(j202_soc_core_memory0_ram_dout0[503]), 
        .B(n21771), .Y(n15296) );
  sky130_fd_sc_hd__nand3_1 U22482 ( .A(n15285), .B(n21738), .C(n15284), .Y(
        n15287) );
  sky130_fd_sc_hd__nor2_1 U22483 ( .A(n15287), .B(n15286), .Y(n15290) );
  sky130_fd_sc_hd__nand4_1 U22484 ( .A(n15291), .B(n15290), .C(n15289), .D(
        n15288), .Y(n15293) );
  sky130_fd_sc_hd__nor2_1 U22485 ( .A(n15293), .B(n15292), .Y(n15295) );
  sky130_fd_sc_hd__nand3_1 U22486 ( .A(n15296), .B(n15295), .C(n15294), .Y(
        n18921) );
  sky130_fd_sc_hd__nor2_1 U22487 ( .A(n15298), .B(n21009), .Y(n15407) );
  sky130_fd_sc_hd__nor2_1 U22488 ( .A(n15299), .B(n15656), .Y(n15300) );
  sky130_fd_sc_hd__xnor2_1 U22489 ( .A(n15301), .B(n15300), .Y(n26069) );
  sky130_fd_sc_hd__nand2_1 U22490 ( .A(n22596), .B(n26069), .Y(n15303) );
  sky130_fd_sc_hd__nand2_1 U22491 ( .A(n22515), .B(n27399), .Y(n15302) );
  sky130_fd_sc_hd__a21oi_1 U22492 ( .A1(n22513), .A2(n16533), .B1(n16554), .Y(
        n15305) );
  sky130_fd_sc_hd__nand2_1 U22493 ( .A(n25176), .B(n12158), .Y(n15306) );
  sky130_fd_sc_hd__nand2_1 U22494 ( .A(j202_soc_core_memory0_ram_dout0[182]), 
        .B(n21590), .Y(n15307) );
  sky130_fd_sc_hd__nand2_1 U22495 ( .A(j202_soc_core_memory0_ram_dout0[470]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n15391) );
  sky130_fd_sc_hd__nand2_1 U22496 ( .A(j202_soc_core_memory0_ram_dout0[438]), 
        .B(n21598), .Y(n15390) );
  sky130_fd_sc_hd__nand2_1 U22497 ( .A(j202_soc_core_memory0_ram_dout0[374]), 
        .B(n21596), .Y(n15389) );
  sky130_fd_sc_hd__a22oi_1 U22498 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[54]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[86]), .Y(n15398) );
  sky130_fd_sc_hd__nand2_1 U22499 ( .A(n21675), .B(j202_soc_core_uart_div1[6]), 
        .Y(n15397) );
  sky130_fd_sc_hd__nand2_1 U22500 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[22]), .Y(n15396) );
  sky130_fd_sc_hd__nand4_1 U22501 ( .A(n15398), .B(n21677), .C(n15397), .D(
        n15396), .Y(n15358) );
  sky130_fd_sc_hd__nand2_1 U22502 ( .A(n15309), .B(n15308), .Y(n15322) );
  sky130_fd_sc_hd__nand2_1 U22503 ( .A(n15340), .B(n15322), .Y(n15311) );
  sky130_fd_sc_hd__nor3_1 U22504 ( .A(n15311), .B(n15365), .C(n15310), .Y(
        n15312) );
  sky130_fd_sc_hd__nand4_1 U22505 ( .A(n15314), .B(n15313), .C(n15312), .D(
        n15560), .Y(n15315) );
  sky130_fd_sc_hd__nand2_1 U22506 ( .A(n15315), .B(n15584), .Y(n15329) );
  sky130_fd_sc_hd__nand2_1 U22507 ( .A(n15316), .B(n16090), .Y(n15328) );
  sky130_fd_sc_hd__nor2_1 U22508 ( .A(n17277), .B(
        j202_soc_core_bootrom_00_address_w[11]), .Y(n19124) );
  sky130_fd_sc_hd__nor4_1 U22509 ( .A(n21207), .B(n15319), .C(n15318), .D(
        n15317), .Y(n15326) );
  sky130_fd_sc_hd__nor2_1 U22510 ( .A(n15321), .B(n15320), .Y(n15345) );
  sky130_fd_sc_hd__nand2_1 U22511 ( .A(n15614), .B(n15322), .Y(n15562) );
  sky130_fd_sc_hd__nor4bb_1 U22512 ( .C_N(n15324), .D_N(n15345), .A(n15323), 
        .B(n15562), .Y(n15325) );
  sky130_fd_sc_hd__nand3_1 U22513 ( .A(n15329), .B(n15328), .C(n15327), .Y(
        n15339) );
  sky130_fd_sc_hd__nor2_1 U22515 ( .A(n15333), .B(n15332), .Y(n15334) );
  sky130_fd_sc_hd__a21oi_1 U22516 ( .A1(n15590), .A2(n15334), .B1(n15384), .Y(
        n15543) );
  sky130_fd_sc_hd__a21oi_1 U22517 ( .A1(n15630), .A2(n15539), .B1(n15543), .Y(
        n15335) );
  sky130_fd_sc_hd__nand3_1 U22518 ( .A(n15337), .B(n15336), .C(n15335), .Y(
        n15338) );
  sky130_fd_sc_hd__a22oi_1 U22519 ( .A1(n15339), .A2(n21697), .B1(n15338), 
        .B2(n13481), .Y(n15401) );
  sky130_fd_sc_hd__nand2_1 U22520 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_duty[10]), .Y(n15400) );
  sky130_fd_sc_hd__nand4_1 U22521 ( .A(n15583), .B(n15342), .C(n15531), .D(
        n15341), .Y(n15343) );
  sky130_fd_sc_hd__nand2_1 U22522 ( .A(n15343), .B(n15584), .Y(n15356) );
  sky130_fd_sc_hd__nand2_1 U22523 ( .A(n15345), .B(n15344), .Y(n15346) );
  sky130_fd_sc_hd__nand2_1 U22524 ( .A(n15346), .B(n15630), .Y(n15355) );
  sky130_fd_sc_hd__nand3_1 U22525 ( .A(n15348), .B(n15577), .C(n16953), .Y(
        n15349) );
  sky130_fd_sc_hd__o21ai_1 U22526 ( .A1(n15349), .A2(n15383), .B1(n17163), .Y(
        n15354) );
  sky130_fd_sc_hd__nand3_1 U22527 ( .A(n15350), .B(n12192), .C(n15533), .Y(
        n15352) );
  sky130_fd_sc_hd__nand4_1 U22529 ( .A(n15356), .B(n15355), .C(n15354), .D(
        n15353), .Y(n15357) );
  sky130_fd_sc_hd__nand2_1 U22530 ( .A(n15357), .B(n21727), .Y(n15399) );
  sky130_fd_sc_hd__nand4b_1 U22531 ( .A_N(n15358), .B(n15401), .C(n15400), .D(
        n15399), .Y(n15387) );
  sky130_fd_sc_hd__nand2_1 U22532 ( .A(n15578), .B(n15359), .Y(n15606) );
  sky130_fd_sc_hd__nor3_1 U22533 ( .A(n15361), .B(n15360), .C(n15606), .Y(
        n15602) );
  sky130_fd_sc_hd__nand4_1 U22534 ( .A(n15602), .B(n15380), .C(n15545), .D(
        n15589), .Y(n15362) );
  sky130_fd_sc_hd__nand2_1 U22535 ( .A(n15362), .B(n15630), .Y(n15378) );
  sky130_fd_sc_hd__nand3_1 U22536 ( .A(n15364), .B(n15363), .C(n15535), .Y(
        n15374) );
  sky130_fd_sc_hd__nand2b_1 U22537 ( .A_N(n15365), .B(n15577), .Y(n15572) );
  sky130_fd_sc_hd__nand3_1 U22538 ( .A(n15601), .B(n15368), .C(n15367), .Y(
        n15607) );
  sky130_fd_sc_hd__nor3_1 U22539 ( .A(n15369), .B(n15572), .C(n15607), .Y(
        n15370) );
  sky130_fd_sc_hd__nand2_1 U22540 ( .A(n15619), .B(n15370), .Y(n15372) );
  sky130_fd_sc_hd__a21oi_1 U22541 ( .A1(n15551), .A2(n15586), .B1(n15384), .Y(
        n15371) );
  sky130_fd_sc_hd__a21oi_1 U22542 ( .A1(n15372), .A2(n17163), .B1(n15371), .Y(
        n15377) );
  sky130_fd_sc_hd__nand2_1 U22543 ( .A(n15373), .B(n15613), .Y(n15375) );
  sky130_fd_sc_hd__o21ai_1 U22544 ( .A1(n15375), .A2(n15374), .B1(n15584), .Y(
        n15376) );
  sky130_fd_sc_hd__nand3_1 U22545 ( .A(n15378), .B(n15377), .C(n15376), .Y(
        n15386) );
  sky130_fd_sc_hd__nor2_1 U22546 ( .A(n15608), .B(n15379), .Y(n15628) );
  sky130_fd_sc_hd__nand4_1 U22547 ( .A(n15381), .B(n15380), .C(n15613), .D(
        n15612), .Y(n15382) );
  sky130_fd_sc_hd__nor2_1 U22548 ( .A(n15383), .B(n15382), .Y(n15385) );
  sky130_fd_sc_hd__a21oi_1 U22549 ( .A1(n15628), .A2(n15385), .B1(n15384), .Y(
        n15620) );
  sky130_fd_sc_hd__o21a_1 U22550 ( .A1(n15386), .A2(n15620), .B1(n20908), .X(
        n15403) );
  sky130_fd_sc_hd__nor2_1 U22551 ( .A(n15387), .B(n15403), .Y(n15388) );
  sky130_fd_sc_hd__nand2_1 U22552 ( .A(j202_soc_core_memory0_ram_dout0[278]), 
        .B(n21605), .Y(n15395) );
  sky130_fd_sc_hd__nand2_1 U22553 ( .A(j202_soc_core_memory0_ram_dout0[406]), 
        .B(n21597), .Y(n15394) );
  sky130_fd_sc_hd__nand2_1 U22554 ( .A(j202_soc_core_memory0_ram_dout0[342]), 
        .B(n21593), .Y(n15393) );
  sky130_fd_sc_hd__nand2_1 U22555 ( .A(j202_soc_core_memory0_ram_dout0[246]), 
        .B(n21735), .Y(n15392) );
  sky130_fd_sc_hd__nand2_1 U22556 ( .A(j202_soc_core_memory0_ram_dout0[502]), 
        .B(n21771), .Y(n15406) );
  sky130_fd_sc_hd__nand4_1 U22557 ( .A(n15398), .B(n21738), .C(n15397), .D(
        n15396), .Y(n15402) );
  sky130_fd_sc_hd__nand4b_1 U22558 ( .A_N(n15402), .B(n15401), .C(n15400), .D(
        n15399), .Y(n15404) );
  sky130_fd_sc_hd__nor2_1 U22559 ( .A(n15404), .B(n15403), .Y(n15405) );
  sky130_fd_sc_hd__nand2_1 U22560 ( .A(n15406), .B(n15405), .Y(n20832) );
  sky130_fd_sc_hd__nand2_1 U22561 ( .A(n15407), .B(
        j202_soc_core_j22_cpu_pc[21]), .Y(n15409) );
  sky130_fd_sc_hd__xor2_1 U22562 ( .A(n15409), .B(n15408), .X(n26111) );
  sky130_fd_sc_hd__nand2_1 U22563 ( .A(n22596), .B(n26111), .Y(n15411) );
  sky130_fd_sc_hd__nand2_1 U22564 ( .A(n22515), .B(n27405), .Y(n15410) );
  sky130_fd_sc_hd__nand2_1 U22565 ( .A(n15771), .B(n15415), .Y(n15659) );
  sky130_fd_sc_hd__nor2_1 U22566 ( .A(n15663), .B(n15659), .Y(n15417) );
  sky130_fd_sc_hd__a21oi_1 U22567 ( .A1(n15770), .A2(n15415), .B1(n15414), .Y(
        n15660) );
  sky130_fd_sc_hd__a22oi_1 U22568 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[50]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[82]), .Y(n15503) );
  sky130_fd_sc_hd__nand2_1 U22569 ( .A(n21675), .B(j202_soc_core_uart_div1[2]), 
        .Y(n15498) );
  sky130_fd_sc_hd__nand2_1 U22570 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[18]), .Y(n15497) );
  sky130_fd_sc_hd__nand4_1 U22571 ( .A(n15503), .B(n21677), .C(n15498), .D(
        n15497), .Y(n15495) );
  sky130_fd_sc_hd__nand2_1 U22572 ( .A(n16171), .B(n19381), .Y(n15438) );
  sky130_fd_sc_hd__nand2_1 U22573 ( .A(n15454), .B(n20787), .Y(n15673) );
  sky130_fd_sc_hd__nand2_1 U22574 ( .A(n15422), .B(n17289), .Y(n15467) );
  sky130_fd_sc_hd__nor2_1 U22575 ( .A(n15438), .B(n15467), .Y(n20606) );
  sky130_fd_sc_hd__nand2_1 U22576 ( .A(n15424), .B(n19354), .Y(n16583) );
  sky130_fd_sc_hd__nor2_1 U22577 ( .A(n16170), .B(n16583), .Y(n20437) );
  sky130_fd_sc_hd__nand2_1 U22578 ( .A(n20437), .B(n15454), .Y(n20669) );
  sky130_fd_sc_hd__nor2_1 U22579 ( .A(j202_soc_core_bootrom_00_address_w[11]), 
        .B(n15454), .Y(n15725) );
  sky130_fd_sc_hd__nand3_1 U22580 ( .A(n15725), .B(n15425), .C(n16171), .Y(
        n20648) );
  sky130_fd_sc_hd__nor2_1 U22581 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .B(n16162), .Y(n20632) );
  sky130_fd_sc_hd__nor3_1 U22582 ( .A(n15705), .B(n15695), .C(n15437), .Y(
        n20479) );
  sky130_fd_sc_hd__nor2_1 U22583 ( .A(n20606), .B(n20678), .Y(n20453) );
  sky130_fd_sc_hd__nand2_1 U22584 ( .A(n20437), .B(
        j202_soc_core_bootrom_00_address_w[9]), .Y(n20582) );
  sky130_fd_sc_hd__nand2_1 U22585 ( .A(n16616), .B(n17274), .Y(n15449) );
  sky130_fd_sc_hd__nor2_1 U22586 ( .A(n15454), .B(n16845), .Y(n15428) );
  sky130_fd_sc_hd__nor2_1 U22587 ( .A(n15449), .B(n15426), .Y(n15741) );
  sky130_fd_sc_hd__nor2_1 U22588 ( .A(n20521), .B(n15741), .Y(n20450) );
  sky130_fd_sc_hd__nor2_1 U22590 ( .A(n15454), .B(n16953), .Y(n20668) );
  sky130_fd_sc_hd__nand2_1 U22591 ( .A(n16171), .B(n17274), .Y(n15431) );
  sky130_fd_sc_hd__nand2_1 U22592 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .B(n13293), .Y(n15427) );
  sky130_fd_sc_hd__nor2_1 U22593 ( .A(n15431), .B(n15427), .Y(n15671) );
  sky130_fd_sc_hd__nor2_1 U22594 ( .A(n15454), .B(n16583), .Y(n15451) );
  sky130_fd_sc_hd__nand2_1 U22595 ( .A(n11994), .B(n17277), .Y(n16159) );
  sky130_fd_sc_hd__nand2_1 U22596 ( .A(n15451), .B(n17161), .Y(n20643) );
  sky130_fd_sc_hd__nand3_1 U22597 ( .A(n16706), .B(n15725), .C(n15458), .Y(
        n20568) );
  sky130_fd_sc_hd__nand2_1 U22598 ( .A(n20643), .B(n20568), .Y(n15720) );
  sky130_fd_sc_hd__nor2_1 U22599 ( .A(n15671), .B(n15720), .Y(n20472) );
  sky130_fd_sc_hd__nand2_1 U22600 ( .A(n15429), .B(n15428), .Y(n20664) );
  sky130_fd_sc_hd__nand2_1 U22601 ( .A(n20472), .B(n20664), .Y(n20466) );
  sky130_fd_sc_hd__nand3_1 U22602 ( .A(n16706), .B(n16616), .C(n15725), .Y(
        n20570) );
  sky130_fd_sc_hd__nand2_1 U22603 ( .A(n13293), .B(n15454), .Y(n15450) );
  sky130_fd_sc_hd__nand2_1 U22604 ( .A(n17161), .B(n17274), .Y(n15434) );
  sky130_fd_sc_hd__nor2_1 U22605 ( .A(n15450), .B(n15434), .Y(n15689) );
  sky130_fd_sc_hd__nor2_1 U22606 ( .A(n20676), .B(n15689), .Y(n20653) );
  sky130_fd_sc_hd__nor4_1 U22607 ( .A(n15716), .B(n20668), .C(n20466), .D(
        n15735), .Y(n15430) );
  sky130_fd_sc_hd__nand2_1 U22608 ( .A(n12137), .B(n20788), .Y(n20681) );
  sky130_fd_sc_hd__a31oi_1 U22609 ( .A1(n20453), .A2(n20450), .A3(n15430), 
        .B1(n20681), .Y(n15446) );
  sky130_fd_sc_hd__nor2_1 U22610 ( .A(n15431), .B(n15450), .Y(n20499) );
  sky130_fd_sc_hd__nor2_1 U22611 ( .A(n20499), .B(n15716), .Y(n15670) );
  sky130_fd_sc_hd__nand2_1 U22612 ( .A(n16616), .B(n19381), .Y(n15703) );
  sky130_fd_sc_hd__nor2_1 U22613 ( .A(n15703), .B(n15467), .Y(n20667) );
  sky130_fd_sc_hd__nor2_1 U22614 ( .A(n20787), .B(n16159), .Y(n17167) );
  sky130_fd_sc_hd__nor3_1 U22615 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .B(n15432), .C(n17164), .Y(n15441) );
  sky130_fd_sc_hd__nand2_1 U22616 ( .A(n15724), .B(n15469), .Y(n15483) );
  sky130_fd_sc_hd__nor4_1 U22617 ( .A(n15741), .B(n20667), .C(n15441), .D(
        n15483), .Y(n15433) );
  sky130_fd_sc_hd__nand2_1 U22618 ( .A(n17175), .B(n20579), .Y(n20651) );
  sky130_fd_sc_hd__a21oi_1 U22619 ( .A1(n15670), .A2(n15433), .B1(n20651), .Y(
        n15445) );
  sky130_fd_sc_hd__nand3_1 U22620 ( .A(n16171), .B(n16706), .C(n15725), .Y(
        n20442) );
  sky130_fd_sc_hd__nor2_1 U22621 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .B(n16845), .Y(n15704) );
  sky130_fd_sc_hd__nor2_1 U22622 ( .A(n15434), .B(n15439), .Y(n20477) );
  sky130_fd_sc_hd__nor2_1 U22623 ( .A(n15716), .B(n20477), .Y(n20672) );
  sky130_fd_sc_hd__nand2_1 U22624 ( .A(n20442), .B(n20672), .Y(n20659) );
  sky130_fd_sc_hd__nand2b_1 U22625 ( .A_N(n20633), .B(n15454), .Y(n15723) );
  sky130_fd_sc_hd__nand2_1 U22626 ( .A(n15723), .B(n20568), .Y(n20495) );
  sky130_fd_sc_hd__nand2_1 U22627 ( .A(n20669), .B(n15738), .Y(n15435) );
  sky130_fd_sc_hd__or4_1 U22628 ( .A(n20499), .B(n20448), .C(n20495), .D(
        n15435), .X(n15436) );
  sky130_fd_sc_hd__nor4_1 U22629 ( .A(n20668), .B(n15437), .C(n20659), .D(
        n15436), .Y(n15443) );
  sky130_fd_sc_hd__nand2_1 U22630 ( .A(n20579), .B(n12137), .Y(n20663) );
  sky130_fd_sc_hd__nor2_1 U22631 ( .A(n15439), .B(n15438), .Y(n20593) );
  sky130_fd_sc_hd__nor2_1 U22632 ( .A(n15705), .B(n20527), .Y(n20585) );
  sky130_fd_sc_hd__nand2_1 U22633 ( .A(n15725), .B(n17289), .Y(n15440) );
  sky130_fd_sc_hd__nor2_1 U22634 ( .A(n15703), .B(n15440), .Y(n20526) );
  sky130_fd_sc_hd__nand2_1 U22635 ( .A(n20585), .B(n20515), .Y(n20650) );
  sky130_fd_sc_hd__or3_1 U22636 ( .A(n20593), .B(n15441), .C(n20650), .X(
        n20446) );
  sky130_fd_sc_hd__nor2_1 U22637 ( .A(n15689), .B(n20668), .Y(n15713) );
  sky130_fd_sc_hd__nand2_1 U22638 ( .A(n15713), .B(n15724), .Y(n20631) );
  sky130_fd_sc_hd__nor4_1 U22639 ( .A(n20592), .B(n20495), .C(n20446), .D(
        n20631), .Y(n15442) );
  sky130_fd_sc_hd__nand2_1 U22640 ( .A(n17175), .B(n20788), .Y(n20683) );
  sky130_fd_sc_hd__o22ai_1 U22641 ( .A1(n15443), .A2(n20663), .B1(n15442), 
        .B2(n20683), .Y(n15444) );
  sky130_fd_sc_hd__nor3_1 U22642 ( .A(n15446), .B(n15445), .C(n15444), .Y(
        n15465) );
  sky130_fd_sc_hd__nand3_1 U22643 ( .A(n19085), .B(n19381), .C(n15454), .Y(
        n15482) );
  sky130_fd_sc_hd__nand2b_1 U22644 ( .A_N(n15482), .B(n17289), .Y(n15718) );
  sky130_fd_sc_hd__nand2_1 U22645 ( .A(n17161), .B(n19381), .Y(n15468) );
  sky130_fd_sc_hd__nor2_1 U22646 ( .A(n15447), .B(n15468), .Y(n20636) );
  sky130_fd_sc_hd__nand2_1 U22647 ( .A(n20636), .B(n17289), .Y(n15696) );
  sky130_fd_sc_hd__nand2_1 U22648 ( .A(n15718), .B(n15696), .Y(n20481) );
  sky130_fd_sc_hd__nand3_1 U22649 ( .A(n15725), .B(n19381), .C(n15458), .Y(
        n20637) );
  sky130_fd_sc_hd__nor4_1 U22650 ( .A(n20668), .B(n20592), .C(n20661), .D(
        n20659), .Y(n15448) );
  sky130_fd_sc_hd__a31oi_1 U22651 ( .A1(n15692), .A2(n20450), .A3(n15448), 
        .B1(n20683), .Y(n15463) );
  sky130_fd_sc_hd__nor2_1 U22652 ( .A(n15450), .B(n15449), .Y(n20518) );
  sky130_fd_sc_hd__nand3_1 U22653 ( .A(n16180), .B(
        j202_soc_core_bootrom_00_address_w[9]), .C(n17161), .Y(n20601) );
  sky130_fd_sc_hd__nor2_1 U22654 ( .A(n20518), .B(n20630), .Y(n15675) );
  sky130_fd_sc_hd__nor2_1 U22655 ( .A(n15716), .B(n20466), .Y(n15453) );
  sky130_fd_sc_hd__nand2_1 U22656 ( .A(n15451), .B(n16616), .Y(n20574) );
  sky130_fd_sc_hd__nand3_1 U22657 ( .A(n16180), .B(n16616), .C(n15454), .Y(
        n20665) );
  sky130_fd_sc_hd__nand2_1 U22658 ( .A(n20574), .B(n20665), .Y(n15677) );
  sky130_fd_sc_hd__nor2_1 U22659 ( .A(n15695), .B(n20592), .Y(n20475) );
  sky130_fd_sc_hd__nand2_1 U22660 ( .A(n20475), .B(n20582), .Y(n20528) );
  sky130_fd_sc_hd__nor3_1 U22661 ( .A(n20477), .B(n15677), .C(n20528), .Y(
        n15452) );
  sky130_fd_sc_hd__a31oi_1 U22662 ( .A1(n15675), .A2(n15453), .A3(n15452), 
        .B1(n20651), .Y(n15462) );
  sky130_fd_sc_hd__nor2_1 U22663 ( .A(n15716), .B(n20526), .Y(n15480) );
  sky130_fd_sc_hd__nand2_1 U22664 ( .A(n15480), .B(n20665), .Y(n15694) );
  sky130_fd_sc_hd__nand2_1 U22665 ( .A(n20442), .B(n15724), .Y(n20514) );
  sky130_fd_sc_hd__nand2_1 U22666 ( .A(n15707), .B(n15723), .Y(n20605) );
  sky130_fd_sc_hd__nand2_1 U22667 ( .A(n15718), .B(n20601), .Y(n15457) );
  sky130_fd_sc_hd__nor2_1 U22668 ( .A(n20605), .B(n15457), .Y(n20613) );
  sky130_fd_sc_hd__nand2b_1 U22669 ( .A_N(n16953), .B(n15454), .Y(n20634) );
  sky130_fd_sc_hd__nand3_1 U22670 ( .A(n20653), .B(n20583), .C(n20634), .Y(
        n20679) );
  sky130_fd_sc_hd__nand4_1 U22671 ( .A(n15470), .B(n20613), .C(n15455), .D(
        n20479), .Y(n15456) );
  sky130_fd_sc_hd__nor2_1 U22672 ( .A(n15694), .B(n15456), .Y(n15460) );
  sky130_fd_sc_hd__nand2_1 U22673 ( .A(n20574), .B(n20570), .Y(n15691) );
  sky130_fd_sc_hd__nand2_1 U22674 ( .A(n20582), .B(n15672), .Y(n20461) );
  sky130_fd_sc_hd__nand2b_1 U22675 ( .A_N(n20461), .B(n20634), .Y(n20504) );
  sky130_fd_sc_hd__nand2_1 U22676 ( .A(n20632), .B(n15458), .Y(n20532) );
  sky130_fd_sc_hd__nand2_1 U22677 ( .A(n15693), .B(n20532), .Y(n20595) );
  sky130_fd_sc_hd__nor4_1 U22678 ( .A(n15705), .B(n15691), .C(n20504), .D(
        n20595), .Y(n15459) );
  sky130_fd_sc_hd__o22ai_1 U22679 ( .A1(n15460), .A2(n20663), .B1(n15459), 
        .B2(n20681), .Y(n15461) );
  sky130_fd_sc_hd__nor3_1 U22680 ( .A(n15463), .B(n15462), .C(n15461), .Y(
        n15464) );
  sky130_fd_sc_hd__mux2i_1 U22681 ( .A0(n15465), .A1(n15464), .S(n20623), .Y(
        n15466) );
  sky130_fd_sc_hd__nand2_1 U22682 ( .A(n15466), .B(n20626), .Y(n15505) );
  sky130_fd_sc_hd__nor2_1 U22683 ( .A(n15468), .B(n15467), .Y(n20476) );
  sky130_fd_sc_hd__nor2_1 U22684 ( .A(n20476), .B(n20667), .Y(n20508) );
  sky130_fd_sc_hd__nand2_1 U22685 ( .A(n15470), .B(n15469), .Y(n15678) );
  sky130_fd_sc_hd__nand2b_1 U22686 ( .A_N(n20637), .B(n17289), .Y(n20502) );
  sky130_fd_sc_hd__nand2_1 U22687 ( .A(n20665), .B(n20502), .Y(n20611) );
  sky130_fd_sc_hd__nand2_1 U22688 ( .A(n15471), .B(n15723), .Y(n20596) );
  sky130_fd_sc_hd__nor4_1 U22689 ( .A(n15678), .B(n20504), .C(n20611), .D(
        n20596), .Y(n15472) );
  sky130_fd_sc_hd__a21oi_1 U22690 ( .A1(n20508), .A2(n15472), .B1(n20663), .Y(
        n15479) );
  sky130_fd_sc_hd__nor2_1 U22691 ( .A(n20636), .B(n20448), .Y(n20517) );
  sky130_fd_sc_hd__nor4_1 U22692 ( .A(n20606), .B(n20605), .C(n20461), .D(
        n15483), .Y(n15473) );
  sky130_fd_sc_hd__a31oi_1 U22693 ( .A1(n20517), .A2(n15473), .A3(n20583), 
        .B1(n20651), .Y(n15478) );
  sky130_fd_sc_hd__nand2_1 U22694 ( .A(n15718), .B(n20634), .Y(n20618) );
  sky130_fd_sc_hd__nor2_1 U22695 ( .A(n20650), .B(n20618), .Y(n20470) );
  sky130_fd_sc_hd__nor3_1 U22696 ( .A(n20476), .B(n15695), .C(n16942), .Y(
        n15474) );
  sky130_fd_sc_hd__a31oi_1 U22697 ( .A1(n20470), .A2(n20516), .A3(n15474), 
        .B1(n20681), .Y(n15477) );
  sky130_fd_sc_hd__nand2_1 U22698 ( .A(n20632), .B(n16159), .Y(n20571) );
  sky130_fd_sc_hd__nand2_1 U22699 ( .A(n20472), .B(n20584), .Y(n20645) );
  sky130_fd_sc_hd__nand2b_1 U22700 ( .A_N(n20518), .B(n20664), .Y(n15740) );
  sky130_fd_sc_hd__nor3_1 U22701 ( .A(n20499), .B(n20521), .C(n15740), .Y(
        n20603) );
  sky130_fd_sc_hd__nor4_1 U22702 ( .A(n15705), .B(n20606), .C(n20645), .D(
        n20674), .Y(n15475) );
  sky130_fd_sc_hd__a31oi_1 U22703 ( .A1(n20458), .A2(n15475), .A3(n20570), 
        .B1(n20683), .Y(n15476) );
  sky130_fd_sc_hd__nor4_1 U22704 ( .A(n15479), .B(n15478), .C(n15477), .D(
        n15476), .Y(n15492) );
  sky130_fd_sc_hd__nand2_1 U22705 ( .A(n20643), .B(n20603), .Y(n20617) );
  sky130_fd_sc_hd__nor2_1 U22706 ( .A(n20647), .B(n15688), .Y(n20652) );
  sky130_fd_sc_hd__a31oi_1 U22707 ( .A1(n20478), .A2(n15480), .A3(n20652), 
        .B1(n20681), .Y(n15490) );
  sky130_fd_sc_hd__nor2_1 U22708 ( .A(n20448), .B(n20618), .Y(n20589) );
  sky130_fd_sc_hd__nand2_1 U22709 ( .A(n15707), .B(n20643), .Y(n20490) );
  sky130_fd_sc_hd__nor4_1 U22710 ( .A(n15671), .B(n20477), .C(n15677), .D(
        n20490), .Y(n15481) );
  sky130_fd_sc_hd__a31oi_1 U22711 ( .A1(n15682), .A2(n20589), .A3(n15481), 
        .B1(n20651), .Y(n15489) );
  sky130_fd_sc_hd__nand2_1 U22712 ( .A(n20636), .B(n17293), .Y(n20473) );
  sky130_fd_sc_hd__nand2_1 U22713 ( .A(n20473), .B(n20442), .Y(n20505) );
  sky130_fd_sc_hd__nor2_1 U22714 ( .A(n20499), .B(n20518), .Y(n20440) );
  sky130_fd_sc_hd__nor2_1 U22715 ( .A(n20505), .B(n20612), .Y(n15736) );
  sky130_fd_sc_hd__nor3_1 U22716 ( .A(n15484), .B(n20495), .C(n15483), .Y(
        n15485) );
  sky130_fd_sc_hd__a21oi_1 U22717 ( .A1(n15736), .A2(n15485), .B1(n20683), .Y(
        n15488) );
  sky130_fd_sc_hd__nor2_1 U22718 ( .A(n15695), .B(n20667), .Y(n20494) );
  sky130_fd_sc_hd__nor4_1 U22719 ( .A(n20513), .B(n20630), .C(n15688), .D(
        n20466), .Y(n15486) );
  sky130_fd_sc_hd__a21oi_1 U22720 ( .A1(n20494), .A2(n15486), .B1(n20663), .Y(
        n15487) );
  sky130_fd_sc_hd__nor4_1 U22721 ( .A(n15490), .B(n15489), .C(n15488), .D(
        n15487), .Y(n15491) );
  sky130_fd_sc_hd__mux2i_1 U22722 ( .A0(n15492), .A1(n15491), .S(n20623), .Y(
        n15494) );
  sky130_fd_sc_hd__nand2_1 U22723 ( .A(n15494), .B(n20693), .Y(n15504) );
  sky130_fd_sc_hd__nand2_1 U22724 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_duty[6]), .Y(n15501) );
  sky130_fd_sc_hd__nand4b_1 U22725 ( .A_N(n15495), .B(n15505), .C(n15504), .D(
        n15501), .Y(n15496) );
  sky130_fd_sc_hd__nand2_1 U22726 ( .A(j202_soc_core_memory0_ram_dout0[498]), 
        .B(n21771), .Y(n15507) );
  sky130_fd_sc_hd__nand2_1 U22727 ( .A(n15497), .B(n21738), .Y(n15500) );
  sky130_fd_sc_hd__nor2_1 U22728 ( .A(n15500), .B(n15499), .Y(n15502) );
  sky130_fd_sc_hd__and4_1 U22729 ( .A(n15504), .B(n15503), .C(n15502), .D(
        n15501), .X(n15506) );
  sky130_fd_sc_hd__nand3_1 U22730 ( .A(n15507), .B(n15506), .C(n15505), .Y(
        n20709) );
  sky130_fd_sc_hd__nor2_1 U22731 ( .A(n21014), .B(n15508), .Y(n15511) );
  sky130_fd_sc_hd__o21ai_0 U22732 ( .A1(n21014), .A2(n15509), .B1(n21015), .Y(
        n15510) );
  sky130_fd_sc_hd__a21oi_1 U22733 ( .A1(n22513), .A2(n15511), .B1(n15510), .Y(
        n15516) );
  sky130_fd_sc_hd__nand2_1 U22734 ( .A(n15514), .B(n15513), .Y(n15515) );
  sky130_fd_sc_hd__xor2_1 U22735 ( .A(n15516), .B(n15515), .X(n24766) );
  sky130_fd_sc_hd__nor2_1 U22736 ( .A(n21008), .B(n21009), .Y(n15517) );
  sky130_fd_sc_hd__xnor2_1 U22737 ( .A(n15518), .B(n15517), .Y(n24799) );
  sky130_fd_sc_hd__o22ai_1 U22738 ( .A1(n15519), .A2(n13603), .B1(n26571), 
        .B2(n11143), .Y(n15520) );
  sky130_fd_sc_hd__a21oi_1 U22739 ( .A1(n17120), .A2(n27432), .B1(n15520), .Y(
        n15522) );
  sky130_fd_sc_hd__nand2b_1 U22740 ( .A_N(n21584), .B(n24799), .Y(n15521) );
  sky130_fd_sc_hd__o211ai_1 U22741 ( .A1(n26572), .A2(n22592), .B1(n15522), 
        .C1(n15521), .Y(n15523) );
  sky130_fd_sc_hd__a21oi_1 U22742 ( .A1(n24766), .A2(n12158), .B1(n15523), .Y(
        n15524) );
  sky130_fd_sc_hd__nand2_1 U22743 ( .A(j202_soc_core_memory0_ram_dout0[181]), 
        .B(n21590), .Y(n15529) );
  sky130_fd_sc_hd__nand2_1 U22744 ( .A(j202_soc_core_memory0_ram_dout0[117]), 
        .B(n21591), .Y(n15528) );
  sky130_fd_sc_hd__nand2_1 U22745 ( .A(j202_soc_core_memory0_ram_dout0[149]), 
        .B(n21592), .Y(n15527) );
  sky130_fd_sc_hd__nand2_1 U22746 ( .A(j202_soc_core_memory0_ram_dout0[341]), 
        .B(n21593), .Y(n15526) );
  sky130_fd_sc_hd__nand2_1 U22747 ( .A(j202_soc_core_memory0_ram_dout0[277]), 
        .B(n21605), .Y(n15641) );
  sky130_fd_sc_hd__nand2_1 U22748 ( .A(j202_soc_core_memory0_ram_dout0[309]), 
        .B(n21603), .Y(n15640) );
  sky130_fd_sc_hd__nand2_1 U22749 ( .A(j202_soc_core_memory0_ram_dout0[53]), 
        .B(n21604), .Y(n15639) );
  sky130_fd_sc_hd__a31oi_1 U22750 ( .A1(n15532), .A2(n15531), .A3(n15530), 
        .B1(n15708), .Y(n15555) );
  sky130_fd_sc_hd__nand4_1 U22751 ( .A(n15535), .B(n15534), .C(n15533), .D(
        n15612), .Y(n15536) );
  sky130_fd_sc_hd__nand2_1 U22752 ( .A(n15578), .B(n15609), .Y(n15544) );
  sky130_fd_sc_hd__nand3_1 U22754 ( .A(n15610), .B(n15538), .C(n15537), .Y(
        n15540) );
  sky130_fd_sc_hd__nand3b_1 U22756 ( .A_N(n15543), .B(n15542), .C(n15541), .Y(
        n15554) );
  sky130_fd_sc_hd__nand2_1 U22757 ( .A(n15612), .B(n15545), .Y(n15546) );
  sky130_fd_sc_hd__nor4b_1 U22758 ( .D_N(n15549), .A(n15548), .B(n15547), .C(
        n15546), .Y(n15552) );
  sky130_fd_sc_hd__a31oi_1 U22759 ( .A1(n15552), .A2(n15551), .A3(n15550), 
        .B1(n15616), .Y(n15553) );
  sky130_fd_sc_hd__o31a_1 U22760 ( .A1(n15555), .A2(n15554), .A3(n15553), .B1(
        n13481), .X(n15652) );
  sky130_fd_sc_hd__a31oi_1 U22761 ( .A1(n15559), .A2(n15558), .A3(n15578), 
        .B1(n15557), .Y(n15567) );
  sky130_fd_sc_hd__nor3_1 U22762 ( .A(n15563), .B(n15562), .C(n15561), .Y(
        n15565) );
  sky130_fd_sc_hd__a31oi_1 U22763 ( .A1(n15565), .A2(n15594), .A3(n15564), 
        .B1(n15708), .Y(n15566) );
  sky130_fd_sc_hd__nor2_1 U22764 ( .A(n15567), .B(n15566), .Y(n15575) );
  sky130_fd_sc_hd__o31ai_1 U22765 ( .A1(n15570), .A2(n15569), .A3(n15568), 
        .B1(n15584), .Y(n15574) );
  sky130_fd_sc_hd__nand3_1 U22767 ( .A(n15575), .B(n15574), .C(n15573), .Y(
        n15576) );
  sky130_fd_sc_hd__nand2_1 U22768 ( .A(n15576), .B(n21697), .Y(n15650) );
  sky130_fd_sc_hd__a22oi_1 U22769 ( .A1(n21675), .A2(
        j202_soc_core_uart_div1[5]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[85]), .Y(n15644) );
  sky130_fd_sc_hd__nand2_1 U22770 ( .A(n21699), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[53]), .Y(n15643) );
  sky130_fd_sc_hd__nand2_1 U22771 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[21]), .Y(n15642) );
  sky130_fd_sc_hd__nand4_1 U22772 ( .A(n15644), .B(n21677), .C(n15643), .D(
        n15642), .Y(n15605) );
  sky130_fd_sc_hd__nand2_1 U22773 ( .A(n15578), .B(n15577), .Y(n15579) );
  sky130_fd_sc_hd__nor3_1 U22774 ( .A(n15581), .B(n15580), .C(n15579), .Y(
        n15582) );
  sky130_fd_sc_hd__nand2_1 U22775 ( .A(n15583), .B(n15582), .Y(n15585) );
  sky130_fd_sc_hd__nand2_1 U22776 ( .A(n15585), .B(n15584), .Y(n15600) );
  sky130_fd_sc_hd__nor2_1 U22777 ( .A(n15588), .B(n15587), .Y(n15617) );
  sky130_fd_sc_hd__nand4_1 U22778 ( .A(n15590), .B(n15617), .C(n15589), .D(
        n15613), .Y(n15591) );
  sky130_fd_sc_hd__nand2_1 U22779 ( .A(n16090), .B(n15591), .Y(n15599) );
  sky130_fd_sc_hd__nand4_1 U22780 ( .A(n15595), .B(n15594), .C(n15593), .D(
        n15592), .Y(n15597) );
  sky130_fd_sc_hd__nand3_1 U22782 ( .A(n15600), .B(n15599), .C(n15598), .Y(
        n15604) );
  sky130_fd_sc_hd__a21oi_1 U22783 ( .A1(n15602), .A2(n15601), .B1(n15708), .Y(
        n15603) );
  sky130_fd_sc_hd__o21a_1 U22784 ( .A1(n15604), .A2(n15603), .B1(n21727), .X(
        n15645) );
  sky130_fd_sc_hd__nor3_1 U22785 ( .A(n15647), .B(n15605), .C(n15645), .Y(
        n15636) );
  sky130_fd_sc_hd__nor3_1 U22786 ( .A(n15608), .B(n15607), .C(n15606), .Y(
        n15611) );
  sky130_fd_sc_hd__and4_1 U22787 ( .A(n15615), .B(n15614), .C(n15613), .D(
        n15612), .X(n15618) );
  sky130_fd_sc_hd__a31oi_1 U22788 ( .A1(n15619), .A2(n15618), .A3(n15617), 
        .B1(n15616), .Y(n15621) );
  sky130_fd_sc_hd__nor2_1 U22789 ( .A(n15621), .B(n15620), .Y(n15633) );
  sky130_fd_sc_hd__nor2_1 U22790 ( .A(n15623), .B(n15622), .Y(n15624) );
  sky130_fd_sc_hd__nand2_1 U22791 ( .A(n18952), .B(n15624), .Y(n15626) );
  sky130_fd_sc_hd__nor2_1 U22792 ( .A(n15626), .B(n15625), .Y(n15627) );
  sky130_fd_sc_hd__nand3_1 U22793 ( .A(n15629), .B(n15628), .C(n15627), .Y(
        n15631) );
  sky130_fd_sc_hd__nand2_1 U22794 ( .A(n15631), .B(n15630), .Y(n15632) );
  sky130_fd_sc_hd__nand3_1 U22795 ( .A(n15634), .B(n15633), .C(n15632), .Y(
        n15635) );
  sky130_fd_sc_hd__nand2_1 U22796 ( .A(n15635), .B(n20908), .Y(n15648) );
  sky130_fd_sc_hd__nand3_1 U22797 ( .A(n15650), .B(n15636), .C(n15648), .Y(
        n15637) );
  sky130_fd_sc_hd__nor2_1 U22798 ( .A(n15652), .B(n15637), .Y(n15638) );
  sky130_fd_sc_hd__nand2_1 U22799 ( .A(j202_soc_core_memory0_ram_dout0[501]), 
        .B(n21771), .Y(n15654) );
  sky130_fd_sc_hd__nand4_1 U22800 ( .A(n15644), .B(n21738), .C(n15643), .D(
        n15642), .Y(n15646) );
  sky130_fd_sc_hd__nor3_1 U22801 ( .A(n15647), .B(n15646), .C(n15645), .Y(
        n15649) );
  sky130_fd_sc_hd__nand3_1 U22802 ( .A(n15650), .B(n15649), .C(n15648), .Y(
        n15651) );
  sky130_fd_sc_hd__nor2_1 U22803 ( .A(n15652), .B(n15651), .Y(n15653) );
  sky130_fd_sc_hd__nand2_1 U22804 ( .A(n15654), .B(n15653), .Y(n21751) );
  sky130_fd_sc_hd__nand2_1 U22805 ( .A(n22515), .B(n27412), .Y(n15658) );
  sky130_fd_sc_hd__xor2_1 U22806 ( .A(n15656), .B(n15655), .X(n25423) );
  sky130_fd_sc_hd__nand2_1 U22807 ( .A(n22596), .B(n25423), .Y(n15657) );
  sky130_fd_sc_hd__a21oi_1 U22808 ( .A1(n22513), .A2(n15662), .B1(n15661), .Y(
        n15667) );
  sky130_fd_sc_hd__nand2_1 U22809 ( .A(n15665), .B(n15664), .Y(n15666) );
  sky130_fd_sc_hd__xor2_1 U22810 ( .A(n15667), .B(n15666), .X(n25412) );
  sky130_fd_sc_hd__nand2_1 U22811 ( .A(n25412), .B(n12158), .Y(n15668) );
  sky130_fd_sc_hd__a22oi_1 U22812 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[51]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[83]), .Y(n15762) );
  sky130_fd_sc_hd__nand2_1 U22813 ( .A(n21675), .B(j202_soc_core_uart_div1[3]), 
        .Y(n15757) );
  sky130_fd_sc_hd__nand2_1 U22814 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[19]), .Y(n15756) );
  sky130_fd_sc_hd__nand4_1 U22815 ( .A(n15762), .B(n21677), .C(n15757), .D(
        n15756), .Y(n15750) );
  sky130_fd_sc_hd__nand2_1 U22816 ( .A(n20632), .B(n17161), .Y(n20602) );
  sky130_fd_sc_hd__nor2_1 U22817 ( .A(n15691), .B(n15733), .Y(n20500) );
  sky130_fd_sc_hd__nand2_1 U22818 ( .A(n15670), .B(n20500), .Y(n20525) );
  sky130_fd_sc_hd__nor2_1 U22819 ( .A(n15671), .B(n20491), .Y(n20498) );
  sky130_fd_sc_hd__nand2_1 U22820 ( .A(n20498), .B(n20669), .Y(n20660) );
  sky130_fd_sc_hd__nor4_1 U22822 ( .A(n20525), .B(n20660), .C(n20481), .D(
        n15732), .Y(n15674) );
  sky130_fd_sc_hd__a31oi_1 U22823 ( .A1(n15675), .A2(n15674), .A3(n15680), 
        .B1(n20681), .Y(n15687) );
  sky130_fd_sc_hd__nor2_1 U22824 ( .A(n20476), .B(n15676), .Y(n15690) );
  sky130_fd_sc_hd__nand2_1 U22825 ( .A(n20517), .B(n15690), .Y(n15717) );
  sky130_fd_sc_hd__nor3_1 U22826 ( .A(n15678), .B(n15677), .C(n15717), .Y(
        n15679) );
  sky130_fd_sc_hd__a31oi_1 U22827 ( .A1(n15679), .A2(n20582), .A3(n20648), 
        .B1(n20663), .Y(n15686) );
  sky130_fd_sc_hd__nor2_1 U22828 ( .A(n15733), .B(n15741), .Y(n20615) );
  sky130_fd_sc_hd__nor4b_1 U22829 ( .D_N(n20615), .A(n20491), .B(n20461), .C(
        n20650), .Y(n15681) );
  sky130_fd_sc_hd__a31oi_1 U22830 ( .A1(n15682), .A2(n15681), .A3(n15680), 
        .B1(n20683), .Y(n15685) );
  sky130_fd_sc_hd__nand2_1 U22831 ( .A(n20508), .B(n15738), .Y(n15714) );
  sky130_fd_sc_hd__nand2_1 U22832 ( .A(n20613), .B(n15722), .Y(n20591) );
  sky130_fd_sc_hd__nor4_1 U22833 ( .A(n20518), .B(n20526), .C(n20466), .D(
        n20591), .Y(n15683) );
  sky130_fd_sc_hd__a31oi_1 U22834 ( .A1(n20516), .A2(n15683), .A3(n15696), 
        .B1(n20651), .Y(n15684) );
  sky130_fd_sc_hd__nor4_1 U22835 ( .A(n15687), .B(n15686), .C(n15685), .D(
        n15684), .Y(n15702) );
  sky130_fd_sc_hd__nor2_1 U22836 ( .A(n15689), .B(n15688), .Y(n20523) );
  sky130_fd_sc_hd__nand2_1 U22837 ( .A(n15690), .B(n20523), .Y(n20675) );
  sky130_fd_sc_hd__nor2_1 U22838 ( .A(n15691), .B(n20675), .Y(n20471) );
  sky130_fd_sc_hd__a31oi_1 U22839 ( .A1(n15692), .A2(n20498), .A3(n20471), 
        .B1(n20681), .Y(n15700) );
  sky130_fd_sc_hd__nand2_1 U22840 ( .A(n15693), .B(n15723), .Y(n20444) );
  sky130_fd_sc_hd__nor4_1 U22841 ( .A(n15720), .B(n20504), .C(n15694), .D(
        n20444), .Y(n15698) );
  sky130_fd_sc_hd__nor3_1 U22842 ( .A(n15695), .B(n20526), .C(n20495), .Y(
        n20671) );
  sky130_fd_sc_hd__nand3_1 U22843 ( .A(n20615), .B(n20458), .C(n20671), .Y(
        n20534) );
  sky130_fd_sc_hd__nand2_1 U22844 ( .A(n20584), .B(n15696), .Y(n20610) );
  sky130_fd_sc_hd__nor4_1 U22845 ( .A(n15705), .B(n20593), .C(n20534), .D(
        n20610), .Y(n15697) );
  sky130_fd_sc_hd__o22ai_1 U22846 ( .A1(n15698), .A2(n20663), .B1(n15697), 
        .B2(n20683), .Y(n15699) );
  sky130_fd_sc_hd__nor2_1 U22847 ( .A(n15700), .B(n15699), .Y(n15701) );
  sky130_fd_sc_hd__mux2_2 U22848 ( .A0(n15702), .A1(n15701), .S(n20687), .X(
        n15711) );
  sky130_fd_sc_hd__nand2b_1 U22849 ( .A_N(n15716), .B(n20602), .Y(n20447) );
  sky130_fd_sc_hd__nand2_1 U22850 ( .A(n15713), .B(n20515), .Y(n20590) );
  sky130_fd_sc_hd__a21oi_1 U22851 ( .A1(n15704), .A2(n15726), .B1(n20590), .Y(
        n20452) );
  sky130_fd_sc_hd__nor2_1 U22852 ( .A(n15706), .B(n15705), .Y(n20609) );
  sky130_fd_sc_hd__nand4b_1 U22853 ( .A_N(n20447), .B(n20452), .C(n20609), .D(
        n15707), .Y(n15709) );
  sky130_fd_sc_hd__nor2_1 U22854 ( .A(n12137), .B(n15708), .Y(n20692) );
  sky130_fd_sc_hd__nand2_1 U22855 ( .A(n15709), .B(n20692), .Y(n15710) );
  sky130_fd_sc_hd__nand2_1 U22856 ( .A(n15711), .B(n15710), .Y(n15712) );
  sky130_fd_sc_hd__nand2_1 U22857 ( .A(n15712), .B(n20626), .Y(n15764) );
  sky130_fd_sc_hd__nor4_1 U22858 ( .A(n15714), .B(n20641), .C(n20528), .D(
        n20447), .Y(n15715) );
  sky130_fd_sc_hd__a31oi_1 U22859 ( .A1(n20440), .A2(n15715), .A3(n15723), 
        .B1(n20683), .Y(n15731) );
  sky130_fd_sc_hd__nor2_1 U22860 ( .A(n15716), .B(n20518), .Y(n20493) );
  sky130_fd_sc_hd__nor3b_1 U22861 ( .C_N(n20493), .A(n20642), .B(n15717), .Y(
        n15719) );
  sky130_fd_sc_hd__a31oi_1 U22862 ( .A1(n20523), .A2(n15719), .A3(n15718), 
        .B1(n20681), .Y(n15730) );
  sky130_fd_sc_hd__nor3_1 U22863 ( .A(n20491), .B(n15720), .C(n20659), .Y(
        n15721) );
  sky130_fd_sc_hd__a31oi_1 U22864 ( .A1(n20479), .A2(n15722), .A3(n15721), 
        .B1(n20651), .Y(n15729) );
  sky130_fd_sc_hd__nor2_1 U22865 ( .A(n20491), .B(n20680), .Y(n20614) );
  sky130_fd_sc_hd__nand2_1 U22866 ( .A(n20614), .B(n15724), .Y(n20480) );
  sky130_fd_sc_hd__nor2_1 U22867 ( .A(n20448), .B(n20480), .Y(n20638) );
  sky130_fd_sc_hd__nor2_1 U22868 ( .A(n16171), .B(n20571), .Y(n20459) );
  sky130_fd_sc_hd__a21oi_1 U22869 ( .A1(n15726), .A2(n15725), .B1(n20459), .Y(
        n15727) );
  sky130_fd_sc_hd__a31oi_1 U22870 ( .A1(n20638), .A2(n20508), .A3(n15727), 
        .B1(n20663), .Y(n15728) );
  sky130_fd_sc_hd__nor4_1 U22871 ( .A(n15731), .B(n15730), .C(n15729), .D(
        n15728), .Y(n15748) );
  sky130_fd_sc_hd__nand2_1 U22872 ( .A(n20601), .B(n20643), .Y(n20646) );
  sky130_fd_sc_hd__nor2_1 U22873 ( .A(n15733), .B(n20646), .Y(n20520) );
  sky130_fd_sc_hd__a31oi_1 U22874 ( .A1(n15734), .A2(n20516), .A3(n20520), 
        .B1(n20663), .Y(n15746) );
  sky130_fd_sc_hd__nor2b_1 U22875 ( .B_N(n20584), .A(n15735), .Y(n20497) );
  sky130_fd_sc_hd__a31oi_1 U22876 ( .A1(n15736), .A2(n20520), .A3(n20497), 
        .B1(n20681), .Y(n15745) );
  sky130_fd_sc_hd__nand4_1 U22877 ( .A(n15738), .B(n20463), .C(n20442), .D(
        n15737), .Y(n15739) );
  sky130_fd_sc_hd__nor3_1 U22878 ( .A(n20521), .B(n15739), .C(n20679), .Y(
        n15743) );
  sky130_fd_sc_hd__nor4_1 U22879 ( .A(n15741), .B(n20481), .C(n20679), .D(
        n15740), .Y(n15742) );
  sky130_fd_sc_hd__o22ai_1 U22880 ( .A1(n15743), .A2(n20651), .B1(n15742), 
        .B2(n20683), .Y(n15744) );
  sky130_fd_sc_hd__nor3_1 U22881 ( .A(n15746), .B(n15745), .C(n15744), .Y(
        n15747) );
  sky130_fd_sc_hd__mux2i_1 U22882 ( .A0(n15748), .A1(n15747), .S(n20623), .Y(
        n15749) );
  sky130_fd_sc_hd__nand2_1 U22883 ( .A(n15749), .B(n20693), .Y(n15763) );
  sky130_fd_sc_hd__nand2_1 U22884 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_duty[7]), .Y(n15760) );
  sky130_fd_sc_hd__nand4b_1 U22885 ( .A_N(n15750), .B(n15764), .C(n15763), .D(
        n15760), .Y(n15751) );
  sky130_fd_sc_hd__a21oi_1 U22886 ( .A1(j202_soc_core_memory0_ram_dout0[147]), 
        .A2(n21592), .B1(n15751), .Y(n15753) );
  sky130_fd_sc_hd__nand4_1 U22887 ( .A(n15755), .B(n15754), .C(n15753), .D(
        n15752), .Y(n20716) );
  sky130_fd_sc_hd__nand2_1 U22888 ( .A(n15756), .B(n21738), .Y(n15759) );
  sky130_fd_sc_hd__nor2_1 U22889 ( .A(n15759), .B(n15758), .Y(n15761) );
  sky130_fd_sc_hd__and4_1 U22890 ( .A(n15763), .B(n15762), .C(n15761), .D(
        n15760), .X(n15765) );
  sky130_fd_sc_hd__xnor2_1 U22891 ( .A(n15767), .B(n15766), .Y(n25669) );
  sky130_fd_sc_hd__nand2_1 U22892 ( .A(n22596), .B(n25669), .Y(n15769) );
  sky130_fd_sc_hd__nand2_1 U22893 ( .A(n22515), .B(n27425), .Y(n15768) );
  sky130_fd_sc_hd__a21oi_1 U22894 ( .A1(n22513), .A2(n15771), .B1(n15770), .Y(
        n15776) );
  sky130_fd_sc_hd__nand2_1 U22895 ( .A(n15774), .B(n15773), .Y(n15775) );
  sky130_fd_sc_hd__xor2_1 U22896 ( .A(n15776), .B(n15775), .X(n24085) );
  sky130_fd_sc_hd__nand2_1 U22897 ( .A(n24085), .B(n12158), .Y(n15777) );
  sky130_fd_sc_hd__a21oi_1 U22898 ( .A1(n19071), .A2(
        j202_soc_core_j22_cpu_memop_MEM__1_), .B1(n23300), .Y(n15779) );
  sky130_fd_sc_hd__mux2i_1 U22899 ( .A0(n15779), .A1(n15778), .S(n24280), .Y(
        n15780) );
  sky130_fd_sc_hd__nand2_1 U22900 ( .A(j202_soc_core_memory0_ram_dout0[26]), 
        .B(n21733), .Y(n15781) );
  sky130_fd_sc_hd__nand2_1 U22901 ( .A(j202_soc_core_memory0_ram_dout0[154]), 
        .B(n21592), .Y(n15785) );
  sky130_fd_sc_hd__nand2_1 U22902 ( .A(j202_soc_core_memory0_ram_dout0[90]), 
        .B(n21734), .Y(n15784) );
  sky130_fd_sc_hd__nand2_1 U22903 ( .A(j202_soc_core_memory0_ram_dout0[218]), 
        .B(n21732), .Y(n15783) );
  sky130_fd_sc_hd__nand2_1 U22904 ( .A(j202_soc_core_memory0_ram_dout0[122]), 
        .B(n21591), .Y(n15782) );
  sky130_fd_sc_hd__a22oi_1 U22905 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[58]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[90]), .Y(n15894) );
  sky130_fd_sc_hd__nand2_1 U22906 ( .A(n21675), .B(j202_soc_core_uart_div0[2]), 
        .Y(n15893) );
  sky130_fd_sc_hd__nand2_1 U22907 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[26]), .Y(n15892) );
  sky130_fd_sc_hd__nand4_1 U22908 ( .A(n15894), .B(n15893), .C(n21677), .D(
        n15892), .Y(n15889) );
  sky130_fd_sc_hd__nand2_1 U22909 ( .A(n15870), .B(n15871), .Y(n15788) );
  sky130_fd_sc_hd__nor2_1 U22910 ( .A(n15786), .B(n15854), .Y(n17027) );
  sky130_fd_sc_hd__nand3_1 U22911 ( .A(n17010), .B(n15788), .C(n15787), .Y(
        n15794) );
  sky130_fd_sc_hd__nand3_1 U22912 ( .A(n15802), .B(n15790), .C(n15789), .Y(
        n15791) );
  sky130_fd_sc_hd__nor2_1 U22913 ( .A(n15794), .B(n15791), .Y(n15792) );
  sky130_fd_sc_hd__nand2_1 U22914 ( .A(n17005), .B(n15792), .Y(n15793) );
  sky130_fd_sc_hd__nand2_1 U22915 ( .A(n15793), .B(n13387), .Y(n15808) );
  sky130_fd_sc_hd__o31ai_1 U22916 ( .A1(n15803), .A2(n15795), .A3(n15794), 
        .B1(n17302), .Y(n15807) );
  sky130_fd_sc_hd__nand2_1 U22917 ( .A(n15796), .B(n17049), .Y(n17016) );
  sky130_fd_sc_hd__nand2_1 U22918 ( .A(n15798), .B(n15797), .Y(n15799) );
  sky130_fd_sc_hd__o21ai_1 U22919 ( .A1(n15800), .A2(n15799), .B1(n17273), .Y(
        n15806) );
  sky130_fd_sc_hd__o21ai_1 U22920 ( .A1(n15804), .A2(n16080), .B1(n13388), .Y(
        n15805) );
  sky130_fd_sc_hd__nand4_1 U22921 ( .A(n15808), .B(n15807), .C(n15806), .D(
        n15805), .Y(n15809) );
  sky130_fd_sc_hd__nor2_1 U22922 ( .A(n15809), .B(n16085), .Y(n15832) );
  sky130_fd_sc_hd__nor2_1 U22923 ( .A(n15810), .B(n16067), .Y(n15812) );
  sky130_fd_sc_hd__nand3_1 U22924 ( .A(n17077), .B(n15812), .C(n15811), .Y(
        n15828) );
  sky130_fd_sc_hd__nor2_1 U22925 ( .A(n17289), .B(n16091), .Y(n15866) );
  sky130_fd_sc_hd__nand4_1 U22926 ( .A(n16059), .B(n15814), .C(n15813), .D(
        n16104), .Y(n15815) );
  sky130_fd_sc_hd__nor4_1 U22927 ( .A(n15817), .B(n15880), .C(n15816), .D(
        n15815), .Y(n15826) );
  sky130_fd_sc_hd__nand4_1 U22928 ( .A(n16058), .B(n16059), .C(n16098), .D(
        n17025), .Y(n15824) );
  sky130_fd_sc_hd__nand2_1 U22929 ( .A(n16564), .B(n15818), .Y(n17024) );
  sky130_fd_sc_hd__nor3_1 U22930 ( .A(n17083), .B(n16101), .C(n15866), .Y(
        n16060) );
  sky130_fd_sc_hd__nor2b_1 U22931 ( .B_N(n16060), .A(n15819), .Y(n15820) );
  sky130_fd_sc_hd__a31oi_1 U22932 ( .A1(n15822), .A2(n15821), .A3(n15820), 
        .B1(n17039), .Y(n15823) );
  sky130_fd_sc_hd__a21oi_1 U22933 ( .A1(n13388), .A2(n15824), .B1(n15823), .Y(
        n15825) );
  sky130_fd_sc_hd__o21ai_1 U22934 ( .A1(n17055), .A2(n15826), .B1(n15825), .Y(
        n15827) );
  sky130_fd_sc_hd__a21oi_1 U22935 ( .A1(n15828), .A2(n17273), .B1(n15827), .Y(
        n15829) );
  sky130_fd_sc_hd__o22ai_1 U22936 ( .A1(n15832), .A2(n15831), .B1(n15830), 
        .B2(n15829), .Y(n15888) );
  sky130_fd_sc_hd__nand3_1 U22937 ( .A(n15834), .B(n17025), .C(n17024), .Y(
        n15835) );
  sky130_fd_sc_hd__nor4_1 U22938 ( .A(n13306), .B(n16095), .C(n15836), .D(
        n15835), .Y(n15843) );
  sky130_fd_sc_hd__nand2_1 U22939 ( .A(n15838), .B(n15837), .Y(n15839) );
  sky130_fd_sc_hd__nand2_1 U22940 ( .A(n15840), .B(n15839), .Y(n15841) );
  sky130_fd_sc_hd__nand2_1 U22941 ( .A(n15841), .B(n13388), .Y(n15842) );
  sky130_fd_sc_hd__o21ai_1 U22942 ( .A1(n17039), .A2(n15843), .B1(n15842), .Y(
        n15862) );
  sky130_fd_sc_hd__or4_1 U22944 ( .A(n16073), .B(n16111), .C(n15848), .D(
        n15847), .X(n16125) );
  sky130_fd_sc_hd__nand2_1 U22945 ( .A(n15850), .B(n15849), .Y(n15851) );
  sky130_fd_sc_hd__nor4_1 U22946 ( .A(n15853), .B(n15852), .C(n16125), .D(
        n15851), .Y(n15860) );
  sky130_fd_sc_hd__nor2_1 U22947 ( .A(n15855), .B(n15854), .Y(n15868) );
  sky130_fd_sc_hd__nor4_1 U22948 ( .A(n15858), .B(n15857), .C(n15868), .D(
        n15856), .Y(n15859) );
  sky130_fd_sc_hd__o22ai_1 U22949 ( .A1(n15860), .A2(n17055), .B1(n15859), 
        .B2(n17037), .Y(n15861) );
  sky130_fd_sc_hd__mux2i_1 U22950 ( .A0(n15862), .A1(n15861), .S(n20787), .Y(
        n15886) );
  sky130_fd_sc_hd__nor4_1 U22951 ( .A(n15867), .B(n15866), .C(n15865), .D(
        n15879), .Y(n15878) );
  sky130_fd_sc_hd__nor3_1 U22952 ( .A(n15869), .B(n15868), .C(n17009), .Y(
        n15876) );
  sky130_fd_sc_hd__nand2_1 U22953 ( .A(n17273), .B(n20787), .Y(n17276) );
  sky130_fd_sc_hd__o21ai_1 U22954 ( .A1(n16126), .A2(n15871), .B1(n15870), .Y(
        n15872) );
  sky130_fd_sc_hd__nand2_1 U22955 ( .A(n17013), .B(n15872), .Y(n15873) );
  sky130_fd_sc_hd__nor3b_1 U22956 ( .C_N(n17048), .A(n15874), .B(n15873), .Y(
        n15875) );
  sky130_fd_sc_hd__o22a_1 U22957 ( .A1(n15876), .A2(n17276), .B1(n15875), .B2(
        n17282), .X(n15877) );
  sky130_fd_sc_hd__nor4_1 U22959 ( .A(n15882), .B(n15881), .C(n15880), .D(
        n15879), .Y(n17072) );
  sky130_fd_sc_hd__a21oi_1 U22960 ( .A1(n17072), .A2(n17028), .B1(n17059), .Y(
        n15883) );
  sky130_fd_sc_hd__nor2_1 U22961 ( .A(n15884), .B(n15883), .Y(n15885) );
  sky130_fd_sc_hd__a21oi_1 U22962 ( .A1(n15886), .A2(n15885), .B1(
        j202_soc_core_bootrom_00_address_w[8]), .Y(n15887) );
  sky130_fd_sc_hd__o21a_1 U22963 ( .A1(n15888), .A2(n15887), .B1(n17098), .X(
        n15896) );
  sky130_fd_sc_hd__nor2_1 U22964 ( .A(n15889), .B(n15896), .Y(n15890) );
  sky130_fd_sc_hd__nand2_1 U22965 ( .A(j202_soc_core_memory0_ram_dout0[506]), 
        .B(n21771), .Y(n15891) );
  sky130_fd_sc_hd__nand4_1 U22966 ( .A(n15894), .B(n15893), .C(n21738), .D(
        n15892), .Y(n15895) );
  sky130_fd_sc_hd__nor2_1 U22967 ( .A(n15896), .B(n15895), .Y(n15897) );
  sky130_fd_sc_hd__nand2_1 U22968 ( .A(n15891), .B(n15897), .Y(n15898) );
  sky130_fd_sc_hd__nor2_1 U22969 ( .A(n15952), .B(n15899), .Y(n16532) );
  sky130_fd_sc_hd__nand2_1 U22970 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[409]), .Y(n15903) );
  sky130_fd_sc_hd__nand2_1 U22971 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[473]), .Y(n15902) );
  sky130_fd_sc_hd__nand2_1 U22972 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[153]), .Y(n15901) );
  sky130_fd_sc_hd__nand2_1 U22973 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[121]), .Y(n15900) );
  sky130_fd_sc_hd__nand4_1 U22974 ( .A(n15903), .B(n15902), .C(n15901), .D(
        n15900), .Y(n15909) );
  sky130_fd_sc_hd__a21oi_1 U22975 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[25]), .B1(n16436), .Y(n15907) );
  sky130_fd_sc_hd__nand2_1 U22976 ( .A(n16431), .B(
        j202_soc_core_j22_cpu_rf_gpr[281]), .Y(n15906) );
  sky130_fd_sc_hd__nand2_1 U22977 ( .A(n11152), .B(
        j202_soc_core_j22_cpu_rf_gpr[57]), .Y(n15905) );
  sky130_fd_sc_hd__nand2_1 U22978 ( .A(n11155), .B(
        j202_soc_core_j22_cpu_rf_gpr[89]), .Y(n15904) );
  sky130_fd_sc_hd__nand4_1 U22979 ( .A(n15907), .B(n15906), .C(n15905), .D(
        n15904), .Y(n15908) );
  sky130_fd_sc_hd__nor2_1 U22980 ( .A(n15909), .B(n15908), .Y(n15921) );
  sky130_fd_sc_hd__nand2_1 U22981 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[249]), .Y(n15913) );
  sky130_fd_sc_hd__nand2_1 U22982 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_rf_gpr[217]), .Y(n15912) );
  sky130_fd_sc_hd__nand2_1 U22983 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[313]), .Y(n15911) );
  sky130_fd_sc_hd__nand2_1 U22984 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[441]), .Y(n15910) );
  sky130_fd_sc_hd__and4_1 U22985 ( .A(n15913), .B(n15912), .C(n15911), .D(
        n15910), .X(n15920) );
  sky130_fd_sc_hd__nand2_1 U22986 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[505]), .Y(n15917) );
  sky130_fd_sc_hd__nand2_1 U22987 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[345]), .Y(n15916) );
  sky130_fd_sc_hd__nand2_1 U22988 ( .A(n15128), .B(
        j202_soc_core_j22_cpu_rf_gpr[185]), .Y(n15915) );
  sky130_fd_sc_hd__nand2_1 U22989 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[377]), .Y(n15914) );
  sky130_fd_sc_hd__nand4_1 U22990 ( .A(n15917), .B(n15916), .C(n15915), .D(
        n15914), .Y(n15918) );
  sky130_fd_sc_hd__a21oi_1 U22991 ( .A1(j202_soc_core_j22_cpu_rf_gpr[25]), 
        .A2(n16285), .B1(n15918), .Y(n15919) );
  sky130_fd_sc_hd__nand3_1 U22992 ( .A(n15921), .B(n15920), .C(n15919), .Y(
        n25137) );
  sky130_fd_sc_hd__inv_2 U22993 ( .A(n25137), .Y(n26706) );
  sky130_fd_sc_hd__o22ai_1 U22994 ( .A1(n16492), .A2(n26706), .B1(n26701), 
        .B2(n13793), .Y(n15954) );
  sky130_fd_sc_hd__nand2_1 U22995 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[185]), .Y(n15925) );
  sky130_fd_sc_hd__nand2_1 U22996 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[249]), .Y(n15924) );
  sky130_fd_sc_hd__nand2_1 U22997 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[505]), .Y(n15923) );
  sky130_fd_sc_hd__nand2_1 U22998 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[441]), .Y(n15922) );
  sky130_fd_sc_hd__nand4_1 U22999 ( .A(n15925), .B(n15924), .C(n15923), .D(
        n15922), .Y(n15931) );
  sky130_fd_sc_hd__nand2_1 U23000 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[25]), .Y(n15929) );
  sky130_fd_sc_hd__nand2_1 U23001 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[57]), .Y(n15928) );
  sky130_fd_sc_hd__nand2_1 U23002 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[121]), .Y(n15927) );
  sky130_fd_sc_hd__nand2_1 U23003 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[409]), .Y(n15926) );
  sky130_fd_sc_hd__nand4_1 U23004 ( .A(n15929), .B(n15928), .C(n15927), .D(
        n15926), .Y(n15930) );
  sky130_fd_sc_hd__nor2_1 U23005 ( .A(n15931), .B(n15930), .Y(n15939) );
  sky130_fd_sc_hd__a22oi_1 U23006 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[313]), .B1(n14724), .B2(
        j202_soc_core_j22_cpu_rf_gpr[473]), .Y(n15938) );
  sky130_fd_sc_hd__a22oi_1 U23007 ( .A1(n23515), .A2(
        j202_soc_core_j22_cpu_rf_gpr[217]), .B1(n16469), .B2(
        j202_soc_core_j22_cpu_rf_gpr[89]), .Y(n15937) );
  sky130_fd_sc_hd__nand2_1 U23008 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[281]), .Y(n15935) );
  sky130_fd_sc_hd__nand2_1 U23009 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[153]), .Y(n15934) );
  sky130_fd_sc_hd__nand2_1 U23010 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[377]), .Y(n15933) );
  sky130_fd_sc_hd__nand2_1 U23011 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[345]), .Y(n15932) );
  sky130_fd_sc_hd__and4_1 U23012 ( .A(n15935), .B(n15934), .C(n15933), .D(
        n15932), .X(n15936) );
  sky130_fd_sc_hd__nand4_1 U23013 ( .A(n15939), .B(n15938), .C(n15937), .D(
        n15936), .Y(n22884) );
  sky130_fd_sc_hd__nand2_1 U23014 ( .A(n22884), .B(n16513), .Y(n15949) );
  sky130_fd_sc_hd__nand2_1 U23015 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[25]), .Y(n15942) );
  sky130_fd_sc_hd__nand2_1 U23016 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[25]), .Y(n15941) );
  sky130_fd_sc_hd__nand2_1 U23017 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[505]), .Y(n15940) );
  sky130_fd_sc_hd__and4_1 U23018 ( .A(n15942), .B(n15941), .C(n16516), .D(
        n15940), .X(n15948) );
  sky130_fd_sc_hd__nand2_1 U23019 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[25]), .Y(n15946) );
  sky130_fd_sc_hd__nand2_1 U23020 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[25]), .Y(n15945) );
  sky130_fd_sc_hd__nand2_1 U23021 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[25]), .Y(n15944) );
  sky130_fd_sc_hd__nand2_1 U23022 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[25]), .Y(n15943) );
  sky130_fd_sc_hd__and4_1 U23023 ( .A(n15946), .B(n15945), .C(n15944), .D(
        n15943), .X(n15947) );
  sky130_fd_sc_hd__nand3_1 U23024 ( .A(n15949), .B(n15948), .C(n15947), .Y(
        n25122) );
  sky130_fd_sc_hd__nand2_1 U23025 ( .A(n25122), .B(n16529), .Y(n15950) );
  sky130_fd_sc_hd__nor2_1 U23027 ( .A(n15954), .B(n15955), .Y(n16531) );
  sky130_fd_sc_hd__nand2_1 U23028 ( .A(n16532), .B(n16152), .Y(n15958) );
  sky130_fd_sc_hd__nor2_1 U23029 ( .A(n15958), .B(n17108), .Y(n15960) );
  sky130_fd_sc_hd__o21ai_1 U23030 ( .A1(n15953), .A2(n15952), .B1(n15951), .Y(
        n16538) );
  sky130_fd_sc_hd__nand2_1 U23031 ( .A(n15955), .B(n15954), .Y(n16536) );
  sky130_fd_sc_hd__a21oi_1 U23032 ( .A1(n16538), .A2(n16152), .B1(n15956), .Y(
        n15957) );
  sky130_fd_sc_hd__o21ai_1 U23033 ( .A1(n15958), .A2(n17110), .B1(n15957), .Y(
        n15959) );
  sky130_fd_sc_hd__a21oi_1 U23034 ( .A1(n22513), .A2(n15960), .B1(n15959), .Y(
        n16026) );
  sky130_fd_sc_hd__nand2_1 U23035 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[410]), .Y(n15964) );
  sky130_fd_sc_hd__nand2_1 U23036 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[474]), .Y(n15963) );
  sky130_fd_sc_hd__nand2_1 U23037 ( .A(n16431), .B(
        j202_soc_core_j22_cpu_rf_gpr[282]), .Y(n15962) );
  sky130_fd_sc_hd__nand2_1 U23038 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[154]), .Y(n15961) );
  sky130_fd_sc_hd__nand4_1 U23039 ( .A(n15964), .B(n15963), .C(n15962), .D(
        n15961), .Y(n15970) );
  sky130_fd_sc_hd__a21oi_1 U23040 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[26]), .B1(n16436), .Y(n15968) );
  sky130_fd_sc_hd__nand2_1 U23041 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[122]), .Y(n15967) );
  sky130_fd_sc_hd__nand2_1 U23042 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[58]), .Y(n15966) );
  sky130_fd_sc_hd__nand2_1 U23043 ( .A(n14204), .B(
        j202_soc_core_j22_cpu_rf_gpr[90]), .Y(n15965) );
  sky130_fd_sc_hd__nand4_1 U23044 ( .A(n15968), .B(n15967), .C(n15966), .D(
        n15965), .Y(n15969) );
  sky130_fd_sc_hd__nor2_1 U23045 ( .A(n15970), .B(n15969), .Y(n15981) );
  sky130_fd_sc_hd__nand2_1 U23046 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[442]), .Y(n15974) );
  sky130_fd_sc_hd__nand2_1 U23047 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[250]), .Y(n15973) );
  sky130_fd_sc_hd__nand2_1 U23048 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[218]), .Y(n15972) );
  sky130_fd_sc_hd__nand2_1 U23049 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[314]), .Y(n15971) );
  sky130_fd_sc_hd__nand2_1 U23050 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[506]), .Y(n15978) );
  sky130_fd_sc_hd__nand2_1 U23051 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[186]), .Y(n15977) );
  sky130_fd_sc_hd__nand2_1 U23052 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[346]), .Y(n15976) );
  sky130_fd_sc_hd__nand2_1 U23053 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[378]), .Y(n15975) );
  sky130_fd_sc_hd__nand4_1 U23054 ( .A(n15978), .B(n15977), .C(n15976), .D(
        n15975), .Y(n15979) );
  sky130_fd_sc_hd__a21oi_1 U23055 ( .A1(j202_soc_core_j22_cpu_rf_gpr[26]), 
        .A2(n16285), .B1(n15979), .Y(n15980) );
  sky130_fd_sc_hd__nand3_1 U23056 ( .A(n15981), .B(n13291), .C(n15980), .Y(
        n26718) );
  sky130_fd_sc_hd__inv_2 U23057 ( .A(n26718), .Y(n26563) );
  sky130_fd_sc_hd__o22ai_1 U23058 ( .A1(n16492), .A2(n26563), .B1(n26706), 
        .B2(n13793), .Y(n16022) );
  sky130_fd_sc_hd__nand2_1 U23059 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[186]), .Y(n15987) );
  sky130_fd_sc_hd__nand2_1 U23060 ( .A(n15982), .B(
        j202_soc_core_j22_cpu_rf_gpr[250]), .Y(n15986) );
  sky130_fd_sc_hd__nand2_1 U23061 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[506]), .Y(n15985) );
  sky130_fd_sc_hd__nand2_1 U23062 ( .A(n15983), .B(
        j202_soc_core_j22_cpu_rf_gpr[442]), .Y(n15984) );
  sky130_fd_sc_hd__nand4_1 U23063 ( .A(n15987), .B(n15986), .C(n15985), .D(
        n15984), .Y(n15993) );
  sky130_fd_sc_hd__nand2_1 U23064 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[26]), .Y(n15991) );
  sky130_fd_sc_hd__nand2_1 U23065 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[58]), .Y(n15990) );
  sky130_fd_sc_hd__nand2_1 U23066 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[122]), .Y(n15989) );
  sky130_fd_sc_hd__nand2_1 U23067 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[410]), .Y(n15988) );
  sky130_fd_sc_hd__nand4_1 U23068 ( .A(n15991), .B(n15990), .C(n15989), .D(
        n15988), .Y(n15992) );
  sky130_fd_sc_hd__nor2_1 U23069 ( .A(n15993), .B(n15992), .Y(n16004) );
  sky130_fd_sc_hd__nand2_1 U23070 ( .A(n16469), .B(
        j202_soc_core_j22_cpu_rf_gpr[90]), .Y(n15997) );
  sky130_fd_sc_hd__nand2_1 U23071 ( .A(n23515), .B(
        j202_soc_core_j22_cpu_rf_gpr[218]), .Y(n15996) );
  sky130_fd_sc_hd__nand2_1 U23072 ( .A(n11160), .B(
        j202_soc_core_j22_cpu_rf_gpr[314]), .Y(n15995) );
  sky130_fd_sc_hd__nand2_1 U23073 ( .A(n14414), .B(
        j202_soc_core_j22_cpu_rf_gpr[474]), .Y(n15994) );
  sky130_fd_sc_hd__and4_1 U23074 ( .A(n15997), .B(n15996), .C(n15995), .D(
        n15994), .X(n16003) );
  sky130_fd_sc_hd__nand2_1 U23075 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[282]), .Y(n16001) );
  sky130_fd_sc_hd__nand2_1 U23076 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[154]), .Y(n16000) );
  sky130_fd_sc_hd__nand2_1 U23077 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[378]), .Y(n15999) );
  sky130_fd_sc_hd__nand2_1 U23078 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[346]), .Y(n15998) );
  sky130_fd_sc_hd__and4_1 U23079 ( .A(n16001), .B(n16000), .C(n15999), .D(
        n15998), .X(n16002) );
  sky130_fd_sc_hd__nand3_1 U23080 ( .A(n16004), .B(n16003), .C(n16002), .Y(
        n22376) );
  sky130_fd_sc_hd__a21oi_1 U23081 ( .A1(n29567), .A2(
        j202_soc_core_j22_cpu_rf_vbr[26]), .B1(n16005), .Y(n16019) );
  sky130_fd_sc_hd__a2bb2oi_1 U23082 ( .B1(j202_soc_core_j22_cpu_rf_gpr[506]), 
        .B2(n29563), .A1_N(n16007), .A2_N(n16006), .Y(n16018) );
  sky130_fd_sc_hd__o22a_1 U23083 ( .A1(n16011), .A2(n16010), .B1(n16009), .B2(
        n16008), .X(n16017) );
  sky130_fd_sc_hd__o22a_1 U23084 ( .A1(n16015), .A2(n16014), .B1(n16013), .B2(
        n11095), .X(n16016) );
  sky130_fd_sc_hd__nand4_1 U23085 ( .A(n16019), .B(n16018), .C(n16017), .D(
        n16016), .Y(n16020) );
  sky130_fd_sc_hd__a21oi_1 U23086 ( .A1(n22376), .A2(n16513), .B1(n16020), .Y(
        n27380) );
  sky130_fd_sc_hd__nand2_1 U23087 ( .A(n27380), .B(n16322), .Y(n16021) );
  sky130_fd_sc_hd__o21ai_1 U23088 ( .A1(n16320), .A2(n27380), .B1(n16021), .Y(
        n16023) );
  sky130_fd_sc_hd__nor2_1 U23089 ( .A(n16022), .B(n16023), .Y(n16535) );
  sky130_fd_sc_hd__nand2_1 U23090 ( .A(n16023), .B(n16022), .Y(n16534) );
  sky130_fd_sc_hd__nand2_1 U23091 ( .A(n16024), .B(n16534), .Y(n16025) );
  sky130_fd_sc_hd__xor2_1 U23092 ( .A(n16026), .B(n16025), .X(n25070) );
  sky130_fd_sc_hd__nand2_1 U23093 ( .A(n25070), .B(n12158), .Y(n16034) );
  sky130_fd_sc_hd__nor2_1 U23094 ( .A(n16028), .B(n16027), .Y(n16030) );
  sky130_fd_sc_hd__o22a_1 U23095 ( .A1(n27380), .A2(n22590), .B1(n26563), .B2(
        n11143), .X(n16031) );
  sky130_fd_sc_hd__a21oi_1 U23097 ( .A1(n25077), .A2(n22596), .B1(n16032), .Y(
        n16033) );
  sky130_fd_sc_hd__nand2_1 U23098 ( .A(n26812), .B(n20428), .Y(n27165) );
  sky130_fd_sc_hd__nor2_1 U23099 ( .A(j202_soc_core_j22_cpu_pc[1]), .B(n24474), 
        .Y(n20548) );
  sky130_fd_sc_hd__a211o_1 U23100 ( .A1(j202_soc_core_j22_cpu_id_opn_v_), .A2(
        n27165), .B1(n20548), .C1(n28965), .X(n16037) );
  sky130_fd_sc_hd__mux2i_1 U23101 ( .A0(n16037), .A1(n16036), .S(n27914), .Y(
        n16053) );
  sky130_fd_sc_hd__nand3_1 U23102 ( .A(n29347), .B(n27955), .C(n27166), .Y(
        n16051) );
  sky130_fd_sc_hd__a2bb2oi_1 U23103 ( .B1(j202_soc_core_intr_level__2_), .B2(
        n21553), .A1_N(n16038), .A2_N(j202_soc_core_j22_cpu_rfuo_sr__i__3_), 
        .Y(n16046) );
  sky130_fd_sc_hd__nand2_1 U23104 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__1_), 
        .B(n16041), .Y(n16039) );
  sky130_fd_sc_hd__nand3_1 U23105 ( .A(n16039), .B(n19451), .C(
        j202_soc_core_intr_level__0_), .Y(n16040) );
  sky130_fd_sc_hd__nand2_1 U23107 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__2_), 
        .B(n16042), .Y(n16043) );
  sky130_fd_sc_hd__nand2_1 U23108 ( .A(n16044), .B(n16043), .Y(n16045) );
  sky130_fd_sc_hd__a2bb2oi_1 U23109 ( .B1(n16046), .B2(n16045), .A1_N(
        j202_soc_core_intr_level__3_), .A2_N(n19043), .Y(n16047) );
  sky130_fd_sc_hd__o21a_1 U23110 ( .A1(j202_soc_core_intr_level__4_), .A2(
        n16047), .B1(j202_soc_core_intr_req_), .X(n27915) );
  sky130_fd_sc_hd__nand2b_1 U23111 ( .A_N(n14849), .B(n27915), .Y(n27906) );
  sky130_fd_sc_hd__nand2_1 U23112 ( .A(n12200), .B(n24474), .Y(n24466) );
  sky130_fd_sc_hd__o211a_2 U23113 ( .A1(n20547), .A2(n24430), .B1(n12142), 
        .C1(n24466), .X(n16050) );
  sky130_fd_sc_hd__nand3_1 U23114 ( .A(n26812), .B(n16054), .C(n20273), .Y(
        n16049) );
  sky130_fd_sc_hd__nand3_1 U23115 ( .A(n27906), .B(n16050), .C(n16049), .Y(
        n23484) );
  sky130_fd_sc_hd__nor2_1 U23116 ( .A(n16051), .B(n23484), .Y(n16052) );
  sky130_fd_sc_hd__nand2_1 U23117 ( .A(n27720), .B(n23299), .Y(n27602) );
  sky130_fd_sc_hd__a22oi_1 U23118 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[57]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[89]), .Y(n16137) );
  sky130_fd_sc_hd__nand2_1 U23119 ( .A(n21675), .B(j202_soc_core_uart_div0[1]), 
        .Y(n16136) );
  sky130_fd_sc_hd__nand2_1 U23120 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[25]), .Y(n16135) );
  sky130_fd_sc_hd__nand4_1 U23121 ( .A(n16137), .B(n21677), .C(n16136), .D(
        n16135), .Y(n16133) );
  sky130_fd_sc_hd__nor3_1 U23122 ( .A(n16056), .B(n16055), .C(n16101), .Y(
        n17063) );
  sky130_fd_sc_hd__a31oi_1 U23123 ( .A1(n16058), .A2(n17063), .A3(n16057), 
        .B1(n17055), .Y(n16071) );
  sky130_fd_sc_hd__nand4_1 U23124 ( .A(n17077), .B(n16064), .C(n16060), .D(
        n16063), .Y(n16061) );
  sky130_fd_sc_hd__o21ai_1 U23125 ( .A1(n16062), .A2(n16061), .B1(n17273), .Y(
        n16070) );
  sky130_fd_sc_hd__nand4b_1 U23126 ( .A_N(n17035), .B(n16065), .C(n16064), .D(
        n16063), .Y(n16066) );
  sky130_fd_sc_hd__nand2_1 U23127 ( .A(n13387), .B(n16066), .Y(n16069) );
  sky130_fd_sc_hd__o21ai_1 U23128 ( .A1(n17031), .A2(n16067), .B1(n13388), .Y(
        n16068) );
  sky130_fd_sc_hd__nand4b_1 U23129 ( .A_N(n16071), .B(n16070), .C(n16069), .D(
        n16068), .Y(n16072) );
  sky130_fd_sc_hd__nand2_1 U23130 ( .A(n16072), .B(n17094), .Y(n16088) );
  sky130_fd_sc_hd__nand2_1 U23131 ( .A(n16074), .B(n13305), .Y(n16076) );
  sky130_fd_sc_hd__nand4_1 U23133 ( .A(n17005), .B(n17007), .C(n16078), .D(
        n16077), .Y(n16079) );
  sky130_fd_sc_hd__nand2_1 U23134 ( .A(n16079), .B(n13387), .Y(n16083) );
  sky130_fd_sc_hd__o21ai_1 U23135 ( .A1(n16081), .A2(n16080), .B1(n13388), .Y(
        n16082) );
  sky130_fd_sc_hd__nand3_1 U23136 ( .A(n16084), .B(n16083), .C(n16082), .Y(
        n16086) );
  sky130_fd_sc_hd__o21ai_1 U23137 ( .A1(n16086), .A2(n16085), .B1(n17021), .Y(
        n16087) );
  sky130_fd_sc_hd__nand2_1 U23138 ( .A(n16088), .B(n16087), .Y(n16089) );
  sky130_fd_sc_hd__nand2_1 U23139 ( .A(n16089), .B(n17098), .Y(n16138) );
  sky130_fd_sc_hd__a21oi_1 U23140 ( .A1(n13294), .A2(n16090), .B1(n16094), .Y(
        n16092) );
  sky130_fd_sc_hd__a31oi_1 U23141 ( .A1(n16093), .A2(n16092), .A3(n16091), 
        .B1(n17037), .Y(n16109) );
  sky130_fd_sc_hd__nor4_1 U23142 ( .A(n13306), .B(n16095), .C(n16094), .D(
        n16101), .Y(n16097) );
  sky130_fd_sc_hd__a31oi_1 U23143 ( .A1(n16097), .A2(n16096), .A3(n16099), 
        .B1(n17039), .Y(n16108) );
  sky130_fd_sc_hd__nand3_1 U23144 ( .A(n16100), .B(n16099), .C(n16098), .Y(
        n17089) );
  sky130_fd_sc_hd__nor3_1 U23145 ( .A(n16102), .B(n16101), .C(n17089), .Y(
        n16103) );
  sky130_fd_sc_hd__a21oi_1 U23146 ( .A1(n17028), .A2(n16103), .B1(n17078), .Y(
        n16107) );
  sky130_fd_sc_hd__a21oi_1 U23147 ( .A1(n16105), .A2(n16104), .B1(n17055), .Y(
        n16106) );
  sky130_fd_sc_hd__nor4_1 U23148 ( .A(n16109), .B(n16108), .C(n16107), .D(
        n16106), .Y(n16131) );
  sky130_fd_sc_hd__nand3b_1 U23149 ( .A_N(n16111), .B(n17014), .C(n16110), .Y(
        n16112) );
  sky130_fd_sc_hd__a31oi_1 U23150 ( .A1(n16115), .A2(n16114), .A3(n16113), 
        .B1(n17078), .Y(n16124) );
  sky130_fd_sc_hd__o31a_1 U23151 ( .A1(n16118), .A2(n16117), .A3(n16116), .B1(
        n13388), .X(n16123) );
  sky130_fd_sc_hd__nor2_1 U23152 ( .A(n16119), .B(n17045), .Y(n16120) );
  sky130_fd_sc_hd__a31oi_1 U23153 ( .A1(n16121), .A2(n17042), .A3(n16120), 
        .B1(n17039), .Y(n16122) );
  sky130_fd_sc_hd__nor3_1 U23154 ( .A(n16124), .B(n16123), .C(n16122), .Y(
        n16129) );
  sky130_fd_sc_hd__a21oi_1 U23155 ( .A1(n16126), .A2(n17301), .B1(n16125), .Y(
        n16127) );
  sky130_fd_sc_hd__a21oi_1 U23156 ( .A1(n16127), .A2(n17049), .B1(n17055), .Y(
        n16128) );
  sky130_fd_sc_hd__nor2b_1 U23157 ( .B_N(n16129), .A(n16128), .Y(n16130) );
  sky130_fd_sc_hd__mux2i_1 U23158 ( .A0(n16131), .A1(n16130), .S(n20787), .Y(
        n16132) );
  sky130_fd_sc_hd__nand2_1 U23159 ( .A(n16132), .B(n20626), .Y(n16141) );
  sky130_fd_sc_hd__nand3b_1 U23160 ( .A_N(n16133), .B(n16138), .C(n16141), .Y(
        n16134) );
  sky130_fd_sc_hd__nand2_1 U23161 ( .A(j202_soc_core_memory0_ram_dout0[505]), 
        .B(n21771), .Y(n16143) );
  sky130_fd_sc_hd__nand4_1 U23162 ( .A(n16137), .B(n21738), .C(n16136), .D(
        n16135), .Y(n16140) );
  sky130_fd_sc_hd__nor2_1 U23163 ( .A(n16140), .B(n16139), .Y(n16142) );
  sky130_fd_sc_hd__nand3_1 U23164 ( .A(n16143), .B(n16142), .C(n16141), .Y(
        n16144) );
  sky130_fd_sc_hd__nand2_1 U23165 ( .A(n22515), .B(n25122), .Y(n16147) );
  sky130_fd_sc_hd__ha_1 U23166 ( .A(n16145), .B(j202_soc_core_j22_cpu_pc[25]), 
        .COUT(n16157), .SUM(n25188) );
  sky130_fd_sc_hd__nand2_1 U23167 ( .A(n22596), .B(n25188), .Y(n16146) );
  sky130_fd_sc_hd__o211a_2 U23168 ( .A1(n26706), .A2(n11143), .B1(n16147), 
        .C1(n16146), .X(n16156) );
  sky130_fd_sc_hd__nor2_1 U23169 ( .A(n16149), .B(n17108), .Y(n16151) );
  sky130_fd_sc_hd__o21ai_1 U23170 ( .A1(n16149), .A2(n17110), .B1(n16148), .Y(
        n16150) );
  sky130_fd_sc_hd__a21oi_1 U23171 ( .A1(n22513), .A2(n16151), .B1(n16150), .Y(
        n16154) );
  sky130_fd_sc_hd__nand2_1 U23172 ( .A(n16152), .B(n16536), .Y(n16153) );
  sky130_fd_sc_hd__xor2_1 U23173 ( .A(n16154), .B(n16153), .X(n25136) );
  sky130_fd_sc_hd__nand2_1 U23174 ( .A(n25136), .B(n12158), .Y(n16155) );
  sky130_fd_sc_hd__ha_1 U23175 ( .A(n16157), .B(j202_soc_core_j22_cpu_pc[26]), 
        .COUT(n17118), .SUM(n25077) );
  sky130_fd_sc_hd__xor2_1 U23176 ( .A(j202_soc_core_j22_cpu_pc[31]), .B(n16158), .X(n26887) );
  sky130_fd_sc_hd__nand2_1 U23177 ( .A(n17175), .B(n20687), .Y(n16964) );
  sky130_fd_sc_hd__nand2_1 U23178 ( .A(n16616), .B(n20579), .Y(n16174) );
  sky130_fd_sc_hd__nand2b_1 U23179 ( .A_N(n16174), .B(n16180), .Y(n16879) );
  sky130_fd_sc_hd__nor2_1 U23180 ( .A(n20579), .B(n16159), .Y(n16615) );
  sky130_fd_sc_hd__nand2b_1 U23181 ( .A_N(n16162), .B(n16615), .Y(n16714) );
  sky130_fd_sc_hd__nand2_1 U23182 ( .A(n16879), .B(n16714), .Y(n16855) );
  sky130_fd_sc_hd__nand2_1 U23183 ( .A(n16180), .B(n16615), .Y(n16577) );
  sky130_fd_sc_hd__nand2_1 U23184 ( .A(n19085), .B(n17301), .Y(n20350) );
  sky130_fd_sc_hd__nand2b_1 U23185 ( .A_N(n20350), .B(n17293), .Y(n16578) );
  sky130_fd_sc_hd__nand2_1 U23186 ( .A(n16577), .B(n16578), .Y(n16787) );
  sky130_fd_sc_hd__nand2_1 U23187 ( .A(n17161), .B(n20579), .Y(n16177) );
  sky130_fd_sc_hd__nand2b_1 U23188 ( .A_N(n16177), .B(n16180), .Y(n16689) );
  sky130_fd_sc_hd__nand2_1 U23189 ( .A(n16616), .B(
        j202_soc_core_bootrom_00_address_w[11]), .Y(n19874) );
  sky130_fd_sc_hd__nand2b_1 U23190 ( .A_N(n19874), .B(n17067), .Y(n16849) );
  sky130_fd_sc_hd__nand2_1 U23191 ( .A(n16689), .B(n16849), .Y(n16620) );
  sky130_fd_sc_hd__nor2_1 U23192 ( .A(n16855), .B(n16715), .Y(n16703) );
  sky130_fd_sc_hd__nand2_1 U23193 ( .A(n20687), .B(n12137), .Y(n16611) );
  sky130_fd_sc_hd__nor2_1 U23194 ( .A(n16160), .B(n16177), .Y(n16858) );
  sky130_fd_sc_hd__nand2_1 U23195 ( .A(n16171), .B(n20788), .Y(n16202) );
  sky130_fd_sc_hd__nand2b_1 U23196 ( .A_N(n16162), .B(n16161), .Y(n16173) );
  sky130_fd_sc_hd__nand2_1 U23197 ( .A(n16182), .B(n20579), .Y(n16770) );
  sky130_fd_sc_hd__nand2_1 U23198 ( .A(n16770), .B(n16578), .Y(n16751) );
  sky130_fd_sc_hd__nor3_1 U23199 ( .A(n16858), .B(n16745), .C(n16751), .Y(
        n16167) );
  sky130_fd_sc_hd__nand2_1 U23200 ( .A(n17044), .B(n17287), .Y(n16691) );
  sky130_fd_sc_hd__nand2_1 U23201 ( .A(n16164), .B(n16163), .Y(n16935) );
  sky130_fd_sc_hd__nand2_1 U23202 ( .A(n16935), .B(n16578), .Y(n16198) );
  sky130_fd_sc_hd__nand2_1 U23203 ( .A(n16691), .B(n16165), .Y(n16215) );
  sky130_fd_sc_hd__nor2_1 U23204 ( .A(n12137), .B(n20687), .Y(n16956) );
  sky130_fd_sc_hd__nand2_1 U23205 ( .A(n16935), .B(n16692), .Y(n16856) );
  sky130_fd_sc_hd__nand2_1 U23206 ( .A(n12137), .B(n20623), .Y(n16596) );
  sky130_fd_sc_hd__a22oi_1 U23207 ( .A1(n16215), .A2(n16956), .B1(n16856), 
        .B2(n16945), .Y(n16166) );
  sky130_fd_sc_hd__o21ai_1 U23208 ( .A1(n16611), .A2(n16167), .B1(n16166), .Y(
        n16168) );
  sky130_fd_sc_hd__o21bai_1 U23209 ( .A1(n16964), .A2(n16703), .B1_N(n16168), 
        .Y(n16169) );
  sky130_fd_sc_hd__nand2_1 U23210 ( .A(n16169), .B(n20908), .Y(n16235) );
  sky130_fd_sc_hd__nor2_1 U23211 ( .A(n20787), .B(n16170), .Y(n17170) );
  sky130_fd_sc_hd__nor2_1 U23212 ( .A(n17289), .B(n21206), .Y(n16882) );
  sky130_fd_sc_hd__nand2_1 U23213 ( .A(n16171), .B(n19354), .Y(n17166) );
  sky130_fd_sc_hd__nand2_1 U23214 ( .A(n16172), .B(n17193), .Y(n16685) );
  sky130_fd_sc_hd__nand2_1 U23215 ( .A(n16202), .B(n16174), .Y(n16846) );
  sky130_fd_sc_hd__nand2_1 U23216 ( .A(n16846), .B(n16180), .Y(n16734) );
  sky130_fd_sc_hd__nand2b_1 U23217 ( .A_N(n16953), .B(n20579), .Y(n16782) );
  sky130_fd_sc_hd__nand4_1 U23218 ( .A(n16173), .B(n16685), .C(n16734), .D(
        n16782), .Y(n16835) );
  sky130_fd_sc_hd__nor4_1 U23219 ( .A(n16882), .B(n16196), .C(n16216), .D(
        n16835), .Y(n16179) );
  sky130_fd_sc_hd__nand3_1 U23220 ( .A(n16564), .B(
        j202_soc_core_bootrom_00_address_w[4]), .C(
        j202_soc_core_bootrom_00_address_w[11]), .Y(n16872) );
  sky130_fd_sc_hd__nand2_1 U23221 ( .A(n16872), .B(n20633), .Y(n16857) );
  sky130_fd_sc_hd__nor2_1 U23222 ( .A(n16583), .B(n16174), .Y(n16773) );
  sky130_fd_sc_hd__nor2b_1 U23223 ( .B_N(n16675), .A(n16773), .Y(n16702) );
  sky130_fd_sc_hd__nor2_1 U23224 ( .A(n16202), .B(n16583), .Y(n16677) );
  sky130_fd_sc_hd__nand2_1 U23225 ( .A(n16840), .B(n20788), .Y(n16844) );
  sky130_fd_sc_hd__nand2b_1 U23226 ( .A_N(n16677), .B(n16844), .Y(n16175) );
  sky130_fd_sc_hd__nand2_1 U23227 ( .A(n16691), .B(n16689), .Y(n16890) );
  sky130_fd_sc_hd__nand2_1 U23228 ( .A(n16615), .B(n16176), .Y(n16880) );
  sky130_fd_sc_hd__nor2_1 U23229 ( .A(n16583), .B(n16177), .Y(n16576) );
  sky130_fd_sc_hd__nor2_1 U23230 ( .A(n16745), .B(n16576), .Y(n16742) );
  sky130_fd_sc_hd__nor2_1 U23231 ( .A(n17293), .B(n21206), .Y(n16891) );
  sky130_fd_sc_hd__nor2_1 U23232 ( .A(n16891), .B(n16881), .Y(n16605) );
  sky130_fd_sc_hd__nand3_1 U23233 ( .A(n16880), .B(n16742), .C(n16605), .Y(
        n16189) );
  sky130_fd_sc_hd__nor4bb_1 U23234 ( .C_N(n16702), .D_N(n16785), .A(n16890), 
        .B(n16189), .Y(n16178) );
  sky130_fd_sc_hd__o22ai_1 U23235 ( .A1(n16179), .A2(n16596), .B1(n16178), 
        .B2(n16964), .Y(n16188) );
  sky130_fd_sc_hd__nor2_1 U23236 ( .A(n16202), .B(n16181), .Y(n16690) );
  sky130_fd_sc_hd__nor2_1 U23237 ( .A(n20788), .B(n20463), .Y(n16911) );
  sky130_fd_sc_hd__nand3b_1 U23238 ( .A_N(n16690), .B(n16578), .C(n16947), .Y(
        n16721) );
  sky130_fd_sc_hd__nand2_1 U23239 ( .A(n16182), .B(n20788), .Y(n16201) );
  sky130_fd_sc_hd__nor2_1 U23240 ( .A(n16677), .B(n16619), .Y(n16566) );
  sky130_fd_sc_hd__nand2_1 U23241 ( .A(n16566), .B(n16685), .Y(n16560) );
  sky130_fd_sc_hd__nand2b_1 U23242 ( .A_N(n16583), .B(n16615), .Y(n16598) );
  sky130_fd_sc_hd__nor2_1 U23243 ( .A(n16560), .B(n16842), .Y(n16191) );
  sky130_fd_sc_hd__nand2b_1 U23244 ( .A_N(n17166), .B(n16564), .Y(n16903) );
  sky130_fd_sc_hd__nand2b_1 U23245 ( .A_N(n17165), .B(n19125), .Y(n20784) );
  sky130_fd_sc_hd__nor2_1 U23246 ( .A(n17289), .B(n20784), .Y(n16905) );
  sky130_fd_sc_hd__nand2b_1 U23247 ( .A_N(n20463), .B(n20788), .Y(n16934) );
  sky130_fd_sc_hd__nand2b_1 U23248 ( .A_N(n16905), .B(n16934), .Y(n16744) );
  sky130_fd_sc_hd__nor2_1 U23249 ( .A(n16735), .B(n16744), .Y(n16688) );
  sky130_fd_sc_hd__nand2b_1 U23250 ( .A_N(n16773), .B(n16577), .Y(n16594) );
  sky130_fd_sc_hd__nor2_1 U23251 ( .A(n16891), .B(n16594), .Y(n16558) );
  sky130_fd_sc_hd__nand2_1 U23252 ( .A(n16688), .B(n16558), .Y(n16853) );
  sky130_fd_sc_hd__nand2_1 U23253 ( .A(n16191), .B(n16183), .Y(n16186) );
  sky130_fd_sc_hd__nand2_1 U23254 ( .A(n16691), .B(n16849), .Y(n16185) );
  sky130_fd_sc_hd__nand2_1 U23255 ( .A(n11994), .B(n20788), .Y(n16184) );
  sky130_fd_sc_hd__nor2_1 U23256 ( .A(n16184), .B(n16583), .Y(n16674) );
  sky130_fd_sc_hd__nand2_1 U23257 ( .A(n16674), .B(n17314), .Y(n16954) );
  sky130_fd_sc_hd__nor2_1 U23258 ( .A(n20788), .B(n16682), .Y(n16769) );
  sky130_fd_sc_hd__nand2_1 U23259 ( .A(n16954), .B(n16778), .Y(n16720) );
  sky130_fd_sc_hd__nor2_1 U23260 ( .A(n16185), .B(n16720), .Y(n16754) );
  sky130_fd_sc_hd__nand2_1 U23261 ( .A(n16754), .B(n16782), .Y(n16960) );
  sky130_fd_sc_hd__o31a_1 U23262 ( .A1(n16721), .A2(n16186), .A3(n16960), .B1(
        n16956), .X(n16187) );
  sky130_fd_sc_hd__o21a_1 U23263 ( .A1(n16188), .A2(n16187), .B1(n13481), .X(
        n16231) );
  sky130_fd_sc_hd__nand2_1 U23264 ( .A(n16688), .B(n16190), .Y(n16870) );
  sky130_fd_sc_hd__nor2_1 U23265 ( .A(n20788), .B(n16722), .Y(n16838) );
  sky130_fd_sc_hd__nor2_1 U23266 ( .A(n16838), .B(n16858), .Y(n16698) );
  sky130_fd_sc_hd__nand3b_1 U23267 ( .A_N(n16870), .B(n16191), .C(n16698), .Y(
        n16192) );
  sky130_fd_sc_hd__nand2_1 U23268 ( .A(n16192), .B(n16937), .Y(n16229) );
  sky130_fd_sc_hd__o2bb2ai_1 U23269 ( .B1(n27043), .B2(n20860), .A1_N(n21676), 
        .A2_N(j202_soc_core_ahblite_interconnect_s_hrdata[31]), .Y(n16193) );
  sky130_fd_sc_hd__a21oi_1 U23270 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[63]), .B1(n16193), .Y(
        n16228) );
  sky130_fd_sc_hd__nand2_1 U23271 ( .A(n21666), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[95]), .Y(n16227) );
  sky130_fd_sc_hd__nand4_1 U23272 ( .A(n16229), .B(n16228), .C(n21677), .D(
        n16227), .Y(n16194) );
  sky130_fd_sc_hd__nor2_1 U23273 ( .A(n16231), .B(n16194), .Y(n16226) );
  sky130_fd_sc_hd__nor2_1 U23274 ( .A(n16911), .B(n16838), .Y(n16915) );
  sky130_fd_sc_hd__nand4_1 U23275 ( .A(n16558), .B(n16915), .C(n16195), .D(
        n16844), .Y(n16199) );
  sky130_fd_sc_hd__nor2_1 U23276 ( .A(n16576), .B(n16882), .Y(n16948) );
  sky130_fd_sc_hd__nor2_1 U23277 ( .A(n16196), .B(n16744), .Y(n16622) );
  sky130_fd_sc_hd__nand2b_1 U23278 ( .A_N(n19121), .B(n16197), .Y(n16740) );
  sky130_fd_sc_hd__nand4b_1 U23279 ( .A_N(n16198), .B(n16948), .C(n16622), .D(
        n16740), .Y(n16614) );
  sky130_fd_sc_hd__o21ai_1 U23280 ( .A1(n16199), .A2(n16614), .B1(n16945), .Y(
        n16212) );
  sky130_fd_sc_hd__nand2_1 U23281 ( .A(n16691), .B(n16685), .Y(n16788) );
  sky130_fd_sc_hd__nor2_1 U23282 ( .A(n16576), .B(n16788), .Y(n16200) );
  sky130_fd_sc_hd__nand3_1 U23283 ( .A(n16201), .B(n16200), .C(n21206), .Y(
        n16204) );
  sky130_fd_sc_hd__o21a_1 U23284 ( .A1(n16202), .A2(n16845), .B1(n16770), .X(
        n16203) );
  sky130_fd_sc_hd__nand3_1 U23285 ( .A(n16915), .B(n16203), .C(n16783), .Y(
        n16617) );
  sky130_fd_sc_hd__o21ai_1 U23286 ( .A1(n16204), .A2(n16617), .B1(n16924), .Y(
        n16211) );
  sky130_fd_sc_hd__nor2_1 U23287 ( .A(n16674), .B(n16882), .Y(n16913) );
  sky130_fd_sc_hd__nand2_1 U23288 ( .A(n16913), .B(n16205), .Y(n16697) );
  sky130_fd_sc_hd__nand2b_1 U23289 ( .A_N(n16891), .B(n16934), .Y(n16914) );
  sky130_fd_sc_hd__nor2_1 U23290 ( .A(n16745), .B(n16594), .Y(n16775) );
  sky130_fd_sc_hd__nand4b_1 U23291 ( .A_N(n16914), .B(n16775), .C(n16562), .D(
        n16880), .Y(n16206) );
  sky130_fd_sc_hd__o21ai_1 U23292 ( .A1(n16697), .A2(n16206), .B1(n16919), .Y(
        n16210) );
  sky130_fd_sc_hd__nor2_1 U23293 ( .A(n16207), .B(n16890), .Y(n16949) );
  sky130_fd_sc_hd__nor2_1 U23294 ( .A(n16745), .B(n16773), .Y(n16612) );
  sky130_fd_sc_hd__nand2_1 U23295 ( .A(n16844), .B(n16740), .Y(n16673) );
  sky130_fd_sc_hd__nand3_1 U23296 ( .A(n16612), .B(n16886), .C(n16904), .Y(
        n16878) );
  sky130_fd_sc_hd__nor2_1 U23297 ( .A(n16764), .B(n16878), .Y(n16717) );
  sky130_fd_sc_hd__nand3_1 U23298 ( .A(n16949), .B(n16699), .C(n16717), .Y(
        n16208) );
  sky130_fd_sc_hd__nand2_1 U23299 ( .A(n16208), .B(n16956), .Y(n16209) );
  sky130_fd_sc_hd__nand4_1 U23300 ( .A(n16212), .B(n16211), .C(n16210), .D(
        n16209), .Y(n16213) );
  sky130_fd_sc_hd__nand2_1 U23301 ( .A(n16213), .B(n21697), .Y(n16234) );
  sky130_fd_sc_hd__nand2b_1 U23302 ( .A_N(n16713), .B(n16577), .Y(n16941) );
  sky130_fd_sc_hd__nor2_1 U23303 ( .A(n16838), .B(n16914), .Y(n16574) );
  sky130_fd_sc_hd__nand4b_1 U23304 ( .A_N(n16941), .B(n16566), .C(n16574), .D(
        n16740), .Y(n16214) );
  sky130_fd_sc_hd__nand4_1 U23306 ( .A(n16754), .B(n16947), .C(n16722), .D(
        n16714), .Y(n16222) );
  sky130_fd_sc_hd__nor2_1 U23307 ( .A(n16216), .B(n16677), .Y(n16746) );
  sky130_fd_sc_hd__nor2b_1 U23308 ( .B_N(n16746), .A(n16576), .Y(n16723) );
  sky130_fd_sc_hd__nand2_1 U23309 ( .A(n16879), .B(n16723), .Y(n16940) );
  sky130_fd_sc_hd__nor4_1 U23310 ( .A(n16735), .B(n16619), .C(n16858), .D(
        n16940), .Y(n16220) );
  sky130_fd_sc_hd__nor2_1 U23311 ( .A(n17290), .B(n17166), .Y(n20863) );
  sky130_fd_sc_hd__nand3_1 U23312 ( .A(n16954), .B(n16873), .C(n16740), .Y(
        n16843) );
  sky130_fd_sc_hd__nand2b_1 U23313 ( .A_N(n16843), .B(n16953), .Y(n16681) );
  sky130_fd_sc_hd__nor4_1 U23314 ( .A(n20863), .B(n16677), .C(n16836), .D(
        n16681), .Y(n16217) );
  sky130_fd_sc_hd__nand2_1 U23315 ( .A(n16689), .B(n16217), .Y(n16218) );
  sky130_fd_sc_hd__nand2_1 U23316 ( .A(n16218), .B(n16924), .Y(n16219) );
  sky130_fd_sc_hd__o21ai_1 U23317 ( .A1(n16220), .A2(n16611), .B1(n16219), .Y(
        n16221) );
  sky130_fd_sc_hd__a21oi_1 U23318 ( .A1(n16222), .A2(n16956), .B1(n16221), .Y(
        n16223) );
  sky130_fd_sc_hd__nand2_1 U23319 ( .A(n16224), .B(n16223), .Y(n16225) );
  sky130_fd_sc_hd__nand2_1 U23320 ( .A(n16225), .B(n21727), .Y(n16232) );
  sky130_fd_sc_hd__nand2_1 U23321 ( .A(j202_soc_core_memory0_ram_dout0[511]), 
        .B(n21771), .Y(n16237) );
  sky130_fd_sc_hd__nand4_1 U23322 ( .A(n16229), .B(n16228), .C(n21738), .D(
        n16227), .Y(n16230) );
  sky130_fd_sc_hd__nor2_1 U23323 ( .A(n16231), .B(n16230), .Y(n16233) );
  sky130_fd_sc_hd__and3_1 U23324 ( .A(n16234), .B(n16233), .C(n16232), .X(
        n16236) );
  sky130_fd_sc_hd__nand3_1 U23325 ( .A(n16237), .B(n16236), .C(n16235), .Y(
        n18981) );
  sky130_fd_sc_hd__nand2_1 U23326 ( .A(n16431), .B(
        j202_soc_core_j22_cpu_rf_gpr[286]), .Y(n16241) );
  sky130_fd_sc_hd__nand2_1 U23327 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[478]), .Y(n16240) );
  sky130_fd_sc_hd__nand2_1 U23328 ( .A(n11150), .B(
        j202_soc_core_j22_cpu_rf_gpr[414]), .Y(n16239) );
  sky130_fd_sc_hd__nand2_1 U23329 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[158]), .Y(n16238) );
  sky130_fd_sc_hd__nand4_1 U23330 ( .A(n16241), .B(n16240), .C(n16239), .D(
        n16238), .Y(n16247) );
  sky130_fd_sc_hd__a21oi_1 U23331 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[30]), .B1(n16436), .Y(n16245) );
  sky130_fd_sc_hd__nand2_1 U23332 ( .A(n11152), .B(
        j202_soc_core_j22_cpu_rf_gpr[62]), .Y(n16244) );
  sky130_fd_sc_hd__nand2_1 U23333 ( .A(n11155), .B(
        j202_soc_core_j22_cpu_rf_gpr[94]), .Y(n16243) );
  sky130_fd_sc_hd__nand2_1 U23334 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[126]), .Y(n16242) );
  sky130_fd_sc_hd__nand4_1 U23335 ( .A(n16245), .B(n16244), .C(n16243), .D(
        n16242), .Y(n16246) );
  sky130_fd_sc_hd__nor2_1 U23336 ( .A(n16247), .B(n16246), .Y(n16260) );
  sky130_fd_sc_hd__nand2_1 U23337 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[446]), .Y(n16252) );
  sky130_fd_sc_hd__nand2_1 U23338 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[318]), .Y(n16251) );
  sky130_fd_sc_hd__nand2_1 U23339 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[254]), .Y(n16250) );
  sky130_fd_sc_hd__nand2_1 U23340 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_rf_gpr[222]), .Y(n16249) );
  sky130_fd_sc_hd__and4_1 U23341 ( .A(n16252), .B(n16251), .C(n16250), .D(
        n16249), .X(n16259) );
  sky130_fd_sc_hd__nand2_1 U23342 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[510]), .Y(n16256) );
  sky130_fd_sc_hd__nand2_1 U23343 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[190]), .Y(n16255) );
  sky130_fd_sc_hd__nand2_1 U23344 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[350]), .Y(n16254) );
  sky130_fd_sc_hd__nand2_1 U23345 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[382]), .Y(n16253) );
  sky130_fd_sc_hd__nand4_1 U23346 ( .A(n16256), .B(n16255), .C(n16254), .D(
        n16253), .Y(n16257) );
  sky130_fd_sc_hd__a21oi_1 U23347 ( .A1(j202_soc_core_j22_cpu_rf_gpr[30]), 
        .A2(n16369), .B1(n16257), .Y(n16258) );
  sky130_fd_sc_hd__nand2_1 U23348 ( .A(n26716), .B(n16261), .Y(n16291) );
  sky130_fd_sc_hd__nand2_1 U23349 ( .A(n11114), .B(
        j202_soc_core_j22_cpu_rf_gpr[415]), .Y(n16266) );
  sky130_fd_sc_hd__nand2_1 U23350 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[479]), .Y(n16265) );
  sky130_fd_sc_hd__nand2_1 U23351 ( .A(n16431), .B(
        j202_soc_core_j22_cpu_rf_gpr[287]), .Y(n16264) );
  sky130_fd_sc_hd__nand2_1 U23352 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[159]), .Y(n16263) );
  sky130_fd_sc_hd__nand4_1 U23353 ( .A(n16266), .B(n16265), .C(n16264), .D(
        n16263), .Y(n16272) );
  sky130_fd_sc_hd__a21oi_1 U23354 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[31]), .B1(n16436), .Y(n16270) );
  sky130_fd_sc_hd__nand2_1 U23355 ( .A(n11116), .B(
        j202_soc_core_j22_cpu_rf_gpr[127]), .Y(n16269) );
  sky130_fd_sc_hd__nand2_1 U23356 ( .A(n11152), .B(
        j202_soc_core_j22_cpu_rf_gpr[63]), .Y(n16268) );
  sky130_fd_sc_hd__nand2_1 U23357 ( .A(n11155), .B(
        j202_soc_core_j22_cpu_rf_gpr[95]), .Y(n16267) );
  sky130_fd_sc_hd__nand4_1 U23358 ( .A(n16270), .B(n16269), .C(n16268), .D(
        n16267), .Y(n16271) );
  sky130_fd_sc_hd__nor2_1 U23359 ( .A(n16272), .B(n16271), .Y(n16288) );
  sky130_fd_sc_hd__nand2_1 U23360 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[447]), .Y(n16277) );
  sky130_fd_sc_hd__nand2_1 U23361 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[255]), .Y(n16276) );
  sky130_fd_sc_hd__nand2_1 U23362 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[223]), .Y(n16275) );
  sky130_fd_sc_hd__nand2_1 U23363 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[319]), .Y(n16274) );
  sky130_fd_sc_hd__and4_1 U23364 ( .A(n16277), .B(n16276), .C(n16275), .D(
        n16274), .X(n16287) );
  sky130_fd_sc_hd__nand2_1 U23365 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[511]), .Y(n16283) );
  sky130_fd_sc_hd__nand2_1 U23366 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[191]), .Y(n16282) );
  sky130_fd_sc_hd__nand2_1 U23367 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[351]), .Y(n16281) );
  sky130_fd_sc_hd__nand2_1 U23368 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[383]), .Y(n16280) );
  sky130_fd_sc_hd__nand4_1 U23369 ( .A(n16283), .B(n16282), .C(n16281), .D(
        n16280), .Y(n16284) );
  sky130_fd_sc_hd__a21oi_1 U23370 ( .A1(j202_soc_core_j22_cpu_rf_gpr[31]), 
        .A2(n13634), .B1(n16284), .Y(n16286) );
  sky130_fd_sc_hd__nand3_1 U23371 ( .A(n16288), .B(n16287), .C(n16286), .Y(
        n26859) );
  sky130_fd_sc_hd__nand2_1 U23372 ( .A(n26859), .B(n16289), .Y(n16290) );
  sky130_fd_sc_hd__nand2_1 U23373 ( .A(n16291), .B(n16290), .Y(n25835) );
  sky130_fd_sc_hd__nand2_1 U23374 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[191]), .Y(n16295) );
  sky130_fd_sc_hd__nand2_1 U23375 ( .A(n13657), .B(
        j202_soc_core_j22_cpu_rf_gpr[255]), .Y(n16294) );
  sky130_fd_sc_hd__nand2_1 U23376 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[511]), .Y(n16293) );
  sky130_fd_sc_hd__nand2_1 U23377 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[447]), .Y(n16292) );
  sky130_fd_sc_hd__nand4_1 U23378 ( .A(n16295), .B(n16294), .C(n16293), .D(
        n16292), .Y(n16301) );
  sky130_fd_sc_hd__nand2_1 U23379 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[31]), .Y(n16299) );
  sky130_fd_sc_hd__nand2_1 U23380 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[63]), .Y(n16298) );
  sky130_fd_sc_hd__nand2_1 U23381 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[127]), .Y(n16297) );
  sky130_fd_sc_hd__nand2_1 U23382 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[415]), .Y(n16296) );
  sky130_fd_sc_hd__nand4_1 U23383 ( .A(n16299), .B(n16298), .C(n16297), .D(
        n16296), .Y(n16300) );
  sky130_fd_sc_hd__nor2_1 U23384 ( .A(n16301), .B(n16300), .Y(n16309) );
  sky130_fd_sc_hd__a22oi_1 U23385 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[319]), .B1(n14414), .B2(
        j202_soc_core_j22_cpu_rf_gpr[479]), .Y(n16308) );
  sky130_fd_sc_hd__a22oi_1 U23386 ( .A1(n23515), .A2(
        j202_soc_core_j22_cpu_rf_gpr[223]), .B1(n16469), .B2(
        j202_soc_core_j22_cpu_rf_gpr[95]), .Y(n16307) );
  sky130_fd_sc_hd__nand2_1 U23387 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[287]), .Y(n16305) );
  sky130_fd_sc_hd__nand2_1 U23388 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[159]), .Y(n16304) );
  sky130_fd_sc_hd__nand2_1 U23389 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[383]), .Y(n16303) );
  sky130_fd_sc_hd__nand2_1 U23390 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[351]), .Y(n16302) );
  sky130_fd_sc_hd__and4_1 U23391 ( .A(n16305), .B(n16304), .C(n16303), .D(
        n16302), .X(n16306) );
  sky130_fd_sc_hd__nand4_1 U23392 ( .A(n16309), .B(n16308), .C(n16307), .D(
        n16306), .Y(n22500) );
  sky130_fd_sc_hd__nand2_1 U23393 ( .A(n22500), .B(n16513), .Y(n16319) );
  sky130_fd_sc_hd__nand2_1 U23394 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[31]), .Y(n16312) );
  sky130_fd_sc_hd__nand2_1 U23395 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[31]), .Y(n16311) );
  sky130_fd_sc_hd__nand2_1 U23396 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[511]), .Y(n16310) );
  sky130_fd_sc_hd__and4_1 U23397 ( .A(n16312), .B(n16311), .C(n16516), .D(
        n16310), .X(n16318) );
  sky130_fd_sc_hd__nand2_1 U23398 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[31]), .Y(n16316) );
  sky130_fd_sc_hd__nand2_1 U23399 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[31]), .Y(n16315) );
  sky130_fd_sc_hd__nand2_1 U23400 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[31]), .Y(n16314) );
  sky130_fd_sc_hd__nand2_1 U23401 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[31]), .Y(n16313) );
  sky130_fd_sc_hd__and4_1 U23402 ( .A(n16316), .B(n16315), .C(n16314), .D(
        n16313), .X(n16317) );
  sky130_fd_sc_hd__nand3_1 U23403 ( .A(n16319), .B(n16318), .C(n16317), .Y(
        n27347) );
  sky130_fd_sc_hd__nand2_1 U23404 ( .A(n27347), .B(n16320), .Y(n16321) );
  sky130_fd_sc_hd__o21a_1 U23405 ( .A1(n27347), .A2(n16322), .B1(n16321), .X(
        n25836) );
  sky130_fd_sc_hd__xor2_1 U23406 ( .A(n25835), .B(n25836), .X(n26610) );
  sky130_fd_sc_hd__nand2_1 U23407 ( .A(n11114), .B(
        j202_soc_core_j22_cpu_rf_gpr[412]), .Y(n16329) );
  sky130_fd_sc_hd__nand2_1 U23408 ( .A(n16323), .B(
        j202_soc_core_j22_cpu_rf_gpr[476]), .Y(n16328) );
  sky130_fd_sc_hd__nand2_1 U23409 ( .A(n16324), .B(
        j202_soc_core_j22_cpu_rf_gpr[284]), .Y(n16327) );
  sky130_fd_sc_hd__nand2_1 U23410 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[156]), .Y(n16326) );
  sky130_fd_sc_hd__nand4_1 U23411 ( .A(n16329), .B(n16328), .C(n16327), .D(
        n16326), .Y(n16335) );
  sky130_fd_sc_hd__a21oi_1 U23412 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[28]), .B1(n16436), .Y(n16333) );
  sky130_fd_sc_hd__nand2_1 U23413 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[124]), .Y(n16332) );
  sky130_fd_sc_hd__nand2_1 U23414 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[60]), .Y(n16331) );
  sky130_fd_sc_hd__nand2_1 U23415 ( .A(n11155), .B(
        j202_soc_core_j22_cpu_rf_gpr[92]), .Y(n16330) );
  sky130_fd_sc_hd__nand4_1 U23416 ( .A(n16333), .B(n16332), .C(n16331), .D(
        n16330), .Y(n16334) );
  sky130_fd_sc_hd__nor2_1 U23417 ( .A(n16335), .B(n16334), .Y(n16346) );
  sky130_fd_sc_hd__nand2_1 U23418 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[444]), .Y(n16339) );
  sky130_fd_sc_hd__nand2_1 U23419 ( .A(n11151), .B(
        j202_soc_core_j22_cpu_rf_gpr[252]), .Y(n16338) );
  sky130_fd_sc_hd__nand2_1 U23420 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_rf_gpr[220]), .Y(n16337) );
  sky130_fd_sc_hd__nand2_1 U23421 ( .A(n14744), .B(
        j202_soc_core_j22_cpu_rf_gpr[316]), .Y(n16336) );
  sky130_fd_sc_hd__nand2_1 U23422 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[508]), .Y(n16343) );
  sky130_fd_sc_hd__nand2_1 U23423 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[188]), .Y(n16342) );
  sky130_fd_sc_hd__nand2_1 U23424 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[348]), .Y(n16341) );
  sky130_fd_sc_hd__nand2_1 U23425 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[380]), .Y(n16340) );
  sky130_fd_sc_hd__nand4_1 U23426 ( .A(n16343), .B(n16342), .C(n16341), .D(
        n16340), .Y(n16344) );
  sky130_fd_sc_hd__a21oi_1 U23427 ( .A1(j202_soc_core_j22_cpu_rf_gpr[28]), 
        .A2(n16285), .B1(n16344), .Y(n16345) );
  sky130_fd_sc_hd__nand3_1 U23428 ( .A(n16346), .B(n13290), .C(n16345), .Y(
        n26414) );
  sky130_fd_sc_hd__inv_2 U23429 ( .A(n26414), .Y(n26705) );
  sky130_fd_sc_hd__nand2_1 U23430 ( .A(n11114), .B(
        j202_soc_core_j22_cpu_rf_gpr[411]), .Y(n16350) );
  sky130_fd_sc_hd__nand2_1 U23431 ( .A(n16262), .B(
        j202_soc_core_j22_cpu_rf_gpr[475]), .Y(n16349) );
  sky130_fd_sc_hd__nand2_1 U23432 ( .A(n16431), .B(
        j202_soc_core_j22_cpu_rf_gpr[283]), .Y(n16348) );
  sky130_fd_sc_hd__nand2_1 U23433 ( .A(n11113), .B(
        j202_soc_core_j22_cpu_rf_gpr[155]), .Y(n16347) );
  sky130_fd_sc_hd__nand4_1 U23434 ( .A(n16350), .B(n16349), .C(n16348), .D(
        n16347), .Y(n16356) );
  sky130_fd_sc_hd__a21oi_1 U23435 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[27]), .B1(n16436), .Y(n16354) );
  sky130_fd_sc_hd__nand2_1 U23436 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[123]), .Y(n16353) );
  sky130_fd_sc_hd__nand2_1 U23437 ( .A(n11152), .B(
        j202_soc_core_j22_cpu_rf_gpr[59]), .Y(n16352) );
  sky130_fd_sc_hd__nand2_1 U23438 ( .A(n11155), .B(
        j202_soc_core_j22_cpu_rf_gpr[91]), .Y(n16351) );
  sky130_fd_sc_hd__nand4_1 U23439 ( .A(n16354), .B(n16353), .C(n16352), .D(
        n16351), .Y(n16355) );
  sky130_fd_sc_hd__nor2_1 U23440 ( .A(n16356), .B(n16355), .Y(n16371) );
  sky130_fd_sc_hd__nand2_1 U23441 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[443]), .Y(n16361) );
  sky130_fd_sc_hd__nand2_1 U23442 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[251]), .Y(n16360) );
  sky130_fd_sc_hd__nand2_1 U23443 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[219]), .Y(n16359) );
  sky130_fd_sc_hd__nand2_1 U23444 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[315]), .Y(n16358) );
  sky130_fd_sc_hd__nand2_1 U23445 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[507]), .Y(n16367) );
  sky130_fd_sc_hd__nand2_1 U23446 ( .A(n16278), .B(
        j202_soc_core_j22_cpu_rf_gpr[187]), .Y(n16366) );
  sky130_fd_sc_hd__nand2_1 U23447 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_rf_gpr[347]), .Y(n16365) );
  sky130_fd_sc_hd__nand2_1 U23448 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_rf_gpr[379]), .Y(n16364) );
  sky130_fd_sc_hd__nand4_1 U23449 ( .A(n16367), .B(n16366), .C(n16365), .D(
        n16364), .Y(n16368) );
  sky130_fd_sc_hd__a21oi_1 U23450 ( .A1(j202_soc_core_j22_cpu_rf_gpr[27]), 
        .A2(n16285), .B1(n16368), .Y(n16370) );
  sky130_fd_sc_hd__nand3_1 U23451 ( .A(n16371), .B(n13341), .C(n16370), .Y(
        n25130) );
  sky130_fd_sc_hd__inv_2 U23452 ( .A(n25130), .Y(n26707) );
  sky130_fd_sc_hd__o22ai_1 U23453 ( .A1(n16492), .A2(n26705), .B1(n26707), 
        .B2(n13793), .Y(n16542) );
  sky130_fd_sc_hd__nand2_1 U23454 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[188]), .Y(n16375) );
  sky130_fd_sc_hd__nand2_1 U23455 ( .A(n15982), .B(
        j202_soc_core_j22_cpu_rf_gpr[252]), .Y(n16374) );
  sky130_fd_sc_hd__nand2_1 U23456 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[508]), .Y(n16373) );
  sky130_fd_sc_hd__nand2_1 U23457 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[444]), .Y(n16372) );
  sky130_fd_sc_hd__nand4_1 U23458 ( .A(n16375), .B(n16374), .C(n16373), .D(
        n16372), .Y(n16381) );
  sky130_fd_sc_hd__nand2_1 U23459 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[28]), .Y(n16379) );
  sky130_fd_sc_hd__nand2_1 U23460 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[60]), .Y(n16378) );
  sky130_fd_sc_hd__nand2_1 U23461 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[124]), .Y(n16377) );
  sky130_fd_sc_hd__nand2_1 U23462 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[412]), .Y(n16376) );
  sky130_fd_sc_hd__nand4_1 U23463 ( .A(n16379), .B(n16378), .C(n16377), .D(
        n16376), .Y(n16380) );
  sky130_fd_sc_hd__nor2_1 U23464 ( .A(n16381), .B(n16380), .Y(n16389) );
  sky130_fd_sc_hd__a22oi_1 U23465 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[316]), .B1(n14414), .B2(
        j202_soc_core_j22_cpu_rf_gpr[476]), .Y(n16388) );
  sky130_fd_sc_hd__a22oi_1 U23466 ( .A1(n23515), .A2(
        j202_soc_core_j22_cpu_rf_gpr[220]), .B1(n23089), .B2(
        j202_soc_core_j22_cpu_rf_gpr[92]), .Y(n16387) );
  sky130_fd_sc_hd__nand2_1 U23467 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[284]), .Y(n16385) );
  sky130_fd_sc_hd__nand2_1 U23468 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[156]), .Y(n16384) );
  sky130_fd_sc_hd__nand2_1 U23469 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[380]), .Y(n16383) );
  sky130_fd_sc_hd__nand2_1 U23470 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[348]), .Y(n16382) );
  sky130_fd_sc_hd__and4_1 U23471 ( .A(n16385), .B(n16384), .C(n16383), .D(
        n16382), .X(n16386) );
  sky130_fd_sc_hd__nand4_1 U23472 ( .A(n16389), .B(n16388), .C(n16387), .D(
        n16386), .Y(n22645) );
  sky130_fd_sc_hd__nand2_1 U23473 ( .A(n22645), .B(n16513), .Y(n16399) );
  sky130_fd_sc_hd__nand2_1 U23474 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[28]), .Y(n16392) );
  sky130_fd_sc_hd__nand2_1 U23475 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[28]), .Y(n16391) );
  sky130_fd_sc_hd__nand2_1 U23476 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[508]), .Y(n16390) );
  sky130_fd_sc_hd__and4_1 U23477 ( .A(n16392), .B(n16391), .C(n16516), .D(
        n16390), .X(n16398) );
  sky130_fd_sc_hd__nand2_1 U23478 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[28]), .Y(n16396) );
  sky130_fd_sc_hd__nand2_1 U23479 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[28]), .Y(n16395) );
  sky130_fd_sc_hd__nand2_1 U23480 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[28]), .Y(n16394) );
  sky130_fd_sc_hd__nand2_1 U23481 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[28]), .Y(n16393) );
  sky130_fd_sc_hd__and4_1 U23482 ( .A(n16396), .B(n16395), .C(n16394), .D(
        n16393), .X(n16397) );
  sky130_fd_sc_hd__nand3_1 U23483 ( .A(n16399), .B(n16398), .C(n16397), .Y(
        n27368) );
  sky130_fd_sc_hd__nand2_1 U23484 ( .A(n27368), .B(n16529), .Y(n16400) );
  sky130_fd_sc_hd__o21ai_1 U23485 ( .A1(n14742), .A2(n27368), .B1(n16400), .Y(
        n16543) );
  sky130_fd_sc_hd__nor2_1 U23486 ( .A(n16542), .B(n16543), .Y(n16657) );
  sky130_fd_sc_hd__o22ai_1 U23487 ( .A1(n16492), .A2(n26707), .B1(n26563), 
        .B2(n13793), .Y(n16540) );
  sky130_fd_sc_hd__nand2_1 U23488 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[187]), .Y(n16404) );
  sky130_fd_sc_hd__nand2_1 U23489 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[251]), .Y(n16403) );
  sky130_fd_sc_hd__nand2_1 U23490 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[507]), .Y(n16402) );
  sky130_fd_sc_hd__nand2_1 U23491 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[443]), .Y(n16401) );
  sky130_fd_sc_hd__nand4_1 U23492 ( .A(n16404), .B(n16403), .C(n16402), .D(
        n16401), .Y(n16410) );
  sky130_fd_sc_hd__nand2_1 U23493 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[27]), .Y(n16408) );
  sky130_fd_sc_hd__nand2_1 U23494 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[59]), .Y(n16407) );
  sky130_fd_sc_hd__nand2_1 U23495 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[123]), .Y(n16406) );
  sky130_fd_sc_hd__nand2_1 U23496 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[411]), .Y(n16405) );
  sky130_fd_sc_hd__nand4_1 U23497 ( .A(n16408), .B(n16407), .C(n16406), .D(
        n16405), .Y(n16409) );
  sky130_fd_sc_hd__nor2_1 U23498 ( .A(n16410), .B(n16409), .Y(n16418) );
  sky130_fd_sc_hd__a22oi_1 U23499 ( .A1(n11160), .A2(
        j202_soc_core_j22_cpu_rf_gpr[315]), .B1(n14724), .B2(
        j202_soc_core_j22_cpu_rf_gpr[475]), .Y(n16417) );
  sky130_fd_sc_hd__a22oi_1 U23500 ( .A1(n16470), .A2(
        j202_soc_core_j22_cpu_rf_gpr[219]), .B1(n16469), .B2(
        j202_soc_core_j22_cpu_rf_gpr[91]), .Y(n16416) );
  sky130_fd_sc_hd__nand2_1 U23501 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[283]), .Y(n16414) );
  sky130_fd_sc_hd__nand2_1 U23502 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[155]), .Y(n16413) );
  sky130_fd_sc_hd__nand2_1 U23503 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[379]), .Y(n16412) );
  sky130_fd_sc_hd__nand2_1 U23504 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[347]), .Y(n16411) );
  sky130_fd_sc_hd__and4_1 U23505 ( .A(n16414), .B(n16413), .C(n16412), .D(
        n16411), .X(n16415) );
  sky130_fd_sc_hd__nand4_1 U23506 ( .A(n16418), .B(n16417), .C(n16416), .D(
        n16415), .Y(n22696) );
  sky130_fd_sc_hd__nand2_1 U23507 ( .A(n22696), .B(n16513), .Y(n16429) );
  sky130_fd_sc_hd__nand2_1 U23508 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[27]), .Y(n16422) );
  sky130_fd_sc_hd__nand2_1 U23509 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[27]), .Y(n16421) );
  sky130_fd_sc_hd__nand2_1 U23510 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[507]), .Y(n16420) );
  sky130_fd_sc_hd__and4_1 U23511 ( .A(n16422), .B(n16421), .C(n16516), .D(
        n16420), .X(n16428) );
  sky130_fd_sc_hd__nand2_1 U23512 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[27]), .Y(n16426) );
  sky130_fd_sc_hd__nand2_1 U23513 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[27]), .Y(n16425) );
  sky130_fd_sc_hd__nand2_1 U23514 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[27]), .Y(n16424) );
  sky130_fd_sc_hd__nand2_1 U23515 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[27]), .Y(n16423) );
  sky130_fd_sc_hd__and4_1 U23516 ( .A(n16426), .B(n16425), .C(n16424), .D(
        n16423), .X(n16427) );
  sky130_fd_sc_hd__nand3_1 U23517 ( .A(n16429), .B(n16428), .C(n16427), .Y(
        n24671) );
  sky130_fd_sc_hd__nand2_1 U23518 ( .A(n24671), .B(n16529), .Y(n16430) );
  sky130_fd_sc_hd__o21ai_1 U23519 ( .A1(n14742), .A2(n24671), .B1(n16430), .Y(
        n16541) );
  sky130_fd_sc_hd__nor2_1 U23520 ( .A(n16540), .B(n16541), .Y(n16651) );
  sky130_fd_sc_hd__nor2_1 U23521 ( .A(n16657), .B(n16651), .Y(n16988) );
  sky130_fd_sc_hd__nand2_1 U23522 ( .A(n16431), .B(
        j202_soc_core_j22_cpu_rf_gpr[285]), .Y(n16435) );
  sky130_fd_sc_hd__nand2_1 U23523 ( .A(n16323), .B(
        j202_soc_core_j22_cpu_rf_gpr[477]), .Y(n16434) );
  sky130_fd_sc_hd__nand2_1 U23524 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_rf_gpr[157]), .Y(n16433) );
  sky130_fd_sc_hd__nand2_1 U23525 ( .A(n11155), .B(
        j202_soc_core_j22_cpu_rf_gpr[93]), .Y(n16432) );
  sky130_fd_sc_hd__nand4_1 U23526 ( .A(n16435), .B(n16434), .C(n16433), .D(
        n16432), .Y(n16442) );
  sky130_fd_sc_hd__a21oi_1 U23527 ( .A1(n13774), .A2(
        j202_soc_core_j22_cpu_rf_tmp[29]), .B1(n16436), .Y(n16440) );
  sky130_fd_sc_hd__nand2_1 U23528 ( .A(n11114), .B(
        j202_soc_core_j22_cpu_rf_gpr[413]), .Y(n16439) );
  sky130_fd_sc_hd__nand2_1 U23529 ( .A(n11094), .B(
        j202_soc_core_j22_cpu_rf_gpr[125]), .Y(n16438) );
  sky130_fd_sc_hd__nand2_1 U23530 ( .A(n11112), .B(
        j202_soc_core_j22_cpu_rf_gpr[61]), .Y(n16437) );
  sky130_fd_sc_hd__nand4_1 U23531 ( .A(n16440), .B(n16439), .C(n16438), .D(
        n16437), .Y(n16441) );
  sky130_fd_sc_hd__nor2_1 U23532 ( .A(n16442), .B(n16441), .Y(n16457) );
  sky130_fd_sc_hd__nand2_1 U23533 ( .A(n11093), .B(
        j202_soc_core_j22_cpu_rf_gpr[445]), .Y(n16447) );
  sky130_fd_sc_hd__nand2_1 U23534 ( .A(n11111), .B(
        j202_soc_core_j22_cpu_rf_gpr[253]), .Y(n16446) );
  sky130_fd_sc_hd__nand2_1 U23535 ( .A(n16443), .B(
        j202_soc_core_j22_cpu_rf_gpr[221]), .Y(n16445) );
  sky130_fd_sc_hd__nand2_1 U23536 ( .A(n16273), .B(
        j202_soc_core_j22_cpu_rf_gpr[317]), .Y(n16444) );
  sky130_fd_sc_hd__and4_1 U23537 ( .A(n16447), .B(n16446), .C(n16445), .D(
        n16444), .X(n16456) );
  sky130_fd_sc_hd__nand2_1 U23538 ( .A(n29564), .B(
        j202_soc_core_j22_cpu_rf_gpr[509]), .Y(n16453) );
  sky130_fd_sc_hd__nand2_1 U23539 ( .A(n16448), .B(
        j202_soc_core_j22_cpu_rf_gpr[349]), .Y(n16452) );
  sky130_fd_sc_hd__nand2_1 U23540 ( .A(n15128), .B(
        j202_soc_core_j22_cpu_rf_gpr[189]), .Y(n16451) );
  sky130_fd_sc_hd__nand2_1 U23541 ( .A(n16449), .B(
        j202_soc_core_j22_cpu_rf_gpr[381]), .Y(n16450) );
  sky130_fd_sc_hd__nand4_1 U23542 ( .A(n16453), .B(n16452), .C(n16451), .D(
        n16450), .Y(n16454) );
  sky130_fd_sc_hd__a21oi_1 U23543 ( .A1(j202_soc_core_j22_cpu_rf_gpr[29]), 
        .A2(n16285), .B1(n16454), .Y(n16455) );
  sky130_fd_sc_hd__o22ai_1 U23544 ( .A1(n16492), .A2(n26702), .B1(n26705), 
        .B2(n13793), .Y(n16544) );
  sky130_fd_sc_hd__nand2_1 U23545 ( .A(n13794), .B(
        j202_soc_core_j22_cpu_rf_gpr[189]), .Y(n16462) );
  sky130_fd_sc_hd__nand2_1 U23546 ( .A(n13657), .B(
        j202_soc_core_j22_cpu_rf_gpr[253]), .Y(n16461) );
  sky130_fd_sc_hd__nand2_1 U23547 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[509]), .Y(n16460) );
  sky130_fd_sc_hd__nand2_1 U23548 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[445]), .Y(n16459) );
  sky130_fd_sc_hd__nand4_1 U23549 ( .A(n16462), .B(n16461), .C(n16460), .D(
        n16459), .Y(n16468) );
  sky130_fd_sc_hd__nand2_1 U23550 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[29]), .Y(n16466) );
  sky130_fd_sc_hd__nand2_1 U23551 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[61]), .Y(n16465) );
  sky130_fd_sc_hd__nand2_1 U23552 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[125]), .Y(n16464) );
  sky130_fd_sc_hd__nand2_1 U23553 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[413]), .Y(n16463) );
  sky130_fd_sc_hd__nand4_1 U23554 ( .A(n16466), .B(n16465), .C(n16464), .D(
        n16463), .Y(n16467) );
  sky130_fd_sc_hd__nor2_1 U23555 ( .A(n16468), .B(n16467), .Y(n16479) );
  sky130_fd_sc_hd__a22oi_1 U23556 ( .A1(n11160), .A2(
        j202_soc_core_j22_cpu_rf_gpr[317]), .B1(n23502), .B2(
        j202_soc_core_j22_cpu_rf_gpr[477]), .Y(n16478) );
  sky130_fd_sc_hd__a22oi_1 U23557 ( .A1(n16470), .A2(
        j202_soc_core_j22_cpu_rf_gpr[221]), .B1(n16469), .B2(
        j202_soc_core_j22_cpu_rf_gpr[93]), .Y(n16477) );
  sky130_fd_sc_hd__nand2_1 U23558 ( .A(n13680), .B(
        j202_soc_core_j22_cpu_rf_gpr[285]), .Y(n16475) );
  sky130_fd_sc_hd__nand2_1 U23559 ( .A(n16471), .B(
        j202_soc_core_j22_cpu_rf_gpr[157]), .Y(n16474) );
  sky130_fd_sc_hd__nand2_1 U23560 ( .A(n13686), .B(
        j202_soc_core_j22_cpu_rf_gpr[381]), .Y(n16473) );
  sky130_fd_sc_hd__nand2_1 U23561 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[349]), .Y(n16472) );
  sky130_fd_sc_hd__and4_1 U23562 ( .A(n16475), .B(n16474), .C(n16473), .D(
        n16472), .X(n16476) );
  sky130_fd_sc_hd__nand4_1 U23563 ( .A(n16479), .B(n16478), .C(n16477), .D(
        n16476), .Y(n22448) );
  sky130_fd_sc_hd__nand2_1 U23564 ( .A(n22448), .B(n16513), .Y(n16490) );
  sky130_fd_sc_hd__nand2_1 U23565 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[29]), .Y(n16483) );
  sky130_fd_sc_hd__nand2_1 U23566 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[29]), .Y(n16482) );
  sky130_fd_sc_hd__nand2_1 U23567 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[509]), .Y(n16481) );
  sky130_fd_sc_hd__and4_1 U23568 ( .A(n16483), .B(n16482), .C(n16516), .D(
        n16481), .X(n16489) );
  sky130_fd_sc_hd__nand2_1 U23569 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[29]), .Y(n16487) );
  sky130_fd_sc_hd__nand2_1 U23570 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[29]), .Y(n16486) );
  sky130_fd_sc_hd__nand2_1 U23571 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[29]), .Y(n16485) );
  sky130_fd_sc_hd__nand2_1 U23572 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[29]), .Y(n16484) );
  sky130_fd_sc_hd__and4_1 U23573 ( .A(n16487), .B(n16486), .C(n16485), .D(
        n16484), .X(n16488) );
  sky130_fd_sc_hd__nand3_1 U23574 ( .A(n16490), .B(n16489), .C(n16488), .Y(
        n24052) );
  sky130_fd_sc_hd__nand2_1 U23575 ( .A(n24052), .B(n16529), .Y(n16491) );
  sky130_fd_sc_hd__o21ai_1 U23576 ( .A1(n14742), .A2(n24052), .B1(n16491), .Y(
        n16545) );
  sky130_fd_sc_hd__nor2_1 U23577 ( .A(n16544), .B(n16545), .Y(n16994) );
  sky130_fd_sc_hd__o22ai_1 U23578 ( .A1(n16492), .A2(n26578), .B1(n26702), 
        .B2(n13793), .Y(n16546) );
  sky130_fd_sc_hd__nand2_1 U23579 ( .A(n23098), .B(
        j202_soc_core_j22_cpu_rf_gpr[190]), .Y(n16497) );
  sky130_fd_sc_hd__nand2_1 U23580 ( .A(n16493), .B(
        j202_soc_core_j22_cpu_rf_gpr[254]), .Y(n16496) );
  sky130_fd_sc_hd__nand2_1 U23581 ( .A(n29566), .B(
        j202_soc_core_j22_cpu_rf_gpr[510]), .Y(n16495) );
  sky130_fd_sc_hd__nand2_1 U23582 ( .A(n15164), .B(
        j202_soc_core_j22_cpu_rf_gpr[446]), .Y(n16494) );
  sky130_fd_sc_hd__nand4_1 U23583 ( .A(n16497), .B(n16496), .C(n16495), .D(
        n16494), .Y(n16504) );
  sky130_fd_sc_hd__nand2_1 U23584 ( .A(n16498), .B(
        j202_soc_core_j22_cpu_rf_gpr[30]), .Y(n16502) );
  sky130_fd_sc_hd__nand2_1 U23585 ( .A(n11165), .B(
        j202_soc_core_j22_cpu_rf_gpr[62]), .Y(n16501) );
  sky130_fd_sc_hd__nand2_1 U23586 ( .A(n11164), .B(
        j202_soc_core_j22_cpu_rf_gpr[126]), .Y(n16500) );
  sky130_fd_sc_hd__nand2_1 U23587 ( .A(n11156), .B(
        j202_soc_core_j22_cpu_rf_gpr[414]), .Y(n16499) );
  sky130_fd_sc_hd__nand4_1 U23588 ( .A(n16502), .B(n16501), .C(n16500), .D(
        n16499), .Y(n16503) );
  sky130_fd_sc_hd__nor2_1 U23589 ( .A(n16504), .B(n16503), .Y(n16512) );
  sky130_fd_sc_hd__a22oi_1 U23590 ( .A1(n11096), .A2(
        j202_soc_core_j22_cpu_rf_gpr[318]), .B1(n23502), .B2(
        j202_soc_core_j22_cpu_rf_gpr[478]), .Y(n16511) );
  sky130_fd_sc_hd__a22oi_1 U23591 ( .A1(n23515), .A2(
        j202_soc_core_j22_cpu_rf_gpr[222]), .B1(n23089), .B2(
        j202_soc_core_j22_cpu_rf_gpr[94]), .Y(n16510) );
  sky130_fd_sc_hd__nand2_1 U23592 ( .A(n11110), .B(
        j202_soc_core_j22_cpu_rf_gpr[286]), .Y(n16508) );
  sky130_fd_sc_hd__nand2_1 U23593 ( .A(n23113), .B(
        j202_soc_core_j22_cpu_rf_gpr[158]), .Y(n16507) );
  sky130_fd_sc_hd__nand2_1 U23594 ( .A(n11115), .B(
        j202_soc_core_j22_cpu_rf_gpr[382]), .Y(n16506) );
  sky130_fd_sc_hd__nand2_1 U23595 ( .A(n23168), .B(
        j202_soc_core_j22_cpu_rf_gpr[350]), .Y(n16505) );
  sky130_fd_sc_hd__and4_1 U23596 ( .A(n16508), .B(n16507), .C(n16506), .D(
        n16505), .X(n16509) );
  sky130_fd_sc_hd__nand4_1 U23597 ( .A(n16512), .B(n16511), .C(n16510), .D(
        n16509), .Y(n22609) );
  sky130_fd_sc_hd__nand2_1 U23598 ( .A(n22609), .B(n16513), .Y(n16528) );
  sky130_fd_sc_hd__nand2_1 U23599 ( .A(n29567), .B(
        j202_soc_core_j22_cpu_rf_vbr[30]), .Y(n16518) );
  sky130_fd_sc_hd__nand2_1 U23600 ( .A(n16514), .B(
        j202_soc_core_j22_cpu_rf_tmp[30]), .Y(n16517) );
  sky130_fd_sc_hd__nand2_1 U23601 ( .A(n29563), .B(
        j202_soc_core_j22_cpu_rf_gpr[510]), .Y(n16515) );
  sky130_fd_sc_hd__and4_1 U23602 ( .A(n16518), .B(n16517), .C(n16516), .D(
        n16515), .X(n16527) );
  sky130_fd_sc_hd__nand2_1 U23603 ( .A(n16519), .B(
        j202_soc_core_j22_cpu_pc[30]), .Y(n16525) );
  sky130_fd_sc_hd__nand2_1 U23604 ( .A(n16520), .B(
        j202_soc_core_j22_cpu_rf_gpr[30]), .Y(n16524) );
  sky130_fd_sc_hd__nand2_1 U23605 ( .A(n16521), .B(
        j202_soc_core_j22_cpu_rf_pr[30]), .Y(n16523) );
  sky130_fd_sc_hd__nand2_1 U23606 ( .A(n16012), .B(
        j202_soc_core_j22_cpu_rf_gbr[30]), .Y(n16522) );
  sky130_fd_sc_hd__and4_1 U23607 ( .A(n16525), .B(n16524), .C(n16523), .D(
        n16522), .X(n16526) );
  sky130_fd_sc_hd__nand3_1 U23608 ( .A(n16528), .B(n16527), .C(n16526), .Y(
        n27357) );
  sky130_fd_sc_hd__nand2_1 U23609 ( .A(n27357), .B(n16529), .Y(n16530) );
  sky130_fd_sc_hd__nor2_1 U23611 ( .A(n16546), .B(n16547), .Y(n16818) );
  sky130_fd_sc_hd__nor2_1 U23612 ( .A(n16994), .B(n16818), .Y(n16549) );
  sky130_fd_sc_hd__nand2_1 U23613 ( .A(n16988), .B(n16549), .Y(n16551) );
  sky130_fd_sc_hd__nor2_1 U23614 ( .A(n16531), .B(n16535), .Y(n16539) );
  sky130_fd_sc_hd__nand2_1 U23615 ( .A(n16532), .B(n16539), .Y(n17111) );
  sky130_fd_sc_hd__nor2_1 U23616 ( .A(n16551), .B(n17111), .Y(n16553) );
  sky130_fd_sc_hd__a21oi_1 U23618 ( .A1(n16539), .A2(n16538), .B1(n16537), .Y(
        n17109) );
  sky130_fd_sc_hd__nand2_1 U23619 ( .A(n16541), .B(n16540), .Y(n17114) );
  sky130_fd_sc_hd__nand2_1 U23620 ( .A(n16543), .B(n16542), .Y(n16658) );
  sky130_fd_sc_hd__o21ai_1 U23621 ( .A1(n17114), .A2(n16657), .B1(n16658), .Y(
        n16987) );
  sky130_fd_sc_hd__nand2_1 U23622 ( .A(n16545), .B(n16544), .Y(n16995) );
  sky130_fd_sc_hd__nand2_1 U23623 ( .A(n16547), .B(n16546), .Y(n16819) );
  sky130_fd_sc_hd__o21ai_1 U23624 ( .A1(n16995), .A2(n16818), .B1(n16819), .Y(
        n16548) );
  sky130_fd_sc_hd__a21oi_1 U23625 ( .A1(n16549), .A2(n16987), .B1(n16548), .Y(
        n16550) );
  sky130_fd_sc_hd__a21oi_1 U23627 ( .A1(n16554), .A2(n16553), .B1(n16552), .Y(
        n16555) );
  sky130_fd_sc_hd__nand2_1 U23628 ( .A(n22510), .B(n26859), .Y(n16557) );
  sky130_fd_sc_hd__nand4_1 U23629 ( .A(n16558), .B(n16742), .C(n16770), .D(
        n16903), .Y(n16559) );
  sky130_fd_sc_hd__nand2_1 U23630 ( .A(n16559), .B(n16945), .Y(n16570) );
  sky130_fd_sc_hd__nand3_1 U23631 ( .A(n16562), .B(n16578), .C(n16561), .Y(
        n16563) );
  sky130_fd_sc_hd__nand2_1 U23632 ( .A(n16954), .B(n16714), .Y(n16833) );
  sky130_fd_sc_hd__o21ai_1 U23633 ( .A1(n16563), .A2(n16833), .B1(n16924), .Y(
        n16569) );
  sky130_fd_sc_hd__nand3b_1 U23634 ( .A_N(n16720), .B(n16934), .C(n16903), .Y(
        n16567) );
  sky130_fd_sc_hd__nand2_1 U23635 ( .A(n16564), .B(n17170), .Y(n16767) );
  sky130_fd_sc_hd__nand2_1 U23636 ( .A(n16947), .B(n16767), .Y(n16719) );
  sky130_fd_sc_hd__nand3_1 U23637 ( .A(n16565), .B(n16593), .C(n16782), .Y(
        n16738) );
  sky130_fd_sc_hd__nand2b_1 U23638 ( .A_N(n16738), .B(n16566), .Y(n16780) );
  sky130_fd_sc_hd__o21ai_1 U23639 ( .A1(n16567), .A2(n16780), .B1(n16956), .Y(
        n16568) );
  sky130_fd_sc_hd__nand3_1 U23640 ( .A(n16570), .B(n16569), .C(n16568), .Y(
        n16571) );
  sky130_fd_sc_hd__nand2_1 U23641 ( .A(n16571), .B(n13481), .Y(n16642) );
  sky130_fd_sc_hd__nand2_1 U23642 ( .A(n21675), .B(j202_soc_core_uart_div0[4]), 
        .Y(n16637) );
  sky130_fd_sc_hd__nand2_1 U23643 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[28]), .Y(n16640) );
  sky130_fd_sc_hd__nand3_1 U23644 ( .A(n16637), .B(n21677), .C(n16640), .Y(
        n16573) );
  sky130_fd_sc_hd__nand2_1 U23645 ( .A(n21699), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[60]), .Y(n16636) );
  sky130_fd_sc_hd__nand2_1 U23646 ( .A(n21666), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[92]), .Y(n16635) );
  sky130_fd_sc_hd__nand2_1 U23647 ( .A(n16636), .B(n16635), .Y(n16572) );
  sky130_fd_sc_hd__nor2_1 U23648 ( .A(n16573), .B(n16572), .Y(n16591) );
  sky130_fd_sc_hd__nor2_1 U23649 ( .A(n16905), .B(n16773), .Y(n16943) );
  sky130_fd_sc_hd__nand2_1 U23650 ( .A(n16935), .B(n16880), .Y(n16875) );
  sky130_fd_sc_hd__nand2b_1 U23651 ( .A_N(n16858), .B(n16598), .Y(n16739) );
  sky130_fd_sc_hd__nor2_1 U23652 ( .A(n16875), .B(n16739), .Y(n16921) );
  sky130_fd_sc_hd__nand4_1 U23653 ( .A(n16943), .B(n16921), .C(n16574), .D(
        n16578), .Y(n16575) );
  sky130_fd_sc_hd__nand2_1 U23654 ( .A(n16575), .B(n16937), .Y(n16641) );
  sky130_fd_sc_hd__nor2b_1 U23655 ( .B_N(n16577), .A(n16576), .Y(n16887) );
  sky130_fd_sc_hd__nand3_1 U23656 ( .A(n16578), .B(n16849), .C(n16903), .Y(
        n16580) );
  sky130_fd_sc_hd__nand2_1 U23657 ( .A(n16598), .B(n16579), .Y(n16711) );
  sky130_fd_sc_hd__nor2_1 U23658 ( .A(n16837), .B(n16711), .Y(n16604) );
  sky130_fd_sc_hd__nand2_1 U23659 ( .A(n16880), .B(n16604), .Y(n16743) );
  sky130_fd_sc_hd__nor3_1 U23660 ( .A(n16580), .B(n16743), .C(n16962), .Y(
        n16581) );
  sky130_fd_sc_hd__nand2_1 U23661 ( .A(n16887), .B(n16581), .Y(n16582) );
  sky130_fd_sc_hd__nand2_1 U23662 ( .A(n16582), .B(n16956), .Y(n16589) );
  sky130_fd_sc_hd__o31a_1 U23663 ( .A1(n16719), .A2(n16856), .A3(n16711), .B1(
        n16924), .X(n16587) );
  sky130_fd_sc_hd__nand2b_1 U23664 ( .A_N(n16583), .B(n11994), .Y(n16686) );
  sky130_fd_sc_hd__nand3b_1 U23665 ( .A_N(n16677), .B(n16782), .C(n16686), .Y(
        n16584) );
  sky130_fd_sc_hd__o21a_1 U23666 ( .A1(n16891), .A2(n16584), .B1(n16945), .X(
        n16918) );
  sky130_fd_sc_hd__nor2_1 U23668 ( .A(n16587), .B(n16586), .Y(n16588) );
  sky130_fd_sc_hd__nand2_1 U23669 ( .A(n16589), .B(n16588), .Y(n16590) );
  sky130_fd_sc_hd__nand2_1 U23670 ( .A(n16590), .B(n20908), .Y(n16638) );
  sky130_fd_sc_hd__nand4_1 U23671 ( .A(n16642), .B(n16591), .C(n16641), .D(
        n16638), .Y(n16609) );
  sky130_fd_sc_hd__nand2_1 U23672 ( .A(n16593), .B(n16592), .Y(n16595) );
  sky130_fd_sc_hd__nand2_1 U23674 ( .A(n16611), .B(n16596), .Y(n16951) );
  sky130_fd_sc_hd__a21oi_1 U23675 ( .A1(n16734), .A2(n20350), .B1(n16964), .Y(
        n16597) );
  sky130_fd_sc_hd__a21oi_1 U23676 ( .A1(n16720), .A2(n16951), .B1(n16597), .Y(
        n16602) );
  sky130_fd_sc_hd__nand3b_1 U23677 ( .A_N(n16905), .B(n16844), .C(n16598), .Y(
        n16917) );
  sky130_fd_sc_hd__nand2_1 U23678 ( .A(n16887), .B(n16599), .Y(n16600) );
  sky130_fd_sc_hd__nand2_1 U23679 ( .A(n16600), .B(n16945), .Y(n16601) );
  sky130_fd_sc_hd__nand3_1 U23680 ( .A(n16603), .B(n16602), .C(n16601), .Y(
        n16608) );
  sky130_fd_sc_hd__nor2_1 U23681 ( .A(n16867), .B(n16735), .Y(n16708) );
  sky130_fd_sc_hd__nand2_1 U23682 ( .A(n16605), .B(n16604), .Y(n16762) );
  sky130_fd_sc_hd__and4b_1 U23683 ( .B(n16746), .C(n16742), .D(n16708), .A_N(
        n16762), .X(n16606) );
  sky130_fd_sc_hd__nor2_1 U23684 ( .A(n20580), .B(n16606), .Y(n16607) );
  sky130_fd_sc_hd__o21a_1 U23685 ( .A1(n16608), .A2(n16607), .B1(n21727), .X(
        n16643) );
  sky130_fd_sc_hd__nor2_1 U23686 ( .A(n16609), .B(n16643), .Y(n16627) );
  sky130_fd_sc_hd__nor3_1 U23687 ( .A(n16858), .B(n16610), .C(n16744), .Y(
        n16613) );
  sky130_fd_sc_hd__a21oi_1 U23688 ( .A1(n16613), .A2(n16612), .B1(n16611), .Y(
        n16750) );
  sky130_fd_sc_hd__a21oi_1 U23689 ( .A1(n16614), .A2(n16945), .B1(n16750), .Y(
        n16731) );
  sky130_fd_sc_hd__a22oi_1 U23690 ( .A1(n19125), .A2(n16616), .B1(n16615), 
        .B2(n19381), .Y(n16618) );
  sky130_fd_sc_hd__o211ai_1 U23691 ( .A1(n16618), .A2(n16845), .B1(n16934), 
        .C1(n16709), .Y(n16624) );
  sky130_fd_sc_hd__nor2_1 U23692 ( .A(n16882), .B(n16619), .Y(n16966) );
  sky130_fd_sc_hd__nor4_1 U23693 ( .A(n16961), .B(n16837), .C(n16620), .D(
        n16673), .Y(n16621) );
  sky130_fd_sc_hd__nand4_1 U23694 ( .A(n16622), .B(n16775), .C(n16966), .D(
        n16621), .Y(n16623) );
  sky130_fd_sc_hd__a22oi_1 U23695 ( .A1(n16924), .A2(n16624), .B1(n16623), 
        .B2(n16956), .Y(n16625) );
  sky130_fd_sc_hd__nand2_1 U23696 ( .A(n16731), .B(n16625), .Y(n16626) );
  sky130_fd_sc_hd__nand2_1 U23697 ( .A(n16626), .B(n21697), .Y(n16646) );
  sky130_fd_sc_hd__nand2_1 U23698 ( .A(j202_soc_core_memory0_ram_dout0[412]), 
        .B(n21597), .Y(n16628) );
  sky130_fd_sc_hd__nand2_1 U23699 ( .A(j202_soc_core_memory0_ram_dout0[124]), 
        .B(n21591), .Y(n16634) );
  sky130_fd_sc_hd__nand2_1 U23701 ( .A(j202_soc_core_memory0_ram_dout0[156]), 
        .B(n21592), .Y(n16632) );
  sky130_fd_sc_hd__nand3_1 U23702 ( .A(n12490), .B(n20965), .C(n20964), .Y(
        n19251) );
  sky130_fd_sc_hd__nand4_1 U23703 ( .A(n16638), .B(n16637), .C(n16636), .D(
        n16635), .Y(n16639) );
  sky130_fd_sc_hd__a21oi_1 U23704 ( .A1(j202_soc_core_memory0_ram_dout0[508]), 
        .A2(n21771), .B1(n16639), .Y(n20970) );
  sky130_fd_sc_hd__and4_1 U23705 ( .A(n16642), .B(n21738), .C(n16641), .D(
        n16640), .X(n16645) );
  sky130_fd_sc_hd__and3_1 U23706 ( .A(n16646), .B(n16645), .C(n16644), .X(
        n20969) );
  sky130_fd_sc_hd__nand2_1 U23707 ( .A(n20970), .B(n20969), .Y(n19250) );
  sky130_fd_sc_hd__ha_1 U23708 ( .A(n16647), .B(j202_soc_core_j22_cpu_pc[28]), 
        .COUT(n16999), .SUM(n26446) );
  sky130_fd_sc_hd__a2bb2oi_1 U23709 ( .B1(n11144), .B2(n26446), .A1_N(n26705), 
        .A2_N(n11143), .Y(n16648) );
  sky130_fd_sc_hd__o21ai_1 U23710 ( .A1(n16649), .A2(n21584), .B1(n16648), .Y(
        n16650) );
  sky130_fd_sc_hd__a21oi_1 U23711 ( .A1(n22515), .A2(n27368), .B1(n16650), .Y(
        n16663) );
  sky130_fd_sc_hd__nand2_1 U23712 ( .A(n16986), .B(n17115), .Y(n16654) );
  sky130_fd_sc_hd__nor2_1 U23713 ( .A(n16654), .B(n17108), .Y(n16656) );
  sky130_fd_sc_hd__a21oi_1 U23714 ( .A1(n16989), .A2(n17115), .B1(n16652), .Y(
        n16653) );
  sky130_fd_sc_hd__o21ai_0 U23715 ( .A1(n16654), .A2(n17110), .B1(n16653), .Y(
        n16655) );
  sky130_fd_sc_hd__a21oi_1 U23716 ( .A1(n22513), .A2(n16656), .B1(n16655), .Y(
        n16661) );
  sky130_fd_sc_hd__nand2_1 U23717 ( .A(n16659), .B(n16658), .Y(n16660) );
  sky130_fd_sc_hd__xor2_1 U23718 ( .A(n16661), .B(n16660), .X(n26410) );
  sky130_fd_sc_hd__nand2_1 U23719 ( .A(n26410), .B(n12158), .Y(n16662) );
  sky130_fd_sc_hd__nand2_1 U23720 ( .A(j202_soc_core_memory0_ram_dout0[382]), 
        .B(n21596), .Y(n16668) );
  sky130_fd_sc_hd__nand2_1 U23721 ( .A(j202_soc_core_memory0_ram_dout0[254]), 
        .B(n21735), .Y(n16667) );
  sky130_fd_sc_hd__nand2_1 U23722 ( .A(j202_soc_core_memory0_ram_dout0[30]), 
        .B(n21733), .Y(n16666) );
  sky130_fd_sc_hd__nand2_1 U23723 ( .A(j202_soc_core_memory0_ram_dout0[318]), 
        .B(n21603), .Y(n16665) );
  sky130_fd_sc_hd__nand2_1 U23724 ( .A(j202_soc_core_memory0_ram_dout0[62]), 
        .B(n21604), .Y(n16672) );
  sky130_fd_sc_hd__nand2_1 U23725 ( .A(j202_soc_core_memory0_ram_dout0[350]), 
        .B(n21593), .Y(n16671) );
  sky130_fd_sc_hd__nand2_1 U23726 ( .A(j202_soc_core_memory0_ram_dout0[286]), 
        .B(n21605), .Y(n16670) );
  sky130_fd_sc_hd__nand2_1 U23727 ( .A(j202_soc_core_memory0_ram_dout0[414]), 
        .B(n21597), .Y(n16669) );
  sky130_fd_sc_hd__nor2_1 U23728 ( .A(n16673), .B(n16914), .Y(n16700) );
  sky130_fd_sc_hd__nand2_1 U23729 ( .A(n16775), .B(n16700), .Y(n16908) );
  sky130_fd_sc_hd__nor2_1 U23730 ( .A(n16908), .B(n16674), .Y(n16676) );
  sky130_fd_sc_hd__nand3_1 U23731 ( .A(n16676), .B(n16675), .C(n16947), .Y(
        n16680) );
  sky130_fd_sc_hd__nor2_1 U23732 ( .A(n16677), .B(n16961), .Y(n16772) );
  sky130_fd_sc_hd__nand3_1 U23733 ( .A(n16772), .B(n16678), .C(n16782), .Y(
        n16679) );
  sky130_fd_sc_hd__nor2_1 U23734 ( .A(n16680), .B(n16679), .Y(n16696) );
  sky130_fd_sc_hd__nand3_1 U23735 ( .A(n16702), .B(n16683), .C(n16682), .Y(
        n16684) );
  sky130_fd_sc_hd__nand2_1 U23736 ( .A(n16684), .B(n16919), .Y(n16928) );
  sky130_fd_sc_hd__nand2_1 U23737 ( .A(n16685), .B(n16714), .Y(n16776) );
  sky130_fd_sc_hd__nand4_1 U23738 ( .A(n16688), .B(n16687), .C(n16953), .D(
        n16686), .Y(n16694) );
  sky130_fd_sc_hd__nand2_1 U23739 ( .A(n16698), .B(n16965), .Y(n16763) );
  sky130_fd_sc_hd__nor2_1 U23740 ( .A(n16690), .B(n16763), .Y(n16693) );
  sky130_fd_sc_hd__nor2b_1 U23741 ( .B_N(n16740), .A(n16769), .Y(n16781) );
  sky130_fd_sc_hd__nand4_1 U23742 ( .A(n16693), .B(n16781), .C(n16692), .D(
        n16691), .Y(n16906) );
  sky130_fd_sc_hd__o211ai_1 U23744 ( .A1(n16696), .A2(n16964), .B1(n16928), 
        .C1(n16695), .Y(n16705) );
  sky130_fd_sc_hd__and4_1 U23745 ( .A(n16894), .B(n16700), .C(n16699), .D(
        n16698), .X(n16701) );
  sky130_fd_sc_hd__a31oi_1 U23746 ( .A1(n16703), .A2(n16702), .A3(n16701), 
        .B1(n20580), .Y(n16704) );
  sky130_fd_sc_hd__o21a_1 U23747 ( .A1(n16705), .A2(n16704), .B1(n20908), .X(
        n16807) );
  sky130_fd_sc_hd__nand2_1 U23748 ( .A(n16706), .B(n17167), .Y(n16707) );
  sky130_fd_sc_hd__nand4_1 U23749 ( .A(n16965), .B(n16879), .C(n16782), .D(
        n16707), .Y(n16852) );
  sky130_fd_sc_hd__nand2_1 U23750 ( .A(n16709), .B(n16708), .Y(n16710) );
  sky130_fd_sc_hd__nor4_1 U23751 ( .A(n16882), .B(n16711), .C(n16852), .D(
        n16710), .Y(n16712) );
  sky130_fd_sc_hd__nand2b_1 U23752 ( .A_N(n16712), .B(n16924), .Y(n16732) );
  sky130_fd_sc_hd__nor2_1 U23753 ( .A(n16713), .B(n16763), .Y(n16936) );
  sky130_fd_sc_hd__nand4_1 U23754 ( .A(n16936), .B(n16754), .C(n16714), .D(
        n16734), .Y(n16729) );
  sky130_fd_sc_hd__nand4b_1 U23755 ( .A_N(n16769), .B(n16717), .C(n16880), .D(
        n16716), .Y(n16718) );
  sky130_fd_sc_hd__nor3_1 U23756 ( .A(n16719), .B(n16718), .C(n16856), .Y(
        n16727) );
  sky130_fd_sc_hd__nand4_1 U23757 ( .A(n16725), .B(n16724), .C(n16723), .D(
        n16722), .Y(n16726) );
  sky130_fd_sc_hd__o2bb2ai_1 U23758 ( .B1(n20580), .B2(n16727), .A1_N(n16919), 
        .A2_N(n16726), .Y(n16728) );
  sky130_fd_sc_hd__a21oi_1 U23759 ( .A1(n16729), .A2(n16945), .B1(n16728), .Y(
        n16730) );
  sky130_fd_sc_hd__nand3_1 U23760 ( .A(n16732), .B(n16731), .C(n16730), .Y(
        n16733) );
  sky130_fd_sc_hd__nand2_1 U23761 ( .A(n16733), .B(n21697), .Y(n16805) );
  sky130_fd_sc_hd__nand2_1 U23762 ( .A(n16770), .B(n16734), .Y(n16874) );
  sky130_fd_sc_hd__nor2_1 U23763 ( .A(n16735), .B(n16874), .Y(n16922) );
  sky130_fd_sc_hd__nand4_1 U23764 ( .A(n16736), .B(n16913), .C(n16785), .D(
        n16922), .Y(n16737) );
  sky130_fd_sc_hd__o21ai_1 U23765 ( .A1(n16737), .A2(n16787), .B1(n16919), .Y(
        n16759) );
  sky130_fd_sc_hd__nor2_1 U23766 ( .A(n16739), .B(n16738), .Y(n16885) );
  sky130_fd_sc_hd__nand2_1 U23767 ( .A(n16849), .B(n16740), .Y(n16868) );
  sky130_fd_sc_hd__nand3_1 U23768 ( .A(n16885), .B(n16742), .C(n16741), .Y(
        n16749) );
  sky130_fd_sc_hd__nor4_1 U23769 ( .A(n16745), .B(n16744), .C(n16856), .D(
        n16743), .Y(n16747) );
  sky130_fd_sc_hd__a21oi_1 U23770 ( .A1(n16747), .A2(n16746), .B1(n20580), .Y(
        n16748) );
  sky130_fd_sc_hd__a21oi_1 U23771 ( .A1(n16749), .A2(n16924), .B1(n16748), .Y(
        n16758) );
  sky130_fd_sc_hd__nand2_1 U23772 ( .A(n20633), .B(n20463), .Y(n16752) );
  sky130_fd_sc_hd__nor2_1 U23773 ( .A(n16752), .B(n16751), .Y(n16753) );
  sky130_fd_sc_hd__nand3_1 U23774 ( .A(n16887), .B(n16754), .C(n16753), .Y(
        n16755) );
  sky130_fd_sc_hd__nand4_1 U23776 ( .A(n16759), .B(n16758), .C(n16757), .D(
        n16756), .Y(n16760) );
  sky130_fd_sc_hd__nand2_1 U23777 ( .A(n16760), .B(n21727), .Y(n16801) );
  sky130_fd_sc_hd__a22oi_1 U23778 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[62]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[94]), .Y(n16799) );
  sky130_fd_sc_hd__nand2_1 U23779 ( .A(n21675), .B(j202_soc_core_uart_div0[6]), 
        .Y(n16798) );
  sky130_fd_sc_hd__nand2_1 U23780 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[30]), .Y(n16797) );
  sky130_fd_sc_hd__nand4_1 U23781 ( .A(n16799), .B(n21677), .C(n16798), .D(
        n16797), .Y(n16761) );
  sky130_fd_sc_hd__nor2b_1 U23782 ( .B_N(n16801), .A(n16761), .Y(n16794) );
  sky130_fd_sc_hd__nor4_1 U23783 ( .A(n16764), .B(n16855), .C(n16763), .D(
        n16762), .Y(n16765) );
  sky130_fd_sc_hd__nand2b_1 U23784 ( .A_N(n16765), .B(n16937), .Y(n16803) );
  sky130_fd_sc_hd__nand2_1 U23785 ( .A(n16767), .B(n16766), .Y(n16768) );
  sky130_fd_sc_hd__nor2_1 U23786 ( .A(n16769), .B(n16768), .Y(n16771) );
  sky130_fd_sc_hd__nand4_1 U23787 ( .A(n16772), .B(n16783), .C(n16771), .D(
        n16770), .Y(n16774) );
  sky130_fd_sc_hd__nor2_1 U23788 ( .A(n16773), .B(n16891), .Y(n16963) );
  sky130_fd_sc_hd__nand2_1 U23789 ( .A(n16913), .B(n16963), .Y(n16786) );
  sky130_fd_sc_hd__o21ai_1 U23790 ( .A1(n16774), .A2(n16786), .B1(n16945), .Y(
        n16792) );
  sky130_fd_sc_hd__nand3b_1 U23791 ( .A_N(n16776), .B(n16775), .C(n16849), .Y(
        n16777) );
  sky130_fd_sc_hd__nor2_1 U23792 ( .A(n16914), .B(n16777), .Y(n16950) );
  sky130_fd_sc_hd__nand2_1 U23793 ( .A(n16950), .B(n16778), .Y(n16779) );
  sky130_fd_sc_hd__nor2_1 U23794 ( .A(n16780), .B(n16779), .Y(n16923) );
  sky130_fd_sc_hd__nand3_1 U23795 ( .A(n16785), .B(n16784), .C(n16783), .Y(
        n16895) );
  sky130_fd_sc_hd__nor4_1 U23796 ( .A(n16788), .B(n16787), .C(n16895), .D(
        n16786), .Y(n16789) );
  sky130_fd_sc_hd__a2bb2oi_1 U23797 ( .B1(n16956), .B2(n16790), .A1_N(n16789), 
        .A2_N(n16964), .Y(n16791) );
  sky130_fd_sc_hd__nand2_1 U23798 ( .A(n16792), .B(n16791), .Y(n16793) );
  sky130_fd_sc_hd__nand2_1 U23799 ( .A(n16793), .B(n13481), .Y(n16802) );
  sky130_fd_sc_hd__nand4_1 U23800 ( .A(n16805), .B(n16794), .C(n16803), .D(
        n16802), .Y(n16795) );
  sky130_fd_sc_hd__nor2_1 U23801 ( .A(n16807), .B(n16795), .Y(n16796) );
  sky130_fd_sc_hd__nand2_1 U23802 ( .A(j202_soc_core_memory0_ram_dout0[510]), 
        .B(n21771), .Y(n16809) );
  sky130_fd_sc_hd__nand4_1 U23803 ( .A(n16799), .B(n21738), .C(n16798), .D(
        n16797), .Y(n16800) );
  sky130_fd_sc_hd__nor2b_1 U23804 ( .B_N(n16801), .A(n16800), .Y(n16804) );
  sky130_fd_sc_hd__nand4_1 U23805 ( .A(n16805), .B(n16804), .C(n16803), .D(
        n16802), .Y(n16806) );
  sky130_fd_sc_hd__nor2_1 U23806 ( .A(n16807), .B(n16806), .Y(n16808) );
  sky130_fd_sc_hd__nand2_1 U23807 ( .A(n16809), .B(n16808), .Y(n21164) );
  sky130_fd_sc_hd__nor2_1 U23808 ( .A(n16994), .B(n16810), .Y(n16813) );
  sky130_fd_sc_hd__nand2_1 U23809 ( .A(n16813), .B(n16986), .Y(n16815) );
  sky130_fd_sc_hd__nor2_1 U23810 ( .A(n16815), .B(n17108), .Y(n16817) );
  sky130_fd_sc_hd__o21ai_0 U23811 ( .A1(n16994), .A2(n16811), .B1(n16995), .Y(
        n16812) );
  sky130_fd_sc_hd__a21oi_1 U23812 ( .A1(n16989), .A2(n16813), .B1(n16812), .Y(
        n16814) );
  sky130_fd_sc_hd__o21ai_0 U23813 ( .A1(n16815), .A2(n17110), .B1(n16814), .Y(
        n16816) );
  sky130_fd_sc_hd__a21oi_1 U23814 ( .A1(n22513), .A2(n16817), .B1(n16816), .Y(
        n16822) );
  sky130_fd_sc_hd__nand2_1 U23815 ( .A(n16820), .B(n16819), .Y(n16821) );
  sky130_fd_sc_hd__xor2_1 U23816 ( .A(n16822), .B(n16821), .X(n24490) );
  sky130_fd_sc_hd__ha_1 U23817 ( .A(n16823), .B(j202_soc_core_j22_cpu_pc[30]), 
        .COUT(n16158), .SUM(n26520) );
  sky130_fd_sc_hd__nand2_1 U23818 ( .A(n26520), .B(n16824), .Y(n16828) );
  sky130_fd_sc_hd__nand2_1 U23819 ( .A(n26520), .B(n11144), .Y(n16827) );
  sky130_fd_sc_hd__nand2_1 U23820 ( .A(n22515), .B(n27357), .Y(n16826) );
  sky130_fd_sc_hd__nand2_1 U23821 ( .A(n22510), .B(n26716), .Y(n16825) );
  sky130_fd_sc_hd__nand4_1 U23822 ( .A(n16828), .B(n16827), .C(n16826), .D(
        n16825), .Y(n16829) );
  sky130_fd_sc_hd__a21oi_1 U23823 ( .A1(n24490), .A2(n12158), .B1(n16829), .Y(
        n16830) );
  sky130_fd_sc_hd__o21a_1 U23824 ( .A1(n17125), .A2(n26538), .B1(n16830), .X(
        n21023) );
  sky130_fd_sc_hd__nand4_1 U23825 ( .A(n12465), .B(n10939), .C(n28919), .D(
        n28920), .Y(n16831) );
  sky130_fd_sc_hd__nand2_1 U23826 ( .A(j202_soc_core_memory0_ram_dout0[189]), 
        .B(n21590), .Y(n16832) );
  sky130_fd_sc_hd__nor4_1 U23827 ( .A(n16941), .B(n16940), .C(n16875), .D(
        n16833), .Y(n16834) );
  sky130_fd_sc_hd__nand2b_1 U23828 ( .A_N(n16834), .B(n16956), .Y(n16865) );
  sky130_fd_sc_hd__nor4_1 U23829 ( .A(n16838), .B(n16837), .C(n16836), .D(
        n16835), .Y(n16839) );
  sky130_fd_sc_hd__nand2b_1 U23830 ( .A_N(n16840), .B(n16839), .Y(n16841) );
  sky130_fd_sc_hd__a22oi_1 U23831 ( .A1(n16842), .A2(n16951), .B1(n16841), 
        .B2(n16945), .Y(n16864) );
  sky130_fd_sc_hd__o21ai_1 U23832 ( .A1(n17274), .A2(n16845), .B1(n16844), .Y(
        n16847) );
  sky130_fd_sc_hd__nand2_1 U23833 ( .A(n16847), .B(n16846), .Y(n16848) );
  sky130_fd_sc_hd__nand4_1 U23834 ( .A(n16966), .B(n16850), .C(n16849), .D(
        n16848), .Y(n16851) );
  sky130_fd_sc_hd__nor3_1 U23835 ( .A(n16853), .B(n16852), .C(n16851), .Y(
        n16854) );
  sky130_fd_sc_hd__nand2b_1 U23836 ( .A_N(n16854), .B(n16924), .Y(n16863) );
  sky130_fd_sc_hd__nor3_1 U23837 ( .A(n16856), .B(n16855), .C(n16895), .Y(
        n16860) );
  sky130_fd_sc_hd__nor2_1 U23838 ( .A(n16858), .B(n16857), .Y(n16859) );
  sky130_fd_sc_hd__nand2_1 U23839 ( .A(n16860), .B(n16859), .Y(n16861) );
  sky130_fd_sc_hd__nand2_1 U23840 ( .A(n16861), .B(n16919), .Y(n16862) );
  sky130_fd_sc_hd__nand4_1 U23841 ( .A(n16865), .B(n16864), .C(n16863), .D(
        n16862), .Y(n16866) );
  sky130_fd_sc_hd__nand2_1 U23842 ( .A(n16866), .B(n21697), .Y(n16979) );
  sky130_fd_sc_hd__nor2_1 U23843 ( .A(n16868), .B(n16867), .Y(n16869) );
  sky130_fd_sc_hd__nand2_1 U23844 ( .A(n16966), .B(n16869), .Y(n16871) );
  sky130_fd_sc_hd__o21ai_1 U23845 ( .A1(n16871), .A2(n16870), .B1(n16956), .Y(
        n16900) );
  sky130_fd_sc_hd__nand4b_1 U23846 ( .A_N(n16874), .B(n20350), .C(n16873), .D(
        n16872), .Y(n16889) );
  sky130_fd_sc_hd__nor3_1 U23847 ( .A(n16911), .B(n16875), .C(n16889), .Y(
        n16876) );
  sky130_fd_sc_hd__nand2b_1 U23848 ( .A_N(n16960), .B(n16876), .Y(n16877) );
  sky130_fd_sc_hd__nand3_1 U23850 ( .A(n16934), .B(n16880), .C(n16879), .Y(
        n16883) );
  sky130_fd_sc_hd__nor3_1 U23851 ( .A(n16883), .B(n16882), .C(n16881), .Y(
        n16884) );
  sky130_fd_sc_hd__nand4_1 U23852 ( .A(n16887), .B(n16886), .C(n16885), .D(
        n16884), .Y(n16888) );
  sky130_fd_sc_hd__nand2_1 U23853 ( .A(n16888), .B(n16924), .Y(n16898) );
  sky130_fd_sc_hd__nor2_1 U23854 ( .A(n16891), .B(n16890), .Y(n16892) );
  sky130_fd_sc_hd__nand4b_1 U23855 ( .A_N(n16895), .B(n16894), .C(n16893), .D(
        n16892), .Y(n16896) );
  sky130_fd_sc_hd__nand2_1 U23856 ( .A(n16896), .B(n16945), .Y(n16897) );
  sky130_fd_sc_hd__nand4_1 U23857 ( .A(n16900), .B(n16899), .C(n16898), .D(
        n16897), .Y(n16901) );
  sky130_fd_sc_hd__nand2_1 U23858 ( .A(n16901), .B(n21727), .Y(n16975) );
  sky130_fd_sc_hd__a22oi_1 U23859 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[61]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[93]), .Y(n16974) );
  sky130_fd_sc_hd__nand2_1 U23860 ( .A(n21675), .B(j202_soc_core_uart_div0[5]), 
        .Y(n16973) );
  sky130_fd_sc_hd__nand2_1 U23861 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[29]), .Y(n16972) );
  sky130_fd_sc_hd__nand4_1 U23862 ( .A(n16974), .B(n21677), .C(n16973), .D(
        n16972), .Y(n16902) );
  sky130_fd_sc_hd__nor2b_1 U23863 ( .B_N(n16975), .A(n16902), .Y(n16939) );
  sky130_fd_sc_hd__nand3b_1 U23864 ( .A_N(n16905), .B(n16904), .C(n16903), .Y(
        n16907) );
  sky130_fd_sc_hd__o21ai_1 U23865 ( .A1(n16907), .A2(n16906), .B1(n16945), .Y(
        n16932) );
  sky130_fd_sc_hd__nand3_1 U23866 ( .A(n16935), .B(n20633), .C(n16909), .Y(
        n16910) );
  sky130_fd_sc_hd__nor3_1 U23867 ( .A(n16911), .B(n16940), .C(n16910), .Y(
        n16912) );
  sky130_fd_sc_hd__nand3_1 U23868 ( .A(n16936), .B(n16913), .C(n16912), .Y(
        n16930) );
  sky130_fd_sc_hd__nand3b_1 U23869 ( .A_N(n16917), .B(n16916), .C(n16915), .Y(
        n16920) );
  sky130_fd_sc_hd__a21oi_1 U23870 ( .A1(n16920), .A2(n16919), .B1(n16918), .Y(
        n16927) );
  sky130_fd_sc_hd__nand3_1 U23871 ( .A(n16923), .B(n16922), .C(n16921), .Y(
        n16925) );
  sky130_fd_sc_hd__nand2_1 U23872 ( .A(n16925), .B(n16924), .Y(n16926) );
  sky130_fd_sc_hd__nand3_1 U23873 ( .A(n16928), .B(n16927), .C(n16926), .Y(
        n16929) );
  sky130_fd_sc_hd__a21oi_1 U23874 ( .A1(n16930), .A2(n16956), .B1(n16929), .Y(
        n16931) );
  sky130_fd_sc_hd__nand2_1 U23875 ( .A(n16932), .B(n16931), .Y(n16933) );
  sky130_fd_sc_hd__nand2_1 U23876 ( .A(n16933), .B(n20908), .Y(n16977) );
  sky130_fd_sc_hd__nand4_1 U23877 ( .A(n16936), .B(n16935), .C(n16934), .D(
        n20633), .Y(n16938) );
  sky130_fd_sc_hd__nand2_1 U23878 ( .A(n16938), .B(n16937), .Y(n16976) );
  sky130_fd_sc_hd__nand4_1 U23879 ( .A(n16979), .B(n16939), .C(n16977), .D(
        n16976), .Y(n16970) );
  sky130_fd_sc_hd__nor3_1 U23880 ( .A(n16942), .B(n16941), .C(n16940), .Y(
        n16944) );
  sky130_fd_sc_hd__nand2_1 U23881 ( .A(n16944), .B(n16943), .Y(n16946) );
  sky130_fd_sc_hd__nand2_1 U23882 ( .A(n16946), .B(n16945), .Y(n16959) );
  sky130_fd_sc_hd__nand4_1 U23883 ( .A(n16950), .B(n16949), .C(n16948), .D(
        n16947), .Y(n16957) );
  sky130_fd_sc_hd__a21oi_1 U23884 ( .A1(n16954), .A2(n16953), .B1(n16952), .Y(
        n16955) );
  sky130_fd_sc_hd__a21oi_1 U23885 ( .A1(n16957), .A2(n16956), .B1(n16955), .Y(
        n16958) );
  sky130_fd_sc_hd__nand2_1 U23886 ( .A(n16959), .B(n16958), .Y(n16969) );
  sky130_fd_sc_hd__nor4b_1 U23887 ( .D_N(n16963), .A(n16962), .B(n16961), .C(
        n16960), .Y(n16967) );
  sky130_fd_sc_hd__a31oi_1 U23888 ( .A1(n16967), .A2(n16966), .A3(n16965), 
        .B1(n16964), .Y(n16968) );
  sky130_fd_sc_hd__o21a_1 U23889 ( .A1(n16969), .A2(n16968), .B1(n13481), .X(
        n16982) );
  sky130_fd_sc_hd__nor2_1 U23890 ( .A(n16970), .B(n16982), .Y(n16971) );
  sky130_fd_sc_hd__nand2_1 U23891 ( .A(j202_soc_core_memory0_ram_dout0[509]), 
        .B(n21771), .Y(n16985) );
  sky130_fd_sc_hd__nand4_1 U23892 ( .A(n16974), .B(n21738), .C(n16973), .D(
        n16972), .Y(n16978) );
  sky130_fd_sc_hd__nand4b_1 U23893 ( .A_N(n16978), .B(n16977), .C(n16976), .D(
        n16975), .Y(n16981) );
  sky130_fd_sc_hd__nor2_1 U23894 ( .A(n16981), .B(n16980), .Y(n16984) );
  sky130_fd_sc_hd__nand3_1 U23895 ( .A(n16985), .B(n16984), .C(n16983), .Y(
        n21814) );
  sky130_fd_sc_hd__nand2_1 U23896 ( .A(n16986), .B(n16988), .Y(n16991) );
  sky130_fd_sc_hd__nor2_1 U23897 ( .A(n16991), .B(n17108), .Y(n16993) );
  sky130_fd_sc_hd__a21oi_1 U23898 ( .A1(n16989), .A2(n16988), .B1(n16987), .Y(
        n16990) );
  sky130_fd_sc_hd__nand2_1 U23899 ( .A(n16996), .B(n16995), .Y(n16997) );
  sky130_fd_sc_hd__xor2_1 U23900 ( .A(n16998), .B(n16997), .X(n24044) );
  sky130_fd_sc_hd__nand2_1 U23901 ( .A(n24044), .B(n12158), .Y(n17002) );
  sky130_fd_sc_hd__ha_1 U23902 ( .A(n16999), .B(j202_soc_core_j22_cpu_pc[29]), 
        .COUT(n16823), .SUM(n26949) );
  sky130_fd_sc_hd__a22oi_1 U23903 ( .A1(n22510), .A2(n26971), .B1(n22596), 
        .B2(n26949), .Y(n17001) );
  sky130_fd_sc_hd__nand2_1 U23904 ( .A(n22515), .B(n24052), .Y(n17000) );
  sky130_fd_sc_hd__nand3_1 U23905 ( .A(n17002), .B(n17001), .C(n17000), .Y(
        n17003) );
  sky130_fd_sc_hd__nand3_1 U23906 ( .A(n17007), .B(n17006), .C(n17005), .Y(
        n17008) );
  sky130_fd_sc_hd__nand3_1 U23909 ( .A(n17014), .B(n17013), .C(n17012), .Y(
        n17015) );
  sky130_fd_sc_hd__nand2_1 U23910 ( .A(n17015), .B(n13388), .Y(n17018) );
  sky130_fd_sc_hd__nand2_1 U23911 ( .A(n17016), .B(n17302), .Y(n17017) );
  sky130_fd_sc_hd__nand4_1 U23912 ( .A(n17020), .B(n17019), .C(n17018), .D(
        n17017), .Y(n17023) );
  sky130_fd_sc_hd__o21ai_1 U23913 ( .A1(n17023), .A2(n17022), .B1(n17021), .Y(
        n17097) );
  sky130_fd_sc_hd__nand2_1 U23914 ( .A(n17025), .B(n17024), .Y(n17026) );
  sky130_fd_sc_hd__nor4b_1 U23915 ( .D_N(n17028), .A(n17071), .B(n17027), .C(
        n17026), .Y(n17060) );
  sky130_fd_sc_hd__o21ai_1 U23916 ( .A1(n17030), .A2(n17029), .B1(n17302), .Y(
        n17041) );
  sky130_fd_sc_hd__nor3_1 U23917 ( .A(n17075), .B(n17032), .C(n17031), .Y(
        n17038) );
  sky130_fd_sc_hd__nor4_1 U23918 ( .A(n17035), .B(n17071), .C(n17034), .D(
        n17033), .Y(n17036) );
  sky130_fd_sc_hd__o22a_1 U23919 ( .A1(n17039), .A2(n17038), .B1(n17037), .B2(
        n17036), .X(n17040) );
  sky130_fd_sc_hd__nand2_1 U23920 ( .A(n17041), .B(n17040), .Y(n17057) );
  sky130_fd_sc_hd__a21oi_1 U23921 ( .A1(n17066), .A2(n17044), .B1(n17043), .Y(
        n17056) );
  sky130_fd_sc_hd__nor2_1 U23922 ( .A(n17047), .B(n17046), .Y(n17050) );
  sky130_fd_sc_hd__nand4_1 U23923 ( .A(n17051), .B(n17050), .C(n17049), .D(
        n17048), .Y(n17052) );
  sky130_fd_sc_hd__nand2_1 U23924 ( .A(n17052), .B(n13387), .Y(n17053) );
  sky130_fd_sc_hd__o21ai_1 U23925 ( .A1(n17060), .A2(n17059), .B1(n17058), .Y(
        n17062) );
  sky130_fd_sc_hd__a211oi_1 U23926 ( .A1(n17067), .A2(n17066), .B1(n17065), 
        .C1(n17064), .Y(n17068) );
  sky130_fd_sc_hd__nand2b_1 U23927 ( .A_N(n17068), .B(n17302), .Y(n17093) );
  sky130_fd_sc_hd__nor4b_1 U23928 ( .D_N(n17072), .A(n17071), .B(n17070), .C(
        n17069), .Y(n17074) );
  sky130_fd_sc_hd__nand3b_1 U23929 ( .A_N(n17075), .B(n17074), .C(n17073), .Y(
        n17080) );
  sky130_fd_sc_hd__nor3b_1 U23930 ( .C_N(n17077), .A(n17076), .B(n17085), .Y(
        n17079) );
  sky130_fd_sc_hd__a2bb2oi_1 U23931 ( .B1(n13387), .B2(n17080), .A1_N(n17079), 
        .A2_N(n17078), .Y(n17092) );
  sky130_fd_sc_hd__nand2_1 U23932 ( .A(n17082), .B(n17081), .Y(n17084) );
  sky130_fd_sc_hd__nor2_1 U23933 ( .A(n17084), .B(n17083), .Y(n17087) );
  sky130_fd_sc_hd__nand3_1 U23934 ( .A(n17088), .B(n17087), .C(n17086), .Y(
        n17090) );
  sky130_fd_sc_hd__o21ai_1 U23935 ( .A1(n17090), .A2(n17089), .B1(n13388), .Y(
        n17091) );
  sky130_fd_sc_hd__nand3_1 U23936 ( .A(n17093), .B(n17092), .C(n17091), .Y(
        n17095) );
  sky130_fd_sc_hd__nand2_1 U23937 ( .A(n17095), .B(n17094), .Y(n17096) );
  sky130_fd_sc_hd__a22oi_1 U23938 ( .A1(n21675), .A2(
        j202_soc_core_uart_div0[3]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[91]), .Y(n17103) );
  sky130_fd_sc_hd__nand2_1 U23939 ( .A(n21699), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[59]), .Y(n17102) );
  sky130_fd_sc_hd__nand4_1 U23940 ( .A(n17104), .B(n17103), .C(n21677), .D(
        n17102), .Y(n17100) );
  sky130_fd_sc_hd__a21oi_1 U23941 ( .A1(j202_soc_core_memory0_ram_dout0[443]), 
        .A2(n21598), .B1(n17100), .Y(n17101) );
  sky130_fd_sc_hd__nand4_1 U23942 ( .A(n17104), .B(n17103), .C(n21738), .D(
        n17102), .Y(n17105) );
  sky130_fd_sc_hd__nor2_1 U23943 ( .A(n17111), .B(n17108), .Y(n17113) );
  sky130_fd_sc_hd__o21ai_1 U23944 ( .A1(n17111), .A2(n17110), .B1(n17109), .Y(
        n17112) );
  sky130_fd_sc_hd__a21oi_1 U23945 ( .A1(n22513), .A2(n17113), .B1(n17112), .Y(
        n17117) );
  sky130_fd_sc_hd__nand2_1 U23946 ( .A(n17115), .B(n17114), .Y(n17116) );
  sky130_fd_sc_hd__xor2_1 U23947 ( .A(n17117), .B(n17116), .X(n23786) );
  sky130_fd_sc_hd__ha_1 U23948 ( .A(n17118), .B(j202_soc_core_j22_cpu_pc[27]), 
        .COUT(n16647), .SUM(n23785) );
  sky130_fd_sc_hd__o22ai_1 U23949 ( .A1(n25151), .A2(n13603), .B1(n26707), 
        .B2(n11143), .Y(n17119) );
  sky130_fd_sc_hd__a21oi_1 U23950 ( .A1(n17120), .A2(n24671), .B1(n17119), .Y(
        n17122) );
  sky130_fd_sc_hd__nand2b_1 U23951 ( .A_N(n21584), .B(n23785), .Y(n17121) );
  sky130_fd_sc_hd__o211ai_1 U23952 ( .A1(n27375), .A2(n22592), .B1(n17122), 
        .C1(n17121), .Y(n17123) );
  sky130_fd_sc_hd__a21oi_1 U23953 ( .A1(n23786), .A2(n12158), .B1(n17123), .Y(
        n17124) );
  sky130_fd_sc_hd__nand2_1 U23954 ( .A(n27823), .B(n29356), .Y(n17143) );
  sky130_fd_sc_hd__inv_1 U23955 ( .A(n17127), .Y(n17128) );
  sky130_fd_sc_hd__nor2_1 U23956 ( .A(n12465), .B(n28919), .Y(n17134) );
  sky130_fd_sc_hd__nor2_1 U23957 ( .A(n28920), .B(n10939), .Y(n17132) );
  sky130_fd_sc_hd__nand4_1 U23959 ( .A(n17135), .B(n17150), .C(n17152), .D(
        n10957), .Y(n17136) );
  sky130_fd_sc_hd__inv_1 U23960 ( .A(n17136), .Y(n17139) );
  sky130_fd_sc_hd__inv_2 U23961 ( .A(n17144), .Y(n17145) );
  sky130_fd_sc_hd__inv_1 U23962 ( .A(n29518), .Y(n17147) );
  sky130_fd_sc_hd__nand3_1 U23963 ( .A(n10957), .B(n21024), .C(n17147), .Y(
        n20978) );
  sky130_fd_sc_hd__nor2_1 U23964 ( .A(n12465), .B(n17149), .Y(n25226) );
  sky130_fd_sc_hd__nand4_1 U23966 ( .A(n25226), .B(n17153), .C(n17152), .D(
        n17151), .Y(n24125) );
  sky130_fd_sc_hd__nor2_1 U23967 ( .A(io_in[14]), .B(n17154), .Y(n20979) );
  sky130_fd_sc_hd__nor2_1 U23968 ( .A(n20979), .B(n17155), .Y(n17156) );
  sky130_fd_sc_hd__mux2i_1 U23969 ( .A0(n24123), .A1(n12400), .S(n17156), .Y(
        n17157) );
  sky130_fd_sc_hd__a21oi_1 U23970 ( .A1(n12400), .A2(n24123), .B1(n17157), .Y(
        n17158) );
  sky130_fd_sc_hd__nand2_1 U23971 ( .A(j202_soc_core_memory0_ram_dout0[322]), 
        .B(n21593), .Y(n17241) );
  sky130_fd_sc_hd__nand2_1 U23972 ( .A(j202_soc_core_memory0_ram_dout0[258]), 
        .B(n21605), .Y(n17240) );
  sky130_fd_sc_hd__nand2_1 U23973 ( .A(j202_soc_core_memory0_ram_dout0[386]), 
        .B(n21597), .Y(n17239) );
  sky130_fd_sc_hd__nand2_1 U23974 ( .A(n17175), .B(n17293), .Y(n20925) );
  sky130_fd_sc_hd__nand2b_1 U23975 ( .A_N(n20784), .B(n20623), .Y(n20306) );
  sky130_fd_sc_hd__nand2_1 U23976 ( .A(n19125), .B(n20623), .Y(n19086) );
  sky130_fd_sc_hd__nand2b_1 U23977 ( .A_N(n17168), .B(n17162), .Y(n20047) );
  sky130_fd_sc_hd__nor2_1 U23978 ( .A(n20011), .B(n20871), .Y(n20207) );
  sky130_fd_sc_hd__nand2_1 U23979 ( .A(n17163), .B(n17170), .Y(n20201) );
  sky130_fd_sc_hd__nor2_1 U23980 ( .A(n20687), .B(n17279), .Y(n17226) );
  sky130_fd_sc_hd__nand2_1 U23981 ( .A(n17167), .B(n17226), .Y(n20885) );
  sky130_fd_sc_hd__nand2_1 U23982 ( .A(n20384), .B(n20885), .Y(n20883) );
  sky130_fd_sc_hd__nand2_1 U23983 ( .A(n17301), .B(n20687), .Y(n17191) );
  sky130_fd_sc_hd__nor2_1 U23984 ( .A(n17164), .B(n17191), .Y(n20094) );
  sky130_fd_sc_hd__nand2_1 U23985 ( .A(n19125), .B(n20687), .Y(n19873) );
  sky130_fd_sc_hd__nand2b_1 U23986 ( .A_N(n17191), .B(n17193), .Y(n20920) );
  sky130_fd_sc_hd__nor2_1 U23988 ( .A(n20094), .B(n20355), .Y(n19119) );
  sky130_fd_sc_hd__nand2_1 U23989 ( .A(n17221), .B(n19119), .Y(n19875) );
  sky130_fd_sc_hd__nor2_1 U23990 ( .A(n17165), .B(n17211), .Y(n20872) );
  sky130_fd_sc_hd__nor2_1 U23991 ( .A(n19121), .B(n17283), .Y(n19841) );
  sky130_fd_sc_hd__nand2_1 U23992 ( .A(n19841), .B(n20687), .Y(n19969) );
  sky130_fd_sc_hd__nor2_1 U23993 ( .A(n20872), .B(n19830), .Y(n20065) );
  sky130_fd_sc_hd__nand2b_1 U23994 ( .A_N(n21206), .B(n20687), .Y(n20842) );
  sky130_fd_sc_hd__nor2_1 U23995 ( .A(n17279), .B(n17166), .Y(n20079) );
  sky130_fd_sc_hd__nand2_1 U23996 ( .A(n20079), .B(n20623), .Y(n20074) );
  sky130_fd_sc_hd__nor2_1 U23997 ( .A(n20687), .B(n17290), .Y(n17192) );
  sky130_fd_sc_hd__nand2b_1 U23998 ( .A_N(n19874), .B(n17192), .Y(n20372) );
  sky130_fd_sc_hd__nand2_1 U23999 ( .A(n20074), .B(n20372), .Y(n17219) );
  sky130_fd_sc_hd__nor2_1 U24000 ( .A(n20924), .B(n17219), .Y(n20013) );
  sky130_fd_sc_hd__nand2_1 U24001 ( .A(n20065), .B(n20013), .Y(n19881) );
  sky130_fd_sc_hd__nor3b_1 U24002 ( .C_N(n20207), .A(n19875), .B(n19881), .Y(
        n17180) );
  sky130_fd_sc_hd__nand2_1 U24003 ( .A(n17175), .B(n17289), .Y(n20906) );
  sky130_fd_sc_hd__nand2b_1 U24004 ( .A_N(n20350), .B(n20687), .Y(n20326) );
  sky130_fd_sc_hd__nand2_1 U24005 ( .A(n19841), .B(n20623), .Y(n20007) );
  sky130_fd_sc_hd__nand2_1 U24006 ( .A(n17271), .B(n20687), .Y(n19120) );
  sky130_fd_sc_hd__nand2b_1 U24007 ( .A_N(n19120), .B(n17193), .Y(n20202) );
  sky130_fd_sc_hd__nand2_1 U24008 ( .A(n20007), .B(n20202), .Y(n20096) );
  sky130_fd_sc_hd__nand2b_1 U24009 ( .A_N(n19120), .B(n17167), .Y(n20118) );
  sky130_fd_sc_hd__nand2_1 U24010 ( .A(n20079), .B(n20687), .Y(n20308) );
  sky130_fd_sc_hd__nor2_1 U24011 ( .A(n20623), .B(n17279), .Y(n17194) );
  sky130_fd_sc_hd__nand2_1 U24012 ( .A(n17167), .B(n17194), .Y(n20376) );
  sky130_fd_sc_hd__nand2_1 U24013 ( .A(n20308), .B(n20376), .Y(n20167) );
  sky130_fd_sc_hd__nor2_1 U24014 ( .A(n19847), .B(n20167), .Y(n19946) );
  sky130_fd_sc_hd__nand2_1 U24015 ( .A(n19946), .B(n20784), .Y(n20225) );
  sky130_fd_sc_hd__nor4_1 U24016 ( .A(n20916), .B(n20110), .C(n20096), .D(
        n20225), .Y(n17178) );
  sky130_fd_sc_hd__nand2_1 U24017 ( .A(n12137), .B(n17289), .Y(n20873) );
  sky130_fd_sc_hd__nand2_1 U24018 ( .A(n17167), .B(n17192), .Y(n20377) );
  sky130_fd_sc_hd__nand2_1 U24019 ( .A(n20885), .B(n20377), .Y(n20082) );
  sky130_fd_sc_hd__nor2_1 U24020 ( .A(n20863), .B(n20011), .Y(n20060) );
  sky130_fd_sc_hd__nand2b_1 U24021 ( .A_N(n20784), .B(n20687), .Y(n20328) );
  sky130_fd_sc_hd__nand2_1 U24022 ( .A(n20328), .B(n20007), .Y(n17171) );
  sky130_fd_sc_hd__nor2_1 U24023 ( .A(n17169), .B(n17168), .Y(n19991) );
  sky130_fd_sc_hd__nand2_1 U24024 ( .A(n19991), .B(n20623), .Y(n20099) );
  sky130_fd_sc_hd__nand2_1 U24025 ( .A(n17192), .B(n17170), .Y(n20375) );
  sky130_fd_sc_hd__nand2_1 U24026 ( .A(n20099), .B(n20375), .Y(n20300) );
  sky130_fd_sc_hd__nand4_1 U24027 ( .A(n17206), .B(n20060), .C(n20378), .D(
        n19995), .Y(n19883) );
  sky130_fd_sc_hd__nand2_1 U24028 ( .A(n20306), .B(n20074), .Y(n20252) );
  sky130_fd_sc_hd__nor2_1 U24029 ( .A(n17171), .B(n20252), .Y(n17174) );
  sky130_fd_sc_hd__nor2b_1 U24030 ( .B_N(n20065), .A(n20863), .Y(n19967) );
  sky130_fd_sc_hd__nand2b_1 U24031 ( .A_N(n19873), .B(n19085), .Y(n20843) );
  sky130_fd_sc_hd__nand2_1 U24032 ( .A(n19971), .B(n20843), .Y(n20887) );
  sky130_fd_sc_hd__nor2_1 U24033 ( .A(n17172), .B(n20887), .Y(n19994) );
  sky130_fd_sc_hd__nand2b_1 U24034 ( .A_N(n17191), .B(n17173), .Y(n20054) );
  sky130_fd_sc_hd__nor2_1 U24035 ( .A(n20110), .B(n20302), .Y(n17190) );
  sky130_fd_sc_hd__nand2b_1 U24036 ( .A_N(n20350), .B(n20623), .Y(n20305) );
  sky130_fd_sc_hd__nand4_1 U24037 ( .A(n17174), .B(n19994), .C(n17190), .D(
        n20305), .Y(n17176) );
  sky130_fd_sc_hd__nor2_1 U24038 ( .A(n17289), .B(n17175), .Y(n20864) );
  sky130_fd_sc_hd__a22oi_1 U24039 ( .A1(n20892), .A2(n19883), .B1(n17176), 
        .B2(n20864), .Y(n17177) );
  sky130_fd_sc_hd__o21a_1 U24040 ( .A1(n20906), .A2(n17178), .B1(n17177), .X(
        n17179) );
  sky130_fd_sc_hd__o21ai_1 U24041 ( .A1(n20925), .A2(n17180), .B1(n17179), .Y(
        n17181) );
  sky130_fd_sc_hd__nand2_1 U24042 ( .A(n17181), .B(n21697), .Y(n17253) );
  sky130_fd_sc_hd__nand2_1 U24043 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_period[2]), .Y(n17249) );
  sky130_fd_sc_hd__nand3_1 U24044 ( .A(n17183), .B(n17182), .C(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[0]), .Y(n17185) );
  sky130_fd_sc_hd__nor2_1 U24045 ( .A(n17185), .B(n17184), .Y(n21698) );
  sky130_fd_sc_hd__a22oi_1 U24046 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[34]), .B1(n21698), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[98]), .Y(n17243) );
  sky130_fd_sc_hd__nor2_1 U24047 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[1]), 
        .B(n27137), .Y(n24376) );
  sky130_fd_sc_hd__nor2_1 U24048 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[0]), 
        .B(j202_soc_core_uart_TOP_rx_fifo_rp[1]), .Y(n21669) );
  sky130_fd_sc_hd__a22oi_1 U24049 ( .A1(n24376), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[18]), .B1(n21669), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[26]), .Y(n17187) );
  sky130_fd_sc_hd__nor2_1 U24050 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[0]), 
        .B(n24378), .Y(n21667) );
  sky130_fd_sc_hd__a22oi_1 U24051 ( .A1(n21667), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[10]), .B1(n21668), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[2]), .Y(n17186) );
  sky130_fd_sc_hd__nand2_1 U24052 ( .A(n17187), .B(n17186), .Y(n17188) );
  sky130_fd_sc_hd__nand2_1 U24053 ( .A(n17188), .B(n21675), .Y(n17244) );
  sky130_fd_sc_hd__nand2_1 U24054 ( .A(n21666), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[66]), .Y(n17247) );
  sky130_fd_sc_hd__nand4_1 U24055 ( .A(n17243), .B(n21677), .C(n17244), .D(
        n17247), .Y(n17189) );
  sky130_fd_sc_hd__nor2b_1 U24056 ( .B_N(n17249), .A(n17189), .Y(n17205) );
  sky130_fd_sc_hd__nor2_1 U24057 ( .A(n19874), .B(n19120), .Y(n20312) );
  sky130_fd_sc_hd__nor3_1 U24058 ( .A(n20312), .B(n20363), .C(n20883), .Y(
        n20006) );
  sky130_fd_sc_hd__nor2_1 U24059 ( .A(n20918), .B(n20871), .Y(n20374) );
  sky130_fd_sc_hd__nor2_1 U24060 ( .A(n20924), .B(n19985), .Y(n19947) );
  sky130_fd_sc_hd__nand2_1 U24061 ( .A(n19947), .B(n13302), .Y(n20251) );
  sky130_fd_sc_hd__o21ai_0 U24062 ( .A1(n19905), .A2(n20251), .B1(n20912), .Y(
        n17198) );
  sky130_fd_sc_hd__nand2b_1 U24063 ( .A_N(n17191), .B(n17287), .Y(n20221) );
  sky130_fd_sc_hd__nand2_1 U24064 ( .A(n20221), .B(n20117), .Y(n20323) );
  sky130_fd_sc_hd__nor2_1 U24065 ( .A(n20924), .B(n19898), .Y(n20361) );
  sky130_fd_sc_hd__nand2b_1 U24066 ( .A_N(n19874), .B(n17194), .Y(n20919) );
  sky130_fd_sc_hd__nand2_1 U24067 ( .A(n20843), .B(n20919), .Y(n20226) );
  sky130_fd_sc_hd__nor2_1 U24068 ( .A(n20871), .B(n20226), .Y(n19952) );
  sky130_fd_sc_hd__nand2_1 U24069 ( .A(n19991), .B(n20687), .Y(n20298) );
  sky130_fd_sc_hd__nand2_1 U24070 ( .A(n20308), .B(n19969), .Y(n20380) );
  sky130_fd_sc_hd__nor2_1 U24071 ( .A(n20313), .B(n20380), .Y(n19986) );
  sky130_fd_sc_hd__nand4_1 U24072 ( .A(n20008), .B(n20361), .C(n19952), .D(
        n19986), .Y(n17195) );
  sky130_fd_sc_hd__nand2_1 U24073 ( .A(n17195), .B(n20335), .Y(n17197) );
  sky130_fd_sc_hd__nand2_1 U24074 ( .A(n19125), .B(n19380), .Y(n17299) );
  sky130_fd_sc_hd__nand2b_1 U24075 ( .A_N(n17299), .B(n20623), .Y(n20214) );
  sky130_fd_sc_hd__nor2_1 U24076 ( .A(n19832), .B(n17228), .Y(n20850) );
  sky130_fd_sc_hd__nand2_1 U24077 ( .A(n20850), .B(n19971), .Y(n19876) );
  sky130_fd_sc_hd__nand4_1 U24079 ( .A(n17199), .B(n17198), .C(n17197), .D(
        n17196), .Y(n17200) );
  sky130_fd_sc_hd__nand2_1 U24080 ( .A(n17200), .B(n13481), .Y(n17251) );
  sky130_fd_sc_hd__nand2_1 U24081 ( .A(n28915), .B(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[2]), .Y(n17202) );
  sky130_fd_sc_hd__nand3_1 U24082 ( .A(n17201), .B(j202_soc_core_aquc_ADR__3_), 
        .C(n20157), .Y(n20154) );
  sky130_fd_sc_hd__nor2_1 U24083 ( .A(n25677), .B(n19858), .Y(n24809) );
  sky130_fd_sc_hd__nand3_1 U24084 ( .A(n24809), .B(n28915), .C(
        j202_soc_core_aquc_ADR__2_), .Y(n20160) );
  sky130_fd_sc_hd__o22ai_1 U24085 ( .A1(n17202), .A2(n20154), .B1(n22996), 
        .B2(n20160), .Y(n17204) );
  sky130_fd_sc_hd__nand2_1 U24086 ( .A(n17204), .B(n20164), .Y(n17250) );
  sky130_fd_sc_hd__nand4_1 U24087 ( .A(n17253), .B(n17205), .C(n17251), .D(
        n17250), .Y(n17237) );
  sky130_fd_sc_hd__nand2_1 U24088 ( .A(n20384), .B(n20117), .Y(n19114) );
  sky130_fd_sc_hd__nand2_1 U24089 ( .A(n17206), .B(n19897), .Y(n19900) );
  sky130_fd_sc_hd__nand3_1 U24090 ( .A(n20018), .B(n20375), .C(n20080), .Y(
        n19845) );
  sky130_fd_sc_hd__nor4b_1 U24091 ( .D_N(n20374), .A(n19832), .B(n19845), .C(
        n20167), .Y(n17207) );
  sky130_fd_sc_hd__nor3_1 U24092 ( .A(n20924), .B(n19848), .C(n19847), .Y(
        n19829) );
  sky130_fd_sc_hd__nand2_1 U24093 ( .A(n17207), .B(n19829), .Y(n17208) );
  sky130_fd_sc_hd__nand2_1 U24094 ( .A(n17208), .B(n20864), .Y(n17216) );
  sky130_fd_sc_hd__nand2_1 U24095 ( .A(n17221), .B(n20214), .Y(n19944) );
  sky130_fd_sc_hd__nor4_1 U24096 ( .A(n20917), .B(n20010), .C(n20301), .D(
        n19944), .Y(n17210) );
  sky130_fd_sc_hd__nand2_1 U24097 ( .A(n20896), .B(n20308), .Y(n20238) );
  sky130_fd_sc_hd__nand2b_1 U24098 ( .A_N(n17219), .B(n20843), .Y(n19973) );
  sky130_fd_sc_hd__o21ai_1 U24099 ( .A1(n20238), .A2(n19973), .B1(n20912), .Y(
        n17209) );
  sky130_fd_sc_hd__nor2_1 U24101 ( .A(n17300), .B(n17211), .Y(n19097) );
  sky130_fd_sc_hd__nand2_1 U24102 ( .A(n20054), .B(n20298), .Y(n20105) );
  sky130_fd_sc_hd__nor4_1 U24103 ( .A(n20010), .B(n19097), .C(n20226), .D(
        n20105), .Y(n17212) );
  sky130_fd_sc_hd__nand2_1 U24104 ( .A(n20884), .B(n20221), .Y(n20904) );
  sky130_fd_sc_hd__a31oi_1 U24105 ( .A1(n17212), .A2(n19135), .A3(n17220), 
        .B1(n20925), .Y(n17213) );
  sky130_fd_sc_hd__nor2_1 U24106 ( .A(n17214), .B(n17213), .Y(n17215) );
  sky130_fd_sc_hd__a21oi_1 U24107 ( .A1(n17216), .A2(n17215), .B1(n19856), .Y(
        n17254) );
  sky130_fd_sc_hd__nand2_1 U24108 ( .A(n20306), .B(n19947), .Y(n20188) );
  sky130_fd_sc_hd__nand2_1 U24109 ( .A(n20202), .B(n20884), .Y(n20349) );
  sky130_fd_sc_hd__nand2_1 U24110 ( .A(n20063), .B(n20328), .Y(n20197) );
  sky130_fd_sc_hd__nand2_1 U24111 ( .A(n20007), .B(n20080), .Y(n17217) );
  sky130_fd_sc_hd__nor4_1 U24112 ( .A(n20188), .B(n20197), .C(n20238), .D(
        n17217), .Y(n17218) );
  sky130_fd_sc_hd__a31oi_1 U24113 ( .A1(n20352), .A2(n17218), .A3(n20326), 
        .B1(n20927), .Y(n17233) );
  sky130_fd_sc_hd__nor2_1 U24114 ( .A(n20917), .B(n17223), .Y(n19831) );
  sky130_fd_sc_hd__nand2_1 U24115 ( .A(n17220), .B(n20054), .Y(n20176) );
  sky130_fd_sc_hd__nand2_1 U24116 ( .A(n17221), .B(n20377), .Y(n20097) );
  sky130_fd_sc_hd__nor4_1 U24117 ( .A(n20058), .B(n20096), .C(n20176), .D(
        n20097), .Y(n17222) );
  sky130_fd_sc_hd__a31oi_1 U24118 ( .A1(n19831), .A2(n20358), .A3(n17222), 
        .B1(n20925), .Y(n17232) );
  sky130_fd_sc_hd__nor2_1 U24119 ( .A(n20180), .B(n19898), .Y(n19836) );
  sky130_fd_sc_hd__nor2_1 U24120 ( .A(n20059), .B(n17223), .Y(n17225) );
  sky130_fd_sc_hd__nand2_1 U24121 ( .A(n20247), .B(n20884), .Y(n19886) );
  sky130_fd_sc_hd__nand3_1 U24122 ( .A(n13302), .B(n20843), .C(n20202), .Y(
        n19833) );
  sky130_fd_sc_hd__nor3_1 U24123 ( .A(n19900), .B(n19886), .C(n19833), .Y(
        n17224) );
  sky130_fd_sc_hd__a31oi_1 U24124 ( .A1(n19836), .A2(n17225), .A3(n17224), 
        .B1(n20873), .Y(n17231) );
  sky130_fd_sc_hd__nand2b_1 U24125 ( .A_N(n19874), .B(n17226), .Y(n20199) );
  sky130_fd_sc_hd__nand2_1 U24126 ( .A(n20376), .B(n20199), .Y(n20219) );
  sky130_fd_sc_hd__nor2_1 U24127 ( .A(n20079), .B(n20219), .Y(n19950) );
  sky130_fd_sc_hd__nand2_1 U24128 ( .A(n20003), .B(n20884), .Y(n20076) );
  sky130_fd_sc_hd__nor2_1 U24129 ( .A(n17227), .B(n20076), .Y(n20232) );
  sky130_fd_sc_hd__nand2_1 U24130 ( .A(n19112), .B(n20298), .Y(n20175) );
  sky130_fd_sc_hd__nand2_1 U24131 ( .A(n20073), .B(n20328), .Y(n20336) );
  sky130_fd_sc_hd__nand2_1 U24132 ( .A(n19951), .B(n20326), .Y(n20388) );
  sky130_fd_sc_hd__nor3_1 U24133 ( .A(n17228), .B(n20175), .C(n20388), .Y(
        n17229) );
  sky130_fd_sc_hd__a31oi_1 U24134 ( .A1(n19950), .A2(n20232), .A3(n17229), 
        .B1(n20906), .Y(n17230) );
  sky130_fd_sc_hd__nor4_1 U24135 ( .A(n17233), .B(n17232), .C(n17231), .D(
        n17230), .Y(n17234) );
  sky130_fd_sc_hd__nand2b_1 U24136 ( .A_N(n17234), .B(n20908), .Y(n17236) );
  sky130_fd_sc_hd__nand2_1 U24137 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[2]), .Y(n17235) );
  sky130_fd_sc_hd__nand2_1 U24138 ( .A(n17236), .B(n17235), .Y(n17242) );
  sky130_fd_sc_hd__nor3_1 U24139 ( .A(n17237), .B(n17254), .C(n17242), .Y(
        n17238) );
  sky130_fd_sc_hd__nand2_1 U24140 ( .A(j202_soc_core_memory0_ram_dout0[482]), 
        .B(n21771), .Y(n17258) );
  sky130_fd_sc_hd__nor2_1 U24141 ( .A(n17246), .B(n17245), .Y(n17248) );
  sky130_fd_sc_hd__and4_1 U24142 ( .A(n17249), .B(n17248), .C(n21738), .D(
        n17247), .X(n17252) );
  sky130_fd_sc_hd__nand4_1 U24143 ( .A(n17253), .B(n17252), .C(n17251), .D(
        n17250), .Y(n17255) );
  sky130_fd_sc_hd__nor2_1 U24144 ( .A(n17255), .B(n17254), .Y(n17256) );
  sky130_fd_sc_hd__nand3_1 U24145 ( .A(n17258), .B(n17257), .C(n17256), .Y(
        n20711) );
  sky130_fd_sc_hd__nand2_1 U24146 ( .A(n20712), .B(n20711), .Y(n23696) );
  sky130_fd_sc_hd__nand2b_1 U24147 ( .A_N(n23696), .B(n22581), .Y(n17270) );
  sky130_fd_sc_hd__nand2_1 U24148 ( .A(n17261), .B(n17260), .Y(n17264) );
  sky130_fd_sc_hd__xnor2_1 U24150 ( .A(n17264), .B(n17263), .Y(n25235) );
  sky130_fd_sc_hd__nand2_1 U24151 ( .A(n25235), .B(n12158), .Y(n17267) );
  sky130_fd_sc_hd__xnor2_1 U24152 ( .A(j202_soc_core_j22_cpu_pc[1]), .B(n19203), .Y(n25244) );
  sky130_fd_sc_hd__nand2_1 U24153 ( .A(n22596), .B(n25244), .Y(n17266) );
  sky130_fd_sc_hd__nand2_1 U24154 ( .A(n22510), .B(n23920), .Y(n17265) );
  sky130_fd_sc_hd__and3_1 U24155 ( .A(n17267), .B(n17266), .C(n17265), .X(
        n17269) );
  sky130_fd_sc_hd__nand2_1 U24156 ( .A(n22515), .B(n27435), .Y(n17268) );
  sky130_fd_sc_hd__nand3_1 U24157 ( .A(n17270), .B(n17269), .C(n17268), .Y(
        n29012) );
  sky130_fd_sc_hd__nand3_1 U24158 ( .A(n13387), .B(n17271), .C(n19354), .Y(
        n19352) );
  sky130_fd_sc_hd__nand2_1 U24159 ( .A(n17284), .B(n17277), .Y(n21613) );
  sky130_fd_sc_hd__nand3_1 U24160 ( .A(n17314), .B(n20788), .C(n19354), .Y(
        n17281) );
  sky130_fd_sc_hd__nand3_1 U24161 ( .A(n13387), .B(n17329), .C(n17274), .Y(
        n20772) );
  sky130_fd_sc_hd__nand2_1 U24162 ( .A(n13388), .B(n19381), .Y(n21169) );
  sky130_fd_sc_hd__nor2_1 U24163 ( .A(n20788), .B(n21170), .Y(n17272) );
  sky130_fd_sc_hd__nand2b_1 U24164 ( .A_N(n21169), .B(n17272), .Y(n21134) );
  sky130_fd_sc_hd__nand2_1 U24165 ( .A(n17273), .B(n17274), .Y(n17330) );
  sky130_fd_sc_hd__nand2b_1 U24166 ( .A_N(n17330), .B(n12181), .Y(n20747) );
  sky130_fd_sc_hd__nand2b_1 U24167 ( .A_N(n20747), .B(n20579), .Y(n21606) );
  sky130_fd_sc_hd__nand3_1 U24168 ( .A(n17328), .B(n21134), .C(n21606), .Y(
        n21713) );
  sky130_fd_sc_hd__nand2_1 U24169 ( .A(n21614), .B(n21221), .Y(n19356) );
  sky130_fd_sc_hd__nand2_1 U24170 ( .A(n13388), .B(n17274), .Y(n17280) );
  sky130_fd_sc_hd__nand2b_1 U24171 ( .A_N(n17280), .B(n12181), .Y(n18927) );
  sky130_fd_sc_hd__a31oi_1 U24172 ( .A1(n20755), .A2(n17275), .A3(n18927), 
        .B1(n21722), .Y(n17297) );
  sky130_fd_sc_hd__nand2b_1 U24173 ( .A_N(n17299), .B(n13387), .Y(n21706) );
  sky130_fd_sc_hd__nand2b_1 U24174 ( .A_N(n18952), .B(n20788), .Y(n21243) );
  sky130_fd_sc_hd__nand2_1 U24175 ( .A(n21243), .B(n21614), .Y(n21714) );
  sky130_fd_sc_hd__nor2_1 U24176 ( .A(n19271), .B(n21714), .Y(n20752) );
  sky130_fd_sc_hd__nand2_1 U24177 ( .A(n21221), .B(n20772), .Y(n21618) );
  sky130_fd_sc_hd__nand2_1 U24178 ( .A(n20778), .B(n17277), .Y(n21246) );
  sky130_fd_sc_hd__nor2_1 U24179 ( .A(n17279), .B(n17278), .Y(n21184) );
  sky130_fd_sc_hd__nand2_1 U24180 ( .A(n21246), .B(n21268), .Y(n21115) );
  sky130_fd_sc_hd__nor2_1 U24181 ( .A(n21618), .B(n21115), .Y(n21708) );
  sky130_fd_sc_hd__nor2_1 U24182 ( .A(n17281), .B(n17280), .Y(n21620) );
  sky130_fd_sc_hd__nor2_1 U24183 ( .A(n17283), .B(n17282), .Y(n21102) );
  sky130_fd_sc_hd__nand2_1 U24184 ( .A(n21102), .B(n17314), .Y(n21685) );
  sky130_fd_sc_hd__nand2_1 U24185 ( .A(n21269), .B(n21685), .Y(n21279) );
  sky130_fd_sc_hd__nand2_1 U24186 ( .A(n17284), .B(n17314), .Y(n21094) );
  sky130_fd_sc_hd__nand3_1 U24187 ( .A(n21708), .B(n19335), .C(n21094), .Y(
        n20734) );
  sky130_fd_sc_hd__a21oi_1 U24188 ( .A1(n17285), .A2(n19125), .B1(n20734), .Y(
        n17286) );
  sky130_fd_sc_hd__a21oi_1 U24189 ( .A1(n20752), .A2(n17286), .B1(n21705), .Y(
        n17296) );
  sky130_fd_sc_hd__nand2_1 U24190 ( .A(n17287), .B(n17301), .Y(n20849) );
  sky130_fd_sc_hd__nand2_1 U24191 ( .A(n13387), .B(n20172), .Y(n21245) );
  sky130_fd_sc_hd__nand2_1 U24192 ( .A(n21184), .B(n13396), .Y(n21287) );
  sky130_fd_sc_hd__nor3_1 U24193 ( .A(n21719), .B(n17288), .C(n21618), .Y(
        n21633) );
  sky130_fd_sc_hd__nand2_1 U24194 ( .A(n20687), .B(n17289), .Y(n21720) );
  sky130_fd_sc_hd__nand2_1 U24195 ( .A(n17302), .B(n19381), .Y(n20790) );
  sky130_fd_sc_hd__nor2_1 U24196 ( .A(n17300), .B(n20790), .Y(n21095) );
  sky130_fd_sc_hd__nand2_1 U24197 ( .A(n21095), .B(n20788), .Y(n21190) );
  sky130_fd_sc_hd__nand2_1 U24198 ( .A(n21207), .B(n20579), .Y(n21628) );
  sky130_fd_sc_hd__nor2_1 U24199 ( .A(n17290), .B(n19874), .Y(n20045) );
  sky130_fd_sc_hd__nand2_1 U24200 ( .A(n20045), .B(n12137), .Y(n21688) );
  sky130_fd_sc_hd__nand3_1 U24201 ( .A(n13387), .B(n19355), .C(n12181), .Y(
        n21631) );
  sky130_fd_sc_hd__nand2_1 U24202 ( .A(n21688), .B(n21631), .Y(n21265) );
  sky130_fd_sc_hd__nand2b_1 U24203 ( .A_N(n18927), .B(n20579), .Y(n21648) );
  sky130_fd_sc_hd__nand2_1 U24204 ( .A(n21648), .B(n20747), .Y(n17291) );
  sky130_fd_sc_hd__nor4_1 U24205 ( .A(n17292), .B(n21126), .C(n21265), .D(
        n17291), .Y(n17294) );
  sky130_fd_sc_hd__nand2_1 U24206 ( .A(n17293), .B(n20623), .Y(n21709) );
  sky130_fd_sc_hd__o22ai_1 U24207 ( .A1(n21633), .A2(n21720), .B1(n17294), 
        .B2(n21709), .Y(n17295) );
  sky130_fd_sc_hd__nor3_1 U24208 ( .A(n17297), .B(n17296), .C(n17295), .Y(
        n17298) );
  sky130_fd_sc_hd__nand2b_1 U24209 ( .A_N(n17298), .B(n21727), .Y(n17350) );
  sky130_fd_sc_hd__nand2b_1 U24210 ( .A_N(n17299), .B(n17302), .Y(n21244) );
  sky130_fd_sc_hd__nand2_1 U24211 ( .A(n21244), .B(n21190), .Y(n21285) );
  sky130_fd_sc_hd__nand2b_1 U24212 ( .A_N(n18952), .B(n20579), .Y(n20736) );
  sky130_fd_sc_hd__nor2_1 U24213 ( .A(n17300), .B(n21169), .Y(n19388) );
  sky130_fd_sc_hd__inv_1 U24214 ( .A(n19388), .Y(n19284) );
  sky130_fd_sc_hd__nand2b_1 U24215 ( .A_N(n21285), .B(n21185), .Y(n17315) );
  sky130_fd_sc_hd__nand2_1 U24216 ( .A(n20908), .B(n21288), .Y(n19272) );
  sky130_fd_sc_hd__nand2_1 U24217 ( .A(n17301), .B(n19380), .Y(n18951) );
  sky130_fd_sc_hd__nand2b_1 U24218 ( .A_N(n18951), .B(n13388), .Y(n21186) );
  sky130_fd_sc_hd__nand2b_1 U24219 ( .A_N(n18951), .B(n17302), .Y(n21267) );
  sky130_fd_sc_hd__nand3_1 U24220 ( .A(n21680), .B(n21256), .C(n21267), .Y(
        n21612) );
  sky130_fd_sc_hd__nand2_1 U24221 ( .A(n21256), .B(n21094), .Y(n21617) );
  sky130_fd_sc_hd__nand2b_1 U24222 ( .A_N(n21617), .B(n17328), .Y(n21626) );
  sky130_fd_sc_hd__a22oi_1 U24223 ( .A1(n13275), .A2(n21612), .B1(n21626), 
        .B2(n21063), .Y(n17303) );
  sky130_fd_sc_hd__nand2_1 U24224 ( .A(n21698), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[103]), .Y(n17341) );
  sky130_fd_sc_hd__nand2_1 U24225 ( .A(n21667), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[15]), .Y(n17307) );
  sky130_fd_sc_hd__nand2_1 U24226 ( .A(n24376), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[23]), .Y(n17306) );
  sky130_fd_sc_hd__nand2_1 U24227 ( .A(n21668), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[7]), .Y(n17305) );
  sky130_fd_sc_hd__nand2_1 U24228 ( .A(n21669), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[31]), .Y(n17304) );
  sky130_fd_sc_hd__nand4_1 U24229 ( .A(n17307), .B(n17306), .C(n17305), .D(
        n17304), .Y(n17308) );
  sky130_fd_sc_hd__nand2_1 U24230 ( .A(n21675), .B(n17308), .Y(n17340) );
  sky130_fd_sc_hd__nand2_1 U24231 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[7]), .Y(n17339) );
  sky130_fd_sc_hd__nand4_1 U24232 ( .A(n17341), .B(n21677), .C(n17340), .D(
        n17339), .Y(n17312) );
  sky130_fd_sc_hd__nand2_1 U24233 ( .A(n21207), .B(n20788), .Y(n21649) );
  sky130_fd_sc_hd__nand2_1 U24234 ( .A(n19943), .B(n21649), .Y(n20733) );
  sky130_fd_sc_hd__nand3_1 U24235 ( .A(n20908), .B(n21636), .C(n20733), .Y(
        n17311) );
  sky130_fd_sc_hd__nand2_1 U24236 ( .A(n21666), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[71]), .Y(n17310) );
  sky130_fd_sc_hd__nand2_1 U24237 ( .A(n21699), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[39]), .Y(n17309) );
  sky130_fd_sc_hd__nand3_1 U24238 ( .A(n17311), .B(n17310), .C(n17309), .Y(
        n17342) );
  sky130_fd_sc_hd__nor2_1 U24239 ( .A(n17312), .B(n17342), .Y(n17318) );
  sky130_fd_sc_hd__nand2_1 U24240 ( .A(n13481), .B(n21251), .Y(n18958) );
  sky130_fd_sc_hd__nor2_1 U24241 ( .A(n20788), .B(n20787), .Y(n20806) );
  sky130_fd_sc_hd__nor2_1 U24242 ( .A(n17313), .B(n17330), .Y(n21203) );
  sky130_fd_sc_hd__nand2_1 U24243 ( .A(n21203), .B(n17314), .Y(n21286) );
  sky130_fd_sc_hd__nand2_1 U24244 ( .A(n21286), .B(n21267), .Y(n21215) );
  sky130_fd_sc_hd__nand2_1 U24245 ( .A(n21095), .B(n20579), .Y(n21632) );
  sky130_fd_sc_hd__nand2_1 U24246 ( .A(n21632), .B(n21648), .Y(n21205) );
  sky130_fd_sc_hd__nor3_1 U24247 ( .A(n17315), .B(n21714), .C(n21205), .Y(
        n17316) );
  sky130_fd_sc_hd__nand3b_1 U24248 ( .A_N(n21215), .B(n17316), .C(n21186), .Y(
        n17317) );
  sky130_fd_sc_hd__nand2_1 U24249 ( .A(n21198), .B(n17317), .Y(n17345) );
  sky130_fd_sc_hd__nand2_1 U24250 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_period[7]), .Y(n17344) );
  sky130_fd_sc_hd__nand4_1 U24251 ( .A(n19398), .B(n17318), .C(n17345), .D(
        n17344), .Y(n17327) );
  sky130_fd_sc_hd__nand2_1 U24252 ( .A(n21244), .B(n21186), .Y(n21098) );
  sky130_fd_sc_hd__nor2_1 U24253 ( .A(n21098), .B(n17319), .Y(n21689) );
  sky130_fd_sc_hd__a31oi_1 U24254 ( .A1(n21689), .A2(n17328), .A3(n21221), 
        .B1(n21709), .Y(n17326) );
  sky130_fd_sc_hd__nand3_1 U24255 ( .A(n13387), .B(n19381), .C(n17329), .Y(
        n20805) );
  sky130_fd_sc_hd__nand4_1 U24256 ( .A(n19284), .B(n21681), .C(n20805), .D(
        n21134), .Y(n17322) );
  sky130_fd_sc_hd__nand2_1 U24257 ( .A(n21614), .B(n21245), .Y(n17320) );
  sky130_fd_sc_hd__nand2_1 U24258 ( .A(n19388), .B(n20579), .Y(n21270) );
  sky130_fd_sc_hd__nand2_1 U24259 ( .A(n21270), .B(n21094), .Y(n21071) );
  sky130_fd_sc_hd__nor2_1 U24260 ( .A(n17320), .B(n21071), .Y(n21687) );
  sky130_fd_sc_hd__nand2_1 U24261 ( .A(n21687), .B(n21221), .Y(n17321) );
  sky130_fd_sc_hd__a22oi_1 U24262 ( .A1(n21235), .A2(n17322), .B1(n17321), 
        .B2(n21288), .Y(n19393) );
  sky130_fd_sc_hd__nand3_1 U24263 ( .A(n13388), .B(
        j202_soc_core_bootrom_00_address_w[11]), .C(n19355), .Y(n19382) );
  sky130_fd_sc_hd__nor2_1 U24264 ( .A(n21719), .B(n21040), .Y(n19366) );
  sky130_fd_sc_hd__nand2_1 U24265 ( .A(n21628), .B(n21631), .Y(n20759) );
  sky130_fd_sc_hd__nand2_1 U24266 ( .A(n21256), .B(n21244), .Y(n19339) );
  sky130_fd_sc_hd__nor4_1 U24267 ( .A(n20778), .B(n19338), .C(n20759), .D(
        n19339), .Y(n17323) );
  sky130_fd_sc_hd__nor2b_1 U24268 ( .B_N(n21251), .A(n17323), .Y(n17324) );
  sky130_fd_sc_hd__o31a_1 U24269 ( .A1(n17326), .A2(n17325), .A3(n17324), .B1(
        n21697), .X(n17347) );
  sky130_fd_sc_hd__nor2_1 U24270 ( .A(n17327), .B(n17347), .Y(n17337) );
  sky130_fd_sc_hd__a21oi_1 U24271 ( .A1(n17328), .A2(n21628), .B1(n21709), .Y(
        n17336) );
  sky130_fd_sc_hd__nand2b_1 U24272 ( .A_N(n18927), .B(n20788), .Y(n21078) );
  sky130_fd_sc_hd__nand2_1 U24273 ( .A(n21078), .B(n21628), .Y(n18925) );
  sky130_fd_sc_hd__nand2_1 U24274 ( .A(n21710), .B(n21646), .Y(n17332) );
  sky130_fd_sc_hd__nand2b_1 U24275 ( .A_N(n17330), .B(n17329), .Y(n21253) );
  sky130_fd_sc_hd__nand2_1 U24276 ( .A(n21246), .B(n21253), .Y(n21201) );
  sky130_fd_sc_hd__nand2_1 U24277 ( .A(n21190), .B(n21268), .Y(n19376) );
  sky130_fd_sc_hd__nand2b_1 U24278 ( .A_N(n21201), .B(n17331), .Y(n18924) );
  sky130_fd_sc_hd__nor4_1 U24279 ( .A(n17333), .B(n21178), .C(n17332), .D(
        n18924), .Y(n17334) );
  sky130_fd_sc_hd__o22ai_1 U24280 ( .A1(n17334), .A2(n21705), .B1(n21720), 
        .B2(n21650), .Y(n17335) );
  sky130_fd_sc_hd__nand2_1 U24282 ( .A(j202_soc_core_memory0_ram_dout0[487]), 
        .B(n21771), .Y(n17352) );
  sky130_fd_sc_hd__nand4_1 U24283 ( .A(n17341), .B(n21738), .C(n17340), .D(
        n17339), .Y(n17343) );
  sky130_fd_sc_hd__nor2_1 U24284 ( .A(n17343), .B(n17342), .Y(n17346) );
  sky130_fd_sc_hd__nand4_1 U24285 ( .A(n19398), .B(n17346), .C(n17345), .D(
        n17344), .Y(n17348) );
  sky130_fd_sc_hd__nor2_1 U24286 ( .A(n17348), .B(n17347), .Y(n17351) );
  sky130_fd_sc_hd__nand4_1 U24287 ( .A(n17352), .B(n17351), .C(n17350), .D(
        n17349), .Y(n17353) );
  sky130_fd_sc_hd__nand2_4 U24288 ( .A(n17358), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .Y(n25219) );
  sky130_fd_sc_hd__nand2_1 U24289 ( .A(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[0]), .Y(n18863) );
  sky130_fd_sc_hd__nand2_1 U24290 ( .A(n17358), .B(n23252), .Y(n17359) );
  sky130_fd_sc_hd__inv_2 U24291 ( .A(n26977), .Y(n17361) );
  sky130_fd_sc_hd__nand2_1 U24292 ( .A(n18867), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .Y(n18861) );
  sky130_fd_sc_hd__a21oi_1 U24293 ( .A1(j202_soc_core_j22_cpu_ml_mach[31]), 
        .A2(n24499), .B1(n17365), .Y(n22054) );
  sky130_fd_sc_hd__o21ai_1 U24294 ( .A1(n12159), .A2(n18296), .B1(n22054), .Y(
        n22061) );
  sky130_fd_sc_hd__xnor2_1 U24295 ( .A(n18687), .B(n22051), .Y(n17362) );
  sky130_fd_sc_hd__buf_6 U24296 ( .A(j202_soc_core_j22_cpu_ml_bufa[31]), .X(
        n22487) );
  sky130_fd_sc_hd__xnor2_1 U24297 ( .A(j202_soc_core_j22_cpu_ml_bufa[30]), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .Y(n17363) );
  sky130_fd_sc_hd__xnor2_1 U24298 ( .A(n18651), .B(n22487), .Y(n17378) );
  sky130_fd_sc_hd__xor2_1 U24299 ( .A(j202_soc_core_j22_cpu_ml_bufa[31]), .B(
        n24505), .X(n17364) );
  sky130_fd_sc_hd__inv_2 U24300 ( .A(n25219), .Y(n26862) );
  sky130_fd_sc_hd__a22oi_1 U24301 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[30]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[14]), .Y(n17367) );
  sky130_fd_sc_hd__nand2_1 U24302 ( .A(n22071), .B(n17367), .Y(n17375) );
  sky130_fd_sc_hd__xnor2_1 U24303 ( .A(n18651), .B(n22051), .Y(n17368) );
  sky130_fd_sc_hd__buf_2 U24304 ( .A(n12767), .X(n18720) );
  sky130_fd_sc_hd__xnor2_1 U24305 ( .A(n22052), .B(n18720), .Y(n17374) );
  sky130_fd_sc_hd__buf_2 U24306 ( .A(n12767), .X(n18672) );
  sky130_fd_sc_hd__xnor2_1 U24307 ( .A(n18651), .B(n18672), .Y(n18622) );
  sky130_fd_sc_hd__xnor2_1 U24308 ( .A(n17370), .B(n12767), .Y(n17372) );
  sky130_fd_sc_hd__nand2_2 U24309 ( .A(n17372), .B(n17371), .Y(n18747) );
  sky130_fd_sc_hd__o22ai_1 U24310 ( .A1(n18750), .A2(n17374), .B1(n18622), 
        .B2(n18747), .Y(n17382) );
  sky130_fd_sc_hd__xnor2_1 U24311 ( .A(n18721), .B(n22051), .Y(n17373) );
  sky130_fd_sc_hd__a21o_1 U24312 ( .A1(n18750), .A2(n18747), .B1(n17374), .X(
        n18615) );
  sky130_fd_sc_hd__fa_1 U24313 ( .A(n17377), .B(n17376), .CIN(n17375), .COUT(
        n22060), .SUM(n18643) );
  sky130_fd_sc_hd__xnor2_1 U24314 ( .A(n18687), .B(n22487), .Y(n17380) );
  sky130_fd_sc_hd__a22oi_1 U24315 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[29]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[13]), .Y(n17379) );
  sky130_fd_sc_hd__nand2_1 U24316 ( .A(n22071), .B(n17379), .Y(n18626) );
  sky130_fd_sc_hd__xnor2_1 U24317 ( .A(n18721), .B(n22487), .Y(n18623) );
  sky130_fd_sc_hd__xnor2_1 U24318 ( .A(n18685), .B(n22051), .Y(n17381) );
  sky130_fd_sc_hd__nor2_1 U24319 ( .A(n17383), .B(n17384), .Y(n22069) );
  sky130_fd_sc_hd__nand2_1 U24320 ( .A(n17384), .B(n17383), .Y(n22183) );
  sky130_fd_sc_hd__nand2_1 U24321 ( .A(n22185), .B(n22183), .Y(n18860) );
  sky130_fd_sc_hd__xnor2_1 U24322 ( .A(j202_soc_core_j22_cpu_ml_bufa[8]), .B(
        j202_soc_core_j22_cpu_ml_bufa[7]), .Y(n17385) );
  sky130_fd_sc_hd__buf_4 U24323 ( .A(n17385), .X(n18067) );
  sky130_fd_sc_hd__xnor2_1 U24324 ( .A(n18685), .B(n22919), .Y(n17487) );
  sky130_fd_sc_hd__xnor2_1 U24325 ( .A(n18673), .B(n22919), .Y(n17415) );
  sky130_fd_sc_hd__o22ai_1 U24326 ( .A1(n18067), .A2(n17487), .B1(n17415), 
        .B2(n10971), .Y(n17516) );
  sky130_fd_sc_hd__nor2b_1 U24327 ( .B_N(n18353), .A(n12140), .Y(n17489) );
  sky130_fd_sc_hd__buf_4 U24328 ( .A(j202_soc_core_j22_cpu_ml_bufa[7]), .X(
        n19012) );
  sky130_fd_sc_hd__xnor2_1 U24329 ( .A(n18687), .B(n19012), .Y(n17505) );
  sky130_fd_sc_hd__xnor2_1 U24330 ( .A(n18721), .B(n19012), .Y(n17405) );
  sky130_fd_sc_hd__xor2_1 U24331 ( .A(j202_soc_core_j22_cpu_ml_bufa[7]), .B(
        j202_soc_core_j22_cpu_ml_bufa[6]), .X(n17388) );
  sky130_fd_sc_hd__o22ai_1 U24332 ( .A1(n17972), .A2(n17505), .B1(n17405), 
        .B2(n11159), .Y(n17488) );
  sky130_fd_sc_hd__xnor2_1 U24333 ( .A(n17489), .B(n17488), .Y(n17515) );
  sky130_fd_sc_hd__xnor2_1 U24334 ( .A(n18426), .B(n18300), .Y(n17419) );
  sky130_fd_sc_hd__xnor2_1 U24335 ( .A(n18367), .B(n18300), .Y(n17444) );
  sky130_fd_sc_hd__xor2_1 U24336 ( .A(j202_soc_core_j22_cpu_ml_bufa[17]), .B(
        j202_soc_core_j22_cpu_ml_bufa[16]), .X(n17391) );
  sky130_fd_sc_hd__o22ai_1 U24337 ( .A1(n18370), .A2(n17419), .B1(n17444), 
        .B2(n17392), .Y(n17463) );
  sky130_fd_sc_hd__xnor2_1 U24338 ( .A(j202_soc_core_j22_cpu_ml_bufa[2]), .B(
        j202_soc_core_j22_cpu_ml_bufa[1]), .Y(n17393) );
  sky130_fd_sc_hd__xnor2_1 U24339 ( .A(n22052), .B(n24132), .Y(n17408) );
  sky130_fd_sc_hd__xnor2_1 U24340 ( .A(n18651), .B(n24132), .Y(n17448) );
  sky130_fd_sc_hd__xor2_1 U24341 ( .A(j202_soc_core_j22_cpu_ml_bufa[3]), .B(
        n11716), .X(n17395) );
  sky130_fd_sc_hd__buf_2 U24342 ( .A(n17393), .X(n17394) );
  sky130_fd_sc_hd__o22ai_1 U24343 ( .A1(n17805), .A2(n17408), .B1(n17448), 
        .B2(n17802), .Y(n17462) );
  sky130_fd_sc_hd__nand2_1 U24344 ( .A(j202_soc_core_j22_cpu_ml_bufa[12]), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .Y(n17398) );
  sky130_fd_sc_hd__nand2_4 U24345 ( .A(n17397), .B(n17398), .Y(n18224) );
  sky130_fd_sc_hd__buf_6 U24346 ( .A(j202_soc_core_j22_cpu_ml_bufa[13]), .X(
        n21887) );
  sky130_fd_sc_hd__xnor2_1 U24347 ( .A(n18667), .B(n21887), .Y(n17412) );
  sky130_fd_sc_hd__xnor2_1 U24348 ( .A(n18511), .B(n21887), .Y(n17428) );
  sky130_fd_sc_hd__nand2_4 U24349 ( .A(n17399), .B(n18224), .Y(n18225) );
  sky130_fd_sc_hd__o22ai_1 U24350 ( .A1(n18224), .A2(n17412), .B1(n17428), 
        .B2(n18225), .Y(n17461) );
  sky130_fd_sc_hd__xnor2_2 U24351 ( .A(j202_soc_core_j22_cpu_ml_bufa[14]), .B(
        n17400), .Y(n18112) );
  sky130_fd_sc_hd__buf_4 U24352 ( .A(j202_soc_core_j22_cpu_ml_bufa[15]), .X(
        n18883) );
  sky130_fd_sc_hd__xnor2_1 U24353 ( .A(n18479), .B(n18883), .Y(n17416) );
  sky130_fd_sc_hd__xnor2_1 U24354 ( .A(n18466), .B(n18883), .Y(n17442) );
  sky130_fd_sc_hd__xor2_1 U24355 ( .A(j202_soc_core_j22_cpu_ml_bufa[15]), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n17401) );
  sky130_fd_sc_hd__o22ai_1 U24356 ( .A1(n18344), .A2(n17416), .B1(n17442), 
        .B2(n17402), .Y(n17460) );
  sky130_fd_sc_hd__xnor2_1 U24357 ( .A(j202_soc_core_j22_cpu_ml_bufa[10]), .B(
        j202_soc_core_j22_cpu_ml_bufa[9]), .Y(n17403) );
  sky130_fd_sc_hd__xnor2_1 U24358 ( .A(n18654), .B(n18147), .Y(n17413) );
  sky130_fd_sc_hd__xnor2_1 U24359 ( .A(n18649), .B(n18147), .Y(n17446) );
  sky130_fd_sc_hd__xor2_1 U24360 ( .A(n12630), .B(n12708), .X(n17404) );
  sky130_fd_sc_hd__nand2_4 U24361 ( .A(n17404), .B(n18151), .Y(n18148) );
  sky130_fd_sc_hd__o22ai_1 U24362 ( .A1(n18151), .A2(n17413), .B1(n17446), 
        .B2(n18148), .Y(n17459) );
  sky130_fd_sc_hd__xnor2_1 U24363 ( .A(n18661), .B(n22919), .Y(n17414) );
  sky130_fd_sc_hd__xnor2_1 U24364 ( .A(n18708), .B(n22919), .Y(n17466) );
  sky130_fd_sc_hd__o22ai_1 U24365 ( .A1(n18067), .A2(n17414), .B1(n17466), 
        .B2(n10971), .Y(n17458) );
  sky130_fd_sc_hd__xnor2_1 U24366 ( .A(n18685), .B(n19012), .Y(n17441) );
  sky130_fd_sc_hd__xnor2_1 U24367 ( .A(j202_soc_core_j22_cpu_ml_bufa[18]), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .Y(n17406) );
  sky130_fd_sc_hd__xnor2_1 U24368 ( .A(n18367), .B(n22951), .Y(n17471) );
  sky130_fd_sc_hd__buf_2 U24369 ( .A(j202_soc_core_j22_cpu_ml_bufb[0]), .X(
        n18226) );
  sky130_fd_sc_hd__xnor2_1 U24370 ( .A(n22951), .B(n18226), .Y(n17407) );
  sky130_fd_sc_hd__nand2_4 U24371 ( .A(n11058), .B(n18469), .Y(n18470) );
  sky130_fd_sc_hd__o22ai_1 U24372 ( .A1(n12367), .A2(n17471), .B1(n17407), 
        .B2(n18470), .Y(n17410) );
  sky130_fd_sc_hd__a21o_1 U24373 ( .A1(n17802), .A2(n17394), .B1(n17408), .X(
        n17409) );
  sky130_fd_sc_hd__fah_1 U24374 ( .A(n17411), .B(n17410), .CI(n17409), .COUT(
        n17486), .SUM(n17430) );
  sky130_fd_sc_hd__xnor2_1 U24375 ( .A(n18649), .B(n21887), .Y(n17468) );
  sky130_fd_sc_hd__o22ai_1 U24376 ( .A1(n18224), .A2(n17468), .B1(n17412), 
        .B2(n18225), .Y(n17422) );
  sky130_fd_sc_hd__xnor2_1 U24377 ( .A(n18708), .B(n18147), .Y(n17470) );
  sky130_fd_sc_hd__o22ai_1 U24378 ( .A1(n18151), .A2(n17470), .B1(n17413), 
        .B2(n18148), .Y(n17421) );
  sky130_fd_sc_hd__o22ai_1 U24379 ( .A1(n18067), .A2(n17415), .B1(n17414), 
        .B2(n10971), .Y(n17420) );
  sky130_fd_sc_hd__xnor2_1 U24380 ( .A(n18511), .B(n18883), .Y(n17473) );
  sky130_fd_sc_hd__o22ai_1 U24381 ( .A1(n18344), .A2(n17473), .B1(n17416), 
        .B2(n17402), .Y(n17425) );
  sky130_fd_sc_hd__nand2b_1 U24382 ( .A_N(n18353), .B(n22951), .Y(n17418) );
  sky130_fd_sc_hd__o22ai_1 U24383 ( .A1(n12367), .A2(n17418), .B1(n17417), 
        .B2(n18470), .Y(n17424) );
  sky130_fd_sc_hd__xnor2_1 U24384 ( .A(n18466), .B(n18300), .Y(n17469) );
  sky130_fd_sc_hd__o22ai_1 U24385 ( .A1(n18370), .A2(n17469), .B1(n17419), 
        .B2(n17392), .Y(n17423) );
  sky130_fd_sc_hd__fah_1 U24386 ( .A(n17425), .B(n17424), .CI(n17423), .COUT(
        n17484), .SUM(n17478) );
  sky130_fd_sc_hd__xnor2_1 U24387 ( .A(n10968), .B(
        j202_soc_core_j22_cpu_ml_bufa[3]), .Y(n17426) );
  sky130_fd_sc_hd__o22ai_1 U24388 ( .A1(n17786), .A2(n17452), .B1(n17464), 
        .B2(n17771), .Y(n17435) );
  sky130_fd_sc_hd__xnor2_1 U24389 ( .A(n18673), .B(n19012), .Y(n17440) );
  sky130_fd_sc_hd__xnor2_1 U24390 ( .A(n18661), .B(n19012), .Y(n17438) );
  sky130_fd_sc_hd__o22ai_1 U24391 ( .A1(n17972), .A2(n17440), .B1(n17438), 
        .B2(n11159), .Y(n17437) );
  sky130_fd_sc_hd__xnor2_1 U24392 ( .A(n18479), .B(n21887), .Y(n17439) );
  sky130_fd_sc_hd__o22ai_1 U24393 ( .A1(n18224), .A2(n17428), .B1(n17439), 
        .B2(n18225), .Y(n17436) );
  sky130_fd_sc_hd__o22ai_1 U24394 ( .A1(n25219), .A2(n17429), .B1(n22198), 
        .B2(n18307), .Y(n17433) );
  sky130_fd_sc_hd__xnor2_1 U24395 ( .A(n17437), .B(n17436), .Y(n17574) );
  sky130_fd_sc_hd__xnor2_1 U24396 ( .A(n18654), .B(n22919), .Y(n17465) );
  sky130_fd_sc_hd__xnor2_1 U24397 ( .A(n18649), .B(n22919), .Y(n17533) );
  sky130_fd_sc_hd__xnor2_1 U24398 ( .A(n18708), .B(n19012), .Y(n17527) );
  sky130_fd_sc_hd__o22ai_1 U24399 ( .A1(n17972), .A2(n17438), .B1(n17527), 
        .B2(n11159), .Y(n17534) );
  sky130_fd_sc_hd__xnor2_1 U24400 ( .A(n18466), .B(n21887), .Y(n17530) );
  sky130_fd_sc_hd__o22ai_1 U24401 ( .A1(n18224), .A2(n17439), .B1(n17530), 
        .B2(n18225), .Y(n17594) );
  sky130_fd_sc_hd__xnor2_1 U24402 ( .A(n18687), .B(n24132), .Y(n17447) );
  sky130_fd_sc_hd__xnor2_1 U24403 ( .A(n18721), .B(n24132), .Y(n17588) );
  sky130_fd_sc_hd__o22ai_1 U24404 ( .A1(n17805), .A2(n17447), .B1(n17588), 
        .B2(n17802), .Y(n17593) );
  sky130_fd_sc_hd__inv_2 U24405 ( .A(j202_soc_core_j22_cpu_ml_bufa[0]), .Y(
        n17812) );
  sky130_fd_sc_hd__buf_6 U24406 ( .A(j202_soc_core_j22_cpu_ml_bufa[1]), .X(
        n22730) );
  sky130_fd_sc_hd__xnor2_1 U24407 ( .A(n22052), .B(n22730), .Y(n17445) );
  sky130_fd_sc_hd__xnor2_1 U24408 ( .A(n18651), .B(n22730), .Y(n17531) );
  sky130_fd_sc_hd__nand2_2 U24409 ( .A(n11749), .B(n17812), .Y(n17801) );
  sky130_fd_sc_hd__o22ai_1 U24410 ( .A1(n17812), .A2(n17445), .B1(n17531), 
        .B2(n17801), .Y(n17592) );
  sky130_fd_sc_hd__o22ai_1 U24411 ( .A1(n17972), .A2(n17441), .B1(n17440), 
        .B2(n11159), .Y(n17453) );
  sky130_fd_sc_hd__xnor2_1 U24412 ( .A(n17454), .B(n17453), .Y(n17457) );
  sky130_fd_sc_hd__xnor2_1 U24413 ( .A(n18426), .B(n18883), .Y(n17542) );
  sky130_fd_sc_hd__o22ai_1 U24414 ( .A1(n18344), .A2(n17442), .B1(n17542), 
        .B2(n17402), .Y(n17551) );
  sky130_fd_sc_hd__xnor2_1 U24415 ( .A(n18300), .B(n18226), .Y(n17443) );
  sky130_fd_sc_hd__o22ai_1 U24416 ( .A1(n18370), .A2(n17444), .B1(n17443), 
        .B2(n17392), .Y(n17550) );
  sky130_fd_sc_hd__a21o_1 U24417 ( .A1(n17801), .A2(n17812), .B1(n17445), .X(
        n17549) );
  sky130_fd_sc_hd__xnor2_1 U24418 ( .A(n18667), .B(n18147), .Y(n17540) );
  sky130_fd_sc_hd__o22ai_1 U24419 ( .A1(n18151), .A2(n17446), .B1(n17540), 
        .B2(n18148), .Y(n17554) );
  sky130_fd_sc_hd__o22ai_1 U24420 ( .A1(n17805), .A2(n17448), .B1(n17447), 
        .B2(n17802), .Y(n17553) );
  sky130_fd_sc_hd__nand2b_1 U24421 ( .A_N(n18353), .B(n18300), .Y(n17449) );
  sky130_fd_sc_hd__o22ai_1 U24422 ( .A1(n18370), .A2(n17449), .B1(n22807), 
        .B2(n17392), .Y(n17552) );
  sky130_fd_sc_hd__o21ai_1 U24423 ( .A1(n17559), .A2(n17560), .B1(n17561), .Y(
        n17451) );
  sky130_fd_sc_hd__nand2_1 U24424 ( .A(n17559), .B(n17560), .Y(n17450) );
  sky130_fd_sc_hd__nand2_1 U24425 ( .A(n17451), .B(n17450), .Y(n17564) );
  sky130_fd_sc_hd__o22ai_1 U24426 ( .A1(n17786), .A2(n17472), .B1(n17452), 
        .B2(n17771), .Y(n17476) );
  sky130_fd_sc_hd__o22ai_1 U24427 ( .A1(n25219), .A2(n17455), .B1(n22953), 
        .B2(n18307), .Y(n17474) );
  sky130_fd_sc_hd__fah_1 U24428 ( .A(n17460), .B(n17459), .CI(n17458), .COUT(
        n17431), .SUM(n17545) );
  sky130_fd_sc_hd__fah_1 U24429 ( .A(n17463), .B(n17462), .CI(n17461), .COUT(
        n17432), .SUM(n17544) );
  sky130_fd_sc_hd__o22ai_1 U24430 ( .A1(n17786), .A2(n17464), .B1(n17538), 
        .B2(n17771), .Y(n17526) );
  sky130_fd_sc_hd__o22ai_1 U24431 ( .A1(n18067), .A2(n17466), .B1(n17465), 
        .B2(n10971), .Y(n17525) );
  sky130_fd_sc_hd__o22ai_1 U24432 ( .A1(n25219), .A2(n17467), .B1(n22806), 
        .B2(n18307), .Y(n17524) );
  sky130_fd_sc_hd__xnor2_1 U24433 ( .A(n18654), .B(n21887), .Y(n17511) );
  sky130_fd_sc_hd__o22ai_1 U24434 ( .A1(n18224), .A2(n17511), .B1(n17468), 
        .B2(n18225), .Y(n17503) );
  sky130_fd_sc_hd__xnor2_1 U24435 ( .A(n18479), .B(n18300), .Y(n17510) );
  sky130_fd_sc_hd__o22ai_1 U24436 ( .A1(n18370), .A2(n17510), .B1(n17469), 
        .B2(n17392), .Y(n17502) );
  sky130_fd_sc_hd__xnor2_1 U24437 ( .A(n18661), .B(n18147), .Y(n17509) );
  sky130_fd_sc_hd__o22ai_1 U24438 ( .A1(n18151), .A2(n17509), .B1(n17470), 
        .B2(n18148), .Y(n17501) );
  sky130_fd_sc_hd__xnor2_1 U24439 ( .A(n18426), .B(n22951), .Y(n17513) );
  sky130_fd_sc_hd__o22ai_1 U24440 ( .A1(n12367), .A2(n17513), .B1(n17471), 
        .B2(n18470), .Y(n17500) );
  sky130_fd_sc_hd__o22ai_1 U24441 ( .A1(n12133), .A2(n17504), .B1(n17472), 
        .B2(n17771), .Y(n17499) );
  sky130_fd_sc_hd__xnor2_1 U24442 ( .A(n18667), .B(n18883), .Y(n17508) );
  sky130_fd_sc_hd__o22ai_1 U24443 ( .A1(n18344), .A2(n17508), .B1(n17473), 
        .B2(n17402), .Y(n17498) );
  sky130_fd_sc_hd__fah_1 U24444 ( .A(n17476), .B(n17475), .CI(n17474), .COUT(
        n17481), .SUM(n17523) );
  sky130_fd_sc_hd__fah_1 U24445 ( .A(n17479), .B(n17478), .CI(n17477), .COUT(
        n17496), .SUM(n17559) );
  sky130_fd_sc_hd__xnor2_1 U24446 ( .A(n17497), .B(n17496), .Y(n17480) );
  sky130_fd_sc_hd__xnor2_1 U24447 ( .A(n17495), .B(n17480), .Y(n17563) );
  sky130_fd_sc_hd__fah_1 U24448 ( .A(n17483), .B(n17482), .CI(n17481), .COUT(
        n17957), .SUM(n17497) );
  sky130_fd_sc_hd__xnor2_1 U24449 ( .A(n18721), .B(n22919), .Y(n17944) );
  sky130_fd_sc_hd__o22ai_1 U24450 ( .A1(n18067), .A2(n17944), .B1(n17487), 
        .B2(n10971), .Y(n17949) );
  sky130_fd_sc_hd__or2_1 U24451 ( .A(n17489), .B(n17488), .X(n17948) );
  sky130_fd_sc_hd__o22ai_1 U24452 ( .A1(n25219), .A2(n17490), .B1(n22113), 
        .B2(n18307), .Y(n17947) );
  sky130_fd_sc_hd__xnor2_1 U24453 ( .A(n17959), .B(n17958), .Y(n17491) );
  sky130_fd_sc_hd__xnor2_1 U24454 ( .A(n17957), .B(n17491), .Y(n18091) );
  sky130_fd_sc_hd__nand2_1 U24455 ( .A(n17493), .B(n17492), .Y(n17494) );
  sky130_fd_sc_hd__xnor2_1 U24456 ( .A(n18651), .B(n19012), .Y(n17940) );
  sky130_fd_sc_hd__o22ai_1 U24457 ( .A1(n17972), .A2(n17940), .B1(n17505), 
        .B2(n11159), .Y(n17931) );
  sky130_fd_sc_hd__buf_6 U24458 ( .A(n12138), .X(n22112) );
  sky130_fd_sc_hd__xnor2_1 U24459 ( .A(n18367), .B(n22112), .Y(n17945) );
  sky130_fd_sc_hd__xnor2_1 U24460 ( .A(n22112), .B(n18226), .Y(n17507) );
  sky130_fd_sc_hd__o22ai_1 U24461 ( .A1(n12140), .A2(n17945), .B1(n17507), 
        .B2(n18424), .Y(n17930) );
  sky130_fd_sc_hd__xnor2_1 U24462 ( .A(n18649), .B(n18883), .Y(n17941) );
  sky130_fd_sc_hd__o22ai_1 U24463 ( .A1(n18344), .A2(n17941), .B1(n17508), 
        .B2(n17402), .Y(n17935) );
  sky130_fd_sc_hd__xnor2_1 U24464 ( .A(n18673), .B(n18147), .Y(n17981) );
  sky130_fd_sc_hd__o22ai_1 U24465 ( .A1(n18151), .A2(n17981), .B1(n17509), 
        .B2(n18148), .Y(n17934) );
  sky130_fd_sc_hd__xnor2_1 U24466 ( .A(n18511), .B(n18300), .Y(n17943) );
  sky130_fd_sc_hd__o22ai_1 U24467 ( .A1(n18370), .A2(n17943), .B1(n17510), 
        .B2(n17392), .Y(n17933) );
  sky130_fd_sc_hd__xnor2_1 U24468 ( .A(n18708), .B(n17400), .Y(n17946) );
  sky130_fd_sc_hd__o22ai_1 U24469 ( .A1(n18224), .A2(n17946), .B1(n17511), 
        .B2(n18225), .Y(n17938) );
  sky130_fd_sc_hd__o22ai_1 U24470 ( .A1(n18514), .A2(n17512), .B1(n22114), 
        .B2(n18515), .Y(n17937) );
  sky130_fd_sc_hd__xnor2_1 U24471 ( .A(n18466), .B(n22951), .Y(n17942) );
  sky130_fd_sc_hd__o22ai_1 U24472 ( .A1(n12367), .A2(n17942), .B1(n17513), 
        .B2(n18470), .Y(n17936) );
  sky130_fd_sc_hd__fah_1 U24473 ( .A(n17516), .B(n17515), .CI(n17514), .COUT(
        n17951), .SUM(n17519) );
  sky130_fd_sc_hd__xnor2_1 U24474 ( .A(n18083), .B(n18084), .Y(n17520) );
  sky130_fd_sc_hd__fah_1 U24475 ( .A(n17519), .B(n17518), .CI(n17517), .COUT(
        n18082), .SUM(n17565) );
  sky130_fd_sc_hd__xnor2_1 U24476 ( .A(n17520), .B(n18082), .Y(n18090) );
  sky130_fd_sc_hd__fah_1 U24477 ( .A(n17526), .B(n17525), .CI(n17524), .COUT(
        n17543), .SUM(n17604) );
  sky130_fd_sc_hd__xnor2_1 U24478 ( .A(n18654), .B(n19012), .Y(n17578) );
  sky130_fd_sc_hd__o22ai_1 U24479 ( .A1(n17972), .A2(n17527), .B1(n17578), 
        .B2(n11159), .Y(n17591) );
  sky130_fd_sc_hd__nand2b_1 U24480 ( .A_N(n18353), .B(n18883), .Y(n17528) );
  sky130_fd_sc_hd__o22ai_1 U24481 ( .A1(n18344), .A2(n17528), .B1(n25264), 
        .B2(n17402), .Y(n17590) );
  sky130_fd_sc_hd__o22ai_1 U24482 ( .A1(n25219), .A2(n17529), .B1(n22530), 
        .B2(n18307), .Y(n17606) );
  sky130_fd_sc_hd__xnor2_1 U24483 ( .A(n18426), .B(n21887), .Y(n17580) );
  sky130_fd_sc_hd__o22ai_1 U24484 ( .A1(n18224), .A2(n17530), .B1(n17580), 
        .B2(n18225), .Y(n17613) );
  sky130_fd_sc_hd__xnor2_1 U24485 ( .A(n18687), .B(n22730), .Y(n17583) );
  sky130_fd_sc_hd__o22ai_1 U24486 ( .A1(n17812), .A2(n17531), .B1(n17583), 
        .B2(n17801), .Y(n17612) );
  sky130_fd_sc_hd__xnor2_1 U24487 ( .A(n18367), .B(n18883), .Y(n17541) );
  sky130_fd_sc_hd__xnor2_1 U24488 ( .A(n18883), .B(n18226), .Y(n17532) );
  sky130_fd_sc_hd__o22ai_1 U24489 ( .A1(n18344), .A2(n17541), .B1(n17532), 
        .B2(n17402), .Y(n17611) );
  sky130_fd_sc_hd__xnor2_1 U24490 ( .A(n18667), .B(n22919), .Y(n17582) );
  sky130_fd_sc_hd__o22ai_1 U24491 ( .A1(n18067), .A2(n17533), .B1(n17582), 
        .B2(n18068), .Y(n17615) );
  sky130_fd_sc_hd__xnor2_1 U24492 ( .A(n18511), .B(n18147), .Y(n17539) );
  sky130_fd_sc_hd__xnor2_1 U24493 ( .A(n18479), .B(n18147), .Y(n17581) );
  sky130_fd_sc_hd__o22ai_1 U24494 ( .A1(n18151), .A2(n17539), .B1(n17581), 
        .B2(n18148), .Y(n17614) );
  sky130_fd_sc_hd__fah_1 U24495 ( .A(n17536), .B(n17535), .CI(n17534), .COUT(
        n17573), .SUM(n17609) );
  sky130_fd_sc_hd__o22ai_1 U24496 ( .A1(n17786), .A2(n17538), .B1(n17537), 
        .B2(n17771), .Y(n17548) );
  sky130_fd_sc_hd__o22ai_1 U24497 ( .A1(n18151), .A2(n17540), .B1(n17539), 
        .B2(n18148), .Y(n17547) );
  sky130_fd_sc_hd__o22ai_1 U24498 ( .A1(n18344), .A2(n17542), .B1(n17541), 
        .B2(n17402), .Y(n17546) );
  sky130_fd_sc_hd__fah_1 U24499 ( .A(n17545), .B(n17544), .CI(n17543), .COUT(
        n17521), .SUM(n17598) );
  sky130_fd_sc_hd__fah_1 U24500 ( .A(n17554), .B(n17553), .CI(n17552), .COUT(
        n17456), .SUM(n17575) );
  sky130_fd_sc_hd__nand2b_1 U24501 ( .A_N(n17598), .B(n17555), .Y(n17556) );
  sky130_fd_sc_hd__nand2_1 U24502 ( .A(n17600), .B(n17556), .Y(n17558) );
  sky130_fd_sc_hd__nand2_1 U24503 ( .A(n17598), .B(n17599), .Y(n17557) );
  sky130_fd_sc_hd__nand2_1 U24504 ( .A(n17558), .B(n17557), .Y(n17567) );
  sky130_fd_sc_hd__xnor2_1 U24505 ( .A(n17560), .B(n17559), .Y(n17562) );
  sky130_fd_sc_hd__xnor2_1 U24506 ( .A(n17562), .B(n17561), .Y(n17566) );
  sky130_fd_sc_hd__fah_1 U24507 ( .A(n17565), .B(n17564), .CI(n17563), .COUT(
        n17928), .SUM(n17927) );
  sky130_fd_sc_hd__fah_1 U24508 ( .A(n17568), .B(n17567), .CI(n17566), .COUT(
        n17926), .SUM(n17925) );
  sky130_fd_sc_hd__fah_1 U24509 ( .A(n17571), .B(n17570), .CI(n17569), .COUT(
        n17561), .SUM(n17623) );
  sky130_fd_sc_hd__fah_1 U24510 ( .A(n17577), .B(n17576), .CI(n17575), .COUT(
        n17599), .SUM(n17620) );
  sky130_fd_sc_hd__xnor2_1 U24511 ( .A(n18649), .B(n19012), .Y(n17584) );
  sky130_fd_sc_hd__o22ai_1 U24512 ( .A1(n17972), .A2(n17578), .B1(n17584), 
        .B2(n11159), .Y(n17625) );
  sky130_fd_sc_hd__o22ai_1 U24513 ( .A1(n17786), .A2(n17579), .B1(n17657), 
        .B2(n17771), .Y(n17624) );
  sky130_fd_sc_hd__xnor2_1 U24514 ( .A(n18367), .B(n21887), .Y(n17653) );
  sky130_fd_sc_hd__o22ai_1 U24515 ( .A1(n18224), .A2(n17580), .B1(n17653), 
        .B2(n18225), .Y(n17629) );
  sky130_fd_sc_hd__xnor2_1 U24516 ( .A(n18466), .B(n18147), .Y(n17659) );
  sky130_fd_sc_hd__o22ai_1 U24517 ( .A1(n18151), .A2(n17581), .B1(n17659), 
        .B2(n18148), .Y(n17628) );
  sky130_fd_sc_hd__xnor2_1 U24518 ( .A(n18511), .B(n22919), .Y(n17649) );
  sky130_fd_sc_hd__o22ai_1 U24519 ( .A1(n18067), .A2(n17582), .B1(n17649), 
        .B2(n10971), .Y(n17627) );
  sky130_fd_sc_hd__xnor2_1 U24520 ( .A(n18721), .B(n22730), .Y(n17651) );
  sky130_fd_sc_hd__o22ai_1 U24521 ( .A1(n17812), .A2(n17583), .B1(n17651), 
        .B2(n17801), .Y(n17632) );
  sky130_fd_sc_hd__xnor2_1 U24522 ( .A(n18685), .B(n24132), .Y(n17587) );
  sky130_fd_sc_hd__xnor2_1 U24523 ( .A(n18673), .B(n24132), .Y(n17655) );
  sky130_fd_sc_hd__o22ai_1 U24524 ( .A1(n17805), .A2(n17587), .B1(n17655), 
        .B2(n17802), .Y(n17631) );
  sky130_fd_sc_hd__xnor2_1 U24525 ( .A(n18667), .B(n19012), .Y(n17637) );
  sky130_fd_sc_hd__o22ai_1 U24526 ( .A1(n17972), .A2(n17584), .B1(n17637), 
        .B2(n11159), .Y(n17634) );
  sky130_fd_sc_hd__o22ai_1 U24527 ( .A1(n17805), .A2(n17588), .B1(n17587), 
        .B2(n17802), .Y(n17618) );
  sky130_fd_sc_hd__inv_2 U24528 ( .A(n26977), .Y(n18882) );
  sky130_fd_sc_hd__ha_1 U24529 ( .A(n17591), .B(n17590), .COUT(n17607), .SUM(
        n17616) );
  sky130_fd_sc_hd__nand2_1 U24530 ( .A(n17902), .B(n17903), .Y(n17596) );
  sky130_fd_sc_hd__nand2_1 U24531 ( .A(n17597), .B(n17596), .Y(n17619) );
  sky130_fd_sc_hd__xnor2_1 U24532 ( .A(n17599), .B(n17598), .Y(n17601) );
  sky130_fd_sc_hd__xnor2_1 U24533 ( .A(n17601), .B(n17600), .Y(n17621) );
  sky130_fd_sc_hd__fah_1 U24534 ( .A(n17607), .B(n17606), .CI(n17605), .COUT(
        n17603), .SUM(n17909) );
  sky130_fd_sc_hd__fah_1 U24535 ( .A(n17610), .B(n17609), .CI(n17608), .COUT(
        n17602), .SUM(n17908) );
  sky130_fd_sc_hd__fah_1 U24536 ( .A(n17613), .B(n17612), .CI(n17611), .COUT(
        n17605), .SUM(n17671) );
  sky130_fd_sc_hd__fah_1 U24537 ( .A(n17618), .B(n17617), .CI(n17616), .COUT(
        n17902), .SUM(n17669) );
  sky130_fd_sc_hd__nor2_1 U24538 ( .A(n17922), .B(n17923), .Y(n19199) );
  sky130_fd_sc_hd__fah_1 U24539 ( .A(n17626), .B(n17625), .CI(n17624), .COUT(
        n17677), .SUM(n17680) );
  sky130_fd_sc_hd__fah_1 U24540 ( .A(n17632), .B(n17631), .CI(n17630), .COUT(
        n17675), .SUM(n17678) );
  sky130_fd_sc_hd__xnor2_1 U24541 ( .A(n18479), .B(n22919), .Y(n17648) );
  sky130_fd_sc_hd__xnor2_1 U24542 ( .A(n18466), .B(n22919), .Y(n17687) );
  sky130_fd_sc_hd__o22ai_1 U24543 ( .A1(n18067), .A2(n17648), .B1(n17687), 
        .B2(n10971), .Y(n17692) );
  sky130_fd_sc_hd__xnor2_1 U24544 ( .A(n18673), .B(n22730), .Y(n17635) );
  sky130_fd_sc_hd__xnor2_1 U24545 ( .A(n18661), .B(n22730), .Y(n17697) );
  sky130_fd_sc_hd__o22ai_1 U24546 ( .A1(n17812), .A2(n17635), .B1(n17697), 
        .B2(n17801), .Y(n17694) );
  sky130_fd_sc_hd__xnor2_1 U24547 ( .A(n18511), .B(n19012), .Y(n17636) );
  sky130_fd_sc_hd__xnor2_1 U24548 ( .A(n18479), .B(n19012), .Y(n17695) );
  sky130_fd_sc_hd__o22ai_1 U24549 ( .A1(n17972), .A2(n17636), .B1(n17695), 
        .B2(n11159), .Y(n17693) );
  sky130_fd_sc_hd__a22o_1 U24550 ( .A1(n23257), .A2(
        j202_soc_core_j22_cpu_ml_macl[28]), .B1(
        j202_soc_core_j22_cpu_ml_macl[12]), .B2(n18183), .X(n17690) );
  sky130_fd_sc_hd__a22o_1 U24551 ( .A1(j202_soc_core_j22_cpu_ml_macl[29]), 
        .A2(n23257), .B1(n18183), .B2(j202_soc_core_j22_cpu_ml_macl[13]), .X(
        n17647) );
  sky130_fd_sc_hd__ha_1 U24552 ( .A(n17634), .B(n17633), .COUT(n17630), .SUM(
        n17646) );
  sky130_fd_sc_hd__nor2b_1 U24553 ( .B_N(n18353), .A(n18224), .Y(n17641) );
  sky130_fd_sc_hd__xnor2_1 U24554 ( .A(n18685), .B(n22730), .Y(n17650) );
  sky130_fd_sc_hd__o22ai_1 U24555 ( .A1(n17812), .A2(n17650), .B1(n17635), 
        .B2(n17801), .Y(n17640) );
  sky130_fd_sc_hd__o22ai_1 U24556 ( .A1(n17972), .A2(n17637), .B1(n17636), 
        .B2(n11159), .Y(n17639) );
  sky130_fd_sc_hd__xnor2_1 U24557 ( .A(n18708), .B(n24132), .Y(n17642) );
  sky130_fd_sc_hd__xnor2_1 U24558 ( .A(n18654), .B(n24132), .Y(n17699) );
  sky130_fd_sc_hd__o22ai_1 U24559 ( .A1(n17805), .A2(n17642), .B1(n17699), 
        .B2(n17802), .Y(n17741) );
  sky130_fd_sc_hd__o22ai_1 U24560 ( .A1(n17786), .A2(n17644), .B1(n17698), 
        .B2(n17771), .Y(n17740) );
  sky130_fd_sc_hd__xnor2_1 U24561 ( .A(n18367), .B(n18147), .Y(n17643) );
  sky130_fd_sc_hd__xnor2_1 U24562 ( .A(n18147), .B(n18226), .Y(n17638) );
  sky130_fd_sc_hd__o22ai_1 U24563 ( .A1(n18151), .A2(n17643), .B1(n17638), 
        .B2(n18148), .Y(n17739) );
  sky130_fd_sc_hd__xnor2_1 U24564 ( .A(n18661), .B(n24132), .Y(n17654) );
  sky130_fd_sc_hd__o22ai_1 U24565 ( .A1(n17805), .A2(n17654), .B1(n17642), 
        .B2(n17802), .Y(n17662) );
  sky130_fd_sc_hd__xnor2_1 U24566 ( .A(n18426), .B(n18147), .Y(n17658) );
  sky130_fd_sc_hd__o22ai_1 U24567 ( .A1(n18151), .A2(n17658), .B1(n17643), 
        .B2(n18148), .Y(n17661) );
  sky130_fd_sc_hd__o22ai_1 U24568 ( .A1(n17786), .A2(n17656), .B1(n17644), 
        .B2(n17771), .Y(n17660) );
  sky130_fd_sc_hd__o22ai_1 U24569 ( .A1(n18882), .A2(n22628), .B1(n23949), 
        .B2(n18307), .Y(n17683) );
  sky130_fd_sc_hd__o22ai_1 U24570 ( .A1(n18067), .A2(n17649), .B1(n17648), 
        .B2(n18068), .Y(n17668) );
  sky130_fd_sc_hd__o22ai_1 U24571 ( .A1(n17812), .A2(n17651), .B1(n17650), 
        .B2(n17801), .Y(n17667) );
  sky130_fd_sc_hd__xnor2_1 U24572 ( .A(n21887), .B(n18226), .Y(n17652) );
  sky130_fd_sc_hd__o22ai_1 U24573 ( .A1(n18224), .A2(n17653), .B1(n17652), 
        .B2(n18225), .Y(n17666) );
  sky130_fd_sc_hd__o22ai_1 U24574 ( .A1(n17805), .A2(n17655), .B1(n17654), 
        .B2(n17802), .Y(n17665) );
  sky130_fd_sc_hd__o22ai_1 U24575 ( .A1(n17786), .A2(n17657), .B1(n17656), 
        .B2(n17771), .Y(n17664) );
  sky130_fd_sc_hd__o22ai_1 U24576 ( .A1(n18151), .A2(n17659), .B1(n17658), 
        .B2(n18148), .Y(n17663) );
  sky130_fd_sc_hd__fah_1 U24577 ( .A(n17671), .B(n17670), .CI(n17669), .COUT(
        n17907), .SUM(n17900) );
  sky130_fd_sc_hd__fah_1 U24578 ( .A(n17674), .B(n17673), .CI(n17672), .COUT(
        n17899), .SUM(n17703) );
  sky130_fd_sc_hd__fa_1 U24580 ( .A(n17684), .B(n17686), .CIN(n17685), .COUT(
        n17672), .SUM(n17887) );
  sky130_fd_sc_hd__xnor2_1 U24581 ( .A(n18426), .B(n22919), .Y(n17696) );
  sky130_fd_sc_hd__o22ai_1 U24582 ( .A1(n18067), .A2(n17687), .B1(n17696), 
        .B2(n10971), .Y(n17744) );
  sky130_fd_sc_hd__nand2b_1 U24583 ( .A_N(n18353), .B(n18147), .Y(n17689) );
  sky130_fd_sc_hd__o22ai_1 U24584 ( .A1(n18151), .A2(n17689), .B1(n17688), 
        .B2(n18148), .Y(n17743) );
  sky130_fd_sc_hd__o22ai_1 U24585 ( .A1(n18882), .A2(n18106), .B1(n23972), 
        .B2(n18307), .Y(n17742) );
  sky130_fd_sc_hd__fah_1 U24586 ( .A(n17692), .B(n17691), .CI(n17690), .COUT(
        n17702), .SUM(n17880) );
  sky130_fd_sc_hd__ha_1 U24587 ( .A(n17694), .B(n17693), .COUT(n17691), .SUM(
        n17735) );
  sky130_fd_sc_hd__xnor2_1 U24588 ( .A(n18466), .B(n19012), .Y(n17708) );
  sky130_fd_sc_hd__xnor2_1 U24589 ( .A(n18367), .B(n22919), .Y(n17713) );
  sky130_fd_sc_hd__o22ai_1 U24590 ( .A1(n18067), .A2(n17696), .B1(n17713), 
        .B2(n10971), .Y(n17723) );
  sky130_fd_sc_hd__xnor2_1 U24591 ( .A(n18708), .B(n22730), .Y(n17707) );
  sky130_fd_sc_hd__o22ai_1 U24592 ( .A1(n17812), .A2(n17697), .B1(n17707), 
        .B2(n17801), .Y(n17728) );
  sky130_fd_sc_hd__o22ai_1 U24593 ( .A1(n17786), .A2(n17698), .B1(n17709), 
        .B2(n17771), .Y(n17727) );
  sky130_fd_sc_hd__xnor2_1 U24594 ( .A(n18649), .B(n24132), .Y(n17730) );
  sky130_fd_sc_hd__o22ai_1 U24595 ( .A1(n17805), .A2(n17699), .B1(n17730), 
        .B2(n17802), .Y(n17726) );
  sky130_fd_sc_hd__fah_1 U24596 ( .A(n17705), .B(n17704), .CI(n17703), .COUT(
        n17895), .SUM(n17894) );
  sky130_fd_sc_hd__nor2_1 U24597 ( .A(n17893), .B(n17894), .Y(n17706) );
  sky130_fd_sc_hd__xnor2_1 U24598 ( .A(n18654), .B(n22730), .Y(n17715) );
  sky130_fd_sc_hd__o22ai_1 U24599 ( .A1(n17812), .A2(n17707), .B1(n17715), 
        .B2(n17801), .Y(n17732) );
  sky130_fd_sc_hd__xnor2_1 U24600 ( .A(n18426), .B(n19012), .Y(n17714) );
  sky130_fd_sc_hd__o22ai_1 U24601 ( .A1(n17972), .A2(n17708), .B1(n17714), 
        .B2(n11159), .Y(n17731) );
  sky130_fd_sc_hd__o22ai_1 U24602 ( .A1(n18882), .A2(n22407), .B1(n19239), 
        .B2(n18307), .Y(n17746) );
  sky130_fd_sc_hd__o22ai_1 U24603 ( .A1(n17786), .A2(n17709), .B1(n17716), 
        .B2(n17771), .Y(n17722) );
  sky130_fd_sc_hd__nand2b_1 U24604 ( .A_N(n18353), .B(n22919), .Y(n17711) );
  sky130_fd_sc_hd__o22ai_1 U24606 ( .A1(n18067), .A2(n17711), .B1(n12569), 
        .B2(n10971), .Y(n17721) );
  sky130_fd_sc_hd__xnor2_1 U24607 ( .A(n22919), .B(n18226), .Y(n17712) );
  sky130_fd_sc_hd__o22ai_1 U24608 ( .A1(n18067), .A2(n17713), .B1(n17712), 
        .B2(n10971), .Y(n17720) );
  sky130_fd_sc_hd__nor2b_1 U24609 ( .B_N(n18353), .A(n18067), .Y(n17757) );
  sky130_fd_sc_hd__xnor2_1 U24610 ( .A(n18367), .B(n19012), .Y(n17754) );
  sky130_fd_sc_hd__o22ai_1 U24611 ( .A1(n17972), .A2(n17714), .B1(n17754), 
        .B2(n11159), .Y(n17756) );
  sky130_fd_sc_hd__xnor2_1 U24612 ( .A(n18649), .B(n22730), .Y(n17717) );
  sky130_fd_sc_hd__o22ai_1 U24613 ( .A1(n17812), .A2(n17715), .B1(n17717), 
        .B2(n17801), .Y(n17755) );
  sky130_fd_sc_hd__xnor2_1 U24614 ( .A(n18667), .B(n24132), .Y(n17729) );
  sky130_fd_sc_hd__xnor2_1 U24615 ( .A(n18511), .B(n24132), .Y(n17752) );
  sky130_fd_sc_hd__o22ai_1 U24616 ( .A1(n17805), .A2(n17729), .B1(n17752), 
        .B2(n17802), .Y(n17847) );
  sky130_fd_sc_hd__o22ai_1 U24617 ( .A1(n17786), .A2(n17716), .B1(n17751), 
        .B2(n17771), .Y(n17846) );
  sky130_fd_sc_hd__xnor2_1 U24618 ( .A(n18667), .B(n22730), .Y(n17770) );
  sky130_fd_sc_hd__o22ai_1 U24619 ( .A1(n17812), .A2(n17717), .B1(n17770), 
        .B2(n17801), .Y(n17781) );
  sky130_fd_sc_hd__nand2b_1 U24620 ( .A_N(n18353), .B(n19012), .Y(n17719) );
  sky130_fd_sc_hd__fah_1 U24621 ( .A(n17725), .B(n17724), .CI(n17723), .COUT(
        n17734), .SUM(n17738) );
  sky130_fd_sc_hd__fah_1 U24622 ( .A(n17728), .B(n17727), .CI(n17726), .COUT(
        n17733), .SUM(n17737) );
  sky130_fd_sc_hd__o22ai_1 U24623 ( .A1(n17805), .A2(n17730), .B1(n17729), 
        .B2(n17802), .Y(n17750) );
  sky130_fd_sc_hd__ha_1 U24624 ( .A(n17732), .B(n17731), .COUT(n17747), .SUM(
        n17748) );
  sky130_fd_sc_hd__fah_1 U24625 ( .A(n17738), .B(n17737), .CI(n17736), .COUT(
        n17871), .SUM(n17761) );
  sky130_fd_sc_hd__fah_1 U24626 ( .A(n17744), .B(n17743), .CI(n17742), .COUT(
        n17881), .SUM(n17877) );
  sky130_fd_sc_hd__fah_1 U24627 ( .A(n17750), .B(n17749), .CI(n17748), .COUT(
        n17736), .SUM(n17859) );
  sky130_fd_sc_hd__a22o_1 U24628 ( .A1(j202_soc_core_j22_cpu_ml_macl[24]), 
        .A2(n26977), .B1(n18183), .B2(j202_soc_core_j22_cpu_ml_macl[8]), .X(
        n17853) );
  sky130_fd_sc_hd__o22ai_1 U24629 ( .A1(n17786), .A2(n17751), .B1(n17765), 
        .B2(n17771), .Y(n17777) );
  sky130_fd_sc_hd__xnor2_1 U24630 ( .A(n18479), .B(n24132), .Y(n17764) );
  sky130_fd_sc_hd__o22ai_1 U24631 ( .A1(n17805), .A2(n17752), .B1(n17764), 
        .B2(n17802), .Y(n17776) );
  sky130_fd_sc_hd__xnor2_1 U24632 ( .A(n19012), .B(n18226), .Y(n17753) );
  sky130_fd_sc_hd__o22ai_1 U24633 ( .A1(n17972), .A2(n17754), .B1(n17753), 
        .B2(n11159), .Y(n17775) );
  sky130_fd_sc_hd__fah_1 U24634 ( .A(n17763), .B(n17762), .CI(n17761), .COUT(
        n17866), .SUM(n17865) );
  sky130_fd_sc_hd__xnor2_1 U24635 ( .A(n18466), .B(n24132), .Y(n17766) );
  sky130_fd_sc_hd__o22ai_1 U24636 ( .A1(n17805), .A2(n17764), .B1(n17766), 
        .B2(n17802), .Y(n17783) );
  sky130_fd_sc_hd__o22ai_1 U24637 ( .A1(n17786), .A2(n17765), .B1(n17768), 
        .B2(n17771), .Y(n17782) );
  sky130_fd_sc_hd__xnor2_1 U24638 ( .A(n18426), .B(n24132), .Y(n17789) );
  sky130_fd_sc_hd__o22ai_1 U24639 ( .A1(n17805), .A2(n17766), .B1(n17802), 
        .B2(n17789), .Y(n17797) );
  sky130_fd_sc_hd__o22ai_1 U24640 ( .A1(n17786), .A2(n17768), .B1(n17767), 
        .B2(n17771), .Y(n17796) );
  sky130_fd_sc_hd__o22ai_1 U24641 ( .A1(n18882), .A2(n22113), .B1(n17769), 
        .B2(n18307), .Y(n17795) );
  sky130_fd_sc_hd__xnor2_1 U24642 ( .A(n18511), .B(n22730), .Y(n17774) );
  sky130_fd_sc_hd__o22ai_1 U24643 ( .A1(n17812), .A2(n17770), .B1(n17774), 
        .B2(n17801), .Y(n17780) );
  sky130_fd_sc_hd__o22ai_1 U24644 ( .A1(n17786), .A2(n29573), .B1(n17772), 
        .B2(n17771), .Y(n17791) );
  sky130_fd_sc_hd__xnor2_1 U24645 ( .A(n18479), .B(n22730), .Y(n17788) );
  sky130_fd_sc_hd__o22ai_1 U24646 ( .A1(n17812), .A2(n17774), .B1(n17788), 
        .B2(n17801), .Y(n17790) );
  sky130_fd_sc_hd__o22ai_1 U24647 ( .A1(n18882), .A2(n22337), .B1(n21537), 
        .B2(n18307), .Y(n17778) );
  sky130_fd_sc_hd__o22ai_1 U24648 ( .A1(n18882), .A2(n22030), .B1(n19008), 
        .B2(n18307), .Y(n17850) );
  sky130_fd_sc_hd__fah_1 U24649 ( .A(n17784), .B(n17783), .CI(n17782), .COUT(
        n17848), .SUM(n17838) );
  sky130_fd_sc_hd__nor2_1 U24650 ( .A(n18993), .B(n18992), .Y(n17842) );
  sky130_fd_sc_hd__nand2b_1 U24651 ( .A_N(n18353), .B(n24132), .Y(n17785) );
  sky130_fd_sc_hd__xnor2_1 U24652 ( .A(n18466), .B(n22730), .Y(n17787) );
  sky130_fd_sc_hd__xnor2_1 U24653 ( .A(n18426), .B(n22730), .Y(n17798) );
  sky130_fd_sc_hd__o22ai_1 U24654 ( .A1(n17812), .A2(n17787), .B1(n17798), 
        .B2(n17801), .Y(n17806) );
  sky130_fd_sc_hd__nor2b_1 U24655 ( .B_N(n18353), .A(n17786), .Y(n17794) );
  sky130_fd_sc_hd__o22ai_1 U24656 ( .A1(n17812), .A2(n17788), .B1(n17787), 
        .B2(n17801), .Y(n17793) );
  sky130_fd_sc_hd__xnor2_1 U24657 ( .A(n18367), .B(n24132), .Y(n17804) );
  sky130_fd_sc_hd__o22ai_1 U24658 ( .A1(n17805), .A2(n17789), .B1(n17804), 
        .B2(n17802), .Y(n17792) );
  sky130_fd_sc_hd__o22ai_1 U24659 ( .A1(n18882), .A2(n22141), .B1(n19428), 
        .B2(n18307), .Y(n17824) );
  sky130_fd_sc_hd__ha_1 U24660 ( .A(n17791), .B(n17790), .COUT(n17779), .SUM(
        n17835) );
  sky130_fd_sc_hd__fah_1 U24661 ( .A(n17794), .B(n17793), .CI(n17792), .COUT(
        n17834), .SUM(n17825) );
  sky130_fd_sc_hd__fah_1 U24662 ( .A(n17797), .B(n17796), .CI(n17795), .COUT(
        n17837), .SUM(n17833) );
  sky130_fd_sc_hd__nor2_1 U24663 ( .A(n17831), .B(n17832), .Y(n21821) );
  sky130_fd_sc_hd__nor2b_1 U24664 ( .B_N(n18353), .A(n17805), .Y(n17811) );
  sky130_fd_sc_hd__xnor2_1 U24665 ( .A(n18367), .B(n22730), .Y(n17799) );
  sky130_fd_sc_hd__o22ai_1 U24666 ( .A1(n17812), .A2(n17798), .B1(n17799), 
        .B2(n17801), .Y(n17810) );
  sky130_fd_sc_hd__o22ai_1 U24667 ( .A1(n17812), .A2(n17799), .B1(n18226), 
        .B2(n17801), .Y(n17814) );
  sky130_fd_sc_hd__nand2b_1 U24668 ( .A_N(n18353), .B(n22730), .Y(n17800) );
  sky130_fd_sc_hd__nand2_1 U24669 ( .A(n17801), .B(n17800), .Y(n17813) );
  sky130_fd_sc_hd__xnor2_1 U24670 ( .A(n24132), .B(n18226), .Y(n17803) );
  sky130_fd_sc_hd__o22ai_1 U24671 ( .A1(n17805), .A2(n17804), .B1(n17803), 
        .B2(n17802), .Y(n17823) );
  sky130_fd_sc_hd__ha_1 U24672 ( .A(n17806), .B(n17807), .COUT(n17826), .SUM(
        n17822) );
  sky130_fd_sc_hd__o22ai_1 U24673 ( .A1(n18882), .A2(n22953), .B1(n17808), 
        .B2(n18307), .Y(n17821) );
  sky130_fd_sc_hd__o22ai_1 U24674 ( .A1(n18882), .A2(n22198), .B1(n19186), 
        .B2(n18307), .Y(n19175) );
  sky130_fd_sc_hd__fah_1 U24675 ( .A(n17811), .B(n17810), .CI(n17809), .COUT(
        n17819), .SUM(n19174) );
  sky130_fd_sc_hd__nor2_1 U24676 ( .A(n19175), .B(n19174), .Y(n17818) );
  sky130_fd_sc_hd__a22o_1 U24677 ( .A1(n23257), .A2(
        j202_soc_core_j22_cpu_ml_macl[16]), .B1(
        j202_soc_core_j22_cpu_ml_macl[0]), .B2(n18183), .X(n21924) );
  sky130_fd_sc_hd__nor2b_1 U24678 ( .B_N(n18353), .A(n17812), .Y(n21925) );
  sky130_fd_sc_hd__nand2_1 U24679 ( .A(n21924), .B(n21925), .Y(n21926) );
  sky130_fd_sc_hd__nand2_1 U24680 ( .A(n17816), .B(n17815), .Y(n22719) );
  sky130_fd_sc_hd__nand2_1 U24681 ( .A(n19174), .B(n19175), .Y(n19176) );
  sky130_fd_sc_hd__nand2_1 U24682 ( .A(n17820), .B(n17819), .Y(n21386) );
  sky130_fd_sc_hd__fah_1 U24683 ( .A(n17823), .B(n17822), .CI(n17821), .COUT(
        n17828), .SUM(n17820) );
  sky130_fd_sc_hd__fah_1 U24684 ( .A(n17826), .B(n17825), .CI(n17824), .COUT(
        n17831), .SUM(n17829) );
  sky130_fd_sc_hd__nor2_1 U24685 ( .A(n17828), .B(n17829), .Y(n17827) );
  sky130_fd_sc_hd__nand2_1 U24686 ( .A(n17829), .B(n17828), .Y(n19424) );
  sky130_fd_sc_hd__nand2_1 U24687 ( .A(n17832), .B(n17831), .Y(n21822) );
  sky130_fd_sc_hd__fah_1 U24688 ( .A(n17835), .B(n17834), .CI(n17833), .COUT(
        n17839), .SUM(n17832) );
  sky130_fd_sc_hd__fah_1 U24689 ( .A(n17837), .B(n17838), .CI(n17836), .COUT(
        n18993), .SUM(n17840) );
  sky130_fd_sc_hd__nand2_1 U24690 ( .A(n17840), .B(n17839), .Y(n21515) );
  sky130_fd_sc_hd__nand2_1 U24691 ( .A(n18992), .B(n18993), .Y(n18994) );
  sky130_fd_sc_hd__fah_1 U24692 ( .A(n17845), .B(n17844), .CI(n17843), .COUT(
        n21969), .SUM(n18992) );
  sky130_fd_sc_hd__fah_1 U24693 ( .A(n17847), .B(n17846), .CI(n11041), .COUT(
        n17759), .SUM(n17856) );
  sky130_fd_sc_hd__fah_1 U24694 ( .A(n17850), .B(n17849), .CI(n17848), .COUT(
        n17855), .SUM(n17843) );
  sky130_fd_sc_hd__fah_1 U24695 ( .A(n17853), .B(n17852), .CI(n17851), .COUT(
        n17858), .SUM(n17854) );
  sky130_fd_sc_hd__nor2_1 U24696 ( .A(n21969), .B(n21968), .Y(n22847) );
  sky130_fd_sc_hd__fah_1 U24697 ( .A(n17856), .B(n17855), .CI(n17854), .COUT(
        n17860), .SUM(n21968) );
  sky130_fd_sc_hd__fah_1 U24698 ( .A(n17859), .B(n17858), .CI(n17857), .COUT(
        n17864), .SUM(n17861) );
  sky130_fd_sc_hd__nor2_1 U24699 ( .A(n22847), .B(n22843), .Y(n17863) );
  sky130_fd_sc_hd__nand2_1 U24700 ( .A(n21968), .B(n21969), .Y(n22845) );
  sky130_fd_sc_hd__nand2_1 U24701 ( .A(n17861), .B(n17860), .Y(n22844) );
  sky130_fd_sc_hd__o21ai_1 U24702 ( .A1(n22845), .A2(n22843), .B1(n22844), .Y(
        n17862) );
  sky130_fd_sc_hd__a21oi_2 U24703 ( .A1(n21967), .A2(n17863), .B1(n17862), .Y(
        n19241) );
  sky130_fd_sc_hd__fah_1 U24704 ( .A(n17872), .B(n17871), .CI(n17870), .COUT(
        n17888), .SUM(n17867) );
  sky130_fd_sc_hd__fah_1 U24705 ( .A(n17875), .B(n17874), .CI(n17873), .COUT(
        n17700), .SUM(n17884) );
  sky130_fd_sc_hd__fah_1 U24706 ( .A(n17878), .B(n17877), .CI(n17876), .COUT(
        n17883), .SUM(n17870) );
  sky130_fd_sc_hd__nor2_1 U24707 ( .A(n17888), .B(n17889), .Y(n21894) );
  sky130_fd_sc_hd__fah_1 U24708 ( .A(n17884), .B(n17883), .CI(n17882), .COUT(
        n17890), .SUM(n17889) );
  sky130_fd_sc_hd__fah_1 U24709 ( .A(n17887), .B(n17886), .CI(n17885), .COUT(
        n17893), .SUM(n17891) );
  sky130_fd_sc_hd__nor2_1 U24710 ( .A(n21894), .B(n21889), .Y(n17892) );
  sky130_fd_sc_hd__nand2_1 U24711 ( .A(n17889), .B(n17888), .Y(n21892) );
  sky130_fd_sc_hd__nand2_1 U24712 ( .A(n17891), .B(n17890), .Y(n21890) );
  sky130_fd_sc_hd__nand2_1 U24713 ( .A(n17894), .B(n17893), .Y(n21504) );
  sky130_fd_sc_hd__nand2_1 U24714 ( .A(n17896), .B(n17895), .Y(n18888) );
  sky130_fd_sc_hd__fah_1 U24715 ( .A(n17900), .B(n17899), .CI(n17898), .COUT(
        n17916), .SUM(n17896) );
  sky130_fd_sc_hd__xor3_1 U24716 ( .A(n17903), .B(n17902), .C(n17901), .X(
        n17912) );
  sky130_fd_sc_hd__fah_1 U24717 ( .A(n17909), .B(n17908), .CI(n17907), .COUT(
        n17914), .SUM(n17910) );
  sky130_fd_sc_hd__nor2_1 U24718 ( .A(n17916), .B(n17917), .Y(n22763) );
  sky130_fd_sc_hd__fah_1 U24719 ( .A(n17912), .B(n17911), .CI(n17910), .COUT(
        n17918), .SUM(n17917) );
  sky130_fd_sc_hd__fah_1 U24720 ( .A(n17915), .B(n17914), .CI(n17913), .COUT(
        n17922), .SUM(n17919) );
  sky130_fd_sc_hd__nand2_1 U24722 ( .A(n17917), .B(n17916), .Y(n22762) );
  sky130_fd_sc_hd__nand2_1 U24723 ( .A(n17919), .B(n17918), .Y(n22760) );
  sky130_fd_sc_hd__nand2_1 U24725 ( .A(n17923), .B(n17922), .Y(n21428) );
  sky130_fd_sc_hd__nand2_1 U24726 ( .A(n17925), .B(n17924), .Y(n21430) );
  sky130_fd_sc_hd__nand2_1 U24727 ( .A(n17927), .B(n17926), .Y(n21803) );
  sky130_fd_sc_hd__nand2_1 U24728 ( .A(n17929), .B(n17928), .Y(n21809) );
  sky130_fd_sc_hd__fah_1 U24729 ( .A(n17932), .B(n17931), .CI(n17930), .COUT(
        n17994), .SUM(n17986) );
  sky130_fd_sc_hd__fah_1 U24730 ( .A(n17938), .B(n17937), .CI(n17936), .COUT(
        n17992), .SUM(n17952) );
  sky130_fd_sc_hd__xnor2_1 U24731 ( .A(n18721), .B(n18147), .Y(n18021) );
  sky130_fd_sc_hd__xnor2_1 U24732 ( .A(n18685), .B(n18147), .Y(n17982) );
  sky130_fd_sc_hd__o22ai_1 U24733 ( .A1(n18151), .A2(n18021), .B1(n17982), 
        .B2(n18148), .Y(n18017) );
  sky130_fd_sc_hd__xnor2_1 U24734 ( .A(j202_soc_core_j22_cpu_ml_bufa[22]), .B(
        j202_soc_core_j22_cpu_ml_bufa[21]), .Y(n17939) );
  sky130_fd_sc_hd__nor2b_1 U24735 ( .B_N(n18353), .A(n18660), .Y(n17985) );
  sky130_fd_sc_hd__xnor2_1 U24736 ( .A(n22052), .B(n19012), .Y(n17971) );
  sky130_fd_sc_hd__o22ai_1 U24737 ( .A1(n17972), .A2(n17971), .B1(n17940), 
        .B2(n11159), .Y(n17984) );
  sky130_fd_sc_hd__o2bb2ai_1 U24738 ( .B1(n22030), .B2(n18307), .A1_N(n26862), 
        .A2_N(j202_soc_core_j22_cpu_ml_mach[7]), .Y(n18015) );
  sky130_fd_sc_hd__xnor2_1 U24739 ( .A(n18654), .B(n18883), .Y(n17968) );
  sky130_fd_sc_hd__o22ai_1 U24740 ( .A1(n18344), .A2(n17968), .B1(n17941), 
        .B2(n17402), .Y(n17967) );
  sky130_fd_sc_hd__xnor2_1 U24741 ( .A(n18479), .B(n22951), .Y(n17979) );
  sky130_fd_sc_hd__o22ai_1 U24742 ( .A1(n12367), .A2(n17979), .B1(n17942), 
        .B2(n18470), .Y(n17966) );
  sky130_fd_sc_hd__xnor2_1 U24743 ( .A(n18667), .B(n18300), .Y(n17980) );
  sky130_fd_sc_hd__o22ai_1 U24744 ( .A1(n18370), .A2(n17980), .B1(n17943), 
        .B2(n17392), .Y(n17965) );
  sky130_fd_sc_hd__xnor2_1 U24745 ( .A(n18687), .B(n22919), .Y(n17978) );
  sky130_fd_sc_hd__xnor2_1 U24746 ( .A(n18426), .B(n22112), .Y(n17974) );
  sky130_fd_sc_hd__o22ai_1 U24747 ( .A1(n18514), .A2(n17974), .B1(n17945), 
        .B2(n18515), .Y(n17963) );
  sky130_fd_sc_hd__xnor2_1 U24748 ( .A(n18661), .B(n21887), .Y(n17977) );
  sky130_fd_sc_hd__o22ai_1 U24749 ( .A1(n18224), .A2(n17977), .B1(n17946), 
        .B2(n18225), .Y(n17962) );
  sky130_fd_sc_hd__xnor2_1 U24750 ( .A(n17950), .B(n18025), .Y(n18077) );
  sky130_fd_sc_hd__fah_1 U24751 ( .A(n17953), .B(n17952), .CI(n17951), .COUT(
        n18089), .SUM(n18084) );
  sky130_fd_sc_hd__fah_1 U24752 ( .A(n17956), .B(n17955), .CI(n17954), .COUT(
        n18025), .SUM(n18088) );
  sky130_fd_sc_hd__o21ai_1 U24753 ( .A1(n17959), .A2(n17958), .B1(n17957), .Y(
        n17961) );
  sky130_fd_sc_hd__nand2_1 U24754 ( .A(n17959), .B(n17958), .Y(n17960) );
  sky130_fd_sc_hd__nand2_1 U24755 ( .A(n17961), .B(n17960), .Y(n18087) );
  sky130_fd_sc_hd__fah_1 U24756 ( .A(n17964), .B(n17963), .CI(n17962), .COUT(
        n18001), .SUM(n17955) );
  sky130_fd_sc_hd__xnor2_1 U24757 ( .A(n18708), .B(n18883), .Y(n18023) );
  sky130_fd_sc_hd__o22ai_1 U24758 ( .A1(n18344), .A2(n18023), .B1(n17968), 
        .B2(n17402), .Y(n18003) );
  sky130_fd_sc_hd__xnor2_1 U24759 ( .A(n18367), .B(n22029), .Y(n18019) );
  sky130_fd_sc_hd__xnor2_1 U24760 ( .A(n22029), .B(n18226), .Y(n17970) );
  sky130_fd_sc_hd__xor2_1 U24761 ( .A(j202_soc_core_j22_cpu_ml_bufa[23]), .B(
        n12725), .X(n17969) );
  sky130_fd_sc_hd__a21o_1 U24762 ( .A1(n11159), .A2(n17972), .B1(n17971), .X(
        n18002) );
  sky130_fd_sc_hd__xnor2_1 U24763 ( .A(n18466), .B(n22112), .Y(n18020) );
  sky130_fd_sc_hd__o22ai_1 U24764 ( .A1(n18514), .A2(n18020), .B1(n17974), 
        .B2(n18515), .Y(n18006) );
  sky130_fd_sc_hd__nand2b_1 U24765 ( .A_N(n18353), .B(n22029), .Y(n17976) );
  sky130_fd_sc_hd__xnor2_1 U24766 ( .A(n18673), .B(n21887), .Y(n17998) );
  sky130_fd_sc_hd__o22ai_1 U24767 ( .A1(n18224), .A2(n17998), .B1(n17977), 
        .B2(n18225), .Y(n18004) );
  sky130_fd_sc_hd__xnor2_1 U24768 ( .A(n18651), .B(n22919), .Y(n18022) );
  sky130_fd_sc_hd__o22ai_1 U24769 ( .A1(n18067), .A2(n18022), .B1(n17978), 
        .B2(n18068), .Y(n18009) );
  sky130_fd_sc_hd__xnor2_1 U24770 ( .A(n18511), .B(n22951), .Y(n17997) );
  sky130_fd_sc_hd__o22ai_1 U24771 ( .A1(n12367), .A2(n17997), .B1(n17979), 
        .B2(n18470), .Y(n18008) );
  sky130_fd_sc_hd__xnor2_1 U24772 ( .A(n18649), .B(n18300), .Y(n18018) );
  sky130_fd_sc_hd__o22ai_1 U24773 ( .A1(n18370), .A2(n18018), .B1(n17980), 
        .B2(n17392), .Y(n18007) );
  sky130_fd_sc_hd__o22ai_1 U24774 ( .A1(n18151), .A2(n17982), .B1(n17981), 
        .B2(n18148), .Y(n17991) );
  sky130_fd_sc_hd__o22ai_1 U24775 ( .A1(n25219), .A2(n17983), .B1(n22337), 
        .B2(n18307), .Y(n17990) );
  sky130_fd_sc_hd__xnor2_1 U24776 ( .A(n17985), .B(n17984), .Y(n17989) );
  sky130_fd_sc_hd__fah_1 U24777 ( .A(n17988), .B(n17987), .CI(n17986), .COUT(
        n18079), .SUM(n18083) );
  sky130_fd_sc_hd__fah_1 U24778 ( .A(n17991), .B(n17990), .CI(n17989), .COUT(
        n18012), .SUM(n18078) );
  sky130_fd_sc_hd__o21ai_1 U24779 ( .A1(n18079), .A2(n18078), .B1(n18081), .Y(
        n17996) );
  sky130_fd_sc_hd__nand2_1 U24780 ( .A(n18079), .B(n18078), .Y(n17995) );
  sky130_fd_sc_hd__xnor2_1 U24781 ( .A(n18667), .B(n22951), .Y(n18063) );
  sky130_fd_sc_hd__o22ai_1 U24782 ( .A1(n12367), .A2(n18063), .B1(n17997), 
        .B2(n18470), .Y(n18071) );
  sky130_fd_sc_hd__nor2b_1 U24783 ( .B_N(n18353), .A(n18711), .Y(n18043) );
  sky130_fd_sc_hd__xnor2_1 U24784 ( .A(n18685), .B(n21887), .Y(n18064) );
  sky130_fd_sc_hd__o22ai_1 U24785 ( .A1(n18224), .A2(n18064), .B1(n17998), 
        .B2(n18225), .Y(n18042) );
  sky130_fd_sc_hd__xnor2_1 U24786 ( .A(n18043), .B(n18042), .Y(n18070) );
  sky130_fd_sc_hd__a22o_1 U24787 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[8]), .B1(n18183), .B2(
        j202_soc_core_j22_cpu_ml_macl[24]), .X(n18069) );
  sky130_fd_sc_hd__fah_1 U24788 ( .A(n18001), .B(n18000), .CI(n17999), .COUT(
        n18073), .SUM(n18011) );
  sky130_fd_sc_hd__fa_1 U24789 ( .A(n18009), .B(n18007), .CIN(n18008), .COUT(
        n18038), .SUM(n18013) );
  sky130_fd_sc_hd__fah_1 U24790 ( .A(n18014), .B(n18013), .CI(n18012), .COUT(
        n18048), .SUM(n18010) );
  sky130_fd_sc_hd__xnor2_1 U24791 ( .A(n18654), .B(n18300), .Y(n18062) );
  sky130_fd_sc_hd__o22ai_1 U24792 ( .A1(n18370), .A2(n18062), .B1(n18018), 
        .B2(n17392), .Y(n18054) );
  sky130_fd_sc_hd__xnor2_1 U24793 ( .A(n18426), .B(n22029), .Y(n18059) );
  sky130_fd_sc_hd__xnor2_1 U24794 ( .A(n18479), .B(n22112), .Y(n18060) );
  sky130_fd_sc_hd__o22ai_1 U24795 ( .A1(n12140), .A2(n18060), .B1(n18020), 
        .B2(n18424), .Y(n18052) );
  sky130_fd_sc_hd__xnor2_1 U24796 ( .A(n18687), .B(n18147), .Y(n18041) );
  sky130_fd_sc_hd__o22ai_1 U24797 ( .A1(n18151), .A2(n18041), .B1(n18021), 
        .B2(n18148), .Y(n18051) );
  sky130_fd_sc_hd__xnor2_1 U24798 ( .A(n22052), .B(n22919), .Y(n18066) );
  sky130_fd_sc_hd__o22ai_1 U24799 ( .A1(n18067), .A2(n18066), .B1(n18022), 
        .B2(n10971), .Y(n18050) );
  sky130_fd_sc_hd__xnor2_1 U24800 ( .A(n18661), .B(n18883), .Y(n18061) );
  sky130_fd_sc_hd__o22ai_1 U24801 ( .A1(n18344), .A2(n18061), .B1(n18023), 
        .B2(n17402), .Y(n18049) );
  sky130_fd_sc_hd__xnor2_1 U24802 ( .A(n18034), .B(n18035), .Y(n18024) );
  sky130_fd_sc_hd__xnor2_1 U24803 ( .A(n18033), .B(n18024), .Y(n18047) );
  sky130_fd_sc_hd__nand2_1 U24804 ( .A(n18027), .B(n18026), .Y(n18028) );
  sky130_fd_sc_hd__nand2_1 U24805 ( .A(n18029), .B(n18028), .Y(n18046) );
  sky130_fd_sc_hd__fah_1 U24806 ( .A(n18032), .B(n18031), .CI(n18030), .COUT(
        n18275), .SUM(n18274) );
  sky130_fd_sc_hd__o21ai_1 U24807 ( .A1(n18034), .A2(n18035), .B1(n18033), .Y(
        n18037) );
  sky130_fd_sc_hd__nand2_1 U24808 ( .A(n18035), .B(n18034), .Y(n18036) );
  sky130_fd_sc_hd__nand2_1 U24809 ( .A(n18037), .B(n18036), .Y(n18126) );
  sky130_fd_sc_hd__fah_1 U24810 ( .A(n18040), .B(n18039), .CI(n18038), .COUT(
        n18128), .SUM(n18072) );
  sky130_fd_sc_hd__xnor2_1 U24811 ( .A(n18651), .B(n18147), .Y(n18149) );
  sky130_fd_sc_hd__o22ai_1 U24812 ( .A1(n18151), .A2(n18149), .B1(n18041), 
        .B2(n18148), .Y(n18118) );
  sky130_fd_sc_hd__o22ai_1 U24814 ( .A1(n25219), .A2(n18044), .B1(n22841), 
        .B2(n18307), .Y(n18116) );
  sky130_fd_sc_hd__xnor2_1 U24815 ( .A(n18128), .B(n18127), .Y(n18045) );
  sky130_fd_sc_hd__xnor2_1 U24816 ( .A(n18126), .B(n18045), .Y(n18179) );
  sky130_fd_sc_hd__fah_1 U24817 ( .A(n18048), .B(n18047), .CI(n18046), .COUT(
        n18178), .SUM(n18030) );
  sky130_fd_sc_hd__fah_1 U24818 ( .A(n18054), .B(n18053), .CI(n18052), .COUT(
        n18159), .SUM(n18034) );
  sky130_fd_sc_hd__buf_4 U24819 ( .A(j202_soc_core_j22_cpu_ml_bufa[25]), .X(
        n18656) );
  sky130_fd_sc_hd__xnor2_1 U24820 ( .A(j202_soc_core_j22_cpu_ml_bufa[25]), .B(
        n24583), .Y(n18055) );
  sky130_fd_sc_hd__nand2_4 U24821 ( .A(n18056), .B(n12131), .Y(n18712) );
  sky130_fd_sc_hd__o22ai_1 U24822 ( .A1(n18711), .A2(n18058), .B1(n18057), 
        .B2(n18712), .Y(n18097) );
  sky130_fd_sc_hd__xnor2_1 U24823 ( .A(n18466), .B(n22029), .Y(n18109) );
  sky130_fd_sc_hd__xnor2_1 U24824 ( .A(n18511), .B(n22112), .Y(n18110) );
  sky130_fd_sc_hd__o22ai_1 U24825 ( .A1(n18514), .A2(n18110), .B1(n18060), 
        .B2(n18515), .Y(n18095) );
  sky130_fd_sc_hd__xnor2_1 U24826 ( .A(n18673), .B(n18883), .Y(n18111) );
  sky130_fd_sc_hd__o22ai_1 U24827 ( .A1(n18344), .A2(n18111), .B1(n18061), 
        .B2(n17402), .Y(n18103) );
  sky130_fd_sc_hd__xnor2_1 U24828 ( .A(n18708), .B(n18300), .Y(n18113) );
  sky130_fd_sc_hd__o22ai_1 U24829 ( .A1(n18370), .A2(n18113), .B1(n18062), 
        .B2(n17392), .Y(n18102) );
  sky130_fd_sc_hd__xnor2_1 U24830 ( .A(n18649), .B(n22951), .Y(n18115) );
  sky130_fd_sc_hd__o22ai_1 U24831 ( .A1(n12367), .A2(n18115), .B1(n18063), 
        .B2(n18470), .Y(n18101) );
  sky130_fd_sc_hd__xnor2_1 U24832 ( .A(n18721), .B(n21887), .Y(n18105) );
  sky130_fd_sc_hd__xnor2_1 U24833 ( .A(n18367), .B(n18656), .Y(n18108) );
  sky130_fd_sc_hd__xnor2_1 U24834 ( .A(n18656), .B(n18353), .Y(n18065) );
  sky130_fd_sc_hd__o22ai_1 U24835 ( .A1(n18711), .A2(n18108), .B1(n18065), 
        .B2(n18712), .Y(n18099) );
  sky130_fd_sc_hd__nor2_1 U24836 ( .A(n21980), .B(n22828), .Y(n18278) );
  sky130_fd_sc_hd__fah_1 U24837 ( .A(n18077), .B(n18076), .CI(n18075), .COUT(
        n18273), .SUM(n18272) );
  sky130_fd_sc_hd__xnor2_1 U24838 ( .A(n18081), .B(n18080), .Y(n18094) );
  sky130_fd_sc_hd__nand2_1 U24839 ( .A(n18084), .B(n18083), .Y(n18085) );
  sky130_fd_sc_hd__fah_1 U24840 ( .A(n18091), .B(n12209), .CI(n18090), .COUT(
        n18269), .SUM(n17929) );
  sky130_fd_sc_hd__fah_1 U24841 ( .A(n18094), .B(n18093), .CI(n18092), .COUT(
        n18271), .SUM(n18270) );
  sky130_fd_sc_hd__nor2_1 U24842 ( .A(n18269), .B(n18270), .Y(n21574) );
  sky130_fd_sc_hd__nand2_1 U24843 ( .A(n18278), .B(n22831), .Y(n19481) );
  sky130_fd_sc_hd__fah_1 U24844 ( .A(n18103), .B(n18102), .CI(n18101), .COUT(
        n18161), .SUM(n18122) );
  sky130_fd_sc_hd__xnor2_1 U24845 ( .A(n18673), .B(n18300), .Y(n18234) );
  sky130_fd_sc_hd__xnor2_1 U24846 ( .A(n18661), .B(n18300), .Y(n18114) );
  sky130_fd_sc_hd__o22ai_1 U24847 ( .A1(n18370), .A2(n18234), .B1(n18114), 
        .B2(n17392), .Y(n18202) );
  sky130_fd_sc_hd__xnor2_1 U24848 ( .A(j202_soc_core_j22_cpu_ml_bufa[26]), .B(
        j202_soc_core_j22_cpu_ml_bufa[25]), .Y(n18104) );
  sky130_fd_sc_hd__buf_2 U24849 ( .A(n18104), .X(n18619) );
  sky130_fd_sc_hd__nor2b_1 U24850 ( .B_N(n18353), .A(n18619), .Y(n18154) );
  sky130_fd_sc_hd__xnor2_1 U24851 ( .A(n18687), .B(n21887), .Y(n18139) );
  sky130_fd_sc_hd__o22ai_1 U24852 ( .A1(n18224), .A2(n18139), .B1(n18105), 
        .B2(n18225), .Y(n18153) );
  sky130_fd_sc_hd__o22ai_1 U24853 ( .A1(n25219), .A2(n18107), .B1(n18106), 
        .B2(n18307), .Y(n18201) );
  sky130_fd_sc_hd__xnor2_1 U24854 ( .A(n18211), .B(n18210), .Y(n18119) );
  sky130_fd_sc_hd__xnor2_1 U24855 ( .A(n18426), .B(n18656), .Y(n18136) );
  sky130_fd_sc_hd__o22ai_1 U24856 ( .A1(n18711), .A2(n18136), .B1(n18108), 
        .B2(n18712), .Y(n18135) );
  sky130_fd_sc_hd__xnor2_1 U24857 ( .A(n18479), .B(n22029), .Y(n18137) );
  sky130_fd_sc_hd__xnor2_1 U24858 ( .A(n18667), .B(n22112), .Y(n18138) );
  sky130_fd_sc_hd__xnor2_1 U24859 ( .A(n18685), .B(n18883), .Y(n18146) );
  sky130_fd_sc_hd__o22ai_1 U24860 ( .A1(n18344), .A2(n18146), .B1(n18111), 
        .B2(n17402), .Y(n18133) );
  sky130_fd_sc_hd__o22ai_1 U24861 ( .A1(n18370), .A2(n18114), .B1(n18113), 
        .B2(n17392), .Y(n18132) );
  sky130_fd_sc_hd__xnor2_1 U24862 ( .A(n18654), .B(n22951), .Y(n18144) );
  sky130_fd_sc_hd__o22ai_1 U24863 ( .A1(n12367), .A2(n18144), .B1(n18115), 
        .B2(n18470), .Y(n18131) );
  sky130_fd_sc_hd__fah_1 U24864 ( .A(n18118), .B(n18117), .CI(n18116), .COUT(
        n18123), .SUM(n18127) );
  sky130_fd_sc_hd__xnor2_1 U24865 ( .A(n18119), .B(n18209), .Y(n18263) );
  sky130_fd_sc_hd__fah_1 U24866 ( .A(n18125), .B(n18124), .CI(n18123), .COUT(
        n18209), .SUM(n18172) );
  sky130_fd_sc_hd__nand2_1 U24867 ( .A(n18128), .B(n18127), .Y(n18129) );
  sky130_fd_sc_hd__nand2_1 U24868 ( .A(n18130), .B(n18129), .Y(n18171) );
  sky130_fd_sc_hd__fah_1 U24869 ( .A(n18133), .B(n18132), .CI(n18131), .COUT(
        n18244), .SUM(n18124) );
  sky130_fd_sc_hd__xnor2_1 U24870 ( .A(n18466), .B(n18656), .Y(n18198) );
  sky130_fd_sc_hd__o22ai_1 U24871 ( .A1(n18711), .A2(n18198), .B1(n18136), 
        .B2(n18712), .Y(n18187) );
  sky130_fd_sc_hd__xnor2_1 U24872 ( .A(n18511), .B(n22029), .Y(n18200) );
  sky130_fd_sc_hd__xnor2_1 U24873 ( .A(n18649), .B(n22112), .Y(n18197) );
  sky130_fd_sc_hd__o22ai_1 U24874 ( .A1(n18514), .A2(n18197), .B1(n18138), 
        .B2(n18424), .Y(n18185) );
  sky130_fd_sc_hd__xnor2_1 U24875 ( .A(n18651), .B(n21887), .Y(n18184) );
  sky130_fd_sc_hd__o22ai_1 U24876 ( .A1(n18224), .A2(n18184), .B1(n18139), 
        .B2(n18225), .Y(n18193) );
  sky130_fd_sc_hd__inv_2 U24877 ( .A(n18140), .Y(n18716) );
  sky130_fd_sc_hd__nand2b_1 U24878 ( .A_N(n18353), .B(n22685), .Y(n18143) );
  sky130_fd_sc_hd__xor2_1 U24879 ( .A(j202_soc_core_j22_cpu_ml_bufa[27]), .B(
        n25085), .X(n18141) );
  sky130_fd_sc_hd__nand2_4 U24880 ( .A(n18141), .B(n18619), .Y(n18713) );
  sky130_fd_sc_hd__o22ai_1 U24881 ( .A1(n18619), .A2(n18143), .B1(n18142), 
        .B2(n18713), .Y(n18192) );
  sky130_fd_sc_hd__xnor2_1 U24882 ( .A(n18708), .B(n22951), .Y(n18195) );
  sky130_fd_sc_hd__o22ai_1 U24883 ( .A1(n12367), .A2(n18195), .B1(n18144), 
        .B2(n18470), .Y(n18191) );
  sky130_fd_sc_hd__xnor2_1 U24884 ( .A(n18367), .B(n22685), .Y(n18199) );
  sky130_fd_sc_hd__xnor2_1 U24885 ( .A(n22685), .B(n18353), .Y(n18145) );
  sky130_fd_sc_hd__o22ai_1 U24886 ( .A1(n18619), .A2(n18199), .B1(n18145), 
        .B2(n18713), .Y(n18190) );
  sky130_fd_sc_hd__xnor2_1 U24887 ( .A(n18721), .B(n18883), .Y(n18194) );
  sky130_fd_sc_hd__o22ai_1 U24888 ( .A1(n18344), .A2(n18194), .B1(n18146), 
        .B2(n17402), .Y(n18189) );
  sky130_fd_sc_hd__xnor2_1 U24889 ( .A(n22052), .B(n18147), .Y(n18150) );
  sky130_fd_sc_hd__o22ai_1 U24890 ( .A1(n18151), .A2(n18150), .B1(n18149), 
        .B2(n18148), .Y(n18157) );
  sky130_fd_sc_hd__o22ai_1 U24891 ( .A1(n25219), .A2(n18152), .B1(n22407), 
        .B2(n18307), .Y(n18156) );
  sky130_fd_sc_hd__xnor2_1 U24892 ( .A(n18154), .B(n18153), .Y(n18155) );
  sky130_fd_sc_hd__fah_1 U24893 ( .A(n18157), .B(n18156), .CI(n18155), .COUT(
        n18206), .SUM(n18166) );
  sky130_fd_sc_hd__fah_1 U24894 ( .A(n18160), .B(n18159), .CI(n18158), .COUT(
        n18170), .SUM(n18176) );
  sky130_fd_sc_hd__fah_1 U24895 ( .A(n18163), .B(n18162), .CI(n18161), .COUT(
        n18211), .SUM(n18167) );
  sky130_fd_sc_hd__nand2_1 U24897 ( .A(n18170), .B(n18166), .Y(n18164) );
  sky130_fd_sc_hd__xnor2_1 U24898 ( .A(n18168), .B(n18167), .Y(n18169) );
  sky130_fd_sc_hd__xor2_1 U24899 ( .A(n18170), .B(n18169), .X(n18182) );
  sky130_fd_sc_hd__fah_1 U24900 ( .A(n18173), .B(n18172), .CI(n18171), .COUT(
        n18262), .SUM(n18181) );
  sky130_fd_sc_hd__fah_1 U24901 ( .A(n18176), .B(n18175), .CI(n18174), .COUT(
        n18180), .SUM(n18177) );
  sky130_fd_sc_hd__nor2_2 U24902 ( .A(n18282), .B(n18281), .Y(n21437) );
  sky130_fd_sc_hd__fah_1 U24903 ( .A(n18179), .B(n18177), .CI(n18178), .COUT(
        n18279), .SUM(n18276) );
  sky130_fd_sc_hd__fah_1 U24904 ( .A(n18182), .B(n18181), .CI(n18180), .COUT(
        n18281), .SUM(n18280) );
  sky130_fd_sc_hd__nor2_1 U24905 ( .A(n18279), .B(n18280), .Y(n19221) );
  sky130_fd_sc_hd__nor2_1 U24906 ( .A(n21437), .B(n19221), .Y(n19482) );
  sky130_fd_sc_hd__xnor2_1 U24907 ( .A(n18673), .B(n22951), .Y(n18313) );
  sky130_fd_sc_hd__xnor2_1 U24908 ( .A(n18661), .B(n22951), .Y(n18196) );
  sky130_fd_sc_hd__o22ai_1 U24909 ( .A1(n12367), .A2(n18313), .B1(n18196), 
        .B2(n18470), .Y(n18323) );
  sky130_fd_sc_hd__nor2b_1 U24910 ( .B_N(n18353), .A(n18750), .Y(n18237) );
  sky130_fd_sc_hd__xnor2_1 U24911 ( .A(n22052), .B(n21887), .Y(n18223) );
  sky130_fd_sc_hd__o22ai_1 U24912 ( .A1(n18224), .A2(n18223), .B1(n18184), 
        .B2(n18225), .Y(n18236) );
  sky130_fd_sc_hd__fah_1 U24913 ( .A(n18187), .B(n18186), .CI(n18185), .COUT(
        n18247), .SUM(n18242) );
  sky130_fd_sc_hd__fah_1 U24914 ( .A(n18190), .B(n18189), .CI(n18188), .COUT(
        n18246), .SUM(n18207) );
  sky130_fd_sc_hd__xnor2_1 U24915 ( .A(n18687), .B(n18883), .Y(n18222) );
  sky130_fd_sc_hd__o22ai_1 U24916 ( .A1(n18344), .A2(n18222), .B1(n18194), 
        .B2(n17402), .Y(n18221) );
  sky130_fd_sc_hd__o22ai_1 U24917 ( .A1(n12367), .A2(n18196), .B1(n18195), 
        .B2(n18470), .Y(n18220) );
  sky130_fd_sc_hd__xnor2_1 U24918 ( .A(n18654), .B(n22112), .Y(n18233) );
  sky130_fd_sc_hd__o22ai_1 U24919 ( .A1(n18514), .A2(n18233), .B1(n18197), 
        .B2(n18515), .Y(n18219) );
  sky130_fd_sc_hd__xnor2_1 U24920 ( .A(n18479), .B(n18656), .Y(n18228) );
  sky130_fd_sc_hd__o22ai_1 U24921 ( .A1(n18711), .A2(n18228), .B1(n18198), 
        .B2(n18712), .Y(n18218) );
  sky130_fd_sc_hd__xnor2_1 U24922 ( .A(n18426), .B(n22685), .Y(n18231) );
  sky130_fd_sc_hd__o22ai_1 U24923 ( .A1(n18619), .A2(n18231), .B1(n18199), 
        .B2(n18713), .Y(n18217) );
  sky130_fd_sc_hd__xnor2_1 U24924 ( .A(n18667), .B(n22029), .Y(n18232) );
  sky130_fd_sc_hd__fah_1 U24925 ( .A(n18205), .B(n18204), .CI(n18203), .COUT(
        n18571), .SUM(n18256) );
  sky130_fd_sc_hd__fah_1 U24926 ( .A(n18208), .B(n18207), .CI(n18206), .COUT(
        n18255), .SUM(n18253) );
  sky130_fd_sc_hd__o21ai_1 U24927 ( .A1(n18211), .A2(n18210), .B1(n18209), .Y(
        n18213) );
  sky130_fd_sc_hd__nand2_1 U24928 ( .A(n18211), .B(n18210), .Y(n18212) );
  sky130_fd_sc_hd__nand2_1 U24929 ( .A(n18213), .B(n18212), .Y(n18258) );
  sky130_fd_sc_hd__o21ai_1 U24930 ( .A1(n18255), .A2(n18256), .B1(n18258), .Y(
        n18215) );
  sky130_fd_sc_hd__nand2_1 U24931 ( .A(n18255), .B(n18256), .Y(n18214) );
  sky130_fd_sc_hd__nand2_1 U24932 ( .A(n18215), .B(n18214), .Y(n18591) );
  sky130_fd_sc_hd__fah_1 U24933 ( .A(n18218), .B(n18217), .CI(n18216), .COUT(
        n18554), .SUM(n18204) );
  sky130_fd_sc_hd__fah_1 U24934 ( .A(n18221), .B(n18219), .CI(n18220), .COUT(
        n18553), .SUM(n18205) );
  sky130_fd_sc_hd__xnor2_1 U24935 ( .A(n18651), .B(n18883), .Y(n18294) );
  sky130_fd_sc_hd__o22ai_1 U24936 ( .A1(n18344), .A2(n18294), .B1(n18222), 
        .B2(n17402), .Y(n18328) );
  sky130_fd_sc_hd__xnor2_1 U24937 ( .A(n18367), .B(n18720), .Y(n18319) );
  sky130_fd_sc_hd__xnor2_1 U24938 ( .A(n18672), .B(n18226), .Y(n18227) );
  sky130_fd_sc_hd__o22ai_1 U24939 ( .A1(n18750), .A2(n18319), .B1(n18227), 
        .B2(n18747), .Y(n18327) );
  sky130_fd_sc_hd__xnor2_1 U24940 ( .A(n18511), .B(n18656), .Y(n18310) );
  sky130_fd_sc_hd__o22ai_1 U24941 ( .A1(n18711), .A2(n18310), .B1(n18228), 
        .B2(n18712), .Y(n18331) );
  sky130_fd_sc_hd__nand2b_1 U24942 ( .A_N(n18353), .B(n18720), .Y(n18230) );
  sky130_fd_sc_hd__xnor2_1 U24943 ( .A(n18466), .B(n22685), .Y(n18317) );
  sky130_fd_sc_hd__o22ai_1 U24944 ( .A1(n18716), .A2(n18317), .B1(n18231), 
        .B2(n18713), .Y(n18329) );
  sky130_fd_sc_hd__xnor2_1 U24945 ( .A(n18721), .B(n18300), .Y(n18311) );
  sky130_fd_sc_hd__xnor2_1 U24946 ( .A(n18685), .B(n18300), .Y(n18235) );
  sky130_fd_sc_hd__o22ai_1 U24947 ( .A1(n18370), .A2(n18311), .B1(n18235), 
        .B2(n17392), .Y(n18334) );
  sky130_fd_sc_hd__xnor2_1 U24948 ( .A(n18649), .B(n22029), .Y(n18305) );
  sky130_fd_sc_hd__xnor2_1 U24949 ( .A(n18708), .B(n22112), .Y(n18315) );
  sky130_fd_sc_hd__o22ai_1 U24950 ( .A1(n18514), .A2(n18315), .B1(n18233), 
        .B2(n18424), .Y(n18332) );
  sky130_fd_sc_hd__o22ai_1 U24951 ( .A1(n18370), .A2(n18235), .B1(n18234), 
        .B2(n17392), .Y(n18241) );
  sky130_fd_sc_hd__xnor2_1 U24952 ( .A(n18237), .B(n18236), .Y(n18240) );
  sky130_fd_sc_hd__o22ai_1 U24953 ( .A1(n25219), .A2(n18238), .B1(n22638), 
        .B2(n18307), .Y(n18239) );
  sky130_fd_sc_hd__fah_1 U24954 ( .A(n18244), .B(n18243), .CI(n18242), .COUT(
        n18252), .SUM(n18254) );
  sky130_fd_sc_hd__nand2_1 U24955 ( .A(n18252), .B(n18250), .Y(n18248) );
  sky130_fd_sc_hd__xnor2_1 U24956 ( .A(n18250), .B(n18249), .Y(n18251) );
  sky130_fd_sc_hd__xnor2_1 U24957 ( .A(n18252), .B(n18251), .Y(n18265) );
  sky130_fd_sc_hd__nand2_1 U24959 ( .A(n18267), .B(n18265), .Y(n18259) );
  sky130_fd_sc_hd__nand2_1 U24960 ( .A(n18260), .B(n18259), .Y(n18285) );
  sky130_fd_sc_hd__nor2_1 U24961 ( .A(n18286), .B(n18285), .Y(n21870) );
  sky130_fd_sc_hd__fah_1 U24962 ( .A(n18262), .B(n18263), .CI(n18261), .COUT(
        n18283), .SUM(n18282) );
  sky130_fd_sc_hd__xnor2_1 U24963 ( .A(n18265), .B(n18264), .Y(n18266) );
  sky130_fd_sc_hd__nor2_1 U24964 ( .A(n21870), .B(n21878), .Y(n18288) );
  sky130_fd_sc_hd__nand2_1 U24965 ( .A(n19482), .B(n18288), .Y(n18290) );
  sky130_fd_sc_hd__nand2_1 U24966 ( .A(n18911), .B(n18268), .Y(n18293) );
  sky130_fd_sc_hd__nand2_1 U24967 ( .A(n18272), .B(n18271), .Y(n18909) );
  sky130_fd_sc_hd__nand2_1 U24968 ( .A(n18274), .B(n18273), .Y(n22832) );
  sky130_fd_sc_hd__nand2_1 U24969 ( .A(n18276), .B(n18275), .Y(n22829) );
  sky130_fd_sc_hd__o21ai_1 U24970 ( .A1(n22832), .A2(n22828), .B1(n22829), .Y(
        n18277) );
  sky130_fd_sc_hd__a21oi_1 U24971 ( .A1(n18278), .A2(n22835), .B1(n18277), .Y(
        n19223) );
  sky130_fd_sc_hd__nand2_1 U24972 ( .A(n18280), .B(n18279), .Y(n19222) );
  sky130_fd_sc_hd__nand2_1 U24973 ( .A(n18281), .B(n18282), .Y(n21438) );
  sky130_fd_sc_hd__nand2_1 U24974 ( .A(n18284), .B(n18283), .Y(n21876) );
  sky130_fd_sc_hd__nand2_1 U24975 ( .A(n18286), .B(n18285), .Y(n21871) );
  sky130_fd_sc_hd__o21ai_1 U24976 ( .A1(n21876), .A2(n21870), .B1(n21871), .Y(
        n18287) );
  sky130_fd_sc_hd__o21ai_1 U24977 ( .A1(n18290), .A2(n19223), .B1(n18289), .Y(
        n18291) );
  sky130_fd_sc_hd__nand2_4 U24978 ( .A(n18293), .B(n18292), .Y(n19249) );
  sky130_fd_sc_hd__xnor2_1 U24979 ( .A(n18687), .B(n22951), .Y(n18373) );
  sky130_fd_sc_hd__xnor2_1 U24980 ( .A(n18721), .B(n22951), .Y(n18298) );
  sky130_fd_sc_hd__o22ai_1 U24981 ( .A1(n12367), .A2(n18373), .B1(n18298), 
        .B2(n18470), .Y(n18364) );
  sky130_fd_sc_hd__xnor2_1 U24982 ( .A(n18479), .B(n18672), .Y(n18371) );
  sky130_fd_sc_hd__xnor2_1 U24983 ( .A(n18466), .B(n18720), .Y(n18304) );
  sky130_fd_sc_hd__o22ai_1 U24984 ( .A1(n18750), .A2(n18371), .B1(n18304), 
        .B2(n18747), .Y(n18363) );
  sky130_fd_sc_hd__xnor2_1 U24985 ( .A(n18661), .B(n22029), .Y(n18351) );
  sky130_fd_sc_hd__xnor2_1 U24986 ( .A(n18708), .B(n22029), .Y(n18299) );
  sky130_fd_sc_hd__xnor2_1 U24987 ( .A(n18426), .B(n22487), .Y(n18374) );
  sky130_fd_sc_hd__xnor2_1 U24988 ( .A(n18367), .B(n22487), .Y(n18342) );
  sky130_fd_sc_hd__xnor2_1 U24989 ( .A(n18667), .B(n22685), .Y(n18372) );
  sky130_fd_sc_hd__xnor2_1 U24990 ( .A(n18511), .B(n22685), .Y(n18297) );
  sky130_fd_sc_hd__o22ai_1 U24991 ( .A1(n18716), .A2(n18372), .B1(n18297), 
        .B2(n18713), .Y(n18360) );
  sky130_fd_sc_hd__xnor2_1 U24992 ( .A(n22052), .B(n18300), .Y(n18369) );
  sky130_fd_sc_hd__xnor2_1 U24993 ( .A(n18651), .B(n18300), .Y(n18301) );
  sky130_fd_sc_hd__o22ai_1 U24994 ( .A1(n18370), .A2(n18369), .B1(n18301), 
        .B2(n17392), .Y(n18359) );
  sky130_fd_sc_hd__xnor2_1 U24995 ( .A(n18673), .B(n22112), .Y(n18376) );
  sky130_fd_sc_hd__xnor2_1 U24996 ( .A(n18661), .B(n22112), .Y(n18316) );
  sky130_fd_sc_hd__o22ai_1 U24997 ( .A1(n12140), .A2(n18376), .B1(n18316), 
        .B2(n18424), .Y(n18326) );
  sky130_fd_sc_hd__nor2b_1 U24998 ( .B_N(n18353), .A(n18719), .Y(n18309) );
  sky130_fd_sc_hd__xnor2_1 U24999 ( .A(n22052), .B(n18883), .Y(n18343) );
  sky130_fd_sc_hd__o22ai_1 U25000 ( .A1(n25219), .A2(n18296), .B1(n18295), 
        .B2(n18307), .Y(n18324) );
  sky130_fd_sc_hd__xnor2_1 U25001 ( .A(n18479), .B(n22685), .Y(n18318) );
  sky130_fd_sc_hd__o22ai_1 U25002 ( .A1(n18619), .A2(n18297), .B1(n18318), 
        .B2(n18713), .Y(n18347) );
  sky130_fd_sc_hd__xnor2_1 U25003 ( .A(n18685), .B(n22951), .Y(n18314) );
  sky130_fd_sc_hd__o22ai_1 U25004 ( .A1(n12367), .A2(n18298), .B1(n18314), 
        .B2(n18470), .Y(n18346) );
  sky130_fd_sc_hd__xnor2_1 U25005 ( .A(n18654), .B(n22029), .Y(n18306) );
  sky130_fd_sc_hd__xnor2_1 U25006 ( .A(n18687), .B(n18300), .Y(n18312) );
  sky130_fd_sc_hd__o22ai_1 U25007 ( .A1(n18370), .A2(n18301), .B1(n18312), 
        .B2(n17392), .Y(n18350) );
  sky130_fd_sc_hd__nand2b_1 U25008 ( .A_N(n18353), .B(n22487), .Y(n18303) );
  sky130_fd_sc_hd__xnor2_1 U25009 ( .A(n18426), .B(n18672), .Y(n18320) );
  sky130_fd_sc_hd__xnor2_1 U25010 ( .A(n18667), .B(n18656), .Y(n18340) );
  sky130_fd_sc_hd__o22ai_1 U25011 ( .A1(n18711), .A2(n18340), .B1(n18310), 
        .B2(n18712), .Y(n18386) );
  sky130_fd_sc_hd__o22ai_1 U25012 ( .A1(n18370), .A2(n18312), .B1(n18311), 
        .B2(n17392), .Y(n18385) );
  sky130_fd_sc_hd__o22ai_1 U25013 ( .A1(n12367), .A2(n18314), .B1(n18313), 
        .B2(n18470), .Y(n18384) );
  sky130_fd_sc_hd__o22ai_1 U25014 ( .A1(n18514), .A2(n18316), .B1(n18315), 
        .B2(n18515), .Y(n18389) );
  sky130_fd_sc_hd__o22ai_1 U25015 ( .A1(n18716), .A2(n18318), .B1(n18317), 
        .B2(n18713), .Y(n18388) );
  sky130_fd_sc_hd__o22ai_1 U25016 ( .A1(n18750), .A2(n18320), .B1(n18319), 
        .B2(n18747), .Y(n18387) );
  sky130_fd_sc_hd__fah_1 U25017 ( .A(n18334), .B(n18333), .CI(n18332), .COUT(
        n18558), .SUM(n18566) );
  sky130_fd_sc_hd__nand2_1 U25018 ( .A(n18578), .B(n18577), .Y(n18335) );
  sky130_fd_sc_hd__nand2_1 U25019 ( .A(n18336), .B(n18335), .Y(n18602) );
  sky130_fd_sc_hd__nand2_1 U25020 ( .A(n18338), .B(n18337), .Y(n18339) );
  sky130_fd_sc_hd__xnor2_1 U25021 ( .A(n18649), .B(n18656), .Y(n18354) );
  sky130_fd_sc_hd__o22ai_1 U25022 ( .A1(n18711), .A2(n18354), .B1(n18340), 
        .B2(n18712), .Y(n18392) );
  sky130_fd_sc_hd__xnor2_1 U25023 ( .A(n22487), .B(n18353), .Y(n18341) );
  sky130_fd_sc_hd__xnor2_1 U25024 ( .A(n18673), .B(n22029), .Y(n18402) );
  sky130_fd_sc_hd__a22oi_1 U25025 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[17]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[1]), .Y(n18352) );
  sky130_fd_sc_hd__xnor2_1 U25027 ( .A(n18654), .B(n18656), .Y(n18365) );
  sky130_fd_sc_hd__o22ai_1 U25028 ( .A1(n18711), .A2(n18365), .B1(n18354), 
        .B2(n18712), .Y(n18378) );
  sky130_fd_sc_hd__or2_0 U25029 ( .A(n18379), .B(n18378), .X(n18430) );
  sky130_fd_sc_hd__xnor2_1 U25030 ( .A(n18419), .B(n18418), .Y(n18358) );
  sky130_fd_sc_hd__xnor2_1 U25031 ( .A(n18358), .B(n18417), .Y(n18605) );
  sky130_fd_sc_hd__nand2_1 U25032 ( .A(n13328), .B(n18605), .Y(n18398) );
  sky130_fd_sc_hd__xnor2_1 U25033 ( .A(n18708), .B(n18656), .Y(n18429) );
  sky130_fd_sc_hd__o22ai_1 U25034 ( .A1(n12131), .A2(n18429), .B1(n18365), 
        .B2(n18712), .Y(n18407) );
  sky130_fd_sc_hd__xnor2_1 U25035 ( .A(n18367), .B(n22051), .Y(n18368) );
  sky130_fd_sc_hd__a21o_1 U25036 ( .A1(n17392), .A2(n18370), .B1(n18369), .X(
        n18405) );
  sky130_fd_sc_hd__xnor2_1 U25037 ( .A(n18721), .B(n22112), .Y(n18425) );
  sky130_fd_sc_hd__xnor2_1 U25038 ( .A(n18685), .B(n22112), .Y(n18377) );
  sky130_fd_sc_hd__o22ai_1 U25039 ( .A1(n12140), .A2(n18425), .B1(n18377), 
        .B2(n18515), .Y(n18413) );
  sky130_fd_sc_hd__xnor2_1 U25040 ( .A(n18511), .B(n18720), .Y(n18428) );
  sky130_fd_sc_hd__o22ai_1 U25041 ( .A1(n18750), .A2(n18428), .B1(n18371), 
        .B2(n18747), .Y(n18412) );
  sky130_fd_sc_hd__xnor2_1 U25042 ( .A(n18649), .B(n22685), .Y(n18403) );
  sky130_fd_sc_hd__o22ai_1 U25043 ( .A1(n18619), .A2(n18403), .B1(n18372), 
        .B2(n18713), .Y(n18411) );
  sky130_fd_sc_hd__xnor2_1 U25044 ( .A(n18651), .B(n22951), .Y(n18422) );
  sky130_fd_sc_hd__o22ai_1 U25045 ( .A1(n12367), .A2(n18422), .B1(n18373), 
        .B2(n18470), .Y(n18410) );
  sky130_fd_sc_hd__xnor2_1 U25046 ( .A(n18466), .B(n22487), .Y(n18423) );
  sky130_fd_sc_hd__xnor2_1 U25047 ( .A(n18379), .B(n18378), .Y(n18382) );
  sky130_fd_sc_hd__a22oi_1 U25048 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[16]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[0]), .Y(n18380) );
  sky130_fd_sc_hd__nand2_1 U25049 ( .A(n22071), .B(n18380), .Y(n18381) );
  sky130_fd_sc_hd__fa_1 U25050 ( .A(n18383), .B(n18382), .CIN(n18381), .COUT(
        n18433), .SUM(n18598) );
  sky130_fd_sc_hd__nand2_1 U25051 ( .A(n13328), .B(n18606), .Y(n18397) );
  sky130_fd_sc_hd__nand2_1 U25052 ( .A(n18605), .B(n18606), .Y(n18396) );
  sky130_fd_sc_hd__nand3_1 U25053 ( .A(n18398), .B(n18397), .C(n18396), .Y(
        n18817) );
  sky130_fd_sc_hd__xnor2_1 U25054 ( .A(n18685), .B(n22029), .Y(n18473) );
  sky130_fd_sc_hd__xnor2_1 U25055 ( .A(n18654), .B(n22685), .Y(n18472) );
  sky130_fd_sc_hd__o22ai_1 U25056 ( .A1(n18716), .A2(n18472), .B1(n18403), 
        .B2(n18713), .Y(n18464) );
  sky130_fd_sc_hd__a22oi_1 U25057 ( .A1(n24499), .A2(
        j202_soc_core_j22_cpu_ml_mach[18]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[2]), .Y(n18404) );
  sky130_fd_sc_hd__nand2_1 U25058 ( .A(n22071), .B(n18404), .Y(n18463) );
  sky130_fd_sc_hd__fah_1 U25059 ( .A(n18416), .B(n18415), .CI(n18414), .COUT(
        n18474), .SUM(n18401) );
  sky130_fd_sc_hd__o21ai_1 U25060 ( .A1(n18419), .A2(n18418), .B1(n18417), .Y(
        n18421) );
  sky130_fd_sc_hd__nand2_1 U25061 ( .A(n18419), .B(n18418), .Y(n18420) );
  sky130_fd_sc_hd__nand2_1 U25062 ( .A(n18421), .B(n18420), .Y(n18455) );
  sky130_fd_sc_hd__xnor2_1 U25063 ( .A(n22052), .B(n22951), .Y(n18468) );
  sky130_fd_sc_hd__o22ai_1 U25064 ( .A1(n12367), .A2(n18468), .B1(n18422), 
        .B2(n18470), .Y(n18454) );
  sky130_fd_sc_hd__xnor2_1 U25065 ( .A(n18479), .B(n22487), .Y(n18446) );
  sky130_fd_sc_hd__xnor2_1 U25066 ( .A(n18687), .B(n22112), .Y(n18471) );
  sky130_fd_sc_hd__o22ai_1 U25067 ( .A1(n12140), .A2(n18471), .B1(n18425), 
        .B2(n18424), .Y(n18452) );
  sky130_fd_sc_hd__xnor2_1 U25068 ( .A(n18426), .B(n22051), .Y(n18427) );
  sky130_fd_sc_hd__xnor2_1 U25069 ( .A(n18667), .B(n18672), .Y(n18447) );
  sky130_fd_sc_hd__xnor2_1 U25070 ( .A(n18661), .B(n18656), .Y(n18445) );
  sky130_fd_sc_hd__o22ai_1 U25071 ( .A1(n18711), .A2(n18445), .B1(n18429), 
        .B2(n18712), .Y(n18489) );
  sky130_fd_sc_hd__inv_1 U25072 ( .A(n18489), .Y(n18449) );
  sky130_fd_sc_hd__xnor2_1 U25074 ( .A(n18455), .B(n18436), .Y(n18437) );
  sky130_fd_sc_hd__nand2_1 U25075 ( .A(n18439), .B(n18438), .Y(n18440) );
  sky130_fd_sc_hd__nand2_1 U25076 ( .A(n18441), .B(n18440), .Y(n18819) );
  sky130_fd_sc_hd__fah_1 U25077 ( .A(n18444), .B(n18443), .CI(n18442), .COUT(
        n18492), .SUM(n18475) );
  sky130_fd_sc_hd__xnor2_1 U25078 ( .A(n18673), .B(n18656), .Y(n18481) );
  sky130_fd_sc_hd__o22ai_1 U25079 ( .A1(n18711), .A2(n18481), .B1(n18445), 
        .B2(n18712), .Y(n18500) );
  sky130_fd_sc_hd__xnor2_1 U25080 ( .A(n18511), .B(n22487), .Y(n18505) );
  sky130_fd_sc_hd__xnor2_1 U25081 ( .A(n18649), .B(n18672), .Y(n18478) );
  sky130_fd_sc_hd__o22ai_1 U25082 ( .A1(n18750), .A2(n18478), .B1(n18447), 
        .B2(n18747), .Y(n18498) );
  sky130_fd_sc_hd__a22oi_1 U25083 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[19]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[3]), .Y(n18448) );
  sky130_fd_sc_hd__nand2_1 U25084 ( .A(n22071), .B(n18448), .Y(n18484) );
  sky130_fd_sc_hd__fah_1 U25085 ( .A(n18451), .B(n18450), .CI(n18449), .COUT(
        n18483), .SUM(n18461) );
  sky130_fd_sc_hd__fah_1 U25086 ( .A(n18454), .B(n18453), .CI(n18452), .COUT(
        n18482), .SUM(n18462) );
  sky130_fd_sc_hd__nor2_1 U25087 ( .A(n18456), .B(n18457), .Y(n18459) );
  sky130_fd_sc_hd__o2bb2ai_1 U25088 ( .B1(n18459), .B2(n18458), .A1_N(n18457), 
        .A2_N(n18456), .Y(n18544) );
  sky130_fd_sc_hd__xnor2_1 U25089 ( .A(n18545), .B(n18544), .Y(n18477) );
  sky130_fd_sc_hd__fah_1 U25090 ( .A(n18462), .B(n18461), .CI(n18460), .COUT(
        n18510), .SUM(n18457) );
  sky130_fd_sc_hd__fah_1 U25091 ( .A(n18465), .B(n18464), .CI(n18463), .COUT(
        n18497), .SUM(n18476) );
  sky130_fd_sc_hd__xnor2_1 U25092 ( .A(n18466), .B(n22051), .Y(n18467) );
  sky130_fd_sc_hd__xnor2_1 U25093 ( .A(n18651), .B(n22112), .Y(n18504) );
  sky130_fd_sc_hd__o22ai_1 U25094 ( .A1(n12140), .A2(n18504), .B1(n18471), 
        .B2(n18515), .Y(n18503) );
  sky130_fd_sc_hd__xnor2_1 U25095 ( .A(n18708), .B(n22685), .Y(n18506) );
  sky130_fd_sc_hd__o22ai_1 U25096 ( .A1(n18716), .A2(n18506), .B1(n18472), 
        .B2(n18713), .Y(n18502) );
  sky130_fd_sc_hd__xnor2_1 U25097 ( .A(n18721), .B(n22029), .Y(n18485) );
  sky130_fd_sc_hd__xnor2_1 U25098 ( .A(n18654), .B(n18720), .Y(n18539) );
  sky130_fd_sc_hd__o22ai_1 U25099 ( .A1(n18750), .A2(n18539), .B1(n18478), 
        .B2(n18747), .Y(n18533) );
  sky130_fd_sc_hd__xnor2_1 U25100 ( .A(n18479), .B(n22051), .Y(n18480) );
  sky130_fd_sc_hd__xnor2_1 U25101 ( .A(n18685), .B(n18656), .Y(n18537) );
  sky130_fd_sc_hd__o22ai_1 U25102 ( .A1(n18711), .A2(n18537), .B1(n18481), 
        .B2(n18712), .Y(n18681) );
  sky130_fd_sc_hd__xnor2_1 U25103 ( .A(n18687), .B(n22029), .Y(n18516) );
  sky130_fd_sc_hd__a22oi_1 U25104 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[20]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[4]), .Y(n18486) );
  sky130_fd_sc_hd__nand2_1 U25105 ( .A(n22071), .B(n18486), .Y(n18521) );
  sky130_fd_sc_hd__fah_1 U25106 ( .A(n18489), .B(n18488), .CI(n18487), .COUT(
        n18520), .SUM(n18496) );
  sky130_fd_sc_hd__nand2_1 U25108 ( .A(n18492), .B(n18491), .Y(n18493) );
  sky130_fd_sc_hd__nand2_1 U25109 ( .A(n18494), .B(n18493), .Y(n18523) );
  sky130_fd_sc_hd__fah_1 U25110 ( .A(n18497), .B(n18496), .CI(n18495), .COUT(
        n18524), .SUM(n18509) );
  sky130_fd_sc_hd__fa_1 U25111 ( .A(n18500), .B(n18499), .CIN(n18498), .COUT(
        n18530), .SUM(n18491) );
  sky130_fd_sc_hd__fa_1 U25112 ( .A(n18501), .B(n18503), .CIN(n18502), .COUT(
        n18529), .SUM(n18495) );
  sky130_fd_sc_hd__xnor2_1 U25113 ( .A(n22052), .B(n22112), .Y(n18513) );
  sky130_fd_sc_hd__o22ai_1 U25114 ( .A1(n12140), .A2(n18513), .B1(n18504), 
        .B2(n18515), .Y(n18536) );
  sky130_fd_sc_hd__xnor2_1 U25115 ( .A(n18667), .B(n22487), .Y(n18538) );
  sky130_fd_sc_hd__xnor2_1 U25116 ( .A(n18661), .B(n22685), .Y(n18517) );
  sky130_fd_sc_hd__o22ai_1 U25117 ( .A1(n18716), .A2(n18517), .B1(n18506), 
        .B2(n18713), .Y(n18534) );
  sky130_fd_sc_hd__fah_1 U25118 ( .A(n18510), .B(n18509), .CI(n18508), .COUT(
        n18549), .SUM(n18546) );
  sky130_fd_sc_hd__xnor2_1 U25119 ( .A(n18511), .B(n22051), .Y(n18512) );
  sky130_fd_sc_hd__a21o_1 U25120 ( .A1(n18515), .A2(n12140), .B1(n18513), .X(
        n18679) );
  sky130_fd_sc_hd__xnor2_1 U25121 ( .A(n18651), .B(n22029), .Y(n18658) );
  sky130_fd_sc_hd__xnor2_1 U25122 ( .A(n18673), .B(n22685), .Y(n18663) );
  sky130_fd_sc_hd__o22ai_1 U25123 ( .A1(n18716), .A2(n18663), .B1(n18517), 
        .B2(n18713), .Y(n18670) );
  sky130_fd_sc_hd__a22oi_1 U25124 ( .A1(n24499), .A2(
        j202_soc_core_j22_cpu_ml_mach[21]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[5]), .Y(n18519) );
  sky130_fd_sc_hd__nand2_1 U25125 ( .A(n22071), .B(n18519), .Y(n18669) );
  sky130_fd_sc_hd__fah_1 U25126 ( .A(n18522), .B(n18521), .CI(n18520), .COUT(
        n18794), .SUM(n18540) );
  sky130_fd_sc_hd__o21ai_1 U25127 ( .A1(n18525), .A2(n18524), .B1(n18523), .Y(
        n18527) );
  sky130_fd_sc_hd__nand2_1 U25128 ( .A(n18525), .B(n18524), .Y(n18526) );
  sky130_fd_sc_hd__nand2_1 U25129 ( .A(n18527), .B(n18526), .Y(n18789) );
  sky130_fd_sc_hd__xnor2_1 U25130 ( .A(n18790), .B(n18789), .Y(n18543) );
  sky130_fd_sc_hd__fah_1 U25131 ( .A(n18530), .B(n18529), .CI(n18528), .COUT(
        n18802), .SUM(n18525) );
  sky130_fd_sc_hd__xnor2_1 U25132 ( .A(n18721), .B(n18656), .Y(n18648) );
  sky130_fd_sc_hd__o22ai_1 U25133 ( .A1(n18711), .A2(n18648), .B1(n18537), 
        .B2(n18712), .Y(n18684) );
  sky130_fd_sc_hd__xnor2_1 U25134 ( .A(n18649), .B(n22487), .Y(n18665) );
  sky130_fd_sc_hd__xnor2_1 U25135 ( .A(n18708), .B(n18720), .Y(n18662) );
  sky130_fd_sc_hd__o22ai_1 U25136 ( .A1(n18750), .A2(n18662), .B1(n18539), 
        .B2(n18747), .Y(n18682) );
  sky130_fd_sc_hd__fah_1 U25137 ( .A(n18542), .B(n18541), .CI(n18540), .COUT(
        n18800), .SUM(n18551) );
  sky130_fd_sc_hd__xnor2_1 U25138 ( .A(n18543), .B(n18791), .Y(n18822) );
  sky130_fd_sc_hd__nand2_1 U25140 ( .A(n18546), .B(n18545), .Y(n18547) );
  sky130_fd_sc_hd__nand2_1 U25141 ( .A(n18548), .B(n18547), .Y(n18820) );
  sky130_fd_sc_hd__fah_1 U25142 ( .A(n18554), .B(n18553), .CI(n18552), .COUT(
        n18588), .SUM(n18564) );
  sky130_fd_sc_hd__fah_1 U25143 ( .A(n18557), .B(n18556), .CI(n18555), .COUT(
        n18583), .SUM(n18587) );
  sky130_fd_sc_hd__fah_1 U25144 ( .A(n18560), .B(n18559), .CI(n18558), .COUT(
        n18578), .SUM(n18586) );
  sky130_fd_sc_hd__xnor2_1 U25145 ( .A(n18561), .B(n18586), .Y(n18562) );
  sky130_fd_sc_hd__fah_1 U25146 ( .A(n18567), .B(n18566), .CI(n18565), .COUT(
        n18576), .SUM(n18563) );
  sky130_fd_sc_hd__fah_1 U25147 ( .A(n18570), .B(n18569), .CI(n18568), .COUT(
        n18579), .SUM(n18575) );
  sky130_fd_sc_hd__xnor2_1 U25148 ( .A(n18578), .B(n18577), .Y(n18580) );
  sky130_fd_sc_hd__xnor2_1 U25149 ( .A(n18580), .B(n18579), .Y(n18609) );
  sky130_fd_sc_hd__fah_1 U25150 ( .A(n18585), .B(n18584), .CI(n18583), .COUT(
        n18600), .SUM(n18603) );
  sky130_fd_sc_hd__nand2_1 U25151 ( .A(n18588), .B(n18587), .Y(n18589) );
  sky130_fd_sc_hd__fah_1 U25152 ( .A(n18592), .B(n18591), .CI(n18590), .COUT(
        n18809), .SUM(n18286) );
  sky130_fd_sc_hd__xnor2_1 U25153 ( .A(n18600), .B(n18599), .Y(n18601) );
  sky130_fd_sc_hd__xnor2_1 U25154 ( .A(n18607), .B(n18606), .Y(n18814) );
  sky130_fd_sc_hd__o21ai_1 U25155 ( .A1(n18610), .A2(n18609), .B1(n18608), .Y(
        n18612) );
  sky130_fd_sc_hd__nand2_1 U25156 ( .A(n18610), .B(n18609), .Y(n18611) );
  sky130_fd_sc_hd__nand2_1 U25157 ( .A(n18612), .B(n18611), .Y(n18812) );
  sky130_fd_sc_hd__fa_1 U25158 ( .A(n18617), .B(n18616), .CIN(n18615), .COUT(
        n18644), .SUM(n18647) );
  sky130_fd_sc_hd__a22oi_1 U25159 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[28]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[12]), .Y(n18618) );
  sky130_fd_sc_hd__nand2_1 U25160 ( .A(n22071), .B(n18618), .Y(n18641) );
  sky130_fd_sc_hd__xnor2_1 U25161 ( .A(n22052), .B(n22685), .Y(n18621) );
  sky130_fd_sc_hd__xnor2_1 U25162 ( .A(n18651), .B(n22685), .Y(n18715) );
  sky130_fd_sc_hd__o22ai_1 U25163 ( .A1(n18619), .A2(n18621), .B1(n18715), 
        .B2(n18713), .Y(n18635) );
  sky130_fd_sc_hd__xnor2_1 U25164 ( .A(n18673), .B(n22051), .Y(n18620) );
  sky130_fd_sc_hd__a21o_1 U25165 ( .A1(n18713), .A2(n18716), .B1(n18621), .X(
        n18633) );
  sky130_fd_sc_hd__xnor2_1 U25166 ( .A(n18687), .B(n18720), .Y(n18749) );
  sky130_fd_sc_hd__o22ai_1 U25167 ( .A1(n18750), .A2(n18622), .B1(n18749), 
        .B2(n18747), .Y(n18638) );
  sky130_fd_sc_hd__xnor2_1 U25168 ( .A(n18685), .B(n22487), .Y(n18631) );
  sky130_fd_sc_hd__a22oi_1 U25169 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[27]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[11]), .Y(n18624) );
  sky130_fd_sc_hd__nand2_1 U25170 ( .A(n22071), .B(n18624), .Y(n18636) );
  sky130_fd_sc_hd__fa_1 U25171 ( .A(n18627), .B(n18626), .CIN(n18625), .COUT(
        n18642), .SUM(n18645) );
  sky130_fd_sc_hd__fah_1 U25172 ( .A(n18630), .B(n18629), .CI(n18628), .COUT(
        n18625), .SUM(n18779) );
  sky130_fd_sc_hd__xnor2_1 U25173 ( .A(n18673), .B(n22487), .Y(n18718) );
  sky130_fd_sc_hd__xnor2_1 U25174 ( .A(n18661), .B(n22051), .Y(n18632) );
  sky130_fd_sc_hd__fah_1 U25175 ( .A(n18638), .B(n18637), .CI(n18636), .COUT(
        n18639), .SUM(n18771) );
  sky130_fd_sc_hd__fa_1 U25176 ( .A(n18641), .B(n18640), .CIN(n18639), .COUT(
        n18646), .SUM(n18777) );
  sky130_fd_sc_hd__nor2_1 U25177 ( .A(n18849), .B(n18850), .Y(n21491) );
  sky130_fd_sc_hd__fa_1 U25178 ( .A(n18644), .B(n18643), .CIN(n18642), .COUT(
        n17384), .SUM(n18851) );
  sky130_fd_sc_hd__nand2_1 U25179 ( .A(n21868), .B(n21490), .Y(n22180) );
  sky130_fd_sc_hd__xnor2_1 U25180 ( .A(n18687), .B(n18656), .Y(n18652) );
  sky130_fd_sc_hd__o22ai_1 U25181 ( .A1(n18711), .A2(n18652), .B1(n18648), 
        .B2(n18712), .Y(n18700) );
  sky130_fd_sc_hd__xnor2_1 U25182 ( .A(n18649), .B(n22051), .Y(n18650) );
  sky130_fd_sc_hd__xnor2_1 U25183 ( .A(n22052), .B(n22029), .Y(n18659) );
  sky130_fd_sc_hd__xnor2_1 U25184 ( .A(n18651), .B(n18656), .Y(n18657) );
  sky130_fd_sc_hd__o22ai_1 U25185 ( .A1(n18711), .A2(n18657), .B1(n18652), 
        .B2(n18712), .Y(n18697) );
  sky130_fd_sc_hd__xnor2_1 U25186 ( .A(n18721), .B(n22685), .Y(n18688) );
  sky130_fd_sc_hd__xnor2_1 U25187 ( .A(n18685), .B(n22685), .Y(n18664) );
  sky130_fd_sc_hd__xnor2_1 U25188 ( .A(n18708), .B(n22487), .Y(n18653) );
  sky130_fd_sc_hd__xnor2_1 U25189 ( .A(n18654), .B(n22487), .Y(n18666) );
  sky130_fd_sc_hd__xnor2_1 U25190 ( .A(n18661), .B(n22487), .Y(n18717) );
  sky130_fd_sc_hd__xnor2_1 U25191 ( .A(n18654), .B(n22051), .Y(n18655) );
  sky130_fd_sc_hd__xnor2_1 U25192 ( .A(n22052), .B(n18656), .Y(n18710) );
  sky130_fd_sc_hd__xnor2_1 U25193 ( .A(n18661), .B(n18672), .Y(n18674) );
  sky130_fd_sc_hd__o22ai_1 U25194 ( .A1(n18750), .A2(n18674), .B1(n18662), 
        .B2(n18747), .Y(n18694) );
  sky130_fd_sc_hd__o22ai_1 U25195 ( .A1(n18716), .A2(n18664), .B1(n18663), 
        .B2(n18713), .Y(n18693) );
  sky130_fd_sc_hd__xnor2_1 U25196 ( .A(n18667), .B(n22051), .Y(n18668) );
  sky130_fd_sc_hd__fah_1 U25197 ( .A(n18671), .B(n18670), .CI(n18669), .COUT(
        n18738), .SUM(n18795) );
  sky130_fd_sc_hd__xnor2_1 U25198 ( .A(n18673), .B(n18672), .Y(n18686) );
  sky130_fd_sc_hd__o22ai_1 U25199 ( .A1(n18750), .A2(n18686), .B1(n18674), 
        .B2(n18747), .Y(n18692) );
  sky130_fd_sc_hd__a22oi_1 U25200 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[23]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[7]), .Y(n18675) );
  sky130_fd_sc_hd__nand2_1 U25201 ( .A(n22071), .B(n18675), .Y(n18691) );
  sky130_fd_sc_hd__a22oi_1 U25202 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[22]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[6]), .Y(n18678) );
  sky130_fd_sc_hd__nand2_1 U25203 ( .A(n22071), .B(n18678), .Y(n18737) );
  sky130_fd_sc_hd__xnor2_1 U25204 ( .A(n18685), .B(n18720), .Y(n18722) );
  sky130_fd_sc_hd__o22ai_1 U25205 ( .A1(n18750), .A2(n18722), .B1(n18686), 
        .B2(n18747), .Y(n18707) );
  sky130_fd_sc_hd__xnor2_1 U25206 ( .A(n18687), .B(n22685), .Y(n18714) );
  sky130_fd_sc_hd__o22ai_1 U25207 ( .A1(n18716), .A2(n18714), .B1(n18688), 
        .B2(n18713), .Y(n18706) );
  sky130_fd_sc_hd__a22oi_1 U25208 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[24]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[8]), .Y(n18689) );
  sky130_fd_sc_hd__nand2_1 U25209 ( .A(n22071), .B(n18689), .Y(n18705) );
  sky130_fd_sc_hd__fah_1 U25210 ( .A(n18692), .B(n18691), .CI(n18690), .COUT(
        n18727), .SUM(n18742) );
  sky130_fd_sc_hd__fah_1 U25211 ( .A(n18695), .B(n18694), .CI(n18693), .COUT(
        n18731), .SUM(n18740) );
  sky130_fd_sc_hd__fah_1 U25212 ( .A(n18700), .B(n18699), .CI(n18698), .COUT(
        n18725), .SUM(n18729) );
  sky130_fd_sc_hd__a22oi_1 U25213 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[25]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[9]), .Y(n18701) );
  sky130_fd_sc_hd__nand2_1 U25214 ( .A(n22071), .B(n18701), .Y(n18767) );
  sky130_fd_sc_hd__xnor2_1 U25215 ( .A(n18708), .B(n22051), .Y(n18709) );
  sky130_fd_sc_hd__a21o_1 U25216 ( .A1(n18712), .A2(n18711), .B1(n18710), .X(
        n18753) );
  sky130_fd_sc_hd__o22ai_1 U25217 ( .A1(n18716), .A2(n18715), .B1(n18714), 
        .B2(n18713), .Y(n18761) );
  sky130_fd_sc_hd__xnor2_1 U25218 ( .A(n18721), .B(n18720), .Y(n18748) );
  sky130_fd_sc_hd__o22ai_1 U25219 ( .A1(n18750), .A2(n18748), .B1(n18722), 
        .B2(n18747), .Y(n18759) );
  sky130_fd_sc_hd__fah_1 U25220 ( .A(n18734), .B(n18733), .CI(n18732), .COUT(
        n18799), .SUM(n18801) );
  sky130_fd_sc_hd__o22ai_1 U25221 ( .A1(n18750), .A2(n18749), .B1(n18748), 
        .B2(n18747), .Y(n18770) );
  sky130_fd_sc_hd__a22oi_1 U25222 ( .A1(n26862), .A2(
        j202_soc_core_j22_cpu_ml_mach[26]), .B1(n18751), .B2(
        j202_soc_core_j22_cpu_ml_mach[10]), .Y(n18752) );
  sky130_fd_sc_hd__nand2_1 U25223 ( .A(n22071), .B(n18752), .Y(n18769) );
  sky130_fd_sc_hd__fa_1 U25224 ( .A(n18761), .B(n18760), .CIN(n18759), .COUT(
        n18776), .SUM(n18757) );
  sky130_fd_sc_hd__fa_1 U25225 ( .A(n18764), .B(n18763), .CIN(n18762), .COUT(
        n18773), .SUM(n18775) );
  sky130_fd_sc_hd__fah_1 U25226 ( .A(n18767), .B(n18766), .CI(n18765), .COUT(
        n18774), .SUM(n18785) );
  sky130_fd_sc_hd__fa_1 U25227 ( .A(n18770), .B(n18769), .CIN(n18768), .COUT(
        n18782), .SUM(n18788) );
  sky130_fd_sc_hd__fah_1 U25228 ( .A(n18776), .B(n18775), .CI(n18774), .COUT(
        n18780), .SUM(n18786) );
  sky130_fd_sc_hd__fah_1 U25229 ( .A(n18782), .B(n18781), .CI(n18780), .COUT(
        n18840), .SUM(n18838) );
  sky130_fd_sc_hd__nor2_1 U25230 ( .A(n18835), .B(n18836), .Y(n19470) );
  sky130_fd_sc_hd__nand2_1 U25232 ( .A(n18791), .B(n18790), .Y(n18792) );
  sky130_fd_sc_hd__nand2_1 U25233 ( .A(n18793), .B(n18792), .Y(n18827) );
  sky130_fd_sc_hd__fa_1 U25234 ( .A(n18796), .B(n18795), .CIN(n18794), .COUT(
        n18804), .SUM(n18790) );
  sky130_fd_sc_hd__inv_2 U25235 ( .A(n18807), .Y(n18902) );
  sky130_fd_sc_hd__nand2_2 U25236 ( .A(n12178), .B(n18902), .Y(n22905) );
  sky130_fd_sc_hd__inv_2 U25237 ( .A(n22471), .Y(n22617) );
  sky130_fd_sc_hd__nor2_1 U25238 ( .A(n22180), .B(n22617), .Y(n18856) );
  sky130_fd_sc_hd__nand2_1 U25239 ( .A(n18811), .B(n18810), .Y(n18873) );
  sky130_fd_sc_hd__nand2_1 U25240 ( .A(n18814), .B(n18813), .Y(n22748) );
  sky130_fd_sc_hd__o21ai_1 U25241 ( .A1(n22751), .A2(n22747), .B1(n22748), .Y(
        n18815) );
  sky130_fd_sc_hd__nand2_1 U25242 ( .A(n18818), .B(n18817), .Y(n21420) );
  sky130_fd_sc_hd__nand2_1 U25243 ( .A(n18822), .B(n18821), .Y(n21786) );
  sky130_fd_sc_hd__o21ai_1 U25244 ( .A1(n21792), .A2(n21785), .B1(n21786), .Y(
        n18823) );
  sky130_fd_sc_hd__o21a_4 U25245 ( .A1(n18826), .A2(n19247), .B1(n18825), .X(
        n21511) );
  sky130_fd_sc_hd__nand2_1 U25246 ( .A(n18828), .B(n18827), .Y(n21510) );
  sky130_fd_sc_hd__nand2_1 U25247 ( .A(n18830), .B(n18829), .Y(n18901) );
  sky130_fd_sc_hd__nand2_1 U25248 ( .A(n12207), .B(n18832), .Y(n22906) );
  sky130_fd_sc_hd__nand2_1 U25249 ( .A(n18834), .B(n18833), .Y(n22903) );
  sky130_fd_sc_hd__o21ai_1 U25250 ( .A1(n22906), .A2(n22902), .B1(n22903), .Y(
        n19228) );
  sky130_fd_sc_hd__nand2_1 U25251 ( .A(n18836), .B(n18835), .Y(n19468) );
  sky130_fd_sc_hd__nand2_1 U25252 ( .A(n18838), .B(n18837), .Y(n21446) );
  sky130_fd_sc_hd__nand2_1 U25253 ( .A(n18840), .B(n18839), .Y(n19466) );
  sky130_fd_sc_hd__a21oi_1 U25254 ( .A1(n18842), .A2(n12166), .B1(n18841), .Y(
        n18843) );
  sky130_fd_sc_hd__nand2_1 U25256 ( .A(n18850), .B(n18849), .Y(n21867) );
  sky130_fd_sc_hd__nand2_1 U25257 ( .A(n18852), .B(n18851), .Y(n21489) );
  sky130_fd_sc_hd__a21oi_2 U25258 ( .A1(n18854), .A2(n21490), .B1(n18853), .Y(
        n22182) );
  sky130_fd_sc_hd__o21ai_1 U25259 ( .A1(n22180), .A2(n22619), .B1(n22182), .Y(
        n18855) );
  sky130_fd_sc_hd__xnor2_2 U25260 ( .A(n18860), .B(n18859), .Y(n23242) );
  sky130_fd_sc_hd__a21oi_1 U25261 ( .A1(n22055), .A2(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[0]), .B1(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .Y(n18862) );
  sky130_fd_sc_hd__o21a_1 U25262 ( .A1(n12763), .A2(n18862), .B1(n18861), .X(
        n18866) );
  sky130_fd_sc_hd__nand3_1 U25263 ( .A(n18865), .B(n18864), .C(n18863), .Y(
        n18892) );
  sky130_fd_sc_hd__o211a_2 U25264 ( .A1(n18869), .A2(n18868), .B1(n18892), 
        .C1(n25824), .X(n18870) );
  sky130_fd_sc_hd__nand2b_1 U25265 ( .A_N(n22936), .B(n12763), .Y(n27271) );
  sky130_fd_sc_hd__nand2_1 U25266 ( .A(n18874), .B(n18873), .Y(n18876) );
  sky130_fd_sc_hd__xnor2_2 U25267 ( .A(n18876), .B(n18875), .Y(n26873) );
  sky130_fd_sc_hd__nand2_1 U25268 ( .A(n26873), .B(n24499), .Y(n18877) );
  sky130_fd_sc_hd__nand2_1 U25269 ( .A(n24138), .B(n26398), .Y(n18897) );
  sky130_fd_sc_hd__nand3_1 U25270 ( .A(n18879), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .C(n24282), .Y(n25338) );
  sky130_fd_sc_hd__nand2_1 U25271 ( .A(n22952), .B(n18882), .Y(n25826) );
  sky130_fd_sc_hd__nand2b_1 U25272 ( .A_N(n22925), .B(
        j202_soc_core_j22_cpu_ml_macl[15]), .Y(n24143) );
  sky130_fd_sc_hd__o2bb2ai_1 U25273 ( .B1(n25264), .B2(n25338), .A1_N(
        j202_soc_core_j22_cpu_ml_mach[15]), .A2_N(n22936), .Y(n24139) );
  sky130_fd_sc_hd__nand2_1 U25274 ( .A(n22923), .B(n18883), .Y(n24142) );
  sky130_fd_sc_hd__a21oi_1 U25275 ( .A1(n24139), .A2(n26398), .B1(n18884), .Y(
        n18885) );
  sky130_fd_sc_hd__nand2_1 U25276 ( .A(n24143), .B(n18885), .Y(n18895) );
  sky130_fd_sc_hd__a21oi_1 U25277 ( .A1(n18886), .A2(n21505), .B1(n18887), .Y(
        n18891) );
  sky130_fd_sc_hd__nand2_1 U25278 ( .A(n18889), .B(n18888), .Y(n18890) );
  sky130_fd_sc_hd__xor2_1 U25279 ( .A(n18891), .B(n18890), .X(n26871) );
  sky130_fd_sc_hd__nor2_4 U25280 ( .A(n26398), .B(n22028), .Y(n22927) );
  sky130_fd_sc_hd__nand2_1 U25281 ( .A(n26871), .B(n22927), .Y(n24159) );
  sky130_fd_sc_hd__nor2_1 U25282 ( .A(n18895), .B(n18894), .Y(n18896) );
  sky130_fd_sc_hd__nand2_1 U25283 ( .A(n18897), .B(n18896), .Y(n18900) );
  sky130_fd_sc_hd__nand2_1 U25284 ( .A(n18900), .B(n22929), .Y(n19075) );
  sky130_fd_sc_hd__inv_2 U25285 ( .A(n21511), .Y(n22661) );
  sky130_fd_sc_hd__nand2_1 U25286 ( .A(n18910), .B(n18909), .Y(n18913) );
  sky130_fd_sc_hd__o21ai_1 U25287 ( .A1(n21574), .A2(n22837), .B1(n21575), .Y(
        n18912) );
  sky130_fd_sc_hd__xnor2_1 U25288 ( .A(n18913), .B(n18912), .Y(n22032) );
  sky130_fd_sc_hd__nand2_1 U25289 ( .A(n22032), .B(n24499), .Y(n18918) );
  sky130_fd_sc_hd__nand2_1 U25290 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[7]), .Y(n18917) );
  sky130_fd_sc_hd__nand2_1 U25291 ( .A(n27721), .B(
        j202_soc_core_j22_cpu_memop_MEM__2_), .Y(n23298) );
  sky130_fd_sc_hd__nand2_1 U25292 ( .A(j202_soc_core_j22_cpu_memop_MEM__3_), 
        .B(j202_soc_core_j22_cpu_memop_MEM__1_), .Y(n19072) );
  sky130_fd_sc_hd__nor2_1 U25293 ( .A(n23298), .B(n18914), .Y(n23573) );
  sky130_fd_sc_hd__nand2b_1 U25294 ( .A_N(n23293), .B(n26802), .Y(n22456) );
  sky130_fd_sc_hd__nand3_1 U25295 ( .A(n18918), .B(n26318), .C(n18917), .Y(
        n22227) );
  sky130_fd_sc_hd__nand3_1 U25296 ( .A(n22228), .B(n22459), .C(n22227), .Y(
        n22507) );
  sky130_fd_sc_hd__nand2_1 U25297 ( .A(j202_soc_core_j22_cpu_ma_M_address[0]), 
        .B(j202_soc_core_j22_cpu_ma_M_address[1]), .Y(n19165) );
  sky130_fd_sc_hd__nor2_1 U25298 ( .A(n18920), .B(n19165), .Y(n18919) );
  sky130_fd_sc_hd__nor2_1 U25299 ( .A(j202_soc_core_j22_cpu_ma_M_address[1]), 
        .B(n18920), .Y(n18980) );
  sky130_fd_sc_hd__nand2_1 U25300 ( .A(n18980), .B(
        j202_soc_core_j22_cpu_ma_M_address[0]), .Y(n19163) );
  sky130_fd_sc_hd__nand3_1 U25301 ( .A(n12419), .B(n18922), .C(n18921), .Y(
        n18984) );
  sky130_fd_sc_hd__nand2_1 U25302 ( .A(n21631), .B(n21078), .Y(n21097) );
  sky130_fd_sc_hd__nand2_1 U25303 ( .A(n21244), .B(n21134), .Y(n18937) );
  sky130_fd_sc_hd__nor4_1 U25304 ( .A(n19271), .B(n21097), .C(n18924), .D(
        n18937), .Y(n18935) );
  sky130_fd_sc_hd__nand2_1 U25305 ( .A(n21190), .B(n21246), .Y(n21615) );
  sky130_fd_sc_hd__nor2_1 U25306 ( .A(n21615), .B(n18925), .Y(n18926) );
  sky130_fd_sc_hd__nand2_1 U25307 ( .A(n21184), .B(n17277), .Y(n21081) );
  sky130_fd_sc_hd__nand2_1 U25308 ( .A(n21221), .B(n21081), .Y(n21053) );
  sky130_fd_sc_hd__nand4_1 U25309 ( .A(n18926), .B(n21608), .C(n21256), .D(
        n21245), .Y(n18933) );
  sky130_fd_sc_hd__nand3_1 U25310 ( .A(n21246), .B(n20747), .C(n21613), .Y(
        n21108) );
  sky130_fd_sc_hd__nor2_1 U25311 ( .A(n21719), .B(n21097), .Y(n21682) );
  sky130_fd_sc_hd__nand3_1 U25312 ( .A(n21243), .B(n21082), .C(n21682), .Y(
        n18928) );
  sky130_fd_sc_hd__o21ai_1 U25313 ( .A1(n21108), .A2(n18928), .B1(n21288), .Y(
        n18931) );
  sky130_fd_sc_hd__nand2_1 U25314 ( .A(n21688), .B(n21613), .Y(n21177) );
  sky130_fd_sc_hd__nand4_1 U25315 ( .A(n21229), .B(n21606), .C(n21245), .D(
        n21219), .Y(n18929) );
  sky130_fd_sc_hd__o21ai_1 U25316 ( .A1(n21177), .A2(n18929), .B1(n21235), .Y(
        n18930) );
  sky130_fd_sc_hd__nand2_1 U25317 ( .A(n18931), .B(n18930), .Y(n18932) );
  sky130_fd_sc_hd__a21oi_1 U25318 ( .A1(n18933), .A2(n21636), .B1(n18932), .Y(
        n18934) );
  sky130_fd_sc_hd__o21ai_1 U25319 ( .A1(n21722), .A2(n18935), .B1(n18934), .Y(
        n18976) );
  sky130_fd_sc_hd__nand2_1 U25320 ( .A(n21245), .B(n21134), .Y(n21114) );
  sky130_fd_sc_hd__nor3_1 U25321 ( .A(n18936), .B(n21126), .C(n21114), .Y(
        n21181) );
  sky130_fd_sc_hd__nor2_1 U25322 ( .A(n21041), .B(n21102), .Y(n21220) );
  sky130_fd_sc_hd__nor2_1 U25323 ( .A(n21226), .B(n19257), .Y(n21077) );
  sky130_fd_sc_hd__nand3_1 U25324 ( .A(n21181), .B(n21220), .C(n21077), .Y(
        n18942) );
  sky130_fd_sc_hd__nand2_1 U25325 ( .A(n21648), .B(n21287), .Y(n21718) );
  sky130_fd_sc_hd__nand2b_1 U25326 ( .A_N(n20759), .B(n21253), .Y(n21247) );
  sky130_fd_sc_hd__nor2_1 U25327 ( .A(n21643), .B(n21046), .Y(n21049) );
  sky130_fd_sc_hd__nand3_1 U25328 ( .A(n21688), .B(n21049), .C(n19352), .Y(
        n21193) );
  sky130_fd_sc_hd__nor3_1 U25329 ( .A(n21718), .B(n21247), .C(n21193), .Y(
        n18940) );
  sky130_fd_sc_hd__nand4_1 U25330 ( .A(n21256), .B(n21688), .C(n21287), .D(
        n19286), .Y(n21224) );
  sky130_fd_sc_hd__nand4_1 U25331 ( .A(n21710), .B(n21084), .C(n21172), .D(
        n21246), .Y(n18938) );
  sky130_fd_sc_hd__nand3_1 U25332 ( .A(n12180), .B(n21632), .C(n21631), .Y(
        n21044) );
  sky130_fd_sc_hd__a21oi_1 U25335 ( .A1(n18942), .A2(n21235), .B1(n18941), .Y(
        n18974) );
  sky130_fd_sc_hd__nand2_1 U25336 ( .A(n21267), .B(n21606), .Y(n21104) );
  sky130_fd_sc_hd__nand3_1 U25337 ( .A(n21706), .B(n21253), .C(n21628), .Y(
        n20791) );
  sky130_fd_sc_hd__nor4_1 U25338 ( .A(n19388), .B(n19257), .C(n21104), .D(
        n20791), .Y(n18943) );
  sky130_fd_sc_hd__nand2_1 U25339 ( .A(n21689), .B(n18943), .Y(n21116) );
  sky130_fd_sc_hd__nand4_1 U25340 ( .A(n21648), .B(n21613), .C(n19382), .D(
        n21270), .Y(n18944) );
  sky130_fd_sc_hd__nor2_1 U25341 ( .A(n21053), .B(n18944), .Y(n21234) );
  sky130_fd_sc_hd__a21oi_1 U25342 ( .A1(n21185), .A2(n21628), .B1(n21709), .Y(
        n18945) );
  sky130_fd_sc_hd__nand2_1 U25343 ( .A(n20908), .B(n18945), .Y(n18949) );
  sky130_fd_sc_hd__a22oi_1 U25344 ( .A1(n21676), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[15]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[79]), .Y(n18948) );
  sky130_fd_sc_hd__nand2_1 U25345 ( .A(n21699), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[47]), .Y(n18947) );
  sky130_fd_sc_hd__nand2_1 U25346 ( .A(n21698), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[111]), .Y(n18946) );
  sky130_fd_sc_hd__nand4_1 U25347 ( .A(n18949), .B(n18948), .C(n18947), .D(
        n18946), .Y(n18955) );
  sky130_fd_sc_hd__nand2b_1 U25348 ( .A_N(n18951), .B(n13387), .Y(n21228) );
  sky130_fd_sc_hd__nand4_1 U25349 ( .A(n18952), .B(n21706), .C(n21228), .D(
        n21245), .Y(n18953) );
  sky130_fd_sc_hd__o2bb2ai_1 U25350 ( .B1(n21220), .B2(n19272), .A1_N(n18953), 
        .A2_N(n13275), .Y(n18954) );
  sky130_fd_sc_hd__nor2_1 U25351 ( .A(n18955), .B(n18954), .Y(n18957) );
  sky130_fd_sc_hd__nand2_1 U25352 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_duty[3]), .Y(n18956) );
  sky130_fd_sc_hd__o211ai_1 U25353 ( .A1(n18958), .A2(n21234), .B1(n18957), 
        .C1(n18956), .Y(n18959) );
  sky130_fd_sc_hd__a21oi_1 U25354 ( .A1(n21116), .A2(n21063), .B1(n18959), .Y(
        n18973) );
  sky130_fd_sc_hd__nand2_1 U25355 ( .A(n21228), .B(n21649), .Y(n21113) );
  sky130_fd_sc_hd__nand2_1 U25356 ( .A(n20736), .B(n21606), .Y(n19297) );
  sky130_fd_sc_hd__nand2_1 U25357 ( .A(n21685), .B(n21253), .Y(n21213) );
  sky130_fd_sc_hd__nand3_1 U25358 ( .A(n21079), .B(n21061), .C(n21287), .Y(
        n18960) );
  sky130_fd_sc_hd__nor3_1 U25359 ( .A(n21113), .B(n19297), .C(n18960), .Y(
        n18970) );
  sky130_fd_sc_hd__nand2_1 U25360 ( .A(n12180), .B(n21632), .Y(n21117) );
  sky130_fd_sc_hd__nand3_1 U25362 ( .A(n21267), .B(n21245), .C(n18961), .Y(
        n18962) );
  sky130_fd_sc_hd__nor2_1 U25363 ( .A(n19388), .B(n18962), .Y(n19294) );
  sky130_fd_sc_hd__nand4_1 U25364 ( .A(n19294), .B(n21243), .C(n21190), .D(
        n21253), .Y(n18965) );
  sky130_fd_sc_hd__nand2_1 U25365 ( .A(n21270), .B(n21613), .Y(n20777) );
  sky130_fd_sc_hd__nand2_1 U25366 ( .A(n21286), .B(n20772), .Y(n18966) );
  sky130_fd_sc_hd__nand2b_1 U25367 ( .A_N(n18966), .B(n21685), .Y(n21039) );
  sky130_fd_sc_hd__nor4b_1 U25368 ( .D_N(n21049), .A(n19351), .B(n21126), .C(
        n21039), .Y(n18963) );
  sky130_fd_sc_hd__nand3b_1 U25369 ( .A_N(n20777), .B(n21082), .C(n18963), .Y(
        n18964) );
  sky130_fd_sc_hd__a22oi_1 U25370 ( .A1(n18965), .A2(n21636), .B1(n18964), 
        .B2(n21251), .Y(n18969) );
  sky130_fd_sc_hd__nand3_1 U25371 ( .A(n21645), .B(n21632), .C(n21094), .Y(
        n19278) );
  sky130_fd_sc_hd__nand2_1 U25372 ( .A(n21244), .B(n20805), .Y(n19300) );
  sky130_fd_sc_hd__nor4_1 U25373 ( .A(n21615), .B(n19278), .C(n21247), .D(
        n19300), .Y(n18967) );
  sky130_fd_sc_hd__nand2b_1 U25374 ( .A_N(n18967), .B(n21235), .Y(n18968) );
  sky130_fd_sc_hd__o211ai_1 U25375 ( .A1(n18970), .A2(n21720), .B1(n18969), 
        .C1(n18968), .Y(n18971) );
  sky130_fd_sc_hd__nand2_1 U25376 ( .A(n18971), .B(n21697), .Y(n18972) );
  sky130_fd_sc_hd__o211ai_1 U25377 ( .A1(n18974), .A2(n21179), .B1(n18973), 
        .C1(n18972), .Y(n18975) );
  sky130_fd_sc_hd__a21oi_1 U25378 ( .A1(n18976), .A2(n21727), .B1(n18975), .Y(
        n18978) );
  sky130_fd_sc_hd__nand2_1 U25379 ( .A(n18978), .B(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n18977) );
  sky130_fd_sc_hd__nand2_1 U25380 ( .A(n18980), .B(n18979), .Y(n21915) );
  sky130_fd_sc_hd__nor2_1 U25381 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[0]), .B(
        n22999), .Y(n18986) );
  sky130_fd_sc_hd__nor2_1 U25382 ( .A(n18986), .B(n26539), .Y(n26314) );
  sky130_fd_sc_hd__nand2_1 U25383 ( .A(n23000), .B(n22999), .Y(n26312) );
  sky130_fd_sc_hd__nand3_1 U25384 ( .A(n26776), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .C(n27910), .Y(n23011) );
  sky130_fd_sc_hd__nand2_1 U25385 ( .A(n23011), .B(n23012), .Y(n24481) );
  sky130_fd_sc_hd__nand2b_1 U25386 ( .A_N(n26682), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n18988) );
  sky130_fd_sc_hd__mux2i_1 U25387 ( .A0(j202_soc_core_j22_cpu_exuop_EXU_[5]), 
        .A1(j202_soc_core_j22_cpu_exuop_EXU_[3]), .S(
        j202_soc_core_j22_cpu_exuop_EXU_[0]), .Y(n18987) );
  sky130_fd_sc_hd__nand2_1 U25388 ( .A(n26690), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[4]), .Y(n26780) );
  sky130_fd_sc_hd__nand3_1 U25389 ( .A(n12382), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[0]), .C(
        j202_soc_core_j22_cpu_exuop_EXU_[5]), .Y(n23927) );
  sky130_fd_sc_hd__nand2_1 U25390 ( .A(n26601), .B(n24785), .Y(n18989) );
  sky130_fd_sc_hd__nand2_1 U25391 ( .A(n18989), .B(n26407), .Y(n18990) );
  sky130_fd_sc_hd__nor2_1 U25392 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[0]), 
        .B(n12382), .Y(n26775) );
  sky130_fd_sc_hd__nand2_1 U25393 ( .A(n26775), .B(n26679), .Y(n19410) );
  sky130_fd_sc_hd__nor2_1 U25394 ( .A(n19410), .B(n24778), .Y(n23940) );
  sky130_fd_sc_hd__nand2_1 U25395 ( .A(n18991), .B(n24494), .Y(n19037) );
  sky130_fd_sc_hd__nand2_1 U25396 ( .A(n18995), .B(n18994), .Y(n18996) );
  sky130_fd_sc_hd__xor2_1 U25397 ( .A(n12789), .B(n18996), .X(n24742) );
  sky130_fd_sc_hd__nand2_1 U25398 ( .A(n24742), .B(n22927), .Y(n22224) );
  sky130_fd_sc_hd__inv_1 U25399 ( .A(n18998), .Y(n22586) );
  sky130_fd_sc_hd__nand2_1 U25400 ( .A(n18999), .B(n22585), .Y(n19000) );
  sky130_fd_sc_hd__xor2_1 U25401 ( .A(n22586), .B(n19000), .X(n23773) );
  sky130_fd_sc_hd__nand2_1 U25402 ( .A(n26603), .B(n26723), .Y(n19001) );
  sky130_fd_sc_hd__nand2_1 U25403 ( .A(n25229), .B(n19001), .Y(n19002) );
  sky130_fd_sc_hd__nand2_1 U25404 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[5]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[3]), .Y(n19025) );
  sky130_fd_sc_hd__nand2_1 U25405 ( .A(n19002), .B(n26747), .Y(n19005) );
  sky130_fd_sc_hd__nor2_1 U25406 ( .A(n26738), .B(n19004), .Y(n23047) );
  sky130_fd_sc_hd__nand2_1 U25407 ( .A(n19005), .B(n23047), .Y(n19006) );
  sky130_fd_sc_hd__nand2_1 U25408 ( .A(n19006), .B(n24785), .Y(n22722) );
  sky130_fd_sc_hd__nand3_1 U25409 ( .A(n26791), .B(n26893), .C(n27429), .Y(
        n19011) );
  sky130_fd_sc_hd__nand2_1 U25410 ( .A(n27455), .B(n19007), .Y(n19026) );
  sky130_fd_sc_hd__nand2b_1 U25411 ( .A_N(n19011), .B(n19027), .Y(n26418) );
  sky130_fd_sc_hd__nor2_1 U25412 ( .A(n19008), .B(n22925), .Y(n22222) );
  sky130_fd_sc_hd__nand2_1 U25413 ( .A(n22222), .B(n26329), .Y(n19010) );
  sky130_fd_sc_hd__nand2_1 U25414 ( .A(n25798), .B(n26790), .Y(n26635) );
  sky130_fd_sc_hd__nor2_1 U25415 ( .A(n27908), .B(n24778), .Y(n26326) );
  sky130_fd_sc_hd__nand2_1 U25416 ( .A(n27402), .B(n26729), .Y(n26634) );
  sky130_fd_sc_hd__nand3_1 U25417 ( .A(n26635), .B(n26326), .C(n26634), .Y(
        n19009) );
  sky130_fd_sc_hd__o211ai_1 U25418 ( .A1(n25788), .A2(n26418), .B1(n19010), 
        .C1(n19009), .Y(n19022) );
  sky130_fd_sc_hd__nor2_1 U25419 ( .A(n23927), .B(n27455), .Y(n23026) );
  sky130_fd_sc_hd__nand2b_1 U25420 ( .A_N(n19011), .B(n23026), .Y(n26419) );
  sky130_fd_sc_hd__nand2_1 U25421 ( .A(n26739), .B(n26727), .Y(n24784) );
  sky130_fd_sc_hd__nor2_1 U25422 ( .A(n24784), .B(n24778), .Y(n25415) );
  sky130_fd_sc_hd__nand2_1 U25423 ( .A(n26790), .B(n25308), .Y(n19016) );
  sky130_fd_sc_hd__nor2_1 U25424 ( .A(j202_soc_core_j22_cpu_macop_MAC_[0]), 
        .B(n25338), .Y(n22965) );
  sky130_fd_sc_hd__nor2_1 U25425 ( .A(n17718), .B(n21972), .Y(n22229) );
  sky130_fd_sc_hd__nor2_1 U25426 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[3]), 
        .B(n19013), .Y(n21548) );
  sky130_fd_sc_hd__nand2_1 U25427 ( .A(n24785), .B(n21548), .Y(n25159) );
  sky130_fd_sc_hd__a21oi_1 U25428 ( .A1(n22229), .A2(n26329), .B1(n26406), .Y(
        n19015) );
  sky130_fd_sc_hd__nor2_1 U25429 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[3]), 
        .B(n12382), .Y(n23020) );
  sky130_fd_sc_hd__nand2_1 U25430 ( .A(n24785), .B(n23020), .Y(n19184) );
  sky130_fd_sc_hd__nand2_1 U25431 ( .A(n26061), .B(n22731), .Y(n19014) );
  sky130_fd_sc_hd__nand3_1 U25432 ( .A(n19016), .B(n19015), .C(n19014), .Y(
        n19017) );
  sky130_fd_sc_hd__a21oi_1 U25433 ( .A1(n19018), .A2(n25415), .B1(n19017), .Y(
        n19020) );
  sky130_fd_sc_hd__nand2_1 U25434 ( .A(n25237), .B(n27429), .Y(n19024) );
  sky130_fd_sc_hd__nand2b_1 U25435 ( .A_N(n19026), .B(n19024), .Y(n26424) );
  sky130_fd_sc_hd__nand2_1 U25436 ( .A(n25063), .B(n26710), .Y(n19019) );
  sky130_fd_sc_hd__o211ai_1 U25437 ( .A1(n26577), .A2(n26419), .B1(n19020), 
        .C1(n19019), .Y(n19021) );
  sky130_fd_sc_hd__nor2_1 U25438 ( .A(n19022), .B(n19021), .Y(n19033) );
  sky130_fd_sc_hd__nand2_1 U25439 ( .A(n26723), .B(n26747), .Y(n23919) );
  sky130_fd_sc_hd__nor2_1 U25440 ( .A(n26603), .B(n23920), .Y(n26714) );
  sky130_fd_sc_hd__nand2_1 U25441 ( .A(n19023), .B(n26714), .Y(n23021) );
  sky130_fd_sc_hd__nor2_1 U25442 ( .A(n24778), .B(n23021), .Y(n26342) );
  sky130_fd_sc_hd__nand2_1 U25443 ( .A(n23026), .B(n19024), .Y(n26427) );
  sky130_fd_sc_hd__nor2_1 U25444 ( .A(n19025), .B(n26723), .Y(n23029) );
  sky130_fd_sc_hd__nand2_1 U25445 ( .A(n23029), .B(n25229), .Y(n23019) );
  sky130_fd_sc_hd__nor2_1 U25446 ( .A(n24778), .B(n23019), .Y(n26338) );
  sky130_fd_sc_hd__nand2_1 U25447 ( .A(n26338), .B(n27354), .Y(n19030) );
  sky130_fd_sc_hd__nand2_1 U25448 ( .A(n27429), .B(n27415), .Y(n23016) );
  sky130_fd_sc_hd__nand2_1 U25449 ( .A(n19028), .B(n19027), .Y(n22729) );
  sky130_fd_sc_hd__o211ai_1 U25450 ( .A1(n11145), .A2(n26427), .B1(n19030), 
        .C1(n19029), .Y(n19031) );
  sky130_fd_sc_hd__a21oi_1 U25451 ( .A1(n26342), .A2(n27399), .B1(n19031), .Y(
        n19032) );
  sky130_fd_sc_hd__o211ai_1 U25452 ( .A1(n26790), .A2(n22722), .B1(n19033), 
        .C1(n19032), .Y(n19034) );
  sky130_fd_sc_hd__a21oi_1 U25453 ( .A1(n23773), .A2(n26409), .B1(n19034), .Y(
        n19035) );
  sky130_fd_sc_hd__o21ai_1 U25454 ( .A1(n18916), .A2(n22224), .B1(n19035), .Y(
        n19036) );
  sky130_fd_sc_hd__a21oi_1 U25455 ( .A1(n19037), .A2(n26729), .B1(n19036), .Y(
        n19038) );
  sky130_fd_sc_hd__nand2_1 U25456 ( .A(n19039), .B(n19038), .Y(n24737) );
  sky130_fd_sc_hd__nand2_1 U25457 ( .A(n24737), .B(n22768), .Y(n22505) );
  sky130_fd_sc_hd__nand2_1 U25458 ( .A(n22507), .B(n22505), .Y(n19040) );
  sky130_fd_sc_hd__nand2_1 U25459 ( .A(n19041), .B(n22873), .Y(n19061) );
  sky130_fd_sc_hd__o22ai_1 U25460 ( .A1(n19043), .A2(n22856), .B1(n19042), 
        .B2(n22854), .Y(n19049) );
  sky130_fd_sc_hd__nand2_1 U25461 ( .A(n19046), .B(n19044), .Y(n22860) );
  sky130_fd_sc_hd__nand2_1 U25462 ( .A(n19046), .B(n19045), .Y(n22858) );
  sky130_fd_sc_hd__o22ai_1 U25463 ( .A1(n19078), .A2(n22860), .B1(n19047), 
        .B2(n22858), .Y(n19048) );
  sky130_fd_sc_hd__nor2_1 U25464 ( .A(n19049), .B(n19048), .Y(n19060) );
  sky130_fd_sc_hd__nor2_1 U25465 ( .A(n19054), .B(n19050), .Y(n22864) );
  sky130_fd_sc_hd__nand2_1 U25466 ( .A(n22864), .B(
        j202_soc_core_j22_cpu_rf_vbr[7]), .Y(n19058) );
  sky130_fd_sc_hd__nand2_1 U25467 ( .A(n19052), .B(n19051), .Y(n22033) );
  sky130_fd_sc_hd__nand2_1 U25468 ( .A(n22867), .B(
        j202_soc_core_j22_cpu_rf_tmp[7]), .Y(n19057) );
  sky130_fd_sc_hd__nand2_1 U25469 ( .A(n22865), .B(
        j202_soc_core_j22_cpu_rf_gpr[487]), .Y(n19056) );
  sky130_fd_sc_hd__nand2_1 U25470 ( .A(n22866), .B(
        j202_soc_core_j22_cpu_rf_gpr[7]), .Y(n19055) );
  sky130_fd_sc_hd__and4_1 U25471 ( .A(n19058), .B(n19057), .C(n19056), .D(
        n19055), .X(n19059) );
  sky130_fd_sc_hd__nand3_1 U25472 ( .A(n19061), .B(n19060), .C(n19059), .Y(
        n22226) );
  sky130_fd_sc_hd__nand3_1 U25473 ( .A(n24279), .B(n27268), .C(
        j202_soc_core_j22_cpu_memop_MEM__3_), .Y(n22545) );
  sky130_fd_sc_hd__nor2_1 U25474 ( .A(j202_soc_core_j22_cpu_memop_MEM__0_), 
        .B(n22545), .Y(n22824) );
  sky130_fd_sc_hd__nand2_1 U25475 ( .A(n22226), .B(n22824), .Y(n22503) );
  sky130_fd_sc_hd__nand2_1 U25476 ( .A(n19062), .B(n22873), .Y(n19070) );
  sky130_fd_sc_hd__o22ai_1 U25477 ( .A1(n19064), .A2(n22854), .B1(n19063), 
        .B2(n22860), .Y(n19065) );
  sky130_fd_sc_hd__a21oi_1 U25478 ( .A1(n22866), .A2(
        j202_soc_core_j22_cpu_rf_gpr[15]), .B1(n19065), .Y(n19069) );
  sky130_fd_sc_hd__a22oi_1 U25479 ( .A1(n21847), .A2(
        j202_soc_core_j22_cpu_rf_gbr[15]), .B1(n22864), .B2(
        j202_soc_core_j22_cpu_rf_vbr[15]), .Y(n19068) );
  sky130_fd_sc_hd__a2bb2oi_1 U25480 ( .B1(j202_soc_core_j22_cpu_rf_gpr[495]), 
        .B2(n22865), .A1_N(n19066), .A2_N(n22033), .Y(n19067) );
  sky130_fd_sc_hd__nand4_1 U25481 ( .A(n19070), .B(n19069), .C(n19068), .D(
        n19067), .Y(n22501) );
  sky130_fd_sc_hd__nor2_1 U25482 ( .A(n19072), .B(n19071), .Y(n22039) );
  sky130_fd_sc_hd__nand2_1 U25483 ( .A(n23574), .B(
        j202_soc_core_j22_cpu_memop_MEM__0_), .Y(n23296) );
  sky130_fd_sc_hd__nand2b_1 U25484 ( .A_N(n22039), .B(n23296), .Y(n22004) );
  sky130_fd_sc_hd__nand2_1 U25485 ( .A(n22501), .B(n22004), .Y(n19073) );
  sky130_fd_sc_hd__nand2_1 U25486 ( .A(j202_soc_core_qspi_wb_wdat[15]), .B(
        n29594), .Y(n28607) );
  sky130_fd_sc_hd__nand2_1 U25487 ( .A(n12727), .B(n22581), .Y(n19083) );
  sky130_fd_sc_hd__nor2_1 U25488 ( .A(n19077), .B(n21762), .Y(n22594) );
  sky130_fd_sc_hd__xnor2_1 U25489 ( .A(n19078), .B(n22594), .Y(n24738) );
  sky130_fd_sc_hd__nor2_1 U25490 ( .A(n23776), .B(n21584), .Y(n19080) );
  sky130_fd_sc_hd__o22ai_1 U25491 ( .A1(n23776), .A2(n13603), .B1(n25798), 
        .B2(n11143), .Y(n19079) );
  sky130_fd_sc_hd__a211oi_1 U25492 ( .A1(n23773), .A2(n12158), .B1(n19080), 
        .C1(n19079), .Y(n19082) );
  sky130_fd_sc_hd__nand2_1 U25493 ( .A(n22515), .B(n27402), .Y(n19081) );
  sky130_fd_sc_hd__nand3_1 U25494 ( .A(n19083), .B(n19082), .C(n19081), .Y(
        n29010) );
  sky130_fd_sc_hd__nand2_1 U25495 ( .A(n20099), .B(n20843), .Y(n20048) );
  sky130_fd_sc_hd__nand2_1 U25496 ( .A(n20384), .B(n20047), .Y(n19974) );
  sky130_fd_sc_hd__nand2_1 U25497 ( .A(n19969), .B(n19112), .Y(n20898) );
  sky130_fd_sc_hd__nand3_1 U25498 ( .A(n20202), .B(n20376), .C(n20326), .Y(
        n20838) );
  sky130_fd_sc_hd__nor4_1 U25499 ( .A(n20048), .B(n19974), .C(n20898), .D(
        n20838), .Y(n19084) );
  sky130_fd_sc_hd__nand2b_1 U25500 ( .A_N(n19084), .B(n13481), .Y(n19091) );
  sky130_fd_sc_hd__nor2_1 U25501 ( .A(n19832), .B(n19985), .Y(n20897) );
  sky130_fd_sc_hd__nand2_1 U25502 ( .A(n20897), .B(n20375), .Y(n20294) );
  sky130_fd_sc_hd__nand2_1 U25503 ( .A(n20919), .B(n20308), .Y(n20116) );
  sky130_fd_sc_hd__nor2_1 U25504 ( .A(n20116), .B(n20898), .Y(n19850) );
  sky130_fd_sc_hd__nand2b_1 U25505 ( .A_N(n19086), .B(n19085), .Y(n20386) );
  sky130_fd_sc_hd__nand2_1 U25506 ( .A(n20298), .B(n20386), .Y(n19113) );
  sky130_fd_sc_hd__nand4_1 U25507 ( .A(n19850), .B(n19970), .C(n20326), .D(
        n20118), .Y(n19087) );
  sky130_fd_sc_hd__o21ai_1 U25508 ( .A1(n20115), .A2(n19087), .B1(n20908), .Y(
        n19090) );
  sky130_fd_sc_hd__nand2_1 U25509 ( .A(n20074), .B(n20008), .Y(n20865) );
  sky130_fd_sc_hd__nand3_1 U25510 ( .A(n20891), .B(n19088), .C(n20298), .Y(
        n20112) );
  sky130_fd_sc_hd__nand2_1 U25511 ( .A(n20112), .B(n21727), .Y(n19089) );
  sky130_fd_sc_hd__nand3_1 U25512 ( .A(n19091), .B(n19090), .C(n19089), .Y(
        n19092) );
  sky130_fd_sc_hd__nand2_1 U25513 ( .A(n19092), .B(n20912), .Y(n19151) );
  sky130_fd_sc_hd__nand2_1 U25514 ( .A(n21699), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[42]), .Y(n19145) );
  sky130_fd_sc_hd__nand2_1 U25515 ( .A(n19145), .B(n21677), .Y(n19096) );
  sky130_fd_sc_hd__nand2_1 U25516 ( .A(n21666), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[74]), .Y(n19095) );
  sky130_fd_sc_hd__nand2_1 U25517 ( .A(n21698), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[106]), .Y(n19094) );
  sky130_fd_sc_hd__nand2_1 U25518 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[10]), .Y(n19093) );
  sky130_fd_sc_hd__nand3_1 U25519 ( .A(n19095), .B(n19094), .C(n19093), .Y(
        n19146) );
  sky130_fd_sc_hd__nor2_1 U25520 ( .A(n19096), .B(n19146), .Y(n19100) );
  sky130_fd_sc_hd__nor4_1 U25521 ( .A(n20917), .B(n19097), .C(n20349), .D(
        n20104), .Y(n19098) );
  sky130_fd_sc_hd__a31oi_1 U25522 ( .A1(n19098), .A2(n20377), .A3(n20074), 
        .B1(n20925), .Y(n19099) );
  sky130_fd_sc_hd__nand2_1 U25523 ( .A(n19099), .B(n20908), .Y(n19149) );
  sky130_fd_sc_hd__nand2_1 U25524 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_period[10]), .Y(n19148) );
  sky130_fd_sc_hd__nand4_1 U25525 ( .A(n19151), .B(n19100), .C(n19149), .D(
        n19148), .Y(n19104) );
  sky130_fd_sc_hd__nand2_1 U25526 ( .A(n20376), .B(n20386), .Y(n20004) );
  sky130_fd_sc_hd__nor2_1 U25527 ( .A(n20180), .B(n19848), .Y(n20327) );
  sky130_fd_sc_hd__nand3_1 U25528 ( .A(n19891), .B(n20327), .C(n20842), .Y(
        n20311) );
  sky130_fd_sc_hd__nor4_1 U25529 ( .A(n20046), .B(n20904), .C(n17217), .D(
        n20311), .Y(n19102) );
  sky130_fd_sc_hd__nor2_1 U25530 ( .A(n20245), .B(n20871), .Y(n20385) );
  sky130_fd_sc_hd__nand4b_1 U25531 ( .A_N(n20105), .B(n20385), .C(n20199), .D(
        n20328), .Y(n20307) );
  sky130_fd_sc_hd__nand2_1 U25532 ( .A(n20919), .B(n20329), .Y(n20083) );
  sky130_fd_sc_hd__nor3_1 U25533 ( .A(n20307), .B(n20294), .C(n20083), .Y(
        n19101) );
  sky130_fd_sc_hd__o22a_1 U25534 ( .A1(n19856), .A2(n19102), .B1(n21179), .B2(
        n19101), .X(n19103) );
  sky130_fd_sc_hd__nor2_1 U25535 ( .A(n20925), .B(n19103), .Y(n19152) );
  sky130_fd_sc_hd__nor2_1 U25536 ( .A(n19104), .B(n19152), .Y(n19143) );
  sky130_fd_sc_hd__nand2_1 U25537 ( .A(n19951), .B(n20117), .Y(n20882) );
  sky130_fd_sc_hd__nor2_1 U25538 ( .A(n19834), .B(n19847), .Y(n20222) );
  sky130_fd_sc_hd__nand3_1 U25539 ( .A(n19891), .B(n20222), .C(n20327), .Y(
        n20353) );
  sky130_fd_sc_hd__nor3_1 U25540 ( .A(n20882), .B(n20353), .C(n20294), .Y(
        n19111) );
  sky130_fd_sc_hd__nand3_1 U25541 ( .A(n12165), .B(n20385), .C(n19971), .Y(
        n20365) );
  sky130_fd_sc_hd__nand2_1 U25542 ( .A(n20054), .B(n20386), .Y(n19997) );
  sky130_fd_sc_hd__a31oi_1 U25543 ( .A1(n19105), .A2(n20241), .A3(n20331), 
        .B1(n21179), .Y(n19109) );
  sky130_fd_sc_hd__nand2_1 U25544 ( .A(n19831), .B(n20080), .Y(n20195) );
  sky130_fd_sc_hd__nand2_1 U25545 ( .A(n20202), .B(n20885), .Y(n20121) );
  sky130_fd_sc_hd__nand2_1 U25546 ( .A(n19106), .B(n20170), .Y(n19107) );
  sky130_fd_sc_hd__nor3_1 U25547 ( .A(n20011), .B(n20180), .C(n19847), .Y(
        n20383) );
  sky130_fd_sc_hd__nand2_1 U25548 ( .A(n20383), .B(n20891), .Y(n20390) );
  sky130_fd_sc_hd__o21a_1 U25549 ( .A1(n19107), .A2(n20390), .B1(n20908), .X(
        n19108) );
  sky130_fd_sc_hd__nor2_1 U25550 ( .A(n19109), .B(n19108), .Y(n19110) );
  sky130_fd_sc_hd__o21ai_1 U25551 ( .A1(n19856), .A2(n19111), .B1(n19110), .Y(
        n19134) );
  sky130_fd_sc_hd__nand3_1 U25552 ( .A(n20384), .B(n20199), .C(n19112), .Y(
        n20190) );
  sky130_fd_sc_hd__nand3_1 U25553 ( .A(n19971), .B(n20306), .C(n20099), .Y(
        n20869) );
  sky130_fd_sc_hd__nor3_1 U25554 ( .A(n20190), .B(n20113), .C(n20869), .Y(
        n19132) );
  sky130_fd_sc_hd__nor2_1 U25555 ( .A(n19114), .B(n19113), .Y(n19116) );
  sky130_fd_sc_hd__nand3_1 U25556 ( .A(n20054), .B(n20843), .C(n20376), .Y(
        n20111) );
  sky130_fd_sc_hd__nor2_1 U25557 ( .A(n20916), .B(n20111), .Y(n19115) );
  sky130_fd_sc_hd__nand4_1 U25558 ( .A(n19850), .B(n19116), .C(n19995), .D(
        n19115), .Y(n19130) );
  sky130_fd_sc_hd__nand2_1 U25559 ( .A(n19891), .B(n20327), .Y(n19117) );
  sky130_fd_sc_hd__nor2_1 U25560 ( .A(n19117), .B(n20048), .Y(n19118) );
  sky130_fd_sc_hd__nand3_1 U25561 ( .A(n19118), .B(n20378), .C(n20358), .Y(
        n19123) );
  sky130_fd_sc_hd__o211ai_1 U25562 ( .A1(n19121), .A2(n19120), .B1(n19119), 
        .C1(n20385), .Y(n19122) );
  sky130_fd_sc_hd__o21ai_1 U25563 ( .A1(n19123), .A2(n19122), .B1(n20335), .Y(
        n19128) );
  sky130_fd_sc_hd__a31o_1 U25564 ( .A1(n19125), .A2(n20623), .A3(n19124), .B1(
        n20872), .X(n19126) );
  sky130_fd_sc_hd__nand2_1 U25565 ( .A(n20326), .B(n20047), .Y(n19998) );
  sky130_fd_sc_hd__nand2_1 U25567 ( .A(n19128), .B(n19127), .Y(n19129) );
  sky130_fd_sc_hd__a21oi_1 U25568 ( .A1(n19130), .A2(n20864), .B1(n19129), .Y(
        n19131) );
  sky130_fd_sc_hd__o21a_1 U25569 ( .A1(n19132), .A2(n20873), .B1(n19131), .X(
        n19133) );
  sky130_fd_sc_hd__a2bb2oi_1 U25570 ( .B1(n20864), .B2(n19134), .A1_N(n21124), 
        .A2_N(n19133), .Y(n19156) );
  sky130_fd_sc_hd__nand3_1 U25571 ( .A(n19135), .B(n20326), .C(n20843), .Y(
        n20379) );
  sky130_fd_sc_hd__nor2_1 U25572 ( .A(n20058), .B(n20379), .Y(n20315) );
  sky130_fd_sc_hd__nand2_1 U25573 ( .A(n20387), .B(n20305), .Y(n20057) );
  sky130_fd_sc_hd__nor4_1 U25574 ( .A(n20872), .B(n20871), .C(n20218), .D(
        n20057), .Y(n19136) );
  sky130_fd_sc_hd__nand2_1 U25575 ( .A(n20315), .B(n19136), .Y(n20078) );
  sky130_fd_sc_hd__nand2_1 U25576 ( .A(n20078), .B(n20908), .Y(n19141) );
  sky130_fd_sc_hd__nand3_1 U25577 ( .A(n20241), .B(n20008), .C(n20007), .Y(
        n19984) );
  sky130_fd_sc_hd__nor4_1 U25578 ( .A(n20312), .B(n20082), .C(n20116), .D(
        n19984), .Y(n19137) );
  sky130_fd_sc_hd__nor2_1 U25579 ( .A(n20918), .B(n19847), .Y(n20016) );
  sky130_fd_sc_hd__nand2_1 U25580 ( .A(n19137), .B(n20016), .Y(n19139) );
  sky130_fd_sc_hd__a21oi_1 U25581 ( .A1(n20850), .A2(n20222), .B1(n19856), .Y(
        n19138) );
  sky130_fd_sc_hd__a21oi_1 U25582 ( .A1(n19139), .A2(n13481), .B1(n19138), .Y(
        n19140) );
  sky130_fd_sc_hd__nand2_1 U25583 ( .A(n19141), .B(n19140), .Y(n19142) );
  sky130_fd_sc_hd__nand2_1 U25584 ( .A(n19142), .B(n20892), .Y(n19154) );
  sky130_fd_sc_hd__nand2_1 U25585 ( .A(j202_soc_core_memory0_ram_dout0[490]), 
        .B(n21771), .Y(n19157) );
  sky130_fd_sc_hd__nand2_1 U25586 ( .A(n19145), .B(n21738), .Y(n19147) );
  sky130_fd_sc_hd__nor2_1 U25587 ( .A(n19147), .B(n19146), .Y(n19150) );
  sky130_fd_sc_hd__nand4_1 U25588 ( .A(n19151), .B(n19150), .C(n19149), .D(
        n19148), .Y(n19153) );
  sky130_fd_sc_hd__nor2_1 U25589 ( .A(n19153), .B(n19152), .Y(n19155) );
  sky130_fd_sc_hd__nand4_1 U25590 ( .A(n19157), .B(n19156), .C(n19155), .D(
        n19154), .Y(n19158) );
  sky130_fd_sc_hd__nand2_1 U25591 ( .A(n21422), .B(n21420), .Y(n19162) );
  sky130_fd_sc_hd__o21ai_2 U25592 ( .A1(n12368), .A2(n22912), .B1(n19160), .Y(
        n19161) );
  sky130_fd_sc_hd__xnor2_2 U25593 ( .A(n19162), .B(n19161), .Y(n23237) );
  sky130_fd_sc_hd__nand2_1 U25594 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[2]), .Y(n25230) );
  sky130_fd_sc_hd__nand2_1 U25595 ( .A(n19163), .B(n26312), .Y(n21813) );
  sky130_fd_sc_hd__nand2_1 U25596 ( .A(n19164), .B(n21813), .Y(n19167) );
  sky130_fd_sc_hd__nand2_1 U25597 ( .A(n26314), .B(n19165), .Y(n22712) );
  sky130_fd_sc_hd__nand2_1 U25598 ( .A(n26606), .B(n26691), .Y(n19169) );
  sky130_fd_sc_hd__nand2_1 U25599 ( .A(n23920), .B(n26323), .Y(n19171) );
  sky130_fd_sc_hd__nand2_1 U25600 ( .A(n19171), .B(n25159), .Y(n19172) );
  sky130_fd_sc_hd__nand2_1 U25601 ( .A(n19177), .B(n19176), .Y(n19178) );
  sky130_fd_sc_hd__xnor2_1 U25602 ( .A(n19179), .B(n19178), .Y(n24805) );
  sky130_fd_sc_hd__nand2_1 U25603 ( .A(n24805), .B(n22927), .Y(n22312) );
  sky130_fd_sc_hd__nand2_1 U25604 ( .A(n26338), .B(n27383), .Y(n19183) );
  sky130_fd_sc_hd__a21oi_1 U25605 ( .A1(n27435), .A2(n25415), .B1(n23940), .Y(
        n19180) );
  sky130_fd_sc_hd__o22ai_1 U25606 ( .A1(n26423), .A2(n27435), .B1(n25229), 
        .B2(n19180), .Y(n19181) );
  sky130_fd_sc_hd__a21oi_1 U25607 ( .A1(n22734), .A2(n26603), .B1(n19181), .Y(
        n19182) );
  sky130_fd_sc_hd__o211ai_1 U25608 ( .A1(n25237), .A2(n22722), .B1(n19183), 
        .C1(n19182), .Y(n19192) );
  sky130_fd_sc_hd__nand2_1 U25609 ( .A(n22729), .B(n19184), .Y(n26341) );
  sky130_fd_sc_hd__a21oi_1 U25610 ( .A1(n26341), .A2(n26728), .B1(n19185), .Y(
        n19190) );
  sky130_fd_sc_hd__nand2_1 U25611 ( .A(n27435), .B(n23920), .Y(n26589) );
  sky130_fd_sc_hd__o21a_1 U25612 ( .A1(n27435), .A2(n23920), .B1(n26589), .X(
        n26638) );
  sky130_fd_sc_hd__o22ai_1 U25613 ( .A1(n21972), .A2(n25231), .B1(n19186), 
        .B2(n22925), .Y(n22313) );
  sky130_fd_sc_hd__a22oi_1 U25614 ( .A1(n26326), .A2(n26638), .B1(n22313), 
        .B2(n26329), .Y(n19189) );
  sky130_fd_sc_hd__o22a_1 U25615 ( .A1(n27007), .A2(n26418), .B1(n25789), .B2(
        n26419), .X(n19188) );
  sky130_fd_sc_hd__nand2_1 U25616 ( .A(n26342), .B(n27432), .Y(n19187) );
  sky130_fd_sc_hd__nand4_1 U25617 ( .A(n19190), .B(n19189), .C(n19188), .D(
        n19187), .Y(n19191) );
  sky130_fd_sc_hd__nor2_1 U25618 ( .A(n19192), .B(n19191), .Y(n19193) );
  sky130_fd_sc_hd__a21oi_1 U25620 ( .A1(n25235), .A2(n26409), .B1(n19194), .Y(
        n19195) );
  sky130_fd_sc_hd__inv_1 U25621 ( .A(n19199), .Y(n21429) );
  sky130_fd_sc_hd__nand2_1 U25622 ( .A(n21429), .B(n21428), .Y(n19201) );
  sky130_fd_sc_hd__xnor2_1 U25623 ( .A(n19201), .B(n19200), .Y(n22197) );
  sky130_fd_sc_hd__nand2_1 U25624 ( .A(n22197), .B(n24499), .Y(n22310) );
  sky130_fd_sc_hd__a22oi_1 U25625 ( .A1(n21847), .A2(
        j202_soc_core_j22_cpu_rf_gbr[2]), .B1(n22864), .B2(
        j202_soc_core_j22_cpu_rf_vbr[2]), .Y(n19208) );
  sky130_fd_sc_hd__o22a_1 U25626 ( .A1(n19203), .A2(n22860), .B1(n19202), .B2(
        n22854), .X(n19207) );
  sky130_fd_sc_hd__a2bb2oi_1 U25627 ( .B1(j202_soc_core_j22_cpu_rf_gpr[482]), 
        .B2(n22865), .A1_N(n19204), .A2_N(n22033), .Y(n19206) );
  sky130_fd_sc_hd__nand2_1 U25628 ( .A(n22866), .B(
        j202_soc_core_j22_cpu_rf_gpr[2]), .Y(n19205) );
  sky130_fd_sc_hd__nand4_1 U25629 ( .A(n19208), .B(n19207), .C(n19206), .D(
        n19205), .Y(n19209) );
  sky130_fd_sc_hd__a21oi_1 U25630 ( .A1(n19210), .A2(n22873), .B1(n19209), .Y(
        n22317) );
  sky130_fd_sc_hd__nand2b_1 U25631 ( .A_N(n22317), .B(n22824), .Y(n19211) );
  sky130_fd_sc_hd__nand2_1 U25632 ( .A(n19212), .B(n22873), .Y(n19220) );
  sky130_fd_sc_hd__o22ai_1 U25633 ( .A1(n19214), .A2(n22854), .B1(n19213), 
        .B2(n22860), .Y(n19215) );
  sky130_fd_sc_hd__a21oi_1 U25634 ( .A1(j202_soc_core_j22_cpu_rf_gpr[10]), 
        .A2(n22866), .B1(n19215), .Y(n19219) );
  sky130_fd_sc_hd__a22oi_1 U25635 ( .A1(n21847), .A2(
        j202_soc_core_j22_cpu_rf_gbr[10]), .B1(n22864), .B2(
        j202_soc_core_j22_cpu_rf_vbr[10]), .Y(n19218) );
  sky130_fd_sc_hd__a2bb2oi_1 U25636 ( .B1(j202_soc_core_j22_cpu_rf_gpr[490]), 
        .B2(n22865), .A1_N(n19216), .A2_N(n22033), .Y(n19217) );
  sky130_fd_sc_hd__nand4_1 U25637 ( .A(n19220), .B(n19219), .C(n19218), .D(
        n19217), .Y(n22382) );
  sky130_fd_sc_hd__nand2_1 U25638 ( .A(n22382), .B(n22004), .Y(n19245) );
  sky130_fd_sc_hd__nand2_1 U25639 ( .A(n21441), .B(n19222), .Y(n19225) );
  sky130_fd_sc_hd__nand2_1 U25641 ( .A(n22410), .B(n24499), .Y(n19236) );
  sky130_fd_sc_hd__a22oi_1 U25642 ( .A1(n12708), .A2(n27187), .B1(n22936), 
        .B2(j202_soc_core_j22_cpu_ml_mach[10]), .Y(n19235) );
  sky130_fd_sc_hd__nand2_1 U25643 ( .A(n19236), .B(n19235), .Y(n25027) );
  sky130_fd_sc_hd__nand2_1 U25644 ( .A(n19226), .B(n19468), .Y(n19234) );
  sky130_fd_sc_hd__nor2_1 U25645 ( .A(n19467), .B(n22905), .Y(n19230) );
  sky130_fd_sc_hd__nand2_1 U25646 ( .A(n22521), .B(n19230), .Y(n19232) );
  sky130_fd_sc_hd__o21ai_1 U25647 ( .A1(n19467), .A2(n22907), .B1(n19469), .Y(
        n19229) );
  sky130_fd_sc_hd__o21ai_2 U25648 ( .A1(n19232), .A2(n22912), .B1(n19231), .Y(
        n19233) );
  sky130_fd_sc_hd__a31oi_1 U25649 ( .A1(n19236), .A2(n26318), .A3(n19235), 
        .B1(n11713), .Y(n19237) );
  sky130_fd_sc_hd__nand2_1 U25650 ( .A(n22923), .B(n12708), .Y(n19238) );
  sky130_fd_sc_hd__o21a_1 U25651 ( .A1(n19239), .A2(n22925), .B1(n19238), .X(
        n25030) );
  sky130_fd_sc_hd__nand2_1 U25652 ( .A(n12208), .B(n19240), .Y(n19242) );
  sky130_fd_sc_hd__inv_1 U25653 ( .A(n19241), .Y(n21461) );
  sky130_fd_sc_hd__xnor2_1 U25654 ( .A(n19242), .B(n21461), .Y(n25049) );
  sky130_fd_sc_hd__nand2_1 U25655 ( .A(n25049), .B(n22927), .Y(n25045) );
  sky130_fd_sc_hd__nand2_1 U25656 ( .A(n19243), .B(n22929), .Y(n19244) );
  sky130_fd_sc_hd__nand2_1 U25657 ( .A(j202_soc_core_qspi_wb_wdat[10]), .B(
        n29594), .Y(n28609) );
  sky130_fd_sc_hd__inv_1 U25658 ( .A(n19246), .Y(n21790) );
  sky130_fd_sc_hd__nand2_2 U25659 ( .A(n23243), .B(n26863), .Y(n24367) );
  sky130_fd_sc_hd__nand2_1 U25660 ( .A(n19251), .B(n19250), .Y(n26311) );
  sky130_fd_sc_hd__nand2b_1 U25661 ( .A_N(n26311), .B(n22714), .Y(n19409) );
  sky130_fd_sc_hd__nand2_1 U25662 ( .A(j202_soc_core_memory0_ram_dout0[396]), 
        .B(n21597), .Y(n19253) );
  sky130_fd_sc_hd__nand2_1 U25663 ( .A(j202_soc_core_memory0_ram_dout0[76]), 
        .B(n21734), .Y(n19252) );
  sky130_fd_sc_hd__nand2_1 U25664 ( .A(j202_soc_core_memory0_ram_dout0[140]), 
        .B(n21592), .Y(n19256) );
  sky130_fd_sc_hd__nand2_1 U25665 ( .A(j202_soc_core_memory0_ram_dout0[204]), 
        .B(n21732), .Y(n19255) );
  sky130_fd_sc_hd__nand2_1 U25666 ( .A(j202_soc_core_memory0_ram_dout0[172]), 
        .B(n21590), .Y(n19254) );
  sky130_fd_sc_hd__nor3_1 U25667 ( .A(n21620), .B(n21201), .C(n19297), .Y(
        n19264) );
  sky130_fd_sc_hd__nor2_1 U25668 ( .A(n19257), .B(n19339), .Y(n20741) );
  sky130_fd_sc_hd__nand2_1 U25669 ( .A(n21081), .B(n21688), .Y(n20810) );
  sky130_fd_sc_hd__nor2_1 U25670 ( .A(n21620), .B(n21201), .Y(n19258) );
  sky130_fd_sc_hd__nand3_1 U25671 ( .A(n21614), .B(n19258), .C(n21094), .Y(
        n19259) );
  sky130_fd_sc_hd__nand3_1 U25673 ( .A(n21632), .B(n21287), .C(n19295), .Y(
        n19260) );
  sky130_fd_sc_hd__o21ai_0 U25674 ( .A1(n19260), .A2(n21617), .B1(n21636), .Y(
        n19261) );
  sky130_fd_sc_hd__o211ai_1 U25675 ( .A1(n21191), .A2(n21705), .B1(n19262), 
        .C1(n19261), .Y(n19263) );
  sky130_fd_sc_hd__o21bai_1 U25676 ( .A1(n21720), .A2(n19264), .B1_N(n19263), 
        .Y(n19265) );
  sky130_fd_sc_hd__nand2_1 U25677 ( .A(n19265), .B(n13481), .Y(n19319) );
  sky130_fd_sc_hd__nand2_1 U25678 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_duty[0]), .Y(n19267) );
  sky130_fd_sc_hd__nand2_1 U25679 ( .A(n21698), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[108]), .Y(n19266) );
  sky130_fd_sc_hd__nand2_1 U25680 ( .A(n19267), .B(n19266), .Y(n19307) );
  sky130_fd_sc_hd__nand3_1 U25681 ( .A(n20736), .B(n21267), .C(n21287), .Y(
        n21070) );
  sky130_fd_sc_hd__nand2_1 U25682 ( .A(n21070), .B(n21235), .Y(n21133) );
  sky130_fd_sc_hd__nand3_1 U25683 ( .A(n21256), .B(n21049), .C(n21206), .Y(
        n19268) );
  sky130_fd_sc_hd__nand2_1 U25684 ( .A(n19268), .B(n21636), .Y(n19269) );
  sky130_fd_sc_hd__nand2_1 U25685 ( .A(n21133), .B(n19269), .Y(n19270) );
  sky130_fd_sc_hd__nand2_1 U25686 ( .A(n19270), .B(n20908), .Y(n19315) );
  sky130_fd_sc_hd__nand2_1 U25687 ( .A(n21666), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[76]), .Y(n19310) );
  sky130_fd_sc_hd__nand2_1 U25688 ( .A(n21699), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[44]), .Y(n19309) );
  sky130_fd_sc_hd__nand2_1 U25689 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[12]), .Y(n19308) );
  sky130_fd_sc_hd__nand4_1 U25690 ( .A(n19310), .B(n19309), .C(n21677), .D(
        n19308), .Y(n19273) );
  sky130_fd_sc_hd__nor2_1 U25691 ( .A(n21620), .B(n19271), .Y(n21068) );
  sky130_fd_sc_hd__nor2_1 U25692 ( .A(n19272), .B(n21068), .Y(n19314) );
  sky130_fd_sc_hd__nor2_1 U25693 ( .A(n19273), .B(n19314), .Y(n19276) );
  sky130_fd_sc_hd__nand3_1 U25694 ( .A(n19274), .B(n21229), .C(n21679), .Y(
        n19275) );
  sky130_fd_sc_hd__nand2_1 U25695 ( .A(n19275), .B(n13275), .Y(n19311) );
  sky130_fd_sc_hd__nand3_1 U25696 ( .A(n19315), .B(n19276), .C(n19311), .Y(
        n19277) );
  sky130_fd_sc_hd__nor2_1 U25697 ( .A(n19307), .B(n19277), .Y(n19293) );
  sky130_fd_sc_hd__nand3_1 U25698 ( .A(n19280), .B(n19279), .C(n21685), .Y(
        n21188) );
  sky130_fd_sc_hd__nand2_1 U25699 ( .A(n21188), .B(n21288), .Y(n19291) );
  sky130_fd_sc_hd__nand2_1 U25700 ( .A(n21221), .B(n21613), .Y(n19299) );
  sky130_fd_sc_hd__nand2_1 U25701 ( .A(n21628), .B(n21688), .Y(n21093) );
  sky130_fd_sc_hd__nor2_1 U25702 ( .A(n19299), .B(n21093), .Y(n19281) );
  sky130_fd_sc_hd__nand3b_1 U25703 ( .A_N(n21039), .B(n21174), .C(n19281), .Y(
        n19282) );
  sky130_fd_sc_hd__nand2_1 U25704 ( .A(n19282), .B(n21251), .Y(n19290) );
  sky130_fd_sc_hd__nand3_1 U25705 ( .A(n21688), .B(n20751), .C(n19283), .Y(
        n21200) );
  sky130_fd_sc_hd__nand3_1 U25706 ( .A(n21614), .B(n21190), .C(n19284), .Y(
        n19285) );
  sky130_fd_sc_hd__nand4_1 U25708 ( .A(n21078), .B(n21220), .C(n21287), .D(
        n19286), .Y(n19287) );
  sky130_fd_sc_hd__nand2_1 U25709 ( .A(n19287), .B(n21636), .Y(n19288) );
  sky130_fd_sc_hd__nand4_1 U25710 ( .A(n19291), .B(n19290), .C(n19289), .D(
        n19288), .Y(n19292) );
  sky130_fd_sc_hd__nand2_1 U25711 ( .A(n19292), .B(n21727), .Y(n19318) );
  sky130_fd_sc_hd__nand3_1 U25712 ( .A(n19319), .B(n19293), .C(n19318), .Y(
        n19305) );
  sky130_fd_sc_hd__nand2_1 U25713 ( .A(n19294), .B(n21286), .Y(n21112) );
  sky130_fd_sc_hd__a21oi_1 U25714 ( .A1(n21270), .A2(n19295), .B1(n21722), .Y(
        n19296) );
  sky130_fd_sc_hd__a21o_1 U25715 ( .A1(n21112), .A2(n21636), .B1(n19296), .X(
        n19304) );
  sky130_fd_sc_hd__nor3_1 U25716 ( .A(n21715), .B(n21042), .C(n19297), .Y(
        n21129) );
  sky130_fd_sc_hd__nand2_1 U25717 ( .A(n21267), .B(n21628), .Y(n21704) );
  sky130_fd_sc_hd__nor4_1 U25718 ( .A(n21095), .B(n21704), .C(n19301), .D(
        n19300), .Y(n19302) );
  sky130_fd_sc_hd__o22ai_1 U25719 ( .A1(n21129), .A2(n21720), .B1(n19302), 
        .B2(n21705), .Y(n19303) );
  sky130_fd_sc_hd__o21a_1 U25720 ( .A1(n19304), .A2(n19303), .B1(n21697), .X(
        n19322) );
  sky130_fd_sc_hd__nor2_1 U25721 ( .A(n19305), .B(n19322), .Y(n19306) );
  sky130_fd_sc_hd__nand2_1 U25722 ( .A(j202_soc_core_memory0_ram_dout0[492]), 
        .B(n21771), .Y(n19325) );
  sky130_fd_sc_hd__nand4_1 U25723 ( .A(n19310), .B(n19309), .C(n21738), .D(
        n19308), .Y(n19313) );
  sky130_fd_sc_hd__nor3_1 U25724 ( .A(n19314), .B(n19313), .C(n19312), .Y(
        n19316) );
  sky130_fd_sc_hd__nand4_1 U25725 ( .A(n19318), .B(n19317), .C(n19316), .D(
        n19315), .Y(n19321) );
  sky130_fd_sc_hd__nor2_1 U25726 ( .A(n19321), .B(n19320), .Y(n19324) );
  sky130_fd_sc_hd__nand3_1 U25727 ( .A(n19325), .B(n19324), .C(n19323), .Y(
        n20973) );
  sky130_fd_sc_hd__nand2_1 U25728 ( .A(n20974), .B(n20973), .Y(n26313) );
  sky130_fd_sc_hd__nand2_1 U25729 ( .A(n26529), .B(n21813), .Y(n19407) );
  sky130_fd_sc_hd__a22oi_1 U25730 ( .A1(j202_soc_core_memory0_ram_dout0[452]), 
        .A2(j202_soc_core_memory0_ram_dout0_sel[14]), .B1(n21596), .B2(
        j202_soc_core_memory0_ram_dout0[356]), .Y(n19329) );
  sky130_fd_sc_hd__nand2_1 U25731 ( .A(j202_soc_core_memory0_ram_dout0[68]), 
        .B(n21734), .Y(n19326) );
  sky130_fd_sc_hd__a22oi_1 U25732 ( .A1(j202_soc_core_memory0_ram_dout0[36]), 
        .A2(n21604), .B1(n21732), .B2(j202_soc_core_memory0_ram_dout0[196]), 
        .Y(n19332) );
  sky130_fd_sc_hd__nand2_1 U25733 ( .A(n21648), .B(n21134), .Y(n21641) );
  sky130_fd_sc_hd__nor4_1 U25734 ( .A(n21207), .B(n21641), .C(n20734), .D(
        n21104), .Y(n19346) );
  sky130_fd_sc_hd__nor2_1 U25735 ( .A(n19350), .B(n19334), .Y(n21711) );
  sky130_fd_sc_hd__nand2_1 U25736 ( .A(n21270), .B(n21134), .Y(n21625) );
  sky130_fd_sc_hd__nor4b_1 U25737 ( .D_N(n19335), .A(n21215), .B(n19347), .C(
        n21625), .Y(n19344) );
  sky130_fd_sc_hd__nand2b_1 U25738 ( .A_N(n21177), .B(n21270), .Y(n21284) );
  sky130_fd_sc_hd__nor2_1 U25739 ( .A(n21113), .B(n21284), .Y(n20750) );
  sky130_fd_sc_hd__nor2_1 U25740 ( .A(n20759), .B(n21615), .Y(n19336) );
  sky130_fd_sc_hd__nand4_1 U25741 ( .A(n20750), .B(n20758), .C(n19336), .D(
        n21685), .Y(n19337) );
  sky130_fd_sc_hd__nand2_1 U25742 ( .A(n19337), .B(n21636), .Y(n19343) );
  sky130_fd_sc_hd__nand2_1 U25743 ( .A(n21190), .B(n21706), .Y(n21045) );
  sky130_fd_sc_hd__nor4_1 U25744 ( .A(n19338), .B(n21641), .C(n21045), .D(
        n21265), .Y(n19340) );
  sky130_fd_sc_hd__nor2_1 U25745 ( .A(n19339), .B(n21115), .Y(n20808) );
  sky130_fd_sc_hd__nand2_1 U25746 ( .A(n19340), .B(n20808), .Y(n19341) );
  sky130_fd_sc_hd__nand2_1 U25747 ( .A(n19341), .B(n21288), .Y(n19342) );
  sky130_fd_sc_hd__o211a_2 U25748 ( .A1(n19344), .A2(n21722), .B1(n19343), 
        .C1(n19342), .X(n19345) );
  sky130_fd_sc_hd__o21a_1 U25749 ( .A1(n21705), .A2(n19346), .B1(n19345), .X(
        n19402) );
  sky130_fd_sc_hd__nand2_1 U25750 ( .A(n21244), .B(n21648), .Y(n21657) );
  sky130_fd_sc_hd__nand2_1 U25751 ( .A(n21256), .B(n21246), .Y(n21684) );
  sky130_fd_sc_hd__nor4_1 U25752 ( .A(n19351), .B(n21657), .C(n19347), .D(
        n21684), .Y(n19348) );
  sky130_fd_sc_hd__nand2_1 U25753 ( .A(n19348), .B(n21079), .Y(n19349) );
  sky130_fd_sc_hd__nand2_1 U25754 ( .A(n19349), .B(n21288), .Y(n19365) );
  sky130_fd_sc_hd__nor2_1 U25755 ( .A(n19351), .B(n19350), .Y(n21630) );
  sky130_fd_sc_hd__nand3_1 U25756 ( .A(n20741), .B(n21173), .C(n21630), .Y(
        n19363) );
  sky130_fd_sc_hd__nand2_1 U25757 ( .A(n21287), .B(n19352), .Y(n21197) );
  sky130_fd_sc_hd__nor2_1 U25758 ( .A(n21641), .B(n21197), .Y(n21609) );
  sky130_fd_sc_hd__nand3_1 U25759 ( .A(n19353), .B(n21245), .C(n20736), .Y(
        n21654) );
  sky130_fd_sc_hd__nand3_1 U25760 ( .A(n19355), .B(n12137), .C(n19354), .Y(
        n21050) );
  sky130_fd_sc_hd__o211ai_1 U25761 ( .A1(n17277), .A2(n21050), .B1(n20739), 
        .C1(n21628), .Y(n19357) );
  sky130_fd_sc_hd__nor2_1 U25762 ( .A(n19357), .B(n19356), .Y(n19358) );
  sky130_fd_sc_hd__nand3_1 U25763 ( .A(n19360), .B(n19359), .C(n19358), .Y(
        n19361) );
  sky130_fd_sc_hd__o2bb2ai_1 U25764 ( .B1(n21609), .B2(n21709), .A1_N(n21251), 
        .A2_N(n19361), .Y(n19362) );
  sky130_fd_sc_hd__a21oi_1 U25765 ( .A1(n19363), .A2(n21235), .B1(n19362), .Y(
        n19364) );
  sky130_fd_sc_hd__nand2_1 U25766 ( .A(n19365), .B(n19364), .Y(n19400) );
  sky130_fd_sc_hd__nand2b_1 U25767 ( .A_N(n21093), .B(n21632), .Y(n21658) );
  sky130_fd_sc_hd__a21oi_1 U25768 ( .A1(n21253), .A2(n20752), .B1(n21709), .Y(
        n19368) );
  sky130_fd_sc_hd__a21oi_1 U25769 ( .A1(n21228), .A2(n19366), .B1(n21705), .Y(
        n19367) );
  sky130_fd_sc_hd__a22oi_1 U25771 ( .A1(n21666), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[68]), .B1(n21698), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[100]), .Y(n19374) );
  sky130_fd_sc_hd__a22oi_1 U25772 ( .A1(n21676), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[4]), .B1(n21699), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[36]), .Y(n19373) );
  sky130_fd_sc_hd__a22oi_1 U25773 ( .A1(n24376), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[20]), .B1(n21669), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[28]), .Y(n19370) );
  sky130_fd_sc_hd__a22oi_1 U25774 ( .A1(n21667), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[12]), .B1(n21668), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[4]), .Y(n19369) );
  sky130_fd_sc_hd__nand2_1 U25775 ( .A(n19370), .B(n19369), .Y(n19371) );
  sky130_fd_sc_hd__nand2_1 U25776 ( .A(n19371), .B(n21675), .Y(n19372) );
  sky130_fd_sc_hd__nand4_1 U25777 ( .A(n19375), .B(n19374), .C(n19373), .D(
        n19372), .Y(n19378) );
  sky130_fd_sc_hd__nand2b_1 U25779 ( .A_N(n19378), .B(n19377), .Y(n19379) );
  sky130_fd_sc_hd__a21oi_1 U25780 ( .A1(n20801), .A2(n21658), .B1(n19379), .Y(
        n19397) );
  sky130_fd_sc_hd__nand2_1 U25781 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_period[4]), .Y(n19396) );
  sky130_fd_sc_hd__nand2_1 U25782 ( .A(n21688), .B(n20772), .Y(n21043) );
  sky130_fd_sc_hd__nor2_1 U25783 ( .A(n21620), .B(n21095), .Y(n20803) );
  sky130_fd_sc_hd__nor2_1 U25784 ( .A(n21178), .B(n21046), .Y(n21651) );
  sky130_fd_sc_hd__nand4_1 U25785 ( .A(n20803), .B(n21651), .C(n21268), .D(
        n21267), .Y(n19384) );
  sky130_fd_sc_hd__a31oi_1 U25786 ( .A1(n21632), .A2(n19382), .A3(n21681), 
        .B1(n21722), .Y(n19383) );
  sky130_fd_sc_hd__a21o_1 U25787 ( .A1(n19384), .A2(n21235), .B1(n19383), .X(
        n19385) );
  sky130_fd_sc_hd__a21oi_1 U25788 ( .A1(n21288), .A2(n19386), .B1(n19385), .Y(
        n19392) );
  sky130_fd_sc_hd__nand4b_1 U25789 ( .A_N(n20759), .B(n21230), .C(n21221), .D(
        n21706), .Y(n21255) );
  sky130_fd_sc_hd__nand2_1 U25790 ( .A(n21255), .B(n21636), .Y(n19391) );
  sky130_fd_sc_hd__nand2_1 U25791 ( .A(n21287), .B(n20784), .Y(n21642) );
  sky130_fd_sc_hd__nor3_1 U25792 ( .A(n19388), .B(n19387), .C(n21642), .Y(
        n19389) );
  sky130_fd_sc_hd__nand2b_1 U25793 ( .A_N(n21654), .B(n19389), .Y(n19390) );
  sky130_fd_sc_hd__nand2_1 U25794 ( .A(n19390), .B(n21636), .Y(n20783) );
  sky130_fd_sc_hd__nand4_1 U25795 ( .A(n19393), .B(n19392), .C(n19391), .D(
        n20783), .Y(n19394) );
  sky130_fd_sc_hd__nand2_1 U25796 ( .A(n19394), .B(n21697), .Y(n19395) );
  sky130_fd_sc_hd__nand4_1 U25797 ( .A(n19398), .B(n19397), .C(n19396), .D(
        n19395), .Y(n19399) );
  sky130_fd_sc_hd__a21oi_1 U25798 ( .A1(n19400), .A2(n13481), .B1(n19399), .Y(
        n19401) );
  sky130_fd_sc_hd__o21a_1 U25799 ( .A1(n19856), .A2(n19402), .B1(n19401), .X(
        n21773) );
  sky130_fd_sc_hd__nor2_1 U25800 ( .A(n21771), .B(n19403), .Y(n21777) );
  sky130_fd_sc_hd__nor2_1 U25801 ( .A(n19404), .B(n21777), .Y(n19405) );
  sky130_fd_sc_hd__nand3_1 U25802 ( .A(n21770), .B(n21773), .C(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n21780) );
  sky130_fd_sc_hd__nand3_1 U25803 ( .A(n21781), .B(n19405), .C(n21780), .Y(
        n19406) );
  sky130_fd_sc_hd__nand2_1 U25804 ( .A(n19410), .B(n23011), .Y(n23022) );
  sky130_fd_sc_hd__nand2b_1 U25805 ( .A_N(n26791), .B(n25415), .Y(n19412) );
  sky130_fd_sc_hd__nand4_1 U25806 ( .A(n27421), .B(n26422), .C(n19413), .D(
        n19412), .Y(n19414) );
  sky130_fd_sc_hd__a21oi_1 U25807 ( .A1(n21531), .A2(n20287), .B1(n19417), .Y(
        n19422) );
  sky130_fd_sc_hd__nand2_1 U25808 ( .A(n19420), .B(n19419), .Y(n19421) );
  sky130_fd_sc_hd__xor2_1 U25809 ( .A(n19422), .B(n19421), .X(n24594) );
  sky130_fd_sc_hd__nand2_1 U25810 ( .A(n19425), .B(n19424), .Y(n19426) );
  sky130_fd_sc_hd__xnor2_1 U25811 ( .A(n19423), .B(n19426), .Y(n24586) );
  sky130_fd_sc_hd__nand2_1 U25812 ( .A(n24586), .B(n22927), .Y(n22265) );
  sky130_fd_sc_hd__o22ai_1 U25813 ( .A1(n25229), .A2(n26419), .B1(n11145), 
        .B2(n26418), .Y(n19427) );
  sky130_fd_sc_hd__a21oi_1 U25814 ( .A1(n26342), .A2(n27419), .B1(n19427), .Y(
        n19437) );
  sky130_fd_sc_hd__nor2_1 U25815 ( .A(n19428), .B(n22925), .Y(n22263) );
  sky130_fd_sc_hd__nand2_1 U25816 ( .A(n22263), .B(n26329), .Y(n19431) );
  sky130_fd_sc_hd__nand2_1 U25817 ( .A(n22923), .B(n10968), .Y(n22260) );
  sky130_fd_sc_hd__o2bb2ai_1 U25818 ( .B1(n18916), .B2(n22260), .A1_N(n22731), 
        .A2_N(n26717), .Y(n19429) );
  sky130_fd_sc_hd__a21oi_1 U25819 ( .A1(n26077), .A2(n26709), .B1(n19429), .Y(
        n19430) );
  sky130_fd_sc_hd__o211ai_1 U25820 ( .A1(n26417), .A2(n22729), .B1(n19431), 
        .C1(n19430), .Y(n19432) );
  sky130_fd_sc_hd__a21oi_1 U25821 ( .A1(n26338), .A2(n27372), .B1(n19432), .Y(
        n19436) );
  sky130_fd_sc_hd__xnor2_1 U25822 ( .A(n26712), .B(n26791), .Y(n26642) );
  sky130_fd_sc_hd__o22ai_1 U25823 ( .A1(n26713), .A2(n26427), .B1(n26577), 
        .B2(n26424), .Y(n19433) );
  sky130_fd_sc_hd__a21oi_1 U25824 ( .A1(n26326), .A2(n26642), .B1(n19433), .Y(
        n19435) );
  sky130_fd_sc_hd__mux2_2 U25825 ( .A0(n26423), .A1(n22722), .S(n27422), .X(
        n19434) );
  sky130_fd_sc_hd__nand4_1 U25826 ( .A(n19437), .B(n19436), .C(n19435), .D(
        n19434), .Y(n19438) );
  sky130_fd_sc_hd__o21bai_1 U25827 ( .A1(n18916), .A2(n22265), .B1_N(n19438), 
        .Y(n19439) );
  sky130_fd_sc_hd__a21oi_1 U25828 ( .A1(n24594), .A2(n26409), .B1(n19439), .Y(
        n19442) );
  sky130_fd_sc_hd__nand3_1 U25829 ( .A(n24481), .B(n23922), .C(n18916), .Y(
        n24792) );
  sky130_fd_sc_hd__o21ai_1 U25830 ( .A1(n24792), .A2(n26712), .B1(n25159), .Y(
        n19440) );
  sky130_fd_sc_hd__a21oi_1 U25831 ( .A1(n19200), .A2(n21802), .B1(n19444), .Y(
        n19447) );
  sky130_fd_sc_hd__nand2_1 U25832 ( .A(n19445), .B(n21803), .Y(n19446) );
  sky130_fd_sc_hd__xor2_1 U25833 ( .A(n19447), .B(n19446), .X(n22144) );
  sky130_fd_sc_hd__nand2_1 U25834 ( .A(n22144), .B(n26862), .Y(n22258) );
  sky130_fd_sc_hd__a22oi_1 U25835 ( .A1(n10968), .A2(n27187), .B1(n22936), 
        .B2(j202_soc_core_j22_cpu_ml_mach[4]), .Y(n22259) );
  sky130_fd_sc_hd__nand2_1 U25836 ( .A(n22258), .B(n22259), .Y(n24368) );
  sky130_fd_sc_hd__nand2_1 U25837 ( .A(n19449), .B(n22873), .Y(n19462) );
  sky130_fd_sc_hd__o22ai_1 U25838 ( .A1(n19451), .A2(n22856), .B1(n19450), 
        .B2(n22854), .Y(n19455) );
  sky130_fd_sc_hd__o22ai_1 U25839 ( .A1(n19453), .A2(n22860), .B1(n19452), 
        .B2(n22858), .Y(n19454) );
  sky130_fd_sc_hd__nor2_1 U25840 ( .A(n19455), .B(n19454), .Y(n19461) );
  sky130_fd_sc_hd__o22ai_1 U25841 ( .A1(n19457), .A2(n22034), .B1(n19456), 
        .B2(n22033), .Y(n19459) );
  sky130_fd_sc_hd__a22o_1 U25842 ( .A1(j202_soc_core_j22_cpu_rf_gpr[484]), 
        .A2(n22865), .B1(n22864), .B2(j202_soc_core_j22_cpu_rf_vbr[4]), .X(
        n19458) );
  sky130_fd_sc_hd__nor2_1 U25843 ( .A(n19459), .B(n19458), .Y(n19460) );
  sky130_fd_sc_hd__nand3_1 U25844 ( .A(n19462), .B(n19461), .C(n19460), .Y(
        n22268) );
  sky130_fd_sc_hd__inv_1 U25845 ( .A(n19463), .Y(n21893) );
  sky130_fd_sc_hd__nand2_1 U25846 ( .A(n19464), .B(n21892), .Y(n19465) );
  sky130_fd_sc_hd__xor2_1 U25847 ( .A(n21893), .B(n19465), .X(n24551) );
  sky130_fd_sc_hd__nand2_1 U25848 ( .A(n24551), .B(n22927), .Y(n26356) );
  sky130_fd_sc_hd__nand2b_1 U25849 ( .A_N(n22925), .B(
        j202_soc_core_j22_cpu_ml_macl[12]), .Y(n26328) );
  sky130_fd_sc_hd__nand2_1 U25850 ( .A(n26356), .B(n26328), .Y(n19493) );
  sky130_fd_sc_hd__nor2_1 U25851 ( .A(n17396), .B(n21972), .Y(n19489) );
  sky130_fd_sc_hd__nand2_1 U25852 ( .A(n26327), .B(n11713), .Y(n19492) );
  sky130_fd_sc_hd__nand2_1 U25853 ( .A(n12166), .B(n19466), .Y(n19479) );
  sky130_fd_sc_hd__nor2_1 U25854 ( .A(n19470), .B(n19467), .Y(n19472) );
  sky130_fd_sc_hd__nand2_1 U25855 ( .A(n21975), .B(n19472), .Y(n21448) );
  sky130_fd_sc_hd__nor2_1 U25856 ( .A(n19473), .B(n21448), .Y(n19475) );
  sky130_fd_sc_hd__a21oi_1 U25858 ( .A1(n21974), .A2(n19472), .B1(n19471), .Y(
        n21449) );
  sky130_fd_sc_hd__o21ai_1 U25859 ( .A1(n19473), .A2(n21449), .B1(n21446), .Y(
        n19474) );
  sky130_fd_sc_hd__xnor2_1 U25860 ( .A(n19479), .B(n19478), .Y(n23249) );
  sky130_fd_sc_hd__nand2_1 U25861 ( .A(n19480), .B(n21876), .Y(n19488) );
  sky130_fd_sc_hd__nand2_1 U25862 ( .A(n21874), .B(n19484), .Y(n19486) );
  sky130_fd_sc_hd__a21oi_1 U25863 ( .A1(n21881), .A2(n19484), .B1(n12578), .Y(
        n19485) );
  sky130_fd_sc_hd__xnor2_1 U25865 ( .A(n19488), .B(n19487), .Y(n22637) );
  sky130_fd_sc_hd__nand2_1 U25866 ( .A(n22637), .B(n26862), .Y(n26319) );
  sky130_fd_sc_hd__nand2_1 U25867 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[12]), .Y(n26317) );
  sky130_fd_sc_hd__nand2_1 U25868 ( .A(n26319), .B(n26317), .Y(n26322) );
  sky130_fd_sc_hd__a21oi_1 U25869 ( .A1(n26321), .A2(n26863), .B1(n26322), .Y(
        n23270) );
  sky130_fd_sc_hd__nor2_1 U25870 ( .A(n19489), .B(n19493), .Y(n19490) );
  sky130_fd_sc_hd__nand2_1 U25871 ( .A(n23270), .B(n19490), .Y(n19491) );
  sky130_fd_sc_hd__nand2_1 U25872 ( .A(n19494), .B(n22873), .Y(n19502) );
  sky130_fd_sc_hd__o22ai_1 U25873 ( .A1(n19496), .A2(n22860), .B1(n22854), 
        .B2(n19495), .Y(n19497) );
  sky130_fd_sc_hd__a21oi_1 U25874 ( .A1(n22866), .A2(
        j202_soc_core_j22_cpu_rf_gpr[12]), .B1(n19497), .Y(n19501) );
  sky130_fd_sc_hd__a22oi_1 U25875 ( .A1(n21847), .A2(
        j202_soc_core_j22_cpu_rf_gbr[12]), .B1(n22864), .B2(
        j202_soc_core_j22_cpu_rf_vbr[12]), .Y(n19500) );
  sky130_fd_sc_hd__a2bb2oi_1 U25876 ( .B1(j202_soc_core_j22_cpu_rf_gpr[492]), 
        .B2(n22865), .A1_N(n19498), .A2_N(n22033), .Y(n19499) );
  sky130_fd_sc_hd__nand4_1 U25877 ( .A(n19502), .B(n19501), .C(n19500), .D(
        n19499), .Y(n22651) );
  sky130_fd_sc_hd__nand2_1 U25878 ( .A(n22651), .B(n22004), .Y(n19503) );
  sky130_fd_sc_hd__nand2_1 U25879 ( .A(j202_soc_core_intc_core_00_in_intreq[7]), .B(j202_soc_core_intc_core_00_rg_itgt[7]), .Y(n19616) );
  sky130_fd_sc_hd__nand2_1 U25880 ( .A(j202_soc_core_intc_core_00_in_intreq[6]), .B(j202_soc_core_intc_core_00_rg_itgt[6]), .Y(n19617) );
  sky130_fd_sc_hd__nand2_1 U25881 ( .A(n19616), .B(n19617), .Y(n19631) );
  sky130_fd_sc_hd__nand2_1 U25882 ( .A(j202_soc_core_intc_core_00_in_intreq[4]), .B(j202_soc_core_intc_core_00_rg_itgt[4]), .Y(n19605) );
  sky130_fd_sc_hd__nand2_1 U25883 ( .A(j202_soc_core_intc_core_00_rg_itgt[5]), 
        .B(j202_soc_core_intc_core_00_in_intreq[5]), .Y(n19606) );
  sky130_fd_sc_hd__nand2_1 U25884 ( .A(n19605), .B(n19606), .Y(n19637) );
  sky130_fd_sc_hd__nor2_1 U25885 ( .A(n19631), .B(n19637), .Y(n19655) );
  sky130_fd_sc_hd__nand2_1 U25886 ( .A(j202_soc_core_intc_core_00_in_intreq[1]), .B(j202_soc_core_intc_core_00_rg_itgt[1]), .Y(n19583) );
  sky130_fd_sc_hd__nand2_1 U25887 ( .A(j202_soc_core_intc_core_00_rg_itgt[0]), 
        .B(j202_soc_core_intc_core_00_in_intreq[0]), .Y(n19582) );
  sky130_fd_sc_hd__nand2_1 U25888 ( .A(n19583), .B(n19582), .Y(n19597) );
  sky130_fd_sc_hd__nand2_1 U25889 ( .A(j202_soc_core_intc_core_00_in_intreq[2]), .B(j202_soc_core_intc_core_00_rg_itgt[2]), .Y(n19572) );
  sky130_fd_sc_hd__nand2_1 U25890 ( .A(j202_soc_core_intc_core_00_in_intreq[3]), .B(j202_soc_core_intc_core_00_rg_itgt[3]), .Y(n19575) );
  sky130_fd_sc_hd__nand2_1 U25891 ( .A(n19572), .B(n19575), .Y(n19595) );
  sky130_fd_sc_hd__nor2_1 U25892 ( .A(n19597), .B(n19595), .Y(n19661) );
  sky130_fd_sc_hd__nand2_1 U25893 ( .A(n19655), .B(n19661), .Y(n19798) );
  sky130_fd_sc_hd__nand2_1 U25894 ( .A(
        j202_soc_core_intc_core_00_in_intreq[10]), .B(
        j202_soc_core_intc_core_00_rg_itgt[10]), .Y(n19674) );
  sky130_fd_sc_hd__nand2_1 U25895 ( .A(
        j202_soc_core_intc_core_00_in_intreq[11]), .B(
        j202_soc_core_intc_core_00_rg_itgt[11]), .Y(n19671) );
  sky130_fd_sc_hd__nand2_1 U25896 ( .A(n19674), .B(n19671), .Y(n19697) );
  sky130_fd_sc_hd__nand2_1 U25897 ( .A(j202_soc_core_intc_core_00_rg_itgt[9]), 
        .B(j202_soc_core_intc_core_00_in_intreq[9]), .Y(n19682) );
  sky130_fd_sc_hd__nand2_1 U25898 ( .A(j202_soc_core_intc_core_00_rg_itgt[8]), 
        .B(j202_soc_core_intc_core_00_in_intreq[8]), .Y(n19681) );
  sky130_fd_sc_hd__nand2_1 U25899 ( .A(n19682), .B(n19681), .Y(n19695) );
  sky130_fd_sc_hd__nor2_1 U25900 ( .A(n19697), .B(n19695), .Y(n19765) );
  sky130_fd_sc_hd__nand2_1 U25901 ( .A(
        j202_soc_core_intc_core_00_in_intreq[15]), .B(
        j202_soc_core_intc_core_00_rg_itgt[15]), .Y(n19705) );
  sky130_fd_sc_hd__nand2_1 U25902 ( .A(
        j202_soc_core_intc_core_00_in_intreq[14]), .B(
        j202_soc_core_intc_core_00_rg_itgt[14]), .Y(n19704) );
  sky130_fd_sc_hd__nand2_1 U25903 ( .A(n19705), .B(n19704), .Y(n19733) );
  sky130_fd_sc_hd__nand2_1 U25904 ( .A(
        j202_soc_core_intc_core_00_in_intreq[12]), .B(
        j202_soc_core_intc_core_00_rg_itgt[12]), .Y(n19715) );
  sky130_fd_sc_hd__nand2_1 U25905 ( .A(
        j202_soc_core_intc_core_00_in_intreq[13]), .B(
        j202_soc_core_intc_core_00_rg_itgt[13]), .Y(n19714) );
  sky130_fd_sc_hd__nand2_1 U25906 ( .A(n19715), .B(n19714), .Y(n19727) );
  sky130_fd_sc_hd__nor2_1 U25907 ( .A(n19733), .B(n19727), .Y(n19762) );
  sky130_fd_sc_hd__nand2_1 U25908 ( .A(n19765), .B(n19762), .Y(n19795) );
  sky130_fd_sc_hd__nor2_1 U25909 ( .A(n19798), .B(n19795), .Y(n19828) );
  sky130_fd_sc_hd__nand2_1 U25910 ( .A(
        j202_soc_core_intc_core_00_in_intreq[18]), .B(
        j202_soc_core_intc_core_00_rg_itgt[18]), .Y(n19516) );
  sky130_fd_sc_hd__nand2_1 U25911 ( .A(
        j202_soc_core_intc_core_00_in_intreq[19]), .B(
        j202_soc_core_intc_core_00_rg_itgt[19]), .Y(n19517) );
  sky130_fd_sc_hd__nand2_1 U25912 ( .A(j202_soc_core_intc_core_00_rg_itgt[16]), 
        .B(j202_soc_core_intc_core_00_in_intreq[16]), .Y(n19509) );
  sky130_fd_sc_hd__nand2_1 U25913 ( .A(
        j202_soc_core_intc_core_00_in_intreq[17]), .B(
        j202_soc_core_intc_core_00_rg_itgt[17]), .Y(n19508) );
  sky130_fd_sc_hd__nand2_1 U25914 ( .A(n19509), .B(n19508), .Y(n19534) );
  sky130_fd_sc_hd__nand2_1 U25915 ( .A(n19529), .B(n19504), .Y(n19564) );
  sky130_fd_sc_hd__nor2_1 U25916 ( .A(n19562), .B(n19564), .Y(n19822) );
  sky130_fd_sc_hd__nand2_1 U25917 ( .A(n19828), .B(n19822), .Y(n25781) );
  sky130_fd_sc_hd__nor2_1 U25918 ( .A(n28590), .B(n25781), .Y(n29059) );
  sky130_fd_sc_hd__nand2_1 U25919 ( .A(n25781), .B(n29594), .Y(n24585) );
  sky130_fd_sc_hd__o22ai_1 U25921 ( .A1(j202_soc_core_intc_core_00_rg_ipr[68]), 
        .A2(n19505), .B1(j202_soc_core_intc_core_00_rg_ipr[69]), .B2(n27665), 
        .Y(n19506) );
  sky130_fd_sc_hd__a222oi_1 U25922 ( .A1(j202_soc_core_intc_core_00_rg_ipr[66]), .A2(n25521), .B1(j202_soc_core_intc_core_00_rg_ipr[66]), .B2(n19506), .C1(
        n25521), .C2(n19506), .Y(n19507) );
  sky130_fd_sc_hd__nand2_1 U25923 ( .A(n26846), .B(
        j202_soc_core_intc_core_00_rg_ipr[66]), .Y(n19512) );
  sky130_fd_sc_hd__o21ai_1 U25924 ( .A1(n25521), .A2(n26846), .B1(n19512), .Y(
        n19538) );
  sky130_fd_sc_hd__a22oi_1 U25925 ( .A1(j202_soc_core_intc_core_00_rg_ipr[73]), 
        .A2(n27805), .B1(j202_soc_core_intc_core_00_rg_ipr[72]), .B2(n26263), 
        .Y(n19514) );
  sky130_fd_sc_hd__o22ai_1 U25926 ( .A1(j202_soc_core_intc_core_00_rg_ipr[73]), 
        .A2(n27805), .B1(j202_soc_core_intc_core_00_rg_ipr[74]), .B2(n27705), 
        .Y(n19513) );
  sky130_fd_sc_hd__o22ai_1 U25927 ( .A1(j202_soc_core_intc_core_00_rg_ipr[78]), 
        .A2(n27283), .B1(n19514), .B2(n19513), .Y(n19515) );
  sky130_fd_sc_hd__a21oi_1 U25928 ( .A1(n19519), .A2(n19518), .B1(n19517), .Y(
        n26850) );
  sky130_fd_sc_hd__nand2_1 U25929 ( .A(n26850), .B(n27705), .Y(n19520) );
  sky130_fd_sc_hd__nand2_1 U25931 ( .A(n26846), .B(n19521), .Y(n19522) );
  sky130_fd_sc_hd__o21ai_1 U25932 ( .A1(j202_soc_core_intc_core_00_rg_ipr[68]), 
        .A2(n26846), .B1(n19522), .Y(n19545) );
  sky130_fd_sc_hd__nand2_1 U25933 ( .A(n26850), .B(n27805), .Y(n19523) );
  sky130_fd_sc_hd__o21ai_1 U25934 ( .A1(j202_soc_core_intc_core_00_rg_ipr[73]), 
        .A2(n26850), .B1(n19523), .Y(n19548) );
  sky130_fd_sc_hd__nand2_1 U25935 ( .A(n26846), .B(
        j202_soc_core_intc_core_00_rg_ipr[65]), .Y(n19524) );
  sky130_fd_sc_hd__o21ai_1 U25936 ( .A1(n26900), .A2(n26846), .B1(n19524), .Y(
        n19549) );
  sky130_fd_sc_hd__nand2_1 U25937 ( .A(n26850), .B(n26263), .Y(n19525) );
  sky130_fd_sc_hd__o21ai_1 U25938 ( .A1(j202_soc_core_intc_core_00_rg_ipr[72]), 
        .A2(n26850), .B1(n19525), .Y(n19544) );
  sky130_fd_sc_hd__o21ai_1 U25939 ( .A1(n19548), .A2(n19549), .B1(n19544), .Y(
        n19526) );
  sky130_fd_sc_hd__o2bb2ai_1 U25940 ( .B1(n19545), .B2(n19526), .A1_N(n19548), 
        .A2_N(n19549), .Y(n19527) );
  sky130_fd_sc_hd__maj3_1 U25941 ( .A(n19536), .B(n19538), .C(n19527), .X(
        n19531) );
  sky130_fd_sc_hd__nand2_1 U25942 ( .A(n26850), .B(n27509), .Y(n19528) );
  sky130_fd_sc_hd__o21ai_1 U25943 ( .A1(j202_soc_core_intc_core_00_rg_ipr[75]), 
        .A2(n26850), .B1(n19528), .Y(n19539) );
  sky130_fd_sc_hd__a21oi_1 U25944 ( .A1(n19531), .A2(n19539), .B1(n19529), .Y(
        n19533) );
  sky130_fd_sc_hd__nand2_1 U25945 ( .A(n26846), .B(
        j202_soc_core_intc_core_00_rg_ipr[67]), .Y(n19530) );
  sky130_fd_sc_hd__o21ai_1 U25947 ( .A1(n19539), .A2(n19531), .B1(n19540), .Y(
        n19532) );
  sky130_fd_sc_hd__nand2_1 U25948 ( .A(n19533), .B(n19532), .Y(n19535) );
  sky130_fd_sc_hd__nand2_1 U25949 ( .A(n26847), .B(n19536), .Y(n19537) );
  sky130_fd_sc_hd__o21ai_1 U25950 ( .A1(n19538), .A2(n26847), .B1(n19537), .Y(
        n19555) );
  sky130_fd_sc_hd__nor2_1 U25951 ( .A(n19541), .B(n26847), .Y(n19542) );
  sky130_fd_sc_hd__a21oi_1 U25952 ( .A1(n19543), .A2(n26847), .B1(n19542), .Y(
        n19817) );
  sky130_fd_sc_hd__nor2_1 U25953 ( .A(n19545), .B(n26847), .Y(n19546) );
  sky130_fd_sc_hd__a21oi_1 U25954 ( .A1(n26847), .A2(n19547), .B1(n19546), .Y(
        n19809) );
  sky130_fd_sc_hd__nand2_1 U25955 ( .A(n26847), .B(n19548), .Y(n19552) );
  sky130_fd_sc_hd__nand2_1 U25956 ( .A(n26849), .B(n19550), .Y(n19551) );
  sky130_fd_sc_hd__nand2_1 U25957 ( .A(n19552), .B(n19551), .Y(n19802) );
  sky130_fd_sc_hd__o22ai_1 U25958 ( .A1(j202_soc_core_intc_core_00_rg_ipr[80]), 
        .A2(n19809), .B1(n19802), .B2(j202_soc_core_intc_core_00_rg_ipr[81]), 
        .Y(n19554) );
  sky130_fd_sc_hd__nand2_1 U25959 ( .A(n19802), .B(
        j202_soc_core_intc_core_00_rg_ipr[81]), .Y(n19553) );
  sky130_fd_sc_hd__nand2_1 U25960 ( .A(n19554), .B(n19553), .Y(n19556) );
  sky130_fd_sc_hd__o21ai_1 U25961 ( .A1(j202_soc_core_intc_core_00_rg_ipr[82]), 
        .A2(n19556), .B1(n19555), .Y(n19558) );
  sky130_fd_sc_hd__nand2_1 U25962 ( .A(n19556), .B(
        j202_soc_core_intc_core_00_rg_ipr[82]), .Y(n19557) );
  sky130_fd_sc_hd__nand2_1 U25963 ( .A(n19558), .B(n19557), .Y(n19559) );
  sky130_fd_sc_hd__o21ai_1 U25964 ( .A1(j202_soc_core_intc_core_00_rg_ipr[83]), 
        .A2(n19817), .B1(n19559), .Y(n19561) );
  sky130_fd_sc_hd__nand2_1 U25965 ( .A(n19817), .B(
        j202_soc_core_intc_core_00_rg_ipr[83]), .Y(n19560) );
  sky130_fd_sc_hd__nand2_1 U25966 ( .A(n19561), .B(n19560), .Y(n19563) );
  sky130_fd_sc_hd__nand2_1 U25967 ( .A(n19563), .B(n19562), .Y(n19565) );
  sky130_fd_sc_hd__nand2_2 U25968 ( .A(n19565), .B(n19564), .Y(n27204) );
  sky130_fd_sc_hd__mux2_2 U25969 ( .A0(n19566), .A1(
        j202_soc_core_intc_core_00_rg_ipr[82]), .S(n27204), .X(n19819) );
  sky130_fd_sc_hd__nand2_1 U25970 ( .A(n24030), .B(
        j202_soc_core_intc_core_00_rg_ipr[13]), .Y(n19567) );
  sky130_fd_sc_hd__o2bb2ai_1 U25971 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[12]), .B2(n25359), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[9]), .A2_N(n25296), .Y(n19568) );
  sky130_fd_sc_hd__nand2_1 U25972 ( .A(n19569), .B(n19568), .Y(n19571) );
  sky130_fd_sc_hd__a2bb2oi_1 U25973 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[11]), .B2(n25277), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[14]), .A2_N(n25349), .Y(n19570) );
  sky130_fd_sc_hd__nand2_1 U25974 ( .A(n19571), .B(n19570), .Y(n19574) );
  sky130_fd_sc_hd__a21oi_1 U25975 ( .A1(n25278), .A2(
        j202_soc_core_intc_core_00_rg_ipr[15]), .B1(n19572), .Y(n19573) );
  sky130_fd_sc_hd__nand2_1 U25976 ( .A(n19574), .B(n19573), .Y(n19577) );
  sky130_fd_sc_hd__mux2i_1 U25977 ( .A0(j202_soc_core_intc_core_00_rg_ipr[14]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[10]), .S(n26839), .Y(n19600) );
  sky130_fd_sc_hd__nand2_1 U25978 ( .A(j202_soc_core_intc_core_00_rg_ipr[5]), 
        .B(n27677), .Y(n19579) );
  sky130_fd_sc_hd__o2bb2ai_1 U25979 ( .B1(j202_soc_core_intc_core_00_rg_ipr[4]), .B2(n24606), .A1_N(j202_soc_core_intc_core_00_rg_ipr[1]), .A2_N(n24056), .Y(
        n19578) );
  sky130_fd_sc_hd__a2bb2oi_1 U25980 ( .B1(j202_soc_core_intc_core_00_rg_ipr[3]), .B2(n24745), .A1_N(j202_soc_core_intc_core_00_rg_ipr[6]), .A2_N(n24987), .Y(
        n19580) );
  sky130_fd_sc_hd__a21oi_1 U25981 ( .A1(n24746), .A2(
        j202_soc_core_intc_core_00_rg_ipr[7]), .B1(n19582), .Y(n19584) );
  sky130_fd_sc_hd__mux2_2 U25982 ( .A0(j202_soc_core_intc_core_00_rg_ipr[2]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[6]), .S(n26842), .X(n19588) );
  sky130_fd_sc_hd__mux2_2 U25983 ( .A0(j202_soc_core_intc_core_00_rg_ipr[1]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[5]), .S(n26842), .X(n19641) );
  sky130_fd_sc_hd__mux2i_1 U25984 ( .A0(j202_soc_core_intc_core_00_rg_ipr[13]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[9]), .S(n26839), .Y(n19643) );
  sky130_fd_sc_hd__mux2_2 U25985 ( .A0(j202_soc_core_intc_core_00_rg_ipr[0]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[4]), .S(n26842), .X(n19647) );
  sky130_fd_sc_hd__mux2i_1 U25986 ( .A0(j202_soc_core_intc_core_00_rg_ipr[12]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[8]), .S(n26839), .Y(n19648) );
  sky130_fd_sc_hd__nand2_1 U25987 ( .A(n19647), .B(n19648), .Y(n19587) );
  sky130_fd_sc_hd__nand2_1 U25988 ( .A(n19641), .B(n19643), .Y(n19586) );
  sky130_fd_sc_hd__o2bb2ai_1 U25989 ( .B1(n19641), .B2(n19643), .A1_N(n19587), 
        .A2_N(n19586), .Y(n19590) );
  sky130_fd_sc_hd__nand2_1 U25990 ( .A(n19588), .B(n19600), .Y(n19589) );
  sky130_fd_sc_hd__nand2_1 U25991 ( .A(n19590), .B(n19589), .Y(n19593) );
  sky130_fd_sc_hd__mux2i_1 U25992 ( .A0(j202_soc_core_intc_core_00_rg_ipr[15]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[11]), .S(n26839), .Y(n19652) );
  sky130_fd_sc_hd__mux2_2 U25993 ( .A0(j202_soc_core_intc_core_00_rg_ipr[3]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[7]), .S(n26842), .X(n19653) );
  sky130_fd_sc_hd__a2bb2oi_1 U25994 ( .B1(n19591), .B2(n19599), .A1_N(n19652), 
        .A2_N(n19653), .Y(n19592) );
  sky130_fd_sc_hd__nand2_1 U25995 ( .A(n19593), .B(n19592), .Y(n19596) );
  sky130_fd_sc_hd__nand2_1 U25996 ( .A(n19653), .B(n19652), .Y(n19594) );
  sky130_fd_sc_hd__nand3_1 U25997 ( .A(n19596), .B(n19595), .C(n19594), .Y(
        n19598) );
  sky130_fd_sc_hd__mux2_2 U25998 ( .A0(n19600), .A1(n19599), .S(n25770), .X(
        n19651) );
  sky130_fd_sc_hd__nand2_1 U25999 ( .A(n25428), .B(
        j202_soc_core_intc_core_00_rg_ipr[21]), .Y(n19602) );
  sky130_fd_sc_hd__o2bb2ai_1 U26000 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[20]), .B2(n25429), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[17]), .A2_N(n19623), .Y(n19601) );
  sky130_fd_sc_hd__o211ai_1 U26001 ( .A1(j202_soc_core_intc_core_00_rg_ipr[18]), .A2(n26499), .B1(n19602), .C1(n19601), .Y(n19604) );
  sky130_fd_sc_hd__a2bb2oi_1 U26002 ( .B1(n26499), .B2(
        j202_soc_core_intc_core_00_rg_ipr[18]), .A1_N(n25431), .A2_N(
        j202_soc_core_intc_core_00_rg_ipr[23]), .Y(n19603) );
  sky130_fd_sc_hd__a21oi_1 U26003 ( .A1(n25431), .A2(
        j202_soc_core_intc_core_00_rg_ipr[23]), .B1(n19605), .Y(n19607) );
  sky130_fd_sc_hd__inv_1 U26004 ( .A(n26837), .Y(n19609) );
  sky130_fd_sc_hd__mux2i_1 U26005 ( .A0(j202_soc_core_intc_core_00_rg_ipr[22]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[18]), .S(n19609), .Y(n19628) );
  sky130_fd_sc_hd__nand2_1 U26006 ( .A(n25196), .B(
        j202_soc_core_intc_core_00_rg_ipr[29]), .Y(n19611) );
  sky130_fd_sc_hd__o2bb2ai_1 U26007 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[28]), .B2(n25863), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[25]), .A2_N(n25446), .Y(n19610) );
  sky130_fd_sc_hd__o211ai_1 U26008 ( .A1(j202_soc_core_intc_core_00_rg_ipr[26]), .A2(n27101), .B1(n19611), .C1(n19610), .Y(n19613) );
  sky130_fd_sc_hd__nand2_1 U26009 ( .A(n27101), .B(
        j202_soc_core_intc_core_00_rg_ipr[26]), .Y(n19612) );
  sky130_fd_sc_hd__nand2_1 U26010 ( .A(n19613), .B(n19612), .Y(n19615) );
  sky130_fd_sc_hd__nand2_1 U26011 ( .A(n25448), .B(
        j202_soc_core_intc_core_00_rg_ipr[31]), .Y(n19614) );
  sky130_fd_sc_hd__nand2_1 U26012 ( .A(n19615), .B(n19614), .Y(n19619) );
  sky130_fd_sc_hd__a21oi_1 U26013 ( .A1(n25447), .A2(
        j202_soc_core_intc_core_00_rg_ipr[27]), .B1(n19616), .Y(n19618) );
  sky130_fd_sc_hd__a21oi_1 U26014 ( .A1(n19619), .A2(n19618), .B1(n19617), .Y(
        n19620) );
  sky130_fd_sc_hd__mux2i_1 U26015 ( .A0(n25088), .A1(n27101), .S(n26838), .Y(
        n19639) );
  sky130_fd_sc_hd__mux2_2 U26016 ( .A0(n25447), .A1(n25448), .S(n19620), .X(
        n19656) );
  sky130_fd_sc_hd__mux2_2 U26017 ( .A0(j202_soc_core_intc_core_00_rg_ipr[19]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[23]), .S(n26837), .X(n19633) );
  sky130_fd_sc_hd__o2bb2ai_1 U26018 ( .B1(n19640), .B2(n19622), .A1_N(n19621), 
        .A2_N(n19657), .Y(n19636) );
  sky130_fd_sc_hd__mux2i_1 U26019 ( .A0(j202_soc_core_intc_core_00_rg_ipr[25]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[29]), .S(n26838), .Y(n19625) );
  sky130_fd_sc_hd__mux2i_1 U26020 ( .A0(n25428), .A1(n19623), .S(n26837), .Y(
        n19650) );
  sky130_fd_sc_hd__nand2_1 U26021 ( .A(n19649), .B(n19624), .Y(n19630) );
  sky130_fd_sc_hd__nand2_1 U26022 ( .A(n19625), .B(n19650), .Y(n19627) );
  sky130_fd_sc_hd__mux2_2 U26023 ( .A0(j202_soc_core_intc_core_00_rg_ipr[16]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[20]), .S(n26837), .X(n19644) );
  sky130_fd_sc_hd__mux2i_1 U26024 ( .A0(j202_soc_core_intc_core_00_rg_ipr[24]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[28]), .S(n26838), .Y(n19645) );
  sky130_fd_sc_hd__nand2_1 U26025 ( .A(n19644), .B(n19645), .Y(n19626) );
  sky130_fd_sc_hd__nand2_1 U26026 ( .A(n19627), .B(n19626), .Y(n19629) );
  sky130_fd_sc_hd__a2bb2oi_1 U26027 ( .B1(n19630), .B2(n19629), .A1_N(n19639), 
        .A2_N(n19628), .Y(n19635) );
  sky130_fd_sc_hd__a21oi_1 U26028 ( .A1(n19656), .A2(n19633), .B1(n19632), .Y(
        n19634) );
  sky130_fd_sc_hd__o21ai_1 U26029 ( .A1(n19636), .A2(n19635), .B1(n19634), .Y(
        n19638) );
  sky130_fd_sc_hd__mux2_2 U26030 ( .A0(n19640), .A1(n19639), .S(n25769), .X(
        n19664) );
  sky130_fd_sc_hd__mux2_2 U26031 ( .A0(n19654), .A1(n19653), .S(n25770), .X(
        n19789) );
  sky130_fd_sc_hd__a21oi_1 U26032 ( .A1(n19658), .A2(n19789), .B1(n19655), .Y(
        n19660) );
  sky130_fd_sc_hd__mux2_2 U26033 ( .A0(n19657), .A1(n19656), .S(n25769), .X(
        n19790) );
  sky130_fd_sc_hd__o21ai_1 U26034 ( .A1(n19789), .A2(n12127), .B1(n19790), .Y(
        n19659) );
  sky130_fd_sc_hd__nand2_1 U26035 ( .A(n19660), .B(n19659), .Y(n19663) );
  sky130_fd_sc_hd__mux2i_1 U26036 ( .A0(n19665), .A1(n19664), .S(n27202), .Y(
        n19785) );
  sky130_fd_sc_hd__nand2_1 U26037 ( .A(n25460), .B(
        j202_soc_core_intc_core_00_rg_ipr[41]), .Y(n19668) );
  sky130_fd_sc_hd__nand2_1 U26038 ( .A(n24027), .B(
        j202_soc_core_intc_core_00_rg_ipr[45]), .Y(n19666) );
  sky130_fd_sc_hd__a2bb2oi_1 U26039 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[47]), .B2(n25463), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[42]), .A2_N(n25450), .Y(n19669) );
  sky130_fd_sc_hd__nand2_1 U26040 ( .A(n19670), .B(n19669), .Y(n19673) );
  sky130_fd_sc_hd__a21oi_1 U26041 ( .A1(n25462), .A2(
        j202_soc_core_intc_core_00_rg_ipr[43]), .B1(n19671), .Y(n19672) );
  sky130_fd_sc_hd__nand2_1 U26042 ( .A(n19673), .B(n19672), .Y(n19676) );
  sky130_fd_sc_hd__inv_2 U26043 ( .A(n19686), .Y(n26826) );
  sky130_fd_sc_hd__mux2_2 U26044 ( .A0(j202_soc_core_intc_core_00_rg_ipr[46]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[42]), .S(n26826), .X(n19699) );
  sky130_fd_sc_hd__nand2_1 U26045 ( .A(n25480), .B(
        j202_soc_core_intc_core_00_rg_ipr[37]), .Y(n19678) );
  sky130_fd_sc_hd__o2bb2ai_1 U26046 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[37]), .B2(n25480), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[32]), .A2_N(n25483), .Y(n19677) );
  sky130_fd_sc_hd__o211ai_1 U26047 ( .A1(j202_soc_core_intc_core_00_rg_ipr[34]), .A2(n25464), .B1(n19678), .C1(n19677), .Y(n19680) );
  sky130_fd_sc_hd__nand2_1 U26048 ( .A(n19680), .B(n19679), .Y(n19684) );
  sky130_fd_sc_hd__a21oi_1 U26049 ( .A1(n25484), .A2(
        j202_soc_core_intc_core_00_rg_ipr[39]), .B1(n19681), .Y(n19683) );
  sky130_fd_sc_hd__a21oi_1 U26050 ( .A1(n19684), .A2(n19683), .B1(n19682), .Y(
        n19685) );
  sky130_fd_sc_hd__mux2i_1 U26051 ( .A0(j202_soc_core_intc_core_00_rg_ipr[38]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[34]), .S(n26823), .Y(n19690) );
  sky130_fd_sc_hd__mux2_2 U26052 ( .A0(j202_soc_core_intc_core_00_rg_ipr[47]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[43]), .S(n26826), .X(n19756) );
  sky130_fd_sc_hd__mux2_2 U26053 ( .A0(j202_soc_core_intc_core_00_rg_ipr[33]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[37]), .S(n19685), .X(n19737) );
  sky130_fd_sc_hd__mux2i_1 U26054 ( .A0(j202_soc_core_intc_core_00_rg_ipr[41]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[45]), .S(n19686), .Y(n19739) );
  sky130_fd_sc_hd__mux2i_1 U26055 ( .A0(j202_soc_core_intc_core_00_rg_ipr[36]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[32]), .S(n26823), .Y(n19744) );
  sky130_fd_sc_hd__nand2_1 U26056 ( .A(n19737), .B(n19739), .Y(n19687) );
  sky130_fd_sc_hd__o21ai_1 U26057 ( .A1(n19737), .A2(n19739), .B1(n19688), .Y(
        n19689) );
  sky130_fd_sc_hd__o21ai_1 U26058 ( .A1(n19699), .A2(n19690), .B1(n19689), .Y(
        n19692) );
  sky130_fd_sc_hd__nand2_1 U26059 ( .A(n19699), .B(n19690), .Y(n19691) );
  sky130_fd_sc_hd__nand2_1 U26060 ( .A(n19692), .B(n19691), .Y(n19693) );
  sky130_fd_sc_hd__mux2i_1 U26061 ( .A0(j202_soc_core_intc_core_00_rg_ipr[39]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[35]), .S(n26823), .Y(n19754) );
  sky130_fd_sc_hd__nand2_1 U26062 ( .A(n19693), .B(n19756), .Y(n19694) );
  sky130_fd_sc_hd__nand2_1 U26063 ( .A(n25195), .B(
        j202_soc_core_intc_core_00_rg_ipr[61]), .Y(n19701) );
  sky130_fd_sc_hd__o2bb2ai_1 U26064 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[60]), .B2(n25854), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[57]), .A2_N(n26952), .Y(n19700) );
  sky130_fd_sc_hd__o211ai_1 U26065 ( .A1(j202_soc_core_intc_core_00_rg_ipr[58]), .A2(n25486), .B1(n19701), .C1(n19700), .Y(n19703) );
  sky130_fd_sc_hd__nand2_1 U26066 ( .A(n19703), .B(n19702), .Y(n19707) );
  sky130_fd_sc_hd__a21oi_1 U26067 ( .A1(n25642), .A2(
        j202_soc_core_intc_core_00_rg_ipr[63]), .B1(n19704), .Y(n19706) );
  sky130_fd_sc_hd__mux2i_1 U26068 ( .A0(j202_soc_core_intc_core_00_rg_ipr[62]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[58]), .S(n26829), .Y(n19736) );
  sky130_fd_sc_hd__nand2_1 U26069 ( .A(n25718), .B(
        j202_soc_core_intc_core_00_rg_ipr[53]), .Y(n19709) );
  sky130_fd_sc_hd__o2bb2ai_1 U26070 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[52]), .B2(n25519), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[49]), .A2_N(n25375), .Y(n19708) );
  sky130_fd_sc_hd__o211ai_1 U26071 ( .A1(j202_soc_core_intc_core_00_rg_ipr[50]), .A2(n25503), .B1(n19709), .C1(n19708), .Y(n19711) );
  sky130_fd_sc_hd__a2bb2oi_1 U26072 ( .B1(
        j202_soc_core_intc_core_00_rg_ipr[51]), .B2(n27020), .A1_N(
        j202_soc_core_intc_core_00_rg_ipr[54]), .A2_N(n25502), .Y(n19710) );
  sky130_fd_sc_hd__nand2_1 U26073 ( .A(n19711), .B(n19710), .Y(n19713) );
  sky130_fd_sc_hd__nand2_1 U26074 ( .A(n25672), .B(
        j202_soc_core_intc_core_00_rg_ipr[55]), .Y(n19712) );
  sky130_fd_sc_hd__nand2_1 U26075 ( .A(n19713), .B(n19712), .Y(n19717) );
  sky130_fd_sc_hd__a21oi_2 U26076 ( .A1(n19717), .A2(n19716), .B1(n19715), .Y(
        n26830) );
  sky130_fd_sc_hd__mux2_2 U26077 ( .A0(j202_soc_core_intc_core_00_rg_ipr[54]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[50]), .S(n26830), .X(n19724) );
  sky130_fd_sc_hd__mux2_2 U26078 ( .A0(n27020), .A1(n25672), .S(n26830), .X(
        n19752) );
  sky130_fd_sc_hd__mux2_2 U26079 ( .A0(j202_soc_core_intc_core_00_rg_ipr[59]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[63]), .S(n19720), .X(n19729) );
  sky130_fd_sc_hd__mux2_2 U26080 ( .A0(n25375), .A1(n25718), .S(n26830), .X(
        n19722) );
  sky130_fd_sc_hd__mux2_2 U26081 ( .A0(j202_soc_core_intc_core_00_rg_ipr[57]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[61]), .S(n19720), .X(n19741) );
  sky130_fd_sc_hd__nand2_1 U26082 ( .A(n19740), .B(n19721), .Y(n19726) );
  sky130_fd_sc_hd__nand2_1 U26083 ( .A(n19722), .B(n19741), .Y(n19723) );
  sky130_fd_sc_hd__mux2_2 U26084 ( .A0(j202_soc_core_intc_core_00_rg_ipr[52]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[48]), .S(n26830), .X(n19747) );
  sky130_fd_sc_hd__mux2i_1 U26085 ( .A0(j202_soc_core_intc_core_00_rg_ipr[60]), 
        .A1(j202_soc_core_intc_core_00_rg_ipr[56]), .S(n26829), .Y(n19749) );
  sky130_fd_sc_hd__nand3_1 U26086 ( .A(n19723), .B(n19747), .C(n19749), .Y(
        n19725) );
  sky130_fd_sc_hd__a2bb2oi_1 U26087 ( .B1(n19726), .B2(n19725), .A1_N(n19724), 
        .A2_N(n19736), .Y(n19731) );
  sky130_fd_sc_hd__a21oi_1 U26088 ( .A1(n19752), .A2(n19729), .B1(n19728), .Y(
        n19730) );
  sky130_fd_sc_hd__o21ai_1 U26089 ( .A1(n19732), .A2(n19731), .B1(n19730), .Y(
        n19734) );
  sky130_fd_sc_hd__mux2_2 U26090 ( .A0(n19736), .A1(n19735), .S(n26827), .X(
        n19767) );
  sky130_fd_sc_hd__mux2_2 U26091 ( .A0(n19739), .A1(n19738), .S(n26824), .X(
        n19780) );
  sky130_fd_sc_hd__mux2_2 U26092 ( .A0(n19741), .A1(n19740), .S(n26827), .X(
        n19778) );
  sky130_fd_sc_hd__nand2_1 U26093 ( .A(n19780), .B(n19778), .Y(n19742) );
  sky130_fd_sc_hd__o21a_1 U26094 ( .A1(n19767), .A2(n19743), .B1(n19742), .X(
        n19751) );
  sky130_fd_sc_hd__mux2_2 U26095 ( .A0(n19746), .A1(n19745), .S(n26824), .X(
        n19774) );
  sky130_fd_sc_hd__mux2_2 U26096 ( .A0(n19749), .A1(n19748), .S(n26827), .X(
        n19772) );
  sky130_fd_sc_hd__o2bb2ai_1 U26097 ( .B1(n19778), .B2(n19780), .A1_N(n19774), 
        .A2_N(n19772), .Y(n19750) );
  sky130_fd_sc_hd__nand2_1 U26098 ( .A(n19751), .B(n19750), .Y(n19759) );
  sky130_fd_sc_hd__mux2_2 U26099 ( .A0(n19753), .A1(n19752), .S(n26827), .X(
        n19786) );
  sky130_fd_sc_hd__nand2_1 U26100 ( .A(n19759), .B(n19758), .Y(n19761) );
  sky130_fd_sc_hd__or2_0 U26101 ( .A(n19786), .B(n19788), .X(n19760) );
  sky130_fd_sc_hd__nand2_1 U26102 ( .A(n19761), .B(n19760), .Y(n19764) );
  sky130_fd_sc_hd__mux2i_1 U26103 ( .A0(n19768), .A1(n19767), .S(n26831), .Y(
        n19800) );
  sky130_fd_sc_hd__mux2i_1 U26104 ( .A0(n19771), .A1(n19770), .S(n27202), .Y(
        n19804) );
  sky130_fd_sc_hd__mux2i_1 U26105 ( .A0(n19774), .A1(n19773), .S(n26831), .Y(
        n19808) );
  sky130_fd_sc_hd__mux2i_1 U26106 ( .A0(n19777), .A1(n19776), .S(n27202), .Y(
        n19807) );
  sky130_fd_sc_hd__nand2_1 U26107 ( .A(n19808), .B(n19807), .Y(n19781) );
  sky130_fd_sc_hd__mux2i_1 U26108 ( .A0(n19780), .A1(n19779), .S(n26831), .Y(
        n19805) );
  sky130_fd_sc_hd__o21ai_1 U26109 ( .A1(n19804), .A2(n19781), .B1(n19805), .Y(
        n19783) );
  sky130_fd_sc_hd__nand2_1 U26110 ( .A(n19781), .B(n19804), .Y(n19782) );
  sky130_fd_sc_hd__nand2_1 U26111 ( .A(n19783), .B(n19782), .Y(n19784) );
  sky130_fd_sc_hd__o21ai_1 U26112 ( .A1(n19785), .A2(n19800), .B1(n19784), .Y(
        n19793) );
  sky130_fd_sc_hd__mux2i_1 U26113 ( .A0(n19788), .A1(n19787), .S(n26831), .Y(
        n19794) );
  sky130_fd_sc_hd__mux2i_1 U26114 ( .A0(n19791), .A1(n19790), .S(n27202), .Y(
        n19816) );
  sky130_fd_sc_hd__nand2_1 U26115 ( .A(n19793), .B(n19792), .Y(n19797) );
  sky130_fd_sc_hd__nand2_4 U26116 ( .A(n19799), .B(n19798), .Y(n26835) );
  sky130_fd_sc_hd__mux2i_1 U26117 ( .A0(n19801), .A1(n19800), .S(n26835), .Y(
        n25524) );
  sky130_fd_sc_hd__mux2_2 U26118 ( .A0(n19803), .A1(
        j202_soc_core_intc_core_00_rg_ipr[81]), .S(n27204), .X(n26901) );
  sky130_fd_sc_hd__mux2i_1 U26119 ( .A0(n19806), .A1(n19805), .S(n26835), .Y(
        n26905) );
  sky130_fd_sc_hd__mux2i_1 U26120 ( .A0(n12126), .A1(n19808), .S(n26835), .Y(
        n25753) );
  sky130_fd_sc_hd__mux2i_1 U26121 ( .A0(n19810), .A1(
        j202_soc_core_intc_core_00_rg_ipr[80]), .S(n27204), .Y(n25754) );
  sky130_fd_sc_hd__nand2_1 U26122 ( .A(n25753), .B(n25754), .Y(n19811) );
  sky130_fd_sc_hd__o21ai_1 U26123 ( .A1(n26901), .A2(n26905), .B1(n19811), .Y(
        n19813) );
  sky130_fd_sc_hd__nand2_1 U26124 ( .A(n26905), .B(n26901), .Y(n19812) );
  sky130_fd_sc_hd__nand2_1 U26125 ( .A(n19813), .B(n19812), .Y(n19814) );
  sky130_fd_sc_hd__o21ai_1 U26126 ( .A1(n19819), .A2(n25524), .B1(n19814), .Y(
        n19827) );
  sky130_fd_sc_hd__mux2i_1 U26127 ( .A0(n19816), .A1(n19815), .S(n26835), .Y(
        n25538) );
  sky130_fd_sc_hd__mux2_2 U26128 ( .A0(n19818), .A1(
        j202_soc_core_intc_core_00_rg_ipr[83]), .S(n27204), .X(n19820) );
  sky130_fd_sc_hd__nand2_1 U26129 ( .A(n25537), .B(n19821), .Y(n19824) );
  sky130_fd_sc_hd__nand2_1 U26130 ( .A(n19824), .B(n19823), .Y(n19825) );
  sky130_fd_sc_hd__nor2_1 U26131 ( .A(n24585), .B(n26851), .Y(n29069) );
  sky130_fd_sc_hd__nor2_1 U26132 ( .A(n20059), .B(n20110), .Y(n20310) );
  sky130_fd_sc_hd__nand2_1 U26133 ( .A(n19829), .B(n20199), .Y(n20179) );
  sky130_fd_sc_hd__a31oi_1 U26134 ( .A1(n20310), .A2(n19893), .A3(n20207), 
        .B1(n20906), .Y(n19840) );
  sky130_fd_sc_hd__a31oi_1 U26135 ( .A1(n19988), .A2(n19994), .A3(n19831), 
        .B1(n20873), .Y(n19839) );
  sky130_fd_sc_hd__nor2_1 U26136 ( .A(n19832), .B(n20114), .Y(n20382) );
  sky130_fd_sc_hd__nor4_1 U26137 ( .A(n19834), .B(n20313), .C(n20188), .D(
        n19833), .Y(n19835) );
  sky130_fd_sc_hd__a31oi_1 U26138 ( .A1(n20382), .A2(n19835), .A3(n20308), 
        .B1(n20927), .Y(n19838) );
  sky130_fd_sc_hd__nor2_1 U26139 ( .A(n20904), .B(n19998), .Y(n20015) );
  sky130_fd_sc_hd__a31oi_1 U26140 ( .A1(n19946), .A2(n20015), .A3(n19836), 
        .B1(n20925), .Y(n19837) );
  sky130_fd_sc_hd__nor4_1 U26141 ( .A(n19840), .B(n19839), .C(n19838), .D(
        n19837), .Y(n19857) );
  sky130_fd_sc_hd__nor2_1 U26142 ( .A(n20363), .B(n20197), .Y(n20174) );
  sky130_fd_sc_hd__nand2_1 U26143 ( .A(n19971), .B(n19842), .Y(n20862) );
  sky130_fd_sc_hd__nand3_1 U26144 ( .A(n20118), .B(n20047), .C(n13279), .Y(
        n19843) );
  sky130_fd_sc_hd__nand2_1 U26145 ( .A(n19992), .B(n20386), .Y(n20189) );
  sky130_fd_sc_hd__nor4_1 U26146 ( .A(n20189), .B(n20240), .C(n20196), .D(
        n20226), .Y(n19844) );
  sky130_fd_sc_hd__a21oi_1 U26147 ( .A1(n20174), .A2(n19844), .B1(n20925), .Y(
        n19854) );
  sky130_fd_sc_hd__nand3_1 U26148 ( .A(n12165), .B(n20073), .C(n20007), .Y(
        n20215) );
  sky130_fd_sc_hd__nor2_1 U26149 ( .A(n20215), .B(n20197), .Y(n20005) );
  sky130_fd_sc_hd__nand2_1 U26150 ( .A(n20052), .B(n20372), .Y(n19945) );
  sky130_fd_sc_hd__nor2_1 U26151 ( .A(n20177), .B(n19945), .Y(n20193) );
  sky130_fd_sc_hd__nor2_1 U26152 ( .A(n20110), .B(n19845), .Y(n19846) );
  sky130_fd_sc_hd__a31oi_1 U26153 ( .A1(n20005), .A2(n20193), .A3(n19846), 
        .B1(n20927), .Y(n19853) );
  sky130_fd_sc_hd__nor2_1 U26154 ( .A(n19848), .B(n19847), .Y(n19849) );
  sky130_fd_sc_hd__nand2_1 U26155 ( .A(n19849), .B(n21206), .Y(n19903) );
  sky130_fd_sc_hd__o31a_1 U26156 ( .A1(n19903), .A2(n20240), .A3(n20312), .B1(
        n20892), .X(n19852) );
  sky130_fd_sc_hd__a31oi_1 U26157 ( .A1(n20170), .A2(n20013), .A3(n19850), 
        .B1(n20906), .Y(n19851) );
  sky130_fd_sc_hd__nor4_1 U26158 ( .A(n19854), .B(n19853), .C(n19852), .D(
        n19851), .Y(n19855) );
  sky130_fd_sc_hd__o22a_1 U26159 ( .A1(n19857), .A2(n19856), .B1(n21179), .B2(
        n19855), .X(n19925) );
  sky130_fd_sc_hd__nand2b_1 U26160 ( .A_N(n19858), .B(n25677), .Y(n20152) );
  sky130_fd_sc_hd__nand2_1 U26161 ( .A(j202_soc_core_bldc_core_00_adc_en), .B(
        n27603), .Y(n19860) );
  sky130_fd_sc_hd__o22ai_1 U26162 ( .A1(n20157), .A2(n19860), .B1(n19859), 
        .B2(n20154), .Y(n19861) );
  sky130_fd_sc_hd__o2bb2ai_1 U26163 ( .B1(n28583), .B2(n20160), .A1_N(n28915), 
        .A2_N(n19861), .Y(n19862) );
  sky130_fd_sc_hd__nand2_1 U26164 ( .A(n19862), .B(n20164), .Y(n19920) );
  sky130_fd_sc_hd__nand2_1 U26165 ( .A(n21666), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[65]), .Y(n19915) );
  sky130_fd_sc_hd__nand2_1 U26166 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[1]), .Y(n19914) );
  sky130_fd_sc_hd__nand3_1 U26167 ( .A(n19915), .B(n21738), .C(n19914), .Y(
        n19871) );
  sky130_fd_sc_hd__nand2_1 U26168 ( .A(n21699), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[33]), .Y(n19870) );
  sky130_fd_sc_hd__nand2_1 U26169 ( .A(n21698), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[97]), .Y(n19869) );
  sky130_fd_sc_hd__nand2_1 U26170 ( .A(n21667), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[9]), .Y(n19866) );
  sky130_fd_sc_hd__nand2_1 U26171 ( .A(n24376), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[17]), .Y(n19865) );
  sky130_fd_sc_hd__nand2_1 U26172 ( .A(n21668), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[1]), .Y(n19864) );
  sky130_fd_sc_hd__nand2_1 U26173 ( .A(n21669), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[25]), .Y(n19863) );
  sky130_fd_sc_hd__nand4_1 U26174 ( .A(n19866), .B(n19865), .C(n19864), .D(
        n19863), .Y(n19867) );
  sky130_fd_sc_hd__nand2_1 U26175 ( .A(n21675), .B(n19867), .Y(n19868) );
  sky130_fd_sc_hd__nand3_1 U26176 ( .A(n19870), .B(n19869), .C(n19868), .Y(
        n19916) );
  sky130_fd_sc_hd__nor2_1 U26177 ( .A(n19871), .B(n19916), .Y(n19872) );
  sky130_fd_sc_hd__nand2_1 U26178 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_period[1]), .Y(n19918) );
  sky130_fd_sc_hd__nand3_1 U26179 ( .A(n19920), .B(n19872), .C(n19918), .Y(
        n19896) );
  sky130_fd_sc_hd__nor2_1 U26180 ( .A(n19874), .B(n19873), .Y(n20356) );
  sky130_fd_sc_hd__nor2_1 U26181 ( .A(n20180), .B(n20215), .Y(n20206) );
  sky130_fd_sc_hd__nand2_1 U26182 ( .A(n19988), .B(n20206), .Y(n20191) );
  sky130_fd_sc_hd__nor4_1 U26183 ( .A(n20356), .B(n19876), .C(n19875), .D(
        n20191), .Y(n19877) );
  sky130_fd_sc_hd__nand2b_1 U26184 ( .A_N(n19877), .B(n20335), .Y(n19890) );
  sky130_fd_sc_hd__and4_1 U26185 ( .A(n20221), .B(n20350), .C(n19879), .D(
        n19878), .X(n19880) );
  sky130_fd_sc_hd__nand4_1 U26186 ( .A(n19880), .B(n20306), .C(n20885), .D(
        n19971), .Y(n19882) );
  sky130_fd_sc_hd__o21ai_1 U26187 ( .A1(n19882), .A2(n19881), .B1(n20912), .Y(
        n19889) );
  sky130_fd_sc_hd__nand2_1 U26188 ( .A(n20214), .B(n20843), .Y(n20198) );
  sky130_fd_sc_hd__nor2_1 U26189 ( .A(n20198), .B(n20313), .Y(n19885) );
  sky130_fd_sc_hd__nand4_1 U26190 ( .A(n19885), .B(n20228), .C(n20384), .D(
        n19884), .Y(n19887) );
  sky130_fd_sc_hd__nand3_1 U26192 ( .A(n19890), .B(n19889), .C(n19888), .Y(
        n19895) );
  sky130_fd_sc_hd__nand2_1 U26193 ( .A(n19891), .B(n20305), .Y(n19976) );
  sky130_fd_sc_hd__nor2_1 U26194 ( .A(n19976), .B(n19901), .Y(n19892) );
  sky130_fd_sc_hd__a31oi_1 U26195 ( .A1(n19893), .A2(n19892), .A3(n20375), 
        .B1(n20873), .Y(n19894) );
  sky130_fd_sc_hd__o21a_1 U26196 ( .A1(n19895), .A2(n19894), .B1(n21697), .X(
        n19921) );
  sky130_fd_sc_hd__nor2_1 U26197 ( .A(n19896), .B(n19921), .Y(n19912) );
  sky130_fd_sc_hd__nand2_1 U26198 ( .A(n19897), .B(n20099), .Y(n20064) );
  sky130_fd_sc_hd__nor2_1 U26199 ( .A(n19898), .B(n20363), .Y(n20050) );
  sky130_fd_sc_hd__nor2_1 U26200 ( .A(n20046), .B(n20114), .Y(n20304) );
  sky130_fd_sc_hd__nand2_1 U26201 ( .A(n20050), .B(n20304), .Y(n20253) );
  sky130_fd_sc_hd__nand2_1 U26202 ( .A(n20328), .B(n20386), .Y(n20049) );
  sky130_fd_sc_hd__nor4_1 U26203 ( .A(n20918), .B(n20064), .C(n20253), .D(
        n20049), .Y(n19899) );
  sky130_fd_sc_hd__a21oi_1 U26204 ( .A1(n20232), .A2(n19899), .B1(n20906), .Y(
        n19910) );
  sky130_fd_sc_hd__nor4_1 U26205 ( .A(n19901), .B(n19900), .C(n20048), .D(
        n20252), .Y(n19902) );
  sky130_fd_sc_hd__a21oi_1 U26206 ( .A1(n20015), .A2(n19902), .B1(n20873), .Y(
        n19909) );
  sky130_fd_sc_hd__nand2_1 U26207 ( .A(n20352), .B(n20306), .Y(n20230) );
  sky130_fd_sc_hd__nor4b_1 U26208 ( .D_N(n20308), .A(n20198), .B(n19903), .C(
        n20230), .Y(n19904) );
  sky130_fd_sc_hd__a31oi_1 U26209 ( .A1(n19904), .A2(n20221), .A3(n20099), 
        .B1(n20927), .Y(n19908) );
  sky130_fd_sc_hd__nor4_1 U26210 ( .A(n20010), .B(n19991), .C(n19974), .D(
        n19905), .Y(n19906) );
  sky130_fd_sc_hd__a21oi_1 U26211 ( .A1(n19950), .A2(n19906), .B1(n20925), .Y(
        n19907) );
  sky130_fd_sc_hd__nor4_1 U26212 ( .A(n19910), .B(n19909), .C(n19908), .D(
        n19907), .Y(n19911) );
  sky130_fd_sc_hd__nand2b_1 U26213 ( .A_N(n19911), .B(n20908), .Y(n19923) );
  sky130_fd_sc_hd__nand3_1 U26214 ( .A(n19925), .B(n19912), .C(n19923), .Y(
        n19913) );
  sky130_fd_sc_hd__nand3_1 U26215 ( .A(n19915), .B(n21677), .C(n19914), .Y(
        n19917) );
  sky130_fd_sc_hd__nor2_1 U26216 ( .A(n19917), .B(n19916), .Y(n19919) );
  sky130_fd_sc_hd__nand3_1 U26217 ( .A(n19920), .B(n19919), .C(n19918), .Y(
        n19922) );
  sky130_fd_sc_hd__nor2_1 U26218 ( .A(n19922), .B(n19921), .Y(n19924) );
  sky130_fd_sc_hd__nand3_1 U26219 ( .A(n19925), .B(n19924), .C(n19923), .Y(
        n19926) );
  sky130_fd_sc_hd__a22oi_1 U26220 ( .A1(j202_soc_core_memory0_ram_dout0[33]), 
        .A2(n21604), .B1(n21591), .B2(j202_soc_core_memory0_ram_dout0[97]), 
        .Y(n19934) );
  sky130_fd_sc_hd__a22oi_1 U26221 ( .A1(j202_soc_core_memory0_ram_dout0[129]), 
        .A2(n21592), .B1(n21734), .B2(j202_soc_core_memory0_ram_dout0[65]), 
        .Y(n19933) );
  sky130_fd_sc_hd__a22oi_1 U26222 ( .A1(j202_soc_core_memory0_ram_dout0[161]), 
        .A2(n21590), .B1(n21733), .B2(j202_soc_core_memory0_ram_dout0[1]), .Y(
        n19932) );
  sky130_fd_sc_hd__a22oi_1 U26223 ( .A1(j202_soc_core_memory0_ram_dout0[193]), 
        .A2(n21732), .B1(n21735), .B2(j202_soc_core_memory0_ram_dout0[225]), 
        .Y(n19931) );
  sky130_fd_sc_hd__nor2_1 U26224 ( .A(n20562), .B(n20707), .Y(n28950) );
  sky130_fd_sc_hd__nand2_1 U26225 ( .A(j202_soc_core_memory0_ram_dout0[67]), 
        .B(n21734), .Y(n19935) );
  sky130_fd_sc_hd__nand2_1 U26226 ( .A(j202_soc_core_memory0_ram_dout0[387]), 
        .B(n21597), .Y(n19941) );
  sky130_fd_sc_hd__nand2_1 U26227 ( .A(j202_soc_core_memory0_ram_dout0[3]), 
        .B(n21733), .Y(n19940) );
  sky130_fd_sc_hd__nand2_1 U26228 ( .A(j202_soc_core_memory0_ram_dout0[227]), 
        .B(n21735), .Y(n19939) );
  sky130_fd_sc_hd__nand2_1 U26229 ( .A(j202_soc_core_memory0_ram_dout0[291]), 
        .B(n21603), .Y(n19938) );
  sky130_fd_sc_hd__nand4_1 U26230 ( .A(n19940), .B(n19941), .C(n19939), .D(
        n19938), .Y(n19942) );
  sky130_fd_sc_hd__nand2_1 U26231 ( .A(n20304), .B(n19943), .Y(n20229) );
  sky130_fd_sc_hd__nor4_1 U26232 ( .A(n20176), .B(n20229), .C(n19944), .D(
        n20057), .Y(n19949) );
  sky130_fd_sc_hd__nor2_1 U26233 ( .A(n20313), .B(n19945), .Y(n19968) );
  sky130_fd_sc_hd__nand4_1 U26234 ( .A(n20247), .B(n19968), .C(n20920), .D(
        n20117), .Y(n20203) );
  sky130_fd_sc_hd__nand2_1 U26235 ( .A(n19946), .B(n20375), .Y(n20903) );
  sky130_fd_sc_hd__nor3b_1 U26236 ( .C_N(n19947), .A(n20203), .B(n20903), .Y(
        n19948) );
  sky130_fd_sc_hd__o22ai_1 U26237 ( .A1(n19949), .A2(n20906), .B1(n19948), 
        .B2(n20925), .Y(n19956) );
  sky130_fd_sc_hd__nand4_1 U26238 ( .A(n20015), .B(n19950), .C(n20327), .D(
        n20377), .Y(n19954) );
  sky130_fd_sc_hd__a31oi_1 U26239 ( .A1(n19952), .A2(n20193), .A3(n19951), 
        .B1(n20873), .Y(n19953) );
  sky130_fd_sc_hd__a21oi_1 U26240 ( .A1(n20864), .A2(n19954), .B1(n19953), .Y(
        n19955) );
  sky130_fd_sc_hd__nand2b_1 U26241 ( .A_N(n19956), .B(n19955), .Y(n19957) );
  sky130_fd_sc_hd__nand2_1 U26242 ( .A(n19957), .B(n21697), .Y(n20041) );
  sky130_fd_sc_hd__nand2_1 U26243 ( .A(n21666), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[67]), .Y(n19959) );
  sky130_fd_sc_hd__nand2_1 U26244 ( .A(n21699), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[35]), .Y(n19958) );
  sky130_fd_sc_hd__nand2_1 U26245 ( .A(n19959), .B(n19958), .Y(n20037) );
  sky130_fd_sc_hd__nand2_1 U26246 ( .A(n21698), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[99]), .Y(n20035) );
  sky130_fd_sc_hd__nand2_1 U26247 ( .A(n21667), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[11]), .Y(n19963) );
  sky130_fd_sc_hd__nand2_1 U26248 ( .A(n24376), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[19]), .Y(n19962) );
  sky130_fd_sc_hd__nand2_1 U26249 ( .A(n21668), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[3]), .Y(n19961) );
  sky130_fd_sc_hd__nand2_1 U26250 ( .A(n21669), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[27]), .Y(n19960) );
  sky130_fd_sc_hd__nand4_1 U26251 ( .A(n19963), .B(n19962), .C(n19961), .D(
        n19960), .Y(n19964) );
  sky130_fd_sc_hd__nand2_1 U26252 ( .A(n21675), .B(n19964), .Y(n20034) );
  sky130_fd_sc_hd__nand2_1 U26253 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[3]), .Y(n20033) );
  sky130_fd_sc_hd__nand4_1 U26254 ( .A(n20035), .B(n21677), .C(n20034), .D(
        n20033), .Y(n19965) );
  sky130_fd_sc_hd__nor2_1 U26255 ( .A(n20037), .B(n19965), .Y(n19983) );
  sky130_fd_sc_hd__nand2_1 U26256 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_period[3]), .Y(n20039) );
  sky130_fd_sc_hd__nor2_1 U26257 ( .A(n20114), .B(n20110), .Y(n19966) );
  sky130_fd_sc_hd__a31oi_1 U26258 ( .A1(n19968), .A2(n19967), .A3(n19966), 
        .B1(n20906), .Y(n19981) );
  sky130_fd_sc_hd__nand2_1 U26259 ( .A(n19970), .B(n19969), .Y(n20243) );
  sky130_fd_sc_hd__nand3_1 U26260 ( .A(n20384), .B(n20842), .C(n20376), .Y(
        n20348) );
  sky130_fd_sc_hd__nand2_1 U26261 ( .A(n20326), .B(n20099), .Y(n20861) );
  sky130_fd_sc_hd__nor4_1 U26262 ( .A(n20872), .B(n20243), .C(n20348), .D(
        n20861), .Y(n19972) );
  sky130_fd_sc_hd__a31oi_1 U26263 ( .A1(n19972), .A2(n19971), .A3(n20372), 
        .B1(n20873), .Y(n19980) );
  sky130_fd_sc_hd__nor4_1 U26264 ( .A(n20096), .B(n19974), .C(n20176), .D(
        n19973), .Y(n19978) );
  sky130_fd_sc_hd__nor2_1 U26265 ( .A(n20059), .B(n20058), .Y(n19975) );
  sky130_fd_sc_hd__nand4_1 U26266 ( .A(n20228), .B(n19975), .C(n20885), .D(
        n20919), .Y(n20217) );
  sky130_fd_sc_hd__nor3_1 U26267 ( .A(n19976), .B(n20300), .C(n20217), .Y(
        n19977) );
  sky130_fd_sc_hd__o22ai_1 U26268 ( .A1(n19978), .A2(n20925), .B1(n19977), 
        .B2(n20927), .Y(n19979) );
  sky130_fd_sc_hd__nor3_1 U26269 ( .A(n19981), .B(n19980), .C(n19979), .Y(
        n19982) );
  sky130_fd_sc_hd__nand2b_1 U26270 ( .A_N(n19982), .B(n21727), .Y(n20038) );
  sky130_fd_sc_hd__nand4_1 U26271 ( .A(n20041), .B(n19983), .C(n20039), .D(
        n20038), .Y(n20026) );
  sky130_fd_sc_hd__nor3_1 U26272 ( .A(n19985), .B(n20918), .C(n19984), .Y(
        n20875) );
  sky130_fd_sc_hd__nand4_1 U26273 ( .A(n19986), .B(n20875), .C(n20099), .D(
        n20080), .Y(n19990) );
  sky130_fd_sc_hd__nor4_1 U26274 ( .A(n20045), .B(n19998), .C(n20219), .D(
        n19997), .Y(n19987) );
  sky130_fd_sc_hd__a31oi_1 U26275 ( .A1(n19988), .A2(n20065), .A3(n19987), 
        .B1(n20873), .Y(n19989) );
  sky130_fd_sc_hd__a21o_1 U26276 ( .A1(n20912), .A2(n19990), .B1(n19989), .X(
        n20002) );
  sky130_fd_sc_hd__nor2_1 U26277 ( .A(n20114), .B(n19991), .Y(n20194) );
  sky130_fd_sc_hd__nand2_1 U26278 ( .A(n19992), .B(n20194), .Y(n20171) );
  sky130_fd_sc_hd__nand2_1 U26279 ( .A(n20919), .B(n20884), .Y(n19993) );
  sky130_fd_sc_hd__nor4_1 U26280 ( .A(n20196), .B(n20171), .C(n19993), .D(
        n20882), .Y(n20000) );
  sky130_fd_sc_hd__nand4_1 U26281 ( .A(n19995), .B(n19994), .C(n20361), .D(
        n20384), .Y(n19996) );
  sky130_fd_sc_hd__nor3_1 U26282 ( .A(n19998), .B(n19997), .C(n19996), .Y(
        n19999) );
  sky130_fd_sc_hd__o22ai_1 U26283 ( .A1(n20000), .A2(n20927), .B1(n19999), 
        .B2(n20925), .Y(n20001) );
  sky130_fd_sc_hd__nand2_1 U26285 ( .A(n20003), .B(n20305), .Y(n20870) );
  sky130_fd_sc_hd__nor2_1 U26286 ( .A(n20004), .B(n20870), .Y(n20332) );
  sky130_fd_sc_hd__a31oi_1 U26287 ( .A1(n20006), .A2(n20005), .A3(n20332), 
        .B1(n20927), .Y(n20022) );
  sky130_fd_sc_hd__nand2_1 U26288 ( .A(n20008), .B(n20007), .Y(n20009) );
  sky130_fd_sc_hd__nor4_1 U26289 ( .A(n20011), .B(n20010), .C(n20105), .D(
        n20009), .Y(n20012) );
  sky130_fd_sc_hd__a21oi_1 U26290 ( .A1(n20013), .A2(n20012), .B1(n20925), .Y(
        n20021) );
  sky130_fd_sc_hd__a31oi_1 U26291 ( .A1(n20016), .A2(n20015), .A3(n20014), 
        .B1(n20906), .Y(n20020) );
  sky130_fd_sc_hd__nor2_1 U26292 ( .A(n20872), .B(n20243), .Y(n20017) );
  sky130_fd_sc_hd__a31oi_1 U26293 ( .A1(n20018), .A2(n20017), .A3(n20306), 
        .B1(n20873), .Y(n20019) );
  sky130_fd_sc_hd__nor4_1 U26294 ( .A(n20022), .B(n20021), .C(n20020), .D(
        n20019), .Y(n20023) );
  sky130_fd_sc_hd__nand2b_1 U26295 ( .A_N(n20023), .B(n20908), .Y(n20024) );
  sky130_fd_sc_hd__nand2_1 U26296 ( .A(n20025), .B(n20024), .Y(n20032) );
  sky130_fd_sc_hd__nor2_1 U26297 ( .A(n20026), .B(n20032), .Y(n20027) );
  sky130_fd_sc_hd__nand2_1 U26298 ( .A(j202_soc_core_memory0_ram_dout0[35]), 
        .B(n21604), .Y(n20030) );
  sky130_fd_sc_hd__nand2_1 U26299 ( .A(j202_soc_core_memory0_ram_dout0[323]), 
        .B(n21593), .Y(n20029) );
  sky130_fd_sc_hd__nand2_1 U26300 ( .A(j202_soc_core_memory0_ram_dout0[259]), 
        .B(n21605), .Y(n20028) );
  sky130_fd_sc_hd__nand3_1 U26301 ( .A(n20030), .B(n20029), .C(n20028), .Y(
        n20031) );
  sky130_fd_sc_hd__nand2_1 U26302 ( .A(j202_soc_core_memory0_ram_dout0[483]), 
        .B(n21771), .Y(n20044) );
  sky130_fd_sc_hd__nand4_1 U26303 ( .A(n20035), .B(n21738), .C(n20034), .D(
        n20033), .Y(n20036) );
  sky130_fd_sc_hd__nor2_1 U26304 ( .A(n20037), .B(n20036), .Y(n20040) );
  sky130_fd_sc_hd__and4_1 U26305 ( .A(n20041), .B(n20040), .C(n20039), .D(
        n20038), .X(n20042) );
  sky130_fd_sc_hd__nor2_1 U26306 ( .A(n20046), .B(n20045), .Y(n20224) );
  sky130_fd_sc_hd__nand4b_1 U26307 ( .A_N(n20048), .B(n20224), .C(n20377), .D(
        n20047), .Y(n20072) );
  sky130_fd_sc_hd__nand2_1 U26308 ( .A(n20383), .B(n20842), .Y(n20902) );
  sky130_fd_sc_hd__nor3_1 U26309 ( .A(n20049), .B(n20072), .C(n20902), .Y(
        n20051) );
  sky130_fd_sc_hd__nand2_1 U26310 ( .A(n20885), .B(n20375), .Y(n20354) );
  sky130_fd_sc_hd__nand2_1 U26311 ( .A(n20052), .B(n20885), .Y(n20053) );
  sky130_fd_sc_hd__nor2_1 U26312 ( .A(n20053), .B(n20072), .Y(n20337) );
  sky130_fd_sc_hd__nand3_1 U26313 ( .A(n20337), .B(n20055), .C(n20054), .Y(
        n20056) );
  sky130_fd_sc_hd__nand2_1 U26314 ( .A(n20056), .B(n20892), .Y(n20070) );
  sky130_fd_sc_hd__nor3_1 U26315 ( .A(n20059), .B(n20058), .C(n20057), .Y(
        n20299) );
  sky130_fd_sc_hd__nand2_1 U26316 ( .A(n20308), .B(n20060), .Y(n20852) );
  sky130_fd_sc_hd__nand4_1 U26317 ( .A(n20299), .B(n20061), .C(n20385), .D(
        n20843), .Y(n20062) );
  sky130_fd_sc_hd__nand2_1 U26318 ( .A(n20062), .B(n20864), .Y(n20069) );
  sky130_fd_sc_hd__nand2_1 U26319 ( .A(n20063), .B(n20386), .Y(n20391) );
  sky130_fd_sc_hd__nor4_1 U26320 ( .A(n20079), .B(n20064), .C(n20391), .D(
        n20111), .Y(n20066) );
  sky130_fd_sc_hd__nand2_1 U26321 ( .A(n20066), .B(n20065), .Y(n20067) );
  sky130_fd_sc_hd__nand2_1 U26322 ( .A(n20067), .B(n20335), .Y(n20068) );
  sky130_fd_sc_hd__nand4_1 U26323 ( .A(n20071), .B(n20070), .C(n20069), .D(
        n20068), .Y(n20092) );
  sky130_fd_sc_hd__nand2b_1 U26324 ( .A_N(n20072), .B(n20305), .Y(n20392) );
  sky130_fd_sc_hd__nand2_1 U26325 ( .A(n20383), .B(n20074), .Y(n20296) );
  sky130_fd_sc_hd__nor3_1 U26326 ( .A(n20882), .B(n20392), .C(n20296), .Y(
        n20090) );
  sky130_fd_sc_hd__nand2_1 U26327 ( .A(n20073), .B(n20375), .Y(n20393) );
  sky130_fd_sc_hd__nor3_1 U26328 ( .A(n20863), .B(n20862), .C(n20393), .Y(
        n20373) );
  sky130_fd_sc_hd__nand2_1 U26329 ( .A(n20075), .B(n20074), .Y(n20324) );
  sky130_fd_sc_hd__nor2_1 U26330 ( .A(n20324), .B(n20076), .Y(n20077) );
  sky130_fd_sc_hd__nand2_1 U26331 ( .A(n20373), .B(n20077), .Y(n20088) );
  sky130_fd_sc_hd__nand4_1 U26332 ( .A(n20841), .B(n20375), .C(n20350), .D(
        n20080), .Y(n20081) );
  sky130_fd_sc_hd__o21ai_0 U26333 ( .A1(n20349), .A2(n20081), .B1(n20335), .Y(
        n20085) );
  sky130_fd_sc_hd__nand2_1 U26334 ( .A(n20221), .B(n20382), .Y(n20845) );
  sky130_fd_sc_hd__o21ai_1 U26335 ( .A1(n20084), .A2(n20845), .B1(n20335), .Y(
        n20877) );
  sky130_fd_sc_hd__o211ai_1 U26336 ( .A1(n20086), .A2(n20927), .B1(n20085), 
        .C1(n20877), .Y(n20087) );
  sky130_fd_sc_hd__a21oi_1 U26337 ( .A1(n20088), .A2(n20912), .B1(n20087), .Y(
        n20089) );
  sky130_fd_sc_hd__o21a_1 U26338 ( .A1(n20873), .A2(n20090), .B1(n20089), .X(
        n20091) );
  sky130_fd_sc_hd__a2bb2oi_1 U26339 ( .B1(n20908), .B2(n20092), .A1_N(n21179), 
        .A2_N(n20091), .Y(n20137) );
  sky130_fd_sc_hd__a22oi_1 U26340 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[43]), .B1(n21698), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[107]), .Y(n20134) );
  sky130_fd_sc_hd__nand2_1 U26341 ( .A(n21666), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[75]), .Y(n20133) );
  sky130_fd_sc_hd__nand2_1 U26342 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[11]), .Y(n20132) );
  sky130_fd_sc_hd__nand4_1 U26343 ( .A(n20134), .B(n21677), .C(n20133), .D(
        n20132), .Y(n20093) );
  sky130_fd_sc_hd__nand2_1 U26344 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_period[11]), .Y(n20135) );
  sky130_fd_sc_hd__nand2b_1 U26345 ( .A_N(n20093), .B(n20135), .Y(n20109) );
  sky130_fd_sc_hd__nor2_1 U26346 ( .A(n20094), .B(n20354), .Y(n20095) );
  sky130_fd_sc_hd__a31oi_1 U26347 ( .A1(n20095), .A2(n20920), .A3(n20919), 
        .B1(n20925), .Y(n20108) );
  sky130_fd_sc_hd__nor3_1 U26348 ( .A(n20916), .B(n20096), .C(n20167), .Y(
        n20103) );
  sky130_fd_sc_hd__nor2_1 U26349 ( .A(n20218), .B(n20097), .Y(n20098) );
  sky130_fd_sc_hd__nand4_1 U26350 ( .A(n20099), .B(n20098), .C(n20386), .D(
        n20202), .Y(n20100) );
  sky130_fd_sc_hd__nand2_1 U26351 ( .A(n20100), .B(n20892), .Y(n20914) );
  sky130_fd_sc_hd__nand3_1 U26352 ( .A(n20306), .B(n20350), .C(n20842), .Y(
        n20101) );
  sky130_fd_sc_hd__o211ai_1 U26354 ( .A1(n20103), .A2(n20906), .B1(n20914), 
        .C1(n20102), .Y(n20107) );
  sky130_fd_sc_hd__nor3_1 U26355 ( .A(n20105), .B(n20104), .C(n20393), .Y(
        n20364) );
  sky130_fd_sc_hd__a31oi_1 U26356 ( .A1(n20364), .A2(n20374), .A3(n20331), 
        .B1(n20927), .Y(n20106) );
  sky130_fd_sc_hd__o31a_1 U26357 ( .A1(n20108), .A2(n20107), .A3(n20106), .B1(
        n21697), .X(n20139) );
  sky130_fd_sc_hd__nor2_1 U26358 ( .A(n20109), .B(n20139), .Y(n20130) );
  sky130_fd_sc_hd__nand2_1 U26359 ( .A(n20228), .B(n20375), .Y(n20922) );
  sky130_fd_sc_hd__nor4_1 U26360 ( .A(n20113), .B(n20112), .C(n20922), .D(
        n20881), .Y(n20128) );
  sky130_fd_sc_hd__nor4_1 U26361 ( .A(n20116), .B(n20336), .C(n20900), .D(
        n20115), .Y(n20126) );
  sky130_fd_sc_hd__nand3_1 U26362 ( .A(n20117), .B(n20118), .C(n20298), .Y(
        n20362) );
  sky130_fd_sc_hd__nor3_1 U26363 ( .A(n20348), .B(n20362), .C(n20845), .Y(
        n20124) );
  sky130_fd_sc_hd__nand2_1 U26364 ( .A(n20118), .B(n20298), .Y(n20119) );
  sky130_fd_sc_hd__nor2_1 U26365 ( .A(n20119), .B(n20348), .Y(n20120) );
  sky130_fd_sc_hd__nand2_1 U26366 ( .A(n20214), .B(n20120), .Y(n20122) );
  sky130_fd_sc_hd__o21a_1 U26368 ( .A1(n20906), .A2(n20124), .B1(n20123), .X(
        n20125) );
  sky130_fd_sc_hd__o21a_1 U26369 ( .A1(n20927), .A2(n20126), .B1(n20125), .X(
        n20127) );
  sky130_fd_sc_hd__nand2_1 U26371 ( .A(n20129), .B(n21727), .Y(n20141) );
  sky130_fd_sc_hd__nand2_1 U26372 ( .A(j202_soc_core_memory0_ram_dout0[491]), 
        .B(n21771), .Y(n20143) );
  sky130_fd_sc_hd__nand4_1 U26373 ( .A(n20134), .B(n21738), .C(n20133), .D(
        n20132), .Y(n20136) );
  sky130_fd_sc_hd__nand2b_1 U26374 ( .A_N(n20136), .B(n20135), .Y(n20140) );
  sky130_fd_sc_hd__nor3_1 U26375 ( .A(n20140), .B(n20139), .C(n20138), .Y(
        n20142) );
  sky130_fd_sc_hd__nand3_1 U26376 ( .A(n20143), .B(n20142), .C(n20141), .Y(
        n20144) );
  sky130_fd_sc_hd__a22oi_1 U26377 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[32]), .B1(n21698), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[96]), .Y(n20263) );
  sky130_fd_sc_hd__nand2_1 U26378 ( .A(n21666), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[64]), .Y(n20262) );
  sky130_fd_sc_hd__nand2_1 U26379 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[0]), .Y(n20261) );
  sky130_fd_sc_hd__nand4_1 U26380 ( .A(n20263), .B(n21738), .C(n20262), .D(
        n20261), .Y(n20166) );
  sky130_fd_sc_hd__nand2b_1 U26381 ( .A_N(n20148), .B(n20147), .Y(n22601) );
  sky130_fd_sc_hd__nand3_1 U26382 ( .A(n20157), .B(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_0_), .C(n25676), .Y(n20150) );
  sky130_fd_sc_hd__nor2_1 U26383 ( .A(n20150), .B(n20149), .Y(n20151) );
  sky130_fd_sc_hd__nand2_1 U26384 ( .A(n25677), .B(n20151), .Y(n25684) );
  sky130_fd_sc_hd__nor2_1 U26385 ( .A(n20152), .B(n28582), .Y(n20153) );
  sky130_fd_sc_hd__a31oi_1 U26386 ( .A1(n25677), .A2(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_), .A3(
        n25676), .B1(n20153), .Y(n20156) );
  sky130_fd_sc_hd__o22ai_1 U26387 ( .A1(n20157), .A2(n20156), .B1(n20155), 
        .B2(n20154), .Y(n20158) );
  sky130_fd_sc_hd__nand2_1 U26388 ( .A(n20158), .B(n28915), .Y(n20159) );
  sky130_fd_sc_hd__o211ai_1 U26389 ( .A1(n28586), .A2(n20160), .B1(n25684), 
        .C1(n20159), .Y(n20165) );
  sky130_fd_sc_hd__a22oi_1 U26390 ( .A1(n21668), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[0]), .B1(n21667), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[8]), .Y(n20162) );
  sky130_fd_sc_hd__a22oi_1 U26391 ( .A1(n21669), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[24]), .B1(n24376), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[16]), .Y(n20161) );
  sky130_fd_sc_hd__a21oi_1 U26392 ( .A1(n20162), .A2(n20161), .B1(n20860), .Y(
        n20163) );
  sky130_fd_sc_hd__a21oi_1 U26393 ( .A1(n20165), .A2(n20164), .B1(n20163), .Y(
        n20265) );
  sky130_fd_sc_hd__nand2_1 U26394 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_period[0]), .Y(n20264) );
  sky130_fd_sc_hd__nand3b_1 U26395 ( .A_N(n20166), .B(n20265), .C(n20264), .Y(
        n20187) );
  sky130_fd_sc_hd__nor4_1 U26396 ( .A(n20168), .B(n20218), .C(n20167), .D(
        n20189), .Y(n20169) );
  sky130_fd_sc_hd__a21oi_1 U26397 ( .A1(n20170), .A2(n20169), .B1(n20925), .Y(
        n20185) );
  sky130_fd_sc_hd__nor4_1 U26398 ( .A(n20180), .B(n20301), .C(n20172), .D(
        n20171), .Y(n20173) );
  sky130_fd_sc_hd__a21oi_1 U26399 ( .A1(n20174), .A2(n20173), .B1(n20927), .Y(
        n20184) );
  sky130_fd_sc_hd__nor4_1 U26400 ( .A(n20180), .B(n20177), .C(n20176), .D(
        n20175), .Y(n20182) );
  sky130_fd_sc_hd__nand2_1 U26401 ( .A(n20376), .B(n20375), .Y(n20178) );
  sky130_fd_sc_hd__nor4_1 U26402 ( .A(n20180), .B(n20301), .C(n20179), .D(
        n20178), .Y(n20181) );
  sky130_fd_sc_hd__o22ai_1 U26403 ( .A1(n20182), .A2(n20906), .B1(n20181), 
        .B2(n20873), .Y(n20183) );
  sky130_fd_sc_hd__nor3_1 U26404 ( .A(n20185), .B(n20184), .C(n20183), .Y(
        n20186) );
  sky130_fd_sc_hd__nor2_1 U26405 ( .A(n21179), .B(n20186), .Y(n20267) );
  sky130_fd_sc_hd__nor2_1 U26406 ( .A(n20187), .B(n20267), .Y(n20259) );
  sky130_fd_sc_hd__nor4_1 U26407 ( .A(n20324), .B(n20190), .C(n20189), .D(
        n20188), .Y(n20212) );
  sky130_fd_sc_hd__nor3_1 U26408 ( .A(n20302), .B(n20198), .C(n20191), .Y(
        n20192) );
  sky130_fd_sc_hd__a31oi_1 U26409 ( .A1(n20194), .A2(n20193), .A3(n20192), 
        .B1(n20873), .Y(n20210) );
  sky130_fd_sc_hd__nor4_1 U26410 ( .A(n20198), .B(n20197), .C(n20196), .D(
        n20195), .Y(n20200) );
  sky130_fd_sc_hd__a31oi_1 U26411 ( .A1(n20200), .A2(n20199), .A3(n20305), 
        .B1(n20927), .Y(n20209) );
  sky130_fd_sc_hd__nand2_1 U26412 ( .A(n20377), .B(n20202), .Y(n20389) );
  sky130_fd_sc_hd__nor3_1 U26413 ( .A(n20204), .B(n20389), .C(n20203), .Y(
        n20205) );
  sky130_fd_sc_hd__a31oi_1 U26414 ( .A1(n20207), .A2(n20206), .A3(n20205), 
        .B1(n20925), .Y(n20208) );
  sky130_fd_sc_hd__nor3_1 U26415 ( .A(n20210), .B(n20209), .C(n20208), .Y(
        n20211) );
  sky130_fd_sc_hd__nand2_1 U26417 ( .A(n20213), .B(n21697), .Y(n20271) );
  sky130_fd_sc_hd__nand2_1 U26418 ( .A(n20326), .B(n20214), .Y(n20216) );
  sky130_fd_sc_hd__nor2_1 U26419 ( .A(n20216), .B(n20215), .Y(n20248) );
  sky130_fd_sc_hd__nor4_1 U26420 ( .A(n20219), .B(n20252), .C(n20218), .D(
        n20217), .Y(n20220) );
  sky130_fd_sc_hd__a21oi_1 U26421 ( .A1(n20248), .A2(n20220), .B1(n20906), .Y(
        n20236) );
  sky130_fd_sc_hd__nand2_1 U26422 ( .A(n20222), .B(n20221), .Y(n20239) );
  sky130_fd_sc_hd__a31oi_1 U26423 ( .A1(n20224), .A2(n20248), .A3(n20223), 
        .B1(n20925), .Y(n20235) );
  sky130_fd_sc_hd__nor4_1 U26424 ( .A(n20226), .B(n20225), .C(n20229), .D(
        n20389), .Y(n20227) );
  sky130_fd_sc_hd__a21oi_1 U26425 ( .A1(n20228), .A2(n20227), .B1(n20873), .Y(
        n20234) );
  sky130_fd_sc_hd__nor2_1 U26426 ( .A(n20230), .B(n20229), .Y(n20231) );
  sky130_fd_sc_hd__a31oi_1 U26427 ( .A1(n13302), .A2(n20232), .A3(n20231), 
        .B1(n20927), .Y(n20233) );
  sky130_fd_sc_hd__nor4_1 U26428 ( .A(n20236), .B(n20235), .C(n20234), .D(
        n20233), .Y(n20237) );
  sky130_fd_sc_hd__nand2b_1 U26429 ( .A_N(n20237), .B(n21727), .Y(n20270) );
  sky130_fd_sc_hd__nor3_1 U26430 ( .A(n20240), .B(n20239), .C(n20238), .Y(
        n20242) );
  sky130_fd_sc_hd__a31oi_1 U26431 ( .A1(n20242), .A2(n20378), .A3(n20241), 
        .B1(n20906), .Y(n20257) );
  sky130_fd_sc_hd__nand4_1 U26432 ( .A(n20844), .B(n20884), .C(n20919), .D(
        n20244), .Y(n20250) );
  sky130_fd_sc_hd__nor3_1 U26433 ( .A(n20245), .B(n20349), .C(n20300), .Y(
        n20246) );
  sky130_fd_sc_hd__nand3_1 U26434 ( .A(n20248), .B(n20247), .C(n20246), .Y(
        n20249) );
  sky130_fd_sc_hd__a22oi_1 U26435 ( .A1(n20892), .A2(n20250), .B1(n20249), 
        .B2(n20864), .Y(n20256) );
  sky130_fd_sc_hd__nor4_1 U26436 ( .A(n20313), .B(n20253), .C(n20252), .D(
        n20251), .Y(n20254) );
  sky130_fd_sc_hd__nand2b_1 U26437 ( .A_N(n20254), .B(n20335), .Y(n20255) );
  sky130_fd_sc_hd__nand3b_1 U26438 ( .A_N(n20257), .B(n20256), .C(n20255), .Y(
        n20258) );
  sky130_fd_sc_hd__nand2_1 U26439 ( .A(n20258), .B(n20908), .Y(n20269) );
  sky130_fd_sc_hd__nand4_1 U26440 ( .A(n20259), .B(n20271), .C(n20270), .D(
        n20269), .Y(n20260) );
  sky130_fd_sc_hd__nand4_1 U26441 ( .A(n20263), .B(n21677), .C(n20262), .D(
        n20261), .Y(n20266) );
  sky130_fd_sc_hd__nand3b_1 U26442 ( .A_N(n20266), .B(n20265), .C(n20264), .Y(
        n20268) );
  sky130_fd_sc_hd__nor2_1 U26443 ( .A(n20268), .B(n20267), .Y(n20272) );
  sky130_fd_sc_hd__nor2_1 U26444 ( .A(n20273), .B(n27914), .Y(n20274) );
  sky130_fd_sc_hd__nand3_1 U26445 ( .A(n27906), .B(n20274), .C(
        j202_soc_core_ahbcs_6__HREADY_), .Y(n27167) );
  sky130_fd_sc_hd__nand2_1 U26446 ( .A(n28950), .B(n22581), .Y(n20283) );
  sky130_fd_sc_hd__nand2_1 U26447 ( .A(n20277), .B(n20276), .Y(n20278) );
  sky130_fd_sc_hd__xor2_1 U26448 ( .A(n20279), .B(n20278), .X(n23781) );
  sky130_fd_sc_hd__o22ai_1 U26449 ( .A1(n25743), .A2(n11143), .B1(
        j202_soc_core_j22_cpu_pc[1]), .B2(n21584), .Y(n20280) );
  sky130_fd_sc_hd__a21oi_1 U26450 ( .A1(n23781), .A2(n12158), .B1(n20280), .Y(
        n20282) );
  sky130_fd_sc_hd__nand2_1 U26451 ( .A(n22515), .B(n27443), .Y(n20281) );
  sky130_fd_sc_hd__nand2_1 U26452 ( .A(n27720), .B(n14849), .Y(n25108) );
  sky130_fd_sc_hd__inv_2 U26453 ( .A(n23305), .Y(n24118) );
  sky130_fd_sc_hd__nor2_1 U26454 ( .A(n29559), .B(n12459), .Y(n28976) );
  sky130_fd_sc_hd__nand2_1 U26455 ( .A(n28921), .B(n22581), .Y(n20293) );
  sky130_fd_sc_hd__xnor2_1 U26456 ( .A(n20285), .B(n21904), .Y(n24651) );
  sky130_fd_sc_hd__o22a_1 U26457 ( .A1(n26713), .A2(n11143), .B1(n26792), .B2(
        n22590), .X(n20290) );
  sky130_fd_sc_hd__nand2_1 U26458 ( .A(n20287), .B(n20286), .Y(n20288) );
  sky130_fd_sc_hd__xnor2_1 U26459 ( .A(n20288), .B(n21531), .Y(n24645) );
  sky130_fd_sc_hd__nand2_1 U26460 ( .A(n24645), .B(n12158), .Y(n20289) );
  sky130_fd_sc_hd__o211ai_1 U26461 ( .A1(n26792), .A2(n22592), .B1(n20290), 
        .C1(n20289), .Y(n20291) );
  sky130_fd_sc_hd__a21oi_1 U26462 ( .A1(n24651), .A2(n22596), .B1(n20291), .Y(
        n20292) );
  sky130_fd_sc_hd__nand2_1 U26463 ( .A(n20293), .B(n20292), .Y(n29013) );
  sky130_fd_sc_hd__a22oi_1 U26464 ( .A1(j202_soc_core_memory0_ram_dout0[392]), 
        .A2(n21597), .B1(n21593), .B2(j202_soc_core_memory0_ram_dout0[328]), 
        .Y(n20404) );
  sky130_fd_sc_hd__nand2_1 U26465 ( .A(n20295), .B(n20841), .Y(n20297) );
  sky130_fd_sc_hd__nor3_1 U26466 ( .A(n20297), .B(n20388), .C(n20296), .Y(
        n20320) );
  sky130_fd_sc_hd__nand3_1 U26467 ( .A(n20299), .B(n21206), .C(n20298), .Y(
        n20839) );
  sky130_fd_sc_hd__nor4_1 U26468 ( .A(n20302), .B(n20301), .C(n20300), .D(
        n20839), .Y(n20303) );
  sky130_fd_sc_hd__a31oi_1 U26469 ( .A1(n20327), .A2(n20304), .A3(n20303), 
        .B1(n20906), .Y(n20318) );
  sky130_fd_sc_hd__nand3_1 U26470 ( .A(n20306), .B(n20377), .C(n20305), .Y(
        n20322) );
  sky130_fd_sc_hd__nor3_1 U26471 ( .A(n20353), .B(n20322), .C(n20307), .Y(
        n20309) );
  sky130_fd_sc_hd__a31oi_1 U26472 ( .A1(n20310), .A2(n20309), .A3(n20308), 
        .B1(n20873), .Y(n20317) );
  sky130_fd_sc_hd__nor4_1 U26473 ( .A(n20918), .B(n20313), .C(n20312), .D(
        n20311), .Y(n20314) );
  sky130_fd_sc_hd__a31oi_1 U26474 ( .A1(n20315), .A2(n20329), .A3(n20314), 
        .B1(n20925), .Y(n20316) );
  sky130_fd_sc_hd__nor3_1 U26475 ( .A(n20318), .B(n20317), .C(n20316), .Y(
        n20319) );
  sky130_fd_sc_hd__nand2_1 U26477 ( .A(n20321), .B(n21727), .Y(n20424) );
  sky130_fd_sc_hd__nor3_1 U26478 ( .A(n20324), .B(n20323), .C(n20322), .Y(
        n20341) );
  sky130_fd_sc_hd__nand4_1 U26479 ( .A(n20841), .B(n20849), .C(n20326), .D(
        n20325), .Y(n20334) );
  sky130_fd_sc_hd__nand2_1 U26480 ( .A(n20328), .B(n20327), .Y(n20366) );
  sky130_fd_sc_hd__nand4_1 U26481 ( .A(n20332), .B(n20331), .C(n20330), .D(
        n20329), .Y(n20333) );
  sky130_fd_sc_hd__a22oi_1 U26482 ( .A1(n20335), .A2(n20334), .B1(n20333), 
        .B2(n20912), .Y(n20340) );
  sky130_fd_sc_hd__nor2_1 U26483 ( .A(n20898), .B(n20336), .Y(n20890) );
  sky130_fd_sc_hd__nand3_1 U26484 ( .A(n20337), .B(n20890), .C(n20384), .Y(
        n20338) );
  sky130_fd_sc_hd__nand2_1 U26485 ( .A(n20338), .B(n20892), .Y(n20339) );
  sky130_fd_sc_hd__o211ai_1 U26486 ( .A1(n20341), .A2(n20927), .B1(n20340), 
        .C1(n20339), .Y(n20342) );
  sky130_fd_sc_hd__nand2_1 U26487 ( .A(n20342), .B(n20908), .Y(n20418) );
  sky130_fd_sc_hd__xnor2_1 U26488 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[1]), 
        .B(j202_soc_core_uart_TOP_rx_fifo_wp[1]), .Y(n27140) );
  sky130_fd_sc_hd__xnor2_1 U26489 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[0]), 
        .B(j202_soc_core_uart_TOP_rx_fifo_wp[0]), .Y(n20343) );
  sky130_fd_sc_hd__nand2_1 U26490 ( .A(n27140), .B(n20343), .Y(n23308) );
  sky130_fd_sc_hd__nor3_1 U26491 ( .A(j202_soc_core_uart_TOP_rx_fifo_gb), .B(
        n20860), .C(n23308), .Y(n20411) );
  sky130_fd_sc_hd__nand2_1 U26492 ( .A(n21699), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[40]), .Y(n20345) );
  sky130_fd_sc_hd__nand2_1 U26493 ( .A(n21666), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[72]), .Y(n20344) );
  sky130_fd_sc_hd__nand2_1 U26494 ( .A(n20345), .B(n20344), .Y(n20416) );
  sky130_fd_sc_hd__nand2_1 U26495 ( .A(n21698), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[104]), .Y(n20414) );
  sky130_fd_sc_hd__nand2_1 U26496 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[8]), .Y(n20412) );
  sky130_fd_sc_hd__nand3_1 U26497 ( .A(n20414), .B(n21677), .C(n20412), .Y(
        n20346) );
  sky130_fd_sc_hd__nor3_1 U26498 ( .A(n20411), .B(n20416), .C(n20346), .Y(
        n20347) );
  sky130_fd_sc_hd__nand2_1 U26499 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_period[8]), .Y(n20417) );
  sky130_fd_sc_hd__nand3_1 U26500 ( .A(n20418), .B(n20347), .C(n20417), .Y(
        n20371) );
  sky130_fd_sc_hd__nor4_1 U26501 ( .A(n20349), .B(n20898), .C(n20348), .D(
        n20869), .Y(n20351) );
  sky130_fd_sc_hd__nand3_1 U26502 ( .A(n20352), .B(n20351), .C(n20350), .Y(
        n20360) );
  sky130_fd_sc_hd__nor4_1 U26503 ( .A(n20356), .B(n20355), .C(n20354), .D(
        n20353), .Y(n20357) );
  sky130_fd_sc_hd__a21oi_1 U26504 ( .A1(n20358), .A2(n20357), .B1(n20925), .Y(
        n20359) );
  sky130_fd_sc_hd__a21o_1 U26505 ( .A1(n20892), .A2(n20360), .B1(n20359), .X(
        n20370) );
  sky130_fd_sc_hd__nand3_1 U26506 ( .A(n20361), .B(n20385), .C(n20372), .Y(
        n20837) );
  sky130_fd_sc_hd__nor4_1 U26507 ( .A(n20363), .B(n20379), .C(n20362), .D(
        n20837), .Y(n20368) );
  sky130_fd_sc_hd__nand2_1 U26508 ( .A(n20364), .B(n20384), .Y(n20915) );
  sky130_fd_sc_hd__nor4_1 U26509 ( .A(n20870), .B(n20366), .C(n20365), .D(
        n20915), .Y(n20367) );
  sky130_fd_sc_hd__o22ai_1 U26510 ( .A1(n20368), .A2(n20906), .B1(n20367), 
        .B2(n20927), .Y(n20369) );
  sky130_fd_sc_hd__o21a_1 U26511 ( .A1(n20370), .A2(n20369), .B1(n21697), .X(
        n20410) );
  sky130_fd_sc_hd__nor2_1 U26512 ( .A(n20371), .B(n20410), .Y(n20400) );
  sky130_fd_sc_hd__a31oi_1 U26513 ( .A1(n20385), .A2(n20373), .A3(n20372), 
        .B1(n20906), .Y(n20398) );
  sky130_fd_sc_hd__nand2_1 U26514 ( .A(n20374), .B(n20885), .Y(n20923) );
  sky130_fd_sc_hd__nand4_1 U26515 ( .A(n20378), .B(n20377), .C(n20376), .D(
        n20375), .Y(n20911) );
  sky130_fd_sc_hd__nor4_1 U26516 ( .A(n20380), .B(n20379), .C(n20923), .D(
        n20911), .Y(n20381) );
  sky130_fd_sc_hd__a31oi_1 U26517 ( .A1(n20383), .A2(n20382), .A3(n20381), 
        .B1(n20925), .Y(n20397) );
  sky130_fd_sc_hd__nand3_1 U26518 ( .A(n12165), .B(n20385), .C(n20384), .Y(
        n20866) );
  sky130_fd_sc_hd__nand2_1 U26519 ( .A(n20387), .B(n20386), .Y(n20901) );
  sky130_fd_sc_hd__nor4_1 U26520 ( .A(n20389), .B(n20388), .C(n20866), .D(
        n20901), .Y(n20395) );
  sky130_fd_sc_hd__nor4_1 U26521 ( .A(n20393), .B(n20392), .C(n20391), .D(
        n20390), .Y(n20394) );
  sky130_fd_sc_hd__o22ai_1 U26522 ( .A1(n20395), .A2(n20927), .B1(n20394), 
        .B2(n20873), .Y(n20396) );
  sky130_fd_sc_hd__nor3_1 U26523 ( .A(n20398), .B(n20397), .C(n20396), .Y(
        n20399) );
  sky130_fd_sc_hd__nand2b_1 U26524 ( .A_N(n20399), .B(n13481), .Y(n20421) );
  sky130_fd_sc_hd__nand3_1 U26525 ( .A(n20424), .B(n20400), .C(n20421), .Y(
        n20401) );
  sky130_fd_sc_hd__a21oi_1 U26526 ( .A1(j202_soc_core_memory0_ram_dout0[424]), 
        .A2(n21598), .B1(n20401), .Y(n20403) );
  sky130_fd_sc_hd__a22oi_1 U26527 ( .A1(j202_soc_core_memory0_ram_dout0[8]), 
        .A2(n21733), .B1(n21605), .B2(j202_soc_core_memory0_ram_dout0[264]), 
        .Y(n20402) );
  sky130_fd_sc_hd__a22oi_1 U26528 ( .A1(j202_soc_core_memory0_ram_dout0[40]), 
        .A2(n21604), .B1(n21735), .B2(j202_soc_core_memory0_ram_dout0[232]), 
        .Y(n20409) );
  sky130_fd_sc_hd__a22oi_1 U26529 ( .A1(j202_soc_core_memory0_ram_dout0[72]), 
        .A2(n21734), .B1(n21603), .B2(j202_soc_core_memory0_ram_dout0[296]), 
        .Y(n20408) );
  sky130_fd_sc_hd__a22oi_1 U26530 ( .A1(j202_soc_core_memory0_ram_dout0[104]), 
        .A2(n21591), .B1(n21592), .B2(j202_soc_core_memory0_ram_dout0[136]), 
        .Y(n20407) );
  sky130_fd_sc_hd__nand2_1 U26531 ( .A(j202_soc_core_memory0_ram_dout0[488]), 
        .B(n21771), .Y(n20426) );
  sky130_fd_sc_hd__nand4_1 U26532 ( .A(n20414), .B(n20413), .C(n21738), .D(
        n20412), .Y(n20415) );
  sky130_fd_sc_hd__nor2_1 U26533 ( .A(n20416), .B(n20415), .Y(n20419) );
  sky130_fd_sc_hd__nand4_1 U26534 ( .A(n20420), .B(n20419), .C(n20418), .D(
        n20417), .Y(n20423) );
  sky130_fd_sc_hd__nor2_1 U26535 ( .A(n20423), .B(n20422), .Y(n20425) );
  sky130_fd_sc_hd__nand3_1 U26536 ( .A(n20426), .B(n20425), .C(n20424), .Y(
        n20427) );
  sky130_fd_sc_hd__a22oi_1 U26537 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__0_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__0_), .Y(n20561) );
  sky130_fd_sc_hd__nand2_1 U26538 ( .A(j202_soc_core_j22_cpu_pc[1]), .B(
        j202_soc_core_j22_cpu_ifetchl), .Y(n20429) );
  sky130_fd_sc_hd__nand2_1 U26539 ( .A(j202_soc_core_memory0_ram_dout0[208]), 
        .B(n21732), .Y(n20432) );
  sky130_fd_sc_hd__nand2_1 U26540 ( .A(j202_soc_core_memory0_ram_dout0[112]), 
        .B(n21591), .Y(n20431) );
  sky130_fd_sc_hd__nand2_1 U26541 ( .A(j202_soc_core_memory0_ram_dout0[400]), 
        .B(n21597), .Y(n20433) );
  sky130_fd_sc_hd__nand2_1 U26542 ( .A(n21666), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[80]), .Y(n20553) );
  sky130_fd_sc_hd__nand2_1 U26543 ( .A(n21675), .B(j202_soc_core_uart_div1[0]), 
        .Y(n20552) );
  sky130_fd_sc_hd__nand2_1 U26544 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[16]), .Y(n20551) );
  sky130_fd_sc_hd__nand4_1 U26545 ( .A(n20553), .B(n21677), .C(n20552), .D(
        n20551), .Y(n20436) );
  sky130_fd_sc_hd__nand2_1 U26546 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_duty[4]), .Y(n20435) );
  sky130_fd_sc_hd__nand2_1 U26547 ( .A(n21699), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[48]), .Y(n20434) );
  sky130_fd_sc_hd__nand2_1 U26548 ( .A(n20435), .B(n20434), .Y(n20550) );
  sky130_fd_sc_hd__nor2_1 U26549 ( .A(n20436), .B(n20550), .Y(n20543) );
  sky130_fd_sc_hd__nor2_1 U26550 ( .A(n20646), .B(n20437), .Y(n20438) );
  sky130_fd_sc_hd__and3_1 U26551 ( .A(n20440), .B(n20439), .C(n20438), .X(
        n20441) );
  sky130_fd_sc_hd__a31oi_1 U26552 ( .A1(n20608), .A2(n20614), .A3(n20441), 
        .B1(n20681), .Y(n20457) );
  sky130_fd_sc_hd__nand2_1 U26553 ( .A(n20442), .B(n20515), .Y(n20443) );
  sky130_fd_sc_hd__nor4_1 U26554 ( .A(n20676), .B(n20444), .C(n20675), .D(
        n20443), .Y(n20445) );
  sky130_fd_sc_hd__a31oi_1 U26555 ( .A1(n20494), .A2(n20445), .A3(n20502), 
        .B1(n20663), .Y(n20456) );
  sky130_fd_sc_hd__nor4_1 U26556 ( .A(n20448), .B(n20447), .C(n20595), .D(
        n20446), .Y(n20449) );
  sky130_fd_sc_hd__a21oi_1 U26557 ( .A1(n20450), .A2(n20449), .B1(n20683), .Y(
        n20455) );
  sky130_fd_sc_hd__nor4_1 U26558 ( .A(n20518), .B(n20667), .C(n20504), .D(
        n20611), .Y(n20451) );
  sky130_fd_sc_hd__a31oi_1 U26559 ( .A1(n20453), .A2(n20452), .A3(n20451), 
        .B1(n20651), .Y(n20454) );
  sky130_fd_sc_hd__nor4_1 U26560 ( .A(n20457), .B(n20456), .C(n20455), .D(
        n20454), .Y(n20488) );
  sky130_fd_sc_hd__nand3_1 U26561 ( .A(n20517), .B(n20458), .C(n20515), .Y(
        n20640) );
  sky130_fd_sc_hd__nor3_1 U26562 ( .A(n20459), .B(n20591), .C(n20640), .Y(
        n20460) );
  sky130_fd_sc_hd__a21oi_1 U26563 ( .A1(n20609), .A2(n20460), .B1(n20651), .Y(
        n20469) );
  sky130_fd_sc_hd__nand2b_1 U26564 ( .A_N(n20476), .B(n20648), .Y(n20462) );
  sky130_fd_sc_hd__nand4_1 U26565 ( .A(n20464), .B(n20584), .C(n20463), .D(
        n20569), .Y(n20467) );
  sky130_fd_sc_hd__o21ai_1 U26566 ( .A1(n20467), .A2(n20466), .B1(n20465), .Y(
        n20468) );
  sky130_fd_sc_hd__nand2b_1 U26567 ( .A_N(n20469), .B(n20468), .Y(n20486) );
  sky130_fd_sc_hd__and3_1 U26568 ( .A(n20472), .B(n20471), .C(n20470), .X(
        n20474) );
  sky130_fd_sc_hd__a31oi_1 U26569 ( .A1(n20475), .A2(n20474), .A3(n20473), 
        .B1(n20683), .Y(n20485) );
  sky130_fd_sc_hd__nor2_1 U26570 ( .A(n20477), .B(n20476), .Y(n20576) );
  sky130_fd_sc_hd__nor2_1 U26571 ( .A(n20676), .B(n20611), .Y(n20483) );
  sky130_fd_sc_hd__nand2_1 U26572 ( .A(n20479), .B(n20478), .Y(n20594) );
  sky130_fd_sc_hd__nor3_1 U26573 ( .A(n20481), .B(n20480), .C(n20594), .Y(
        n20482) );
  sky130_fd_sc_hd__a31oi_1 U26574 ( .A1(n20576), .A2(n20483), .A3(n20482), 
        .B1(n20681), .Y(n20484) );
  sky130_fd_sc_hd__nor3_1 U26575 ( .A(n20486), .B(n20485), .C(n20484), .Y(
        n20487) );
  sky130_fd_sc_hd__mux2i_1 U26576 ( .A0(n20488), .A1(n20487), .S(n20623), .Y(
        n20489) );
  sky130_fd_sc_hd__nand2_1 U26577 ( .A(n20489), .B(n20626), .Y(n20557) );
  sky130_fd_sc_hd__nor4_1 U26578 ( .A(n20491), .B(n20596), .C(n20631), .D(
        n20490), .Y(n20492) );
  sky130_fd_sc_hd__a31oi_1 U26579 ( .A1(n20494), .A2(n20493), .A3(n20492), 
        .B1(n20683), .Y(n20512) );
  sky130_fd_sc_hd__nor2_1 U26580 ( .A(n20518), .B(n20495), .Y(n20496) );
  sky130_fd_sc_hd__a31oi_1 U26581 ( .A1(n20498), .A2(n20497), .A3(n20496), 
        .B1(n20663), .Y(n20511) );
  sky130_fd_sc_hd__nor2b_1 U26582 ( .B_N(n20517), .A(n20499), .Y(n20501) );
  sky130_fd_sc_hd__a31oi_1 U26583 ( .A1(n20501), .A2(n20500), .A3(n20665), 
        .B1(n20681), .Y(n20510) );
  sky130_fd_sc_hd__nand2_1 U26584 ( .A(n20615), .B(n20601), .Y(n20503) );
  sky130_fd_sc_hd__nor4_1 U26585 ( .A(n20506), .B(n20505), .C(n20504), .D(
        n20503), .Y(n20507) );
  sky130_fd_sc_hd__a31oi_1 U26586 ( .A1(n20584), .A2(n20508), .A3(n20507), 
        .B1(n20651), .Y(n20509) );
  sky130_fd_sc_hd__nor4_1 U26587 ( .A(n20512), .B(n20511), .C(n20510), .D(
        n20509), .Y(n20541) );
  sky130_fd_sc_hd__nor2_1 U26588 ( .A(n20514), .B(n20513), .Y(n20573) );
  sky130_fd_sc_hd__nand3_1 U26589 ( .A(n20517), .B(n20516), .C(n20515), .Y(
        n20677) );
  sky130_fd_sc_hd__nor4b_1 U26590 ( .D_N(n20672), .A(n20518), .B(n20667), .C(
        n20677), .Y(n20519) );
  sky130_fd_sc_hd__a31oi_1 U26591 ( .A1(n20573), .A2(n20520), .A3(n20519), 
        .B1(n20663), .Y(n20539) );
  sky130_fd_sc_hd__nor2_1 U26592 ( .A(n20660), .B(n20659), .Y(n20524) );
  sky130_fd_sc_hd__nor2_1 U26593 ( .A(n20632), .B(n20521), .Y(n20522) );
  sky130_fd_sc_hd__a31oi_1 U26594 ( .A1(n20524), .A2(n20523), .A3(n20522), 
        .B1(n20681), .Y(n20537) );
  sky130_fd_sc_hd__nor3_1 U26595 ( .A(n20527), .B(n20526), .C(n20525), .Y(
        n20639) );
  sky130_fd_sc_hd__nor4_1 U26596 ( .A(n20647), .B(n20662), .C(n20646), .D(
        n20528), .Y(n20529) );
  sky130_fd_sc_hd__nand4_1 U26597 ( .A(n20532), .B(n20570), .C(n20531), .D(
        n20583), .Y(n20535) );
  sky130_fd_sc_hd__o21ai_1 U26598 ( .A1(n20535), .A2(n20534), .B1(n20533), .Y(
        n20536) );
  sky130_fd_sc_hd__nand3b_1 U26599 ( .A_N(n20537), .B(n20530), .C(n20536), .Y(
        n20538) );
  sky130_fd_sc_hd__nor2_1 U26600 ( .A(n20539), .B(n20538), .Y(n20540) );
  sky130_fd_sc_hd__mux2i_1 U26601 ( .A0(n20541), .A1(n20540), .S(n20623), .Y(
        n20542) );
  sky130_fd_sc_hd__nand2_1 U26602 ( .A(n20542), .B(n20693), .Y(n20556) );
  sky130_fd_sc_hd__nand2_1 U26603 ( .A(j202_soc_core_memory0_ram_dout0[16]), 
        .B(n21733), .Y(n20546) );
  sky130_fd_sc_hd__nand2_1 U26604 ( .A(j202_soc_core_memory0_ram_dout0[48]), 
        .B(n21604), .Y(n20545) );
  sky130_fd_sc_hd__nand2_1 U26605 ( .A(j202_soc_core_memory0_ram_dout0[304]), 
        .B(n21603), .Y(n20544) );
  sky130_fd_sc_hd__nand2_1 U26606 ( .A(n20549), .B(n20548), .Y(n20967) );
  sky130_fd_sc_hd__nand2_1 U26607 ( .A(j202_soc_core_memory0_ram_dout0[496]), 
        .B(n21771), .Y(n20559) );
  sky130_fd_sc_hd__and4_1 U26608 ( .A(n20553), .B(n21738), .C(n20552), .D(
        n20551), .X(n20554) );
  sky130_fd_sc_hd__and3_1 U26609 ( .A(n20556), .B(n20555), .C(n20554), .X(
        n20558) );
  sky130_fd_sc_hd__nand3_1 U26610 ( .A(n20559), .B(n20558), .C(n20557), .Y(
        n20987) );
  sky130_fd_sc_hd__nand2_1 U26611 ( .A(j202_soc_core_memory0_ram_dout0[305]), 
        .B(n21603), .Y(n20563) );
  sky130_fd_sc_hd__nand2_1 U26612 ( .A(j202_soc_core_memory0_ram_dout0[49]), 
        .B(n21604), .Y(n20567) );
  sky130_fd_sc_hd__nand2_1 U26613 ( .A(j202_soc_core_memory0_ram_dout0[337]), 
        .B(n21593), .Y(n20566) );
  sky130_fd_sc_hd__nand2_1 U26614 ( .A(j202_soc_core_memory0_ram_dout0[273]), 
        .B(n21605), .Y(n20565) );
  sky130_fd_sc_hd__nand2_1 U26615 ( .A(j202_soc_core_memory0_ram_dout0[401]), 
        .B(n21597), .Y(n20564) );
  sky130_fd_sc_hd__nand2_1 U26616 ( .A(j202_soc_core_memory0_ram_dout0[177]), 
        .B(n21590), .Y(n20696) );
  sky130_fd_sc_hd__a22oi_1 U26617 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[49]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[81]), .Y(n20700) );
  sky130_fd_sc_hd__nand2_1 U26618 ( .A(n21675), .B(j202_soc_core_uart_div1[1]), 
        .Y(n20699) );
  sky130_fd_sc_hd__nand2_1 U26619 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[17]), .Y(n20698) );
  sky130_fd_sc_hd__nand4_1 U26620 ( .A(n20700), .B(n21677), .C(n20699), .D(
        n20698), .Y(n20629) );
  sky130_fd_sc_hd__nand4_1 U26621 ( .A(n20571), .B(n20570), .C(n20569), .D(
        n20568), .Y(n20572) );
  sky130_fd_sc_hd__nor2b_1 U26622 ( .B_N(n20573), .A(n20572), .Y(n20581) );
  sky130_fd_sc_hd__nor4_1 U26623 ( .A(n20612), .B(n20678), .C(n20611), .D(
        n20631), .Y(n20575) );
  sky130_fd_sc_hd__nand4_1 U26624 ( .A(n20589), .B(n20576), .C(n20575), .D(
        n20574), .Y(n20577) );
  sky130_fd_sc_hd__nand2_1 U26625 ( .A(n20577), .B(n20692), .Y(n20578) );
  sky130_fd_sc_hd__o31ai_1 U26626 ( .A1(n20581), .A2(n20580), .A3(n20579), 
        .B1(n20578), .Y(n20628) );
  sky130_fd_sc_hd__nand2_1 U26627 ( .A(n20583), .B(n20582), .Y(n20587) );
  sky130_fd_sc_hd__nand4_1 U26628 ( .A(n20585), .B(n20615), .C(n20584), .D(
        n20614), .Y(n20586) );
  sky130_fd_sc_hd__nor4_1 U26629 ( .A(n20668), .B(n20667), .C(n20587), .D(
        n20586), .Y(n20588) );
  sky130_fd_sc_hd__a21oi_1 U26630 ( .A1(n20589), .A2(n20588), .B1(n20681), .Y(
        n20600) );
  sky130_fd_sc_hd__nor4_1 U26631 ( .A(n20593), .B(n20592), .C(n20591), .D(
        n20590), .Y(n20598) );
  sky130_fd_sc_hd__nor4_1 U26632 ( .A(n20668), .B(n20596), .C(n20595), .D(
        n20594), .Y(n20597) );
  sky130_fd_sc_hd__o22ai_1 U26633 ( .A1(n20598), .A2(n20683), .B1(n20597), 
        .B2(n20663), .Y(n20599) );
  sky130_fd_sc_hd__nor2_1 U26634 ( .A(n20600), .B(n20599), .Y(n20625) );
  sky130_fd_sc_hd__nand4_1 U26635 ( .A(n20603), .B(n20602), .C(n20601), .D(
        n20648), .Y(n20604) );
  sky130_fd_sc_hd__nor4_1 U26636 ( .A(n20606), .B(n20605), .C(n20618), .D(
        n20604), .Y(n20607) );
  sky130_fd_sc_hd__a31oi_1 U26637 ( .A1(n20609), .A2(n20608), .A3(n20607), 
        .B1(n20663), .Y(n20622) );
  sky130_fd_sc_hd__nor4b_1 U26638 ( .D_N(n20613), .A(n20612), .B(n20611), .C(
        n20610), .Y(n20620) );
  sky130_fd_sc_hd__nand2_1 U26639 ( .A(n20615), .B(n20614), .Y(n20616) );
  sky130_fd_sc_hd__nor4_1 U26640 ( .A(n20667), .B(n20618), .C(n20617), .D(
        n20616), .Y(n20619) );
  sky130_fd_sc_hd__o22ai_1 U26641 ( .A1(n20620), .A2(n20651), .B1(n20619), 
        .B2(n20681), .Y(n20621) );
  sky130_fd_sc_hd__nor2_1 U26642 ( .A(n20622), .B(n20621), .Y(n20624) );
  sky130_fd_sc_hd__mux2i_1 U26643 ( .A0(n20625), .A1(n20624), .S(n20623), .Y(
        n20627) );
  sky130_fd_sc_hd__o21a_1 U26644 ( .A1(n20628), .A2(n20627), .B1(n20626), .X(
        n20701) );
  sky130_fd_sc_hd__nor3_1 U26645 ( .A(n20703), .B(n20629), .C(n20701), .Y(
        n20695) );
  sky130_fd_sc_hd__a211oi_1 U26646 ( .A1(n20632), .A2(
        j202_soc_core_bootrom_00_address_w[4]), .B1(n20631), .C1(n20630), .Y(
        n20635) );
  sky130_fd_sc_hd__nand4b_1 U26647 ( .A_N(n20636), .B(n20635), .C(n20634), .D(
        n20633), .Y(n20691) );
  sky130_fd_sc_hd__a31oi_1 U26648 ( .A1(n20639), .A2(n20638), .A3(n20637), 
        .B1(n20683), .Y(n20658) );
  sky130_fd_sc_hd__nor3_1 U26649 ( .A(n20642), .B(n20641), .C(n20640), .Y(
        n20644) );
  sky130_fd_sc_hd__a31oi_1 U26650 ( .A1(n20672), .A2(n20644), .A3(n20643), 
        .B1(n20681), .Y(n20657) );
  sky130_fd_sc_hd__nor4_1 U26651 ( .A(n20647), .B(n20650), .C(n20646), .D(
        n20645), .Y(n20649) );
  sky130_fd_sc_hd__a21oi_1 U26652 ( .A1(n20649), .A2(n20648), .B1(n20663), .Y(
        n20656) );
  sky130_fd_sc_hd__a31oi_1 U26653 ( .A1(n20654), .A2(n20653), .A3(n20652), 
        .B1(n20651), .Y(n20655) );
  sky130_fd_sc_hd__nor4_1 U26654 ( .A(n20658), .B(n20657), .C(n20656), .D(
        n20655), .Y(n20689) );
  sky130_fd_sc_hd__nor4_1 U26655 ( .A(n20662), .B(n20661), .C(n20660), .D(
        n20659), .Y(n20666) );
  sky130_fd_sc_hd__a31oi_1 U26656 ( .A1(n20666), .A2(n20665), .A3(n20664), 
        .B1(n20663), .Y(n20686) );
  sky130_fd_sc_hd__nor2_1 U26657 ( .A(n20668), .B(n20667), .Y(n20670) );
  sky130_fd_sc_hd__nand4_1 U26658 ( .A(n20672), .B(n20671), .C(n20670), .D(
        n20669), .Y(n20673) );
  sky130_fd_sc_hd__nor4_1 U26659 ( .A(n20676), .B(n20675), .C(n20674), .D(
        n20673), .Y(n20684) );
  sky130_fd_sc_hd__nor4_1 U26660 ( .A(n20680), .B(n20679), .C(n20678), .D(
        n20677), .Y(n20682) );
  sky130_fd_sc_hd__o22ai_1 U26661 ( .A1(n20684), .A2(n20683), .B1(n20682), 
        .B2(n20681), .Y(n20685) );
  sky130_fd_sc_hd__nor2_1 U26662 ( .A(n20686), .B(n20685), .Y(n20688) );
  sky130_fd_sc_hd__mux2i_1 U26663 ( .A0(n20689), .A1(n20688), .S(n20687), .Y(
        n20690) );
  sky130_fd_sc_hd__a21o_1 U26664 ( .A1(n20692), .A2(n20691), .B1(n20690), .X(
        n20694) );
  sky130_fd_sc_hd__nand2_1 U26665 ( .A(n20694), .B(n20693), .Y(n20704) );
  sky130_fd_sc_hd__nand2_1 U26666 ( .A(j202_soc_core_memory0_ram_dout0[81]), 
        .B(n21734), .Y(n20697) );
  sky130_fd_sc_hd__nand2_1 U26667 ( .A(j202_soc_core_memory0_ram_dout0[497]), 
        .B(n21771), .Y(n20706) );
  sky130_fd_sc_hd__nand4_1 U26668 ( .A(n20700), .B(n21738), .C(n20699), .D(
        n20698), .Y(n20702) );
  sky130_fd_sc_hd__nor3_1 U26669 ( .A(n20703), .B(n20702), .C(n20701), .Y(
        n20705) );
  sky130_fd_sc_hd__nand3_1 U26670 ( .A(n20706), .B(n20705), .C(n20704), .Y(
        n21006) );
  sky130_fd_sc_hd__a22oi_1 U26671 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__1_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__1_), .Y(n20708) );
  sky130_fd_sc_hd__buf_2 U26672 ( .A(n22277), .X(n29071) );
  sky130_fd_sc_hd__a22oi_1 U26673 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__2_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__2_), .Y(n20713) );
  sky130_fd_sc_hd__a22oi_1 U26674 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__3_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__3_), .Y(n20722) );
  sky130_fd_sc_hd__nand2_1 U26675 ( .A(n20716), .B(n29572), .Y(n20721) );
  sky130_fd_sc_hd__a22oi_1 U26676 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__6_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__6_), .Y(n20834) );
  sky130_fd_sc_hd__nand2_1 U26677 ( .A(j202_soc_core_memory0_ram_dout0[134]), 
        .B(n21592), .Y(n20726) );
  sky130_fd_sc_hd__nand2_1 U26678 ( .A(j202_soc_core_memory0_ram_dout0[70]), 
        .B(n21734), .Y(n20725) );
  sky130_fd_sc_hd__nand2_1 U26679 ( .A(j202_soc_core_memory0_ram_dout0[166]), 
        .B(n21590), .Y(n20724) );
  sky130_fd_sc_hd__nand2_1 U26680 ( .A(j202_soc_core_memory0_ram_dout0[326]), 
        .B(n21593), .Y(n20723) );
  sky130_fd_sc_hd__nand4_1 U26681 ( .A(n20726), .B(n20725), .C(n20724), .D(
        n20723), .Y(n20732) );
  sky130_fd_sc_hd__nand2_1 U26682 ( .A(j202_soc_core_memory0_ram_dout0[358]), 
        .B(n21596), .Y(n20730) );
  sky130_fd_sc_hd__nand2_1 U26683 ( .A(j202_soc_core_memory0_ram_dout0[390]), 
        .B(n21597), .Y(n20729) );
  sky130_fd_sc_hd__nand2_1 U26684 ( .A(j202_soc_core_memory0_ram_dout0[454]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n20728) );
  sky130_fd_sc_hd__nand2_1 U26685 ( .A(j202_soc_core_memory0_ram_dout0[422]), 
        .B(n21598), .Y(n20727) );
  sky130_fd_sc_hd__nand4_1 U26686 ( .A(n20730), .B(n20729), .C(n20728), .D(
        n20727), .Y(n20731) );
  sky130_fd_sc_hd__nor2_1 U26687 ( .A(n20732), .B(n20731), .Y(n20827) );
  sky130_fd_sc_hd__nand2_1 U26688 ( .A(j202_soc_core_memory0_ram_dout0[262]), 
        .B(n21605), .Y(n20821) );
  sky130_fd_sc_hd__nand2_1 U26689 ( .A(j202_soc_core_memory0_ram_dout0[294]), 
        .B(n21603), .Y(n20820) );
  sky130_fd_sc_hd__nand2_1 U26690 ( .A(j202_soc_core_memory0_ram_dout0[38]), 
        .B(n21604), .Y(n20819) );
  sky130_fd_sc_hd__nand2_1 U26691 ( .A(n20736), .B(n21228), .Y(n21655) );
  sky130_fd_sc_hd__nor4_1 U26692 ( .A(n21285), .B(n20734), .C(n21655), .D(
        n20733), .Y(n20735) );
  sky130_fd_sc_hd__a31oi_1 U26693 ( .A1(n20735), .A2(n21706), .A3(n21270), 
        .B1(n21705), .Y(n20745) );
  sky130_fd_sc_hd__nor2_1 U26694 ( .A(n21715), .B(n21716), .Y(n20738) );
  sky130_fd_sc_hd__nor2_1 U26695 ( .A(n21627), .B(n21625), .Y(n20737) );
  sky130_fd_sc_hd__nand2_1 U26696 ( .A(n20736), .B(n21649), .Y(n20773) );
  sky130_fd_sc_hd__a31oi_1 U26697 ( .A1(n20738), .A2(n20737), .A3(n21132), 
        .B1(n21722), .Y(n20744) );
  sky130_fd_sc_hd__and3_1 U26698 ( .A(n21628), .B(n21613), .C(n20739), .X(
        n20740) );
  sky130_fd_sc_hd__a31oi_1 U26699 ( .A1(n20803), .A2(n20740), .A3(n21243), 
        .B1(n21709), .Y(n20743) );
  sky130_fd_sc_hd__a31oi_1 U26700 ( .A1(n20741), .A2(n21245), .A3(n21134), 
        .B1(n21720), .Y(n20742) );
  sky130_fd_sc_hd__nor4_1 U26701 ( .A(n20745), .B(n20744), .C(n20743), .D(
        n20742), .Y(n20746) );
  sky130_fd_sc_hd__nand2b_1 U26702 ( .A_N(n20746), .B(n21727), .Y(n20817) );
  sky130_fd_sc_hd__nand4_1 U26703 ( .A(n21243), .B(n21256), .C(n20747), .D(
        n21269), .Y(n20748) );
  sky130_fd_sc_hd__nor2_1 U26704 ( .A(n21618), .B(n20748), .Y(n20749) );
  sky130_fd_sc_hd__nand2_1 U26705 ( .A(n20750), .B(n20749), .Y(n20802) );
  sky130_fd_sc_hd__nand4_1 U26706 ( .A(n21648), .B(n20752), .C(n21081), .D(
        n20751), .Y(n20753) );
  sky130_fd_sc_hd__nor2_1 U26707 ( .A(n21201), .B(n20753), .Y(n21634) );
  sky130_fd_sc_hd__nand2_1 U26708 ( .A(n21634), .B(n21607), .Y(n20754) );
  sky130_fd_sc_hd__o2bb2ai_1 U26709 ( .B1(n20755), .B2(n21179), .A1_N(n20908), 
        .A2_N(n20754), .Y(n20756) );
  sky130_fd_sc_hd__nand2_1 U26710 ( .A(n20756), .B(n21636), .Y(n20771) );
  sky130_fd_sc_hd__nor2_1 U26711 ( .A(n20811), .B(n21207), .Y(n20757) );
  sky130_fd_sc_hd__nand4_1 U26712 ( .A(n20758), .B(n21258), .C(n20757), .D(
        n21270), .Y(n20768) );
  sky130_fd_sc_hd__nand3_1 U26713 ( .A(n20759), .B(n21288), .C(n13481), .Y(
        n20766) );
  sky130_fd_sc_hd__a22oi_1 U26714 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[38]), .B1(n21698), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[102]), .Y(n20765) );
  sky130_fd_sc_hd__a22oi_1 U26715 ( .A1(n21676), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[6]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[70]), .Y(n20764) );
  sky130_fd_sc_hd__a22oi_1 U26716 ( .A1(n24376), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[22]), .B1(n21669), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[30]), .Y(n20761) );
  sky130_fd_sc_hd__a22oi_1 U26717 ( .A1(n21667), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[14]), .B1(n21668), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[6]), .Y(n20760) );
  sky130_fd_sc_hd__nand2_1 U26718 ( .A(n20761), .B(n20760), .Y(n20762) );
  sky130_fd_sc_hd__nand2_1 U26719 ( .A(n20762), .B(n21675), .Y(n20763) );
  sky130_fd_sc_hd__nand4_1 U26720 ( .A(n20766), .B(n20765), .C(n20764), .D(
        n20763), .Y(n20767) );
  sky130_fd_sc_hd__a21oi_1 U26721 ( .A1(n20768), .A2(n21198), .B1(n20767), .Y(
        n20770) );
  sky130_fd_sc_hd__nand2_1 U26722 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_period[6]), .Y(n20769) );
  sky130_fd_sc_hd__nand3_1 U26723 ( .A(n20771), .B(n20770), .C(n20769), .Y(
        n20799) );
  sky130_fd_sc_hd__nand3_1 U26724 ( .A(n21081), .B(n20784), .C(n20772), .Y(
        n20774) );
  sky130_fd_sc_hd__nor2_1 U26725 ( .A(n20774), .B(n20773), .Y(n20775) );
  sky130_fd_sc_hd__nand2_1 U26726 ( .A(n20775), .B(n21687), .Y(n20776) );
  sky130_fd_sc_hd__nand2_1 U26727 ( .A(n20776), .B(n21288), .Y(n20782) );
  sky130_fd_sc_hd__nor2_1 U26728 ( .A(n20778), .B(n20777), .Y(n20779) );
  sky130_fd_sc_hd__nand3_1 U26729 ( .A(n12180), .B(n21710), .C(n20779), .Y(
        n20780) );
  sky130_fd_sc_hd__nand2_1 U26730 ( .A(n20780), .B(n21251), .Y(n20781) );
  sky130_fd_sc_hd__a31oi_1 U26731 ( .A1(n20783), .A2(n20782), .A3(n20781), 
        .B1(n21124), .Y(n20798) );
  sky130_fd_sc_hd__nand3_1 U26732 ( .A(n20785), .B(n21608), .C(n20784), .Y(
        n20786) );
  sky130_fd_sc_hd__o21ai_0 U26733 ( .A1(n21626), .A2(n20786), .B1(n21235), .Y(
        n20796) );
  sky130_fd_sc_hd__nand2_1 U26734 ( .A(n20788), .B(n20787), .Y(n20789) );
  sky130_fd_sc_hd__nor2_1 U26736 ( .A(n20791), .B(n21717), .Y(n20792) );
  sky130_fd_sc_hd__nand2_1 U26737 ( .A(n21082), .B(n20792), .Y(n20793) );
  sky130_fd_sc_hd__o21ai_0 U26738 ( .A1(n20793), .A2(n21626), .B1(n21251), .Y(
        n20795) );
  sky130_fd_sc_hd__a21oi_1 U26739 ( .A1(n20796), .A2(n20795), .B1(n20794), .Y(
        n20797) );
  sky130_fd_sc_hd__nor3_1 U26740 ( .A(n20799), .B(n20798), .C(n20797), .Y(
        n20800) );
  sky130_fd_sc_hd__nand3_1 U26741 ( .A(n20803), .B(n21614), .C(n21681), .Y(
        n21624) );
  sky130_fd_sc_hd__a21bo_2 U26742 ( .A1(n20806), .A2(n20807), .B1_N(n20805), 
        .X(n21264) );
  sky130_fd_sc_hd__a21oi_1 U26743 ( .A1(n20807), .A2(n12181), .B1(n21264), .Y(
        n21101) );
  sky130_fd_sc_hd__nand2_1 U26744 ( .A(n20808), .B(n21101), .Y(n20809) );
  sky130_fd_sc_hd__o21ai_1 U26745 ( .A1(n21624), .A2(n20809), .B1(n21697), .Y(
        n20813) );
  sky130_fd_sc_hd__o21ai_1 U26746 ( .A1(n20811), .A2(n20810), .B1(n13481), .Y(
        n20812) );
  sky130_fd_sc_hd__nand2_1 U26747 ( .A(n20813), .B(n20812), .Y(n20814) );
  sky130_fd_sc_hd__nand2_1 U26748 ( .A(n20814), .B(n21235), .Y(n20815) );
  sky130_fd_sc_hd__nand3_1 U26749 ( .A(n20817), .B(n20816), .C(n20815), .Y(
        n20828) );
  sky130_fd_sc_hd__nor2_1 U26750 ( .A(j202_soc_core_memory0_ram_dout0_sel[15]), 
        .B(n20828), .Y(n20818) );
  sky130_fd_sc_hd__and4_1 U26751 ( .A(n20821), .B(n20820), .C(n20819), .D(
        n20818), .X(n20826) );
  sky130_fd_sc_hd__nand2_1 U26752 ( .A(j202_soc_core_memory0_ram_dout0[198]), 
        .B(n21732), .Y(n20825) );
  sky130_fd_sc_hd__nand2_1 U26753 ( .A(j202_soc_core_memory0_ram_dout0[230]), 
        .B(n21735), .Y(n20824) );
  sky130_fd_sc_hd__nand2_1 U26754 ( .A(j202_soc_core_memory0_ram_dout0[6]), 
        .B(n21733), .Y(n20823) );
  sky130_fd_sc_hd__nand2_1 U26755 ( .A(j202_soc_core_memory0_ram_dout0[102]), 
        .B(n21591), .Y(n20822) );
  sky130_fd_sc_hd__nand2_1 U26756 ( .A(n20831), .B(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n20829) );
  sky130_fd_sc_hd__a2bb2oi_1 U26757 ( .B1(n20831), .B2(n20830), .A1_N(n20829), 
        .A2_N(j202_soc_core_memory0_ram_dout0[486]), .Y(n21520) );
  sky130_fd_sc_hd__a22oi_1 U26758 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__8_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__8_), .Y(n20836) );
  sky130_fd_sc_hd__a22oi_1 U26759 ( .A1(j202_soc_core_memory0_ram_dout0[329]), 
        .A2(n21593), .B1(n21605), .B2(j202_soc_core_memory0_ram_dout0[265]), 
        .Y(n20935) );
  sky130_fd_sc_hd__nor3_1 U26760 ( .A(n20838), .B(n20870), .C(n20837), .Y(
        n20856) );
  sky130_fd_sc_hd__nor3_1 U26761 ( .A(n20898), .B(n20869), .C(n20839), .Y(
        n20840) );
  sky130_fd_sc_hd__a21oi_1 U26762 ( .A1(n20841), .A2(n20840), .B1(n20925), .Y(
        n20848) );
  sky130_fd_sc_hd__nand3_1 U26763 ( .A(n20844), .B(n20843), .C(n20842), .Y(
        n20846) );
  sky130_fd_sc_hd__o21a_1 U26764 ( .A1(n20846), .A2(n20845), .B1(n20912), .X(
        n20847) );
  sky130_fd_sc_hd__nor2_1 U26765 ( .A(n20848), .B(n20847), .Y(n20855) );
  sky130_fd_sc_hd__nand2_1 U26766 ( .A(n20850), .B(n20849), .Y(n20851) );
  sky130_fd_sc_hd__nor4_1 U26767 ( .A(n20898), .B(n20911), .C(n20852), .D(
        n20851), .Y(n20853) );
  sky130_fd_sc_hd__nand2b_1 U26768 ( .A_N(n20853), .B(n20864), .Y(n20854) );
  sky130_fd_sc_hd__o211ai_1 U26769 ( .A1(n20856), .A2(n20873), .B1(n20855), 
        .C1(n20854), .Y(n20857) );
  sky130_fd_sc_hd__nand2_1 U26770 ( .A(n20857), .B(n21727), .Y(n20949) );
  sky130_fd_sc_hd__nor2_1 U26771 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[0]), 
        .B(n28753), .Y(n20858) );
  sky130_fd_sc_hd__xor2_1 U26772 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[1]), 
        .B(j202_soc_core_uart_TOP_tx_fifo_wp[1]), .X(n24698) );
  sky130_fd_sc_hd__nor2_1 U26773 ( .A(n20858), .B(n24698), .Y(n27993) );
  sky130_fd_sc_hd__nand2_1 U26774 ( .A(n28753), .B(
        j202_soc_core_uart_TOP_tx_fifo_wp[0]), .Y(n27991) );
  sky130_fd_sc_hd__nand3_1 U26775 ( .A(n27993), .B(
        j202_soc_core_uart_TOP_tx_fifo_gb), .C(n27991), .Y(n20859) );
  sky130_fd_sc_hd__a2bb2oi_1 U26776 ( .B1(
        j202_soc_core_ahblite_interconnect_s_hrdata[105]), .B2(n21698), .A1_N(
        n20860), .A2_N(n20859), .Y(n20945) );
  sky130_fd_sc_hd__a22oi_1 U26777 ( .A1(n21676), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[9]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[73]), .Y(n20944) );
  sky130_fd_sc_hd__nand2_1 U26778 ( .A(n21699), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[41]), .Y(n20943) );
  sky130_fd_sc_hd__and4_1 U26779 ( .A(n20945), .B(n20944), .C(n21677), .D(
        n20943), .X(n20880) );
  sky130_fd_sc_hd__nor4_1 U26780 ( .A(n20863), .B(n20862), .C(n20861), .D(
        n20923), .Y(n20868) );
  sky130_fd_sc_hd__o21ai_0 U26782 ( .A1(n20868), .A2(n20906), .B1(n20867), .Y(
        n20878) );
  sky130_fd_sc_hd__nor4_1 U26783 ( .A(n20872), .B(n20871), .C(n20870), .D(
        n20869), .Y(n20874) );
  sky130_fd_sc_hd__a21o_1 U26784 ( .A1(n20875), .A2(n20874), .B1(n20873), .X(
        n20876) );
  sky130_fd_sc_hd__nand3b_1 U26785 ( .A_N(n20878), .B(n20877), .C(n20876), .Y(
        n20879) );
  sky130_fd_sc_hd__nand2_1 U26786 ( .A(n20879), .B(n13481), .Y(n20947) );
  sky130_fd_sc_hd__nand2_1 U26787 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_period[9]), .Y(n20946) );
  sky130_fd_sc_hd__nand4_1 U26788 ( .A(n20949), .B(n20880), .C(n20947), .D(
        n20946), .Y(n20931) );
  sky130_fd_sc_hd__nor4_1 U26789 ( .A(n20883), .B(n20904), .C(n20882), .D(
        n20881), .Y(n20895) );
  sky130_fd_sc_hd__nand2_1 U26790 ( .A(n20885), .B(n20919), .Y(n20886) );
  sky130_fd_sc_hd__nor4_1 U26791 ( .A(n20916), .B(n20888), .C(n20887), .D(
        n20886), .Y(n20889) );
  sky130_fd_sc_hd__nand4_1 U26792 ( .A(n13302), .B(n20891), .C(n20890), .D(
        n20889), .Y(n20893) );
  sky130_fd_sc_hd__nand2_1 U26793 ( .A(n20893), .B(n20892), .Y(n20894) );
  sky130_fd_sc_hd__nand3b_1 U26795 ( .A_N(n20898), .B(n20897), .C(n20896), .Y(
        n20899) );
  sky130_fd_sc_hd__nor4_1 U26796 ( .A(n20901), .B(n20923), .C(n20900), .D(
        n20899), .Y(n20907) );
  sky130_fd_sc_hd__nor3_1 U26797 ( .A(n20904), .B(n20903), .C(n20902), .Y(
        n20905) );
  sky130_fd_sc_hd__o22ai_1 U26798 ( .A1(n20907), .A2(n20906), .B1(n20905), 
        .B2(n20927), .Y(n20909) );
  sky130_fd_sc_hd__o21a_1 U26799 ( .A1(n20910), .A2(n20909), .B1(n20908), .X(
        n20951) );
  sky130_fd_sc_hd__nand2_1 U26800 ( .A(n20912), .B(n20911), .Y(n20913) );
  sky130_fd_sc_hd__nand2_1 U26801 ( .A(n20914), .B(n20913), .Y(n20930) );
  sky130_fd_sc_hd__nor4_1 U26802 ( .A(n20918), .B(n20917), .C(n20916), .D(
        n20915), .Y(n20928) );
  sky130_fd_sc_hd__nand2_1 U26803 ( .A(n20920), .B(n20919), .Y(n20921) );
  sky130_fd_sc_hd__nor4_1 U26804 ( .A(n20924), .B(n20923), .C(n20922), .D(
        n20921), .Y(n20926) );
  sky130_fd_sc_hd__o22ai_1 U26805 ( .A1(n20928), .A2(n20927), .B1(n20926), 
        .B2(n20925), .Y(n20929) );
  sky130_fd_sc_hd__o21a_1 U26806 ( .A1(n20930), .A2(n20929), .B1(n21697), .X(
        n20950) );
  sky130_fd_sc_hd__nor3_1 U26807 ( .A(n20931), .B(n20951), .C(n20950), .Y(
        n20932) );
  sky130_fd_sc_hd__nand4_1 U26808 ( .A(n20935), .B(n20936), .C(n20934), .D(
        n20933), .Y(n20937) );
  sky130_fd_sc_hd__inv_1 U26809 ( .A(n20937), .Y(n20956) );
  sky130_fd_sc_hd__a22oi_1 U26810 ( .A1(j202_soc_core_memory0_ram_dout0[9]), 
        .A2(n21733), .B1(n21603), .B2(j202_soc_core_memory0_ram_dout0[297]), 
        .Y(n20941) );
  sky130_fd_sc_hd__a22oi_1 U26811 ( .A1(j202_soc_core_memory0_ram_dout0[41]), 
        .A2(n21604), .B1(n21590), .B2(j202_soc_core_memory0_ram_dout0[169]), 
        .Y(n20940) );
  sky130_fd_sc_hd__nand4_1 U26812 ( .A(n20941), .B(n20940), .C(n20939), .D(
        n20938), .Y(n20942) );
  sky130_fd_sc_hd__nand2_1 U26813 ( .A(j202_soc_core_memory0_ram_dout0[489]), 
        .B(n21771), .Y(n20954) );
  sky130_fd_sc_hd__and4_1 U26814 ( .A(n20945), .B(n20944), .C(n21738), .D(
        n20943), .X(n20948) );
  sky130_fd_sc_hd__nand4_1 U26815 ( .A(n20949), .B(n20948), .C(n20947), .D(
        n20946), .Y(n20952) );
  sky130_fd_sc_hd__nor3_1 U26816 ( .A(n20952), .B(n20951), .C(n20950), .Y(
        n20953) );
  sky130_fd_sc_hd__nand2_1 U26817 ( .A(n28970), .B(n21750), .Y(n20959) );
  sky130_fd_sc_hd__a22oi_1 U26818 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__9_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__9_), .Y(n20958) );
  sky130_fd_sc_hd__nand2_1 U26819 ( .A(n12743), .B(n21776), .Y(n20957) );
  sky130_fd_sc_hd__a22oi_1 U26820 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__10_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__10_), .Y(n20961) );
  sky130_fd_sc_hd__a22oi_1 U26821 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__11_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__11_), .Y(n20963) );
  sky130_fd_sc_hd__nand2_1 U26822 ( .A(j202_soc_core_j22_cpu_id_op2_v_), .B(
        j202_soc_core_j22_cpu_id_op2_inst__12_), .Y(n20968) );
  sky130_fd_sc_hd__nand2_1 U26823 ( .A(n20967), .B(n20968), .Y(n20971) );
  sky130_fd_sc_hd__nand2_1 U26824 ( .A(n21775), .B(
        j202_soc_core_j22_cpu_id_opn_inst__12_), .Y(n20975) );
  sky130_fd_sc_hd__nor3_1 U26825 ( .A(n25881), .B(n24123), .C(n20978), .Y(
        n20981) );
  sky130_fd_sc_hd__xnor2_1 U26826 ( .A(n20979), .B(n12400), .Y(n25224) );
  sky130_fd_sc_hd__and3_1 U26827 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[2]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_sck), .C(n12142), .X(n28642) );
  sky130_fd_sc_hd__nand2_1 U26828 ( .A(n28642), .B(
        j202_soc_core_wbqspiflash_00_lldriver_state[0]), .Y(n28747) );
  sky130_fd_sc_hd__nand3_1 U26829 ( .A(n28642), .B(n20984), .C(n26261), .Y(
        n26225) );
  sky130_fd_sc_hd__nand2_1 U26830 ( .A(n25944), .B(
        j202_soc_core_wbqspiflash_00_spi_wr), .Y(n26198) );
  sky130_fd_sc_hd__nor2_1 U26831 ( .A(n28649), .B(n26198), .Y(n28637) );
  sky130_fd_sc_hd__nand2_1 U26832 ( .A(n23907), .B(n20984), .Y(n26260) );
  sky130_fd_sc_hd__nor2_1 U26833 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[2]), .B(n20984), .Y(n28638) );
  sky130_fd_sc_hd__nand3_1 U26834 ( .A(n28638), .B(n12142), .C(n26261), .Y(
        n26202) );
  sky130_fd_sc_hd__o211ai_1 U26835 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .A2(n28747), .B1(
        n20985), .C1(n26209), .Y(n29091) );
  sky130_fd_sc_hd__nand3_1 U26836 ( .A(n24814), .B(n20986), .C(
        j202_soc_core_ahb2apb_00_state[1]), .Y(n24818) );
  sky130_fd_sc_hd__nand2_1 U26837 ( .A(n24817), .B(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[0]), .Y(n24810) );
  sky130_fd_sc_hd__nor2_1 U26838 ( .A(n24818), .B(n24810), .Y(n28969) );
  sky130_fd_sc_hd__nand2_1 U26840 ( .A(n22321), .B(n20990), .Y(n21319) );
  sky130_fd_sc_hd__nand2_1 U26841 ( .A(n21341), .B(n20992), .Y(n22509) );
  sky130_fd_sc_hd__nor2_1 U26842 ( .A(n19063), .B(n22509), .Y(n20993) );
  sky130_fd_sc_hd__xnor2_1 U26843 ( .A(n20994), .B(n20993), .Y(n25261) );
  sky130_fd_sc_hd__nand2_1 U26844 ( .A(n22596), .B(n25261), .Y(n20996) );
  sky130_fd_sc_hd__nand2_1 U26845 ( .A(n22515), .B(n27447), .Y(n20995) );
  sky130_fd_sc_hd__a21oi_1 U26846 ( .A1(n22513), .A2(n22512), .B1(n20998), .Y(
        n21003) );
  sky130_fd_sc_hd__nand2_1 U26847 ( .A(n21001), .B(n21000), .Y(n21002) );
  sky130_fd_sc_hd__xor2_1 U26848 ( .A(n21003), .B(n21002), .X(n23996) );
  sky130_fd_sc_hd__nand2_1 U26849 ( .A(n23996), .B(n12158), .Y(n21004) );
  sky130_fd_sc_hd__nand3_1 U26850 ( .A(n21005), .B(n12213), .C(n21004), .Y(
        n28946) );
  sky130_fd_sc_hd__nand2b_1 U26851 ( .A_N(n26524), .B(n22581), .Y(n21021) );
  sky130_fd_sc_hd__xor2_1 U26852 ( .A(n21009), .B(n21008), .X(n25715) );
  sky130_fd_sc_hd__nand2_1 U26853 ( .A(n22596), .B(n25715), .Y(n21011) );
  sky130_fd_sc_hd__nand2_1 U26854 ( .A(n22515), .B(n24613), .Y(n21010) );
  sky130_fd_sc_hd__o211a_2 U26855 ( .A1(n25128), .A2(n11143), .B1(n21011), 
        .C1(n21010), .X(n21020) );
  sky130_fd_sc_hd__a21oi_1 U26856 ( .A1(n22513), .A2(n21013), .B1(n21012), .Y(
        n21018) );
  sky130_fd_sc_hd__nand2_1 U26857 ( .A(n21016), .B(n21015), .Y(n21017) );
  sky130_fd_sc_hd__xor2_1 U26858 ( .A(n21018), .B(n21017), .X(n24626) );
  sky130_fd_sc_hd__nand2_1 U26859 ( .A(n24626), .B(n12158), .Y(n21019) );
  sky130_fd_sc_hd__nand3_1 U26860 ( .A(n21021), .B(n21020), .C(n21019), .Y(
        n28922) );
  sky130_fd_sc_hd__nand4_1 U26861 ( .A(n21025), .B(n28919), .C(n21024), .D(
        n21023), .Y(n21029) );
  sky130_fd_sc_hd__nand2_1 U26862 ( .A(n21027), .B(n21026), .Y(n21028) );
  sky130_fd_sc_hd__nand3_1 U26863 ( .A(n22672), .B(n22671), .C(n28946), .Y(
        n21030) );
  sky130_fd_sc_hd__nor2_1 U26864 ( .A(j202_soc_core_wbqspiflash_00_state[3]), 
        .B(j202_soc_core_wbqspiflash_00_state[1]), .Y(n25916) );
  sky130_fd_sc_hd__nand2_1 U26865 ( .A(j202_soc_core_wbqspiflash_00_state[2]), 
        .B(j202_soc_core_wbqspiflash_00_state[4]), .Y(n25928) );
  sky130_fd_sc_hd__nand2_1 U26866 ( .A(n25916), .B(n26161), .Y(n28232) );
  sky130_fd_sc_hd__nand2_1 U26867 ( .A(n28232), .B(n29594), .Y(n28968) );
  sky130_fd_sc_hd__nand2_1 U26868 ( .A(j202_soc_core_memory0_ram_dout0[366]), 
        .B(n21596), .Y(n21034) );
  sky130_fd_sc_hd__nand2_1 U26869 ( .A(j202_soc_core_memory0_ram_dout0[334]), 
        .B(n21593), .Y(n21033) );
  sky130_fd_sc_hd__nand2_1 U26870 ( .A(j202_soc_core_memory0_ram_dout0[270]), 
        .B(n21605), .Y(n21032) );
  sky130_fd_sc_hd__nand2_1 U26871 ( .A(j202_soc_core_memory0_ram_dout0[398]), 
        .B(n21597), .Y(n21031) );
  sky130_fd_sc_hd__nand2_1 U26872 ( .A(j202_soc_core_memory0_ram_dout0[238]), 
        .B(n21735), .Y(n21038) );
  sky130_fd_sc_hd__nand2_1 U26873 ( .A(j202_soc_core_memory0_ram_dout0[14]), 
        .B(n21733), .Y(n21037) );
  sky130_fd_sc_hd__nand2_1 U26874 ( .A(j202_soc_core_memory0_ram_dout0[302]), 
        .B(n21603), .Y(n21036) );
  sky130_fd_sc_hd__nand2_1 U26875 ( .A(j202_soc_core_memory0_ram_dout0[46]), 
        .B(n21604), .Y(n21035) );
  sky130_fd_sc_hd__nand2_1 U26876 ( .A(j202_soc_core_memory0_ram_dout0[174]), 
        .B(n21590), .Y(n21143) );
  sky130_fd_sc_hd__nor4_1 U26877 ( .A(n21041), .B(n21040), .C(n21108), .D(
        n21039), .Y(n21048) );
  sky130_fd_sc_hd__nand2_1 U26878 ( .A(n21243), .B(n21228), .Y(n21176) );
  sky130_fd_sc_hd__nand2_1 U26879 ( .A(n21094), .B(n21267), .Y(n21227) );
  sky130_fd_sc_hd__nor4b_1 U26880 ( .D_N(n21136), .A(n21046), .B(n21045), .C(
        n21044), .Y(n21047) );
  sky130_fd_sc_hd__o22ai_1 U26881 ( .A1(n21048), .A2(n21722), .B1(n21047), 
        .B2(n21705), .Y(n21059) );
  sky130_fd_sc_hd__nand4_1 U26882 ( .A(n21050), .B(n21187), .C(n21049), .D(
        n21229), .Y(n21057) );
  sky130_fd_sc_hd__nor2_1 U26883 ( .A(n21051), .B(n21070), .Y(n21211) );
  sky130_fd_sc_hd__nand4_1 U26884 ( .A(n21190), .B(n21094), .C(n21286), .D(
        n21228), .Y(n21052) );
  sky130_fd_sc_hd__nor4_1 U26885 ( .A(n21054), .B(n21715), .C(n21053), .D(
        n21052), .Y(n21055) );
  sky130_fd_sc_hd__a31oi_1 U26886 ( .A1(n21211), .A2(n21191), .A3(n21055), 
        .B1(n21709), .Y(n21056) );
  sky130_fd_sc_hd__a21oi_1 U26887 ( .A1(n21288), .A2(n21057), .B1(n21056), .Y(
        n21058) );
  sky130_fd_sc_hd__nand2b_1 U26888 ( .A_N(n21059), .B(n21058), .Y(n21060) );
  sky130_fd_sc_hd__nand2_1 U26889 ( .A(n21060), .B(n13481), .Y(n21158) );
  sky130_fd_sc_hd__a22oi_1 U26890 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[46]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[78]), .Y(n21152) );
  sky130_fd_sc_hd__nand2_1 U26891 ( .A(n21698), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[110]), .Y(n21151) );
  sky130_fd_sc_hd__nand2_1 U26892 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[14]), .Y(n21150) );
  sky130_fd_sc_hd__nand4_1 U26893 ( .A(n21152), .B(n21677), .C(n21151), .D(
        n21150), .Y(n21065) );
  sky130_fd_sc_hd__nand2_1 U26894 ( .A(n21228), .B(n21650), .Y(n21062) );
  sky130_fd_sc_hd__nand2_1 U26895 ( .A(n21081), .B(n21186), .Y(n21653) );
  sky130_fd_sc_hd__nor2_1 U26896 ( .A(n21062), .B(n21653), .Y(n21064) );
  sky130_fd_sc_hd__nor2_1 U26897 ( .A(n21065), .B(n21153), .Y(n21092) );
  sky130_fd_sc_hd__nand3_1 U26898 ( .A(n21068), .B(n21221), .C(n21649), .Y(
        n21066) );
  sky130_fd_sc_hd__nor2_1 U26899 ( .A(n21224), .B(n21066), .Y(n21217) );
  sky130_fd_sc_hd__o21ai_0 U26900 ( .A1(n21188), .A2(n21067), .B1(n21288), .Y(
        n21090) );
  sky130_fd_sc_hd__nor2_1 U26901 ( .A(n21108), .B(n21069), .Y(n21135) );
  sky130_fd_sc_hd__nor2_1 U26902 ( .A(n21071), .B(n21070), .Y(n21074) );
  sky130_fd_sc_hd__nand2_1 U26903 ( .A(n21206), .B(n21219), .Y(n21072) );
  sky130_fd_sc_hd__nor2_1 U26904 ( .A(n21072), .B(n21207), .Y(n21073) );
  sky130_fd_sc_hd__nand4_1 U26905 ( .A(n21135), .B(n21075), .C(n21074), .D(
        n21073), .Y(n21076) );
  sky130_fd_sc_hd__nand2_1 U26906 ( .A(n21076), .B(n21251), .Y(n21089) );
  sky130_fd_sc_hd__and3_1 U26907 ( .A(n21078), .B(n21077), .C(n21287), .X(
        n21647) );
  sky130_fd_sc_hd__nor2_1 U26908 ( .A(n21176), .B(n21620), .Y(n21223) );
  sky130_fd_sc_hd__nand4_1 U26909 ( .A(n21647), .B(n21079), .C(n21223), .D(
        n21221), .Y(n21080) );
  sky130_fd_sc_hd__nand2_1 U26910 ( .A(n21080), .B(n21636), .Y(n21088) );
  sky130_fd_sc_hd__nand4_1 U26911 ( .A(n21229), .B(n21606), .C(n21681), .D(
        n21081), .Y(n21083) );
  sky130_fd_sc_hd__nand2_1 U26912 ( .A(n21082), .B(n21228), .Y(n21131) );
  sky130_fd_sc_hd__nor2_1 U26913 ( .A(n21083), .B(n21131), .Y(n21085) );
  sky130_fd_sc_hd__nand2_1 U26914 ( .A(n21085), .B(n21084), .Y(n21086) );
  sky130_fd_sc_hd__nand2_1 U26915 ( .A(n21086), .B(n21235), .Y(n21087) );
  sky130_fd_sc_hd__nand4_1 U26916 ( .A(n21090), .B(n21089), .C(n21088), .D(
        n21087), .Y(n21091) );
  sky130_fd_sc_hd__nand2_1 U26917 ( .A(n21091), .B(n21727), .Y(n21156) );
  sky130_fd_sc_hd__nand2_1 U26918 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_duty[2]), .Y(n21155) );
  sky130_fd_sc_hd__nand4_1 U26919 ( .A(n21158), .B(n21092), .C(n21156), .D(
        n21155), .Y(n21125) );
  sky130_fd_sc_hd__nand2b_1 U26920 ( .A_N(n21095), .B(n21094), .Y(n21214) );
  sky130_fd_sc_hd__nor4_1 U26921 ( .A(n21098), .B(n21097), .C(n21096), .D(
        n21214), .Y(n21099) );
  sky130_fd_sc_hd__a31oi_1 U26922 ( .A1(n21101), .A2(n21100), .A3(n21099), 
        .B1(n21705), .Y(n21122) );
  sky130_fd_sc_hd__nor2_1 U26923 ( .A(n21715), .B(n21653), .Y(n21107) );
  sky130_fd_sc_hd__nand3_1 U26924 ( .A(n21687), .B(n21688), .C(n21103), .Y(
        n21259) );
  sky130_fd_sc_hd__nor4_1 U26925 ( .A(n21207), .B(n21643), .C(n21104), .D(
        n21201), .Y(n21105) );
  sky130_fd_sc_hd__a31oi_1 U26926 ( .A1(n21107), .A2(n21106), .A3(n21105), 
        .B1(n21720), .Y(n21121) );
  sky130_fd_sc_hd__nor2_1 U26927 ( .A(n21109), .B(n21620), .Y(n21110) );
  sky130_fd_sc_hd__nand3_1 U26928 ( .A(n21111), .B(n21110), .C(n21221), .Y(
        n21289) );
  sky130_fd_sc_hd__nor4_1 U26929 ( .A(n21657), .B(n21113), .C(n21289), .D(
        n21112), .Y(n21119) );
  sky130_fd_sc_hd__nor3_1 U26930 ( .A(n21714), .B(n21115), .C(n21114), .Y(
        n21128) );
  sky130_fd_sc_hd__nor4b_1 U26931 ( .D_N(n21128), .A(n21265), .B(n21117), .C(
        n21116), .Y(n21118) );
  sky130_fd_sc_hd__o22ai_1 U26932 ( .A1(n21119), .A2(n21722), .B1(n21118), 
        .B2(n21709), .Y(n21120) );
  sky130_fd_sc_hd__nor3_1 U26933 ( .A(n21122), .B(n21121), .C(n21120), .Y(
        n21123) );
  sky130_fd_sc_hd__nor2_1 U26934 ( .A(n21124), .B(n21123), .Y(n21159) );
  sky130_fd_sc_hd__nor2_1 U26935 ( .A(n21125), .B(n21159), .Y(n21142) );
  sky130_fd_sc_hd__nor3_1 U26936 ( .A(n21126), .B(n21618), .C(n21131), .Y(
        n21127) );
  sky130_fd_sc_hd__a31oi_1 U26937 ( .A1(n21129), .A2(n21128), .A3(n21127), 
        .B1(n21709), .Y(n21140) );
  sky130_fd_sc_hd__nand2_1 U26938 ( .A(n21630), .B(n21631), .Y(n21611) );
  sky130_fd_sc_hd__a31oi_1 U26939 ( .A1(n21132), .A2(n21281), .A3(n21134), 
        .B1(n21722), .Y(n21139) );
  sky130_fd_sc_hd__nand2_1 U26940 ( .A(n21253), .B(n21134), .Y(n21656) );
  sky130_fd_sc_hd__a31oi_1 U26941 ( .A1(n21136), .A2(n21257), .A3(n21135), 
        .B1(n21720), .Y(n21137) );
  sky130_fd_sc_hd__nor4_1 U26942 ( .A(n21140), .B(n21139), .C(n21138), .D(
        n21137), .Y(n21141) );
  sky130_fd_sc_hd__nand2_1 U26943 ( .A(j202_soc_core_memory0_ram_dout0[142]), 
        .B(n21592), .Y(n21145) );
  sky130_fd_sc_hd__nand2_1 U26944 ( .A(j202_soc_core_memory0_ram_dout0[78]), 
        .B(n21734), .Y(n21144) );
  sky130_fd_sc_hd__nand2_1 U26945 ( .A(j202_soc_core_memory0_ram_dout0[206]), 
        .B(n21732), .Y(n21149) );
  sky130_fd_sc_hd__nand2_1 U26946 ( .A(j202_soc_core_memory0_ram_dout0[110]), 
        .B(n21591), .Y(n21148) );
  sky130_fd_sc_hd__nand2_1 U26947 ( .A(j202_soc_core_memory0_ram_dout0[462]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n21147) );
  sky130_fd_sc_hd__nand2_1 U26948 ( .A(j202_soc_core_memory0_ram_dout0[430]), 
        .B(n21598), .Y(n21146) );
  sky130_fd_sc_hd__nand2_1 U26949 ( .A(j202_soc_core_memory0_ram_dout0[494]), 
        .B(n21771), .Y(n21163) );
  sky130_fd_sc_hd__nand4_1 U26950 ( .A(n21152), .B(n21738), .C(n21151), .D(
        n21150), .Y(n21154) );
  sky130_fd_sc_hd__nor2_1 U26951 ( .A(n21154), .B(n21153), .Y(n21157) );
  sky130_fd_sc_hd__nand4_1 U26952 ( .A(n21158), .B(n21157), .C(n21156), .D(
        n21155), .Y(n21160) );
  sky130_fd_sc_hd__nor2_1 U26953 ( .A(n21160), .B(n21159), .Y(n21162) );
  sky130_fd_sc_hd__nand3_1 U26954 ( .A(n21163), .B(n21162), .C(n21161), .Y(
        n21317) );
  sky130_fd_sc_hd__a22oi_1 U26955 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__13_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__13_), .Y(n21316) );
  sky130_fd_sc_hd__nand2_1 U26956 ( .A(j202_soc_core_memory0_ram_dout0[365]), 
        .B(n21596), .Y(n21168) );
  sky130_fd_sc_hd__nand2_1 U26957 ( .A(j202_soc_core_memory0_ram_dout0[397]), 
        .B(n21597), .Y(n21167) );
  sky130_fd_sc_hd__nand2_1 U26958 ( .A(j202_soc_core_memory0_ram_dout0[333]), 
        .B(n21593), .Y(n21295) );
  sky130_fd_sc_hd__o21a_1 U26959 ( .A1(n21170), .A2(n21169), .B1(n21606), .X(
        n21171) );
  sky130_fd_sc_hd__nand4_1 U26960 ( .A(n21172), .B(n21645), .C(n21171), .D(
        n21649), .Y(n21175) );
  sky130_fd_sc_hd__nand3b_1 U26961 ( .A_N(n21247), .B(n21174), .C(n21173), .Y(
        n21283) );
  sky130_fd_sc_hd__o21a_1 U26962 ( .A1(n21175), .A2(n21283), .B1(n20908), .X(
        n21183) );
  sky130_fd_sc_hd__nor4_1 U26963 ( .A(n21178), .B(n21177), .C(n21201), .D(
        n21176), .Y(n21180) );
  sky130_fd_sc_hd__a21oi_1 U26964 ( .A1(n21181), .A2(n21180), .B1(n21179), .Y(
        n21182) );
  sky130_fd_sc_hd__o21a_1 U26965 ( .A1(n21183), .A2(n21182), .B1(n21636), .X(
        n21310) );
  sky130_fd_sc_hd__nor2_1 U26966 ( .A(n21184), .B(n21719), .Y(n21278) );
  sky130_fd_sc_hd__nand4_1 U26967 ( .A(n21187), .B(n21278), .C(n21186), .D(
        n21185), .Y(n21189) );
  sky130_fd_sc_hd__nand4_1 U26969 ( .A(n21223), .B(n21191), .C(n21681), .D(
        n21190), .Y(n21192) );
  sky130_fd_sc_hd__o21ai_0 U26970 ( .A1(n21193), .A2(n21192), .B1(n21288), .Y(
        n21194) );
  sky130_fd_sc_hd__nand2_1 U26971 ( .A(n21195), .B(n21194), .Y(n21196) );
  sky130_fd_sc_hd__nand2_1 U26972 ( .A(n21196), .B(n20908), .Y(n21307) );
  sky130_fd_sc_hd__a22oi_1 U26973 ( .A1(n21699), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[45]), .B1(n21666), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[77]), .Y(n21301) );
  sky130_fd_sc_hd__nand2_1 U26974 ( .A(n21698), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[109]), .Y(n21300) );
  sky130_fd_sc_hd__nand2_1 U26975 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[13]), .Y(n21299) );
  sky130_fd_sc_hd__nand4_1 U26976 ( .A(n21301), .B(n21677), .C(n21300), .D(
        n21299), .Y(n21202) );
  sky130_fd_sc_hd__nand2b_1 U26977 ( .A_N(n21197), .B(n21685), .Y(n21199) );
  sky130_fd_sc_hd__o31a_1 U26978 ( .A1(n21201), .A2(n21200), .A3(n21199), .B1(
        n21198), .X(n21302) );
  sky130_fd_sc_hd__nor2_1 U26979 ( .A(n21202), .B(n21302), .Y(n21242) );
  sky130_fd_sc_hd__nand2_1 U26980 ( .A(n21233), .B(n21223), .Y(n21204) );
  sky130_fd_sc_hd__nor3_1 U26981 ( .A(n21205), .B(n21204), .C(n21203), .Y(
        n21210) );
  sky130_fd_sc_hd__nor2_1 U26982 ( .A(n21208), .B(n21207), .Y(n21209) );
  sky130_fd_sc_hd__nand4_1 U26983 ( .A(n21211), .B(n21210), .C(n21209), .D(
        n21688), .Y(n21212) );
  sky130_fd_sc_hd__nand2_1 U26984 ( .A(n21212), .B(n21251), .Y(n21240) );
  sky130_fd_sc_hd__nor3_1 U26985 ( .A(n21215), .B(n21214), .C(n21213), .Y(
        n21216) );
  sky130_fd_sc_hd__nand2_1 U26986 ( .A(n21217), .B(n21216), .Y(n21218) );
  sky130_fd_sc_hd__nand2_1 U26987 ( .A(n21218), .B(n21288), .Y(n21239) );
  sky130_fd_sc_hd__and4_1 U26988 ( .A(n21245), .B(n21631), .C(n21220), .D(
        n21219), .X(n21222) );
  sky130_fd_sc_hd__nand3_1 U26989 ( .A(n21223), .B(n21222), .C(n21221), .Y(
        n21225) );
  sky130_fd_sc_hd__o21ai_0 U26990 ( .A1(n21225), .A2(n21224), .B1(n21636), .Y(
        n21238) );
  sky130_fd_sc_hd__nor2_1 U26991 ( .A(n21227), .B(n21226), .Y(n21232) );
  sky130_fd_sc_hd__and4_1 U26992 ( .A(n21230), .B(n21229), .C(n21287), .D(
        n21228), .X(n21231) );
  sky130_fd_sc_hd__nand4_1 U26993 ( .A(n21234), .B(n21233), .C(n21232), .D(
        n21231), .Y(n21236) );
  sky130_fd_sc_hd__nand2_1 U26994 ( .A(n21236), .B(n21235), .Y(n21237) );
  sky130_fd_sc_hd__nand4_1 U26995 ( .A(n21240), .B(n21239), .C(n21238), .D(
        n21237), .Y(n21241) );
  sky130_fd_sc_hd__nand2_1 U26996 ( .A(n21241), .B(n21727), .Y(n21305) );
  sky130_fd_sc_hd__nand2_1 U26997 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_duty[1]), .Y(n21304) );
  sky130_fd_sc_hd__nand4_1 U26998 ( .A(n21307), .B(n21242), .C(n21305), .D(
        n21304), .Y(n21277) );
  sky130_fd_sc_hd__nand4_1 U26999 ( .A(n21246), .B(n21269), .C(n21245), .D(
        n21244), .Y(n21248) );
  sky130_fd_sc_hd__nor3_1 U27000 ( .A(n21249), .B(n21248), .C(n21247), .Y(
        n21250) );
  sky130_fd_sc_hd__nand2_1 U27001 ( .A(n21274), .B(n21250), .Y(n21252) );
  sky130_fd_sc_hd__nand2_1 U27002 ( .A(n21252), .B(n21251), .Y(n21263) );
  sky130_fd_sc_hd__nand3_1 U27003 ( .A(n21258), .B(n21253), .C(n21287), .Y(
        n21254) );
  sky130_fd_sc_hd__o21ai_1 U27004 ( .A1(n21255), .A2(n21254), .B1(n21636), .Y(
        n21262) );
  sky130_fd_sc_hd__nand4_1 U27005 ( .A(n21258), .B(n21608), .C(n21257), .D(
        n21256), .Y(n21260) );
  sky130_fd_sc_hd__o21ai_1 U27006 ( .A1(n21260), .A2(n21259), .B1(n21288), .Y(
        n21261) );
  sky130_fd_sc_hd__nand3_1 U27007 ( .A(n21263), .B(n21262), .C(n21261), .Y(
        n21276) );
  sky130_fd_sc_hd__nor2_1 U27008 ( .A(n21641), .B(n21264), .Y(n21678) );
  sky130_fd_sc_hd__nand4_1 U27009 ( .A(n21269), .B(n21268), .C(n21267), .D(
        n21266), .Y(n21272) );
  sky130_fd_sc_hd__nand2_1 U27010 ( .A(n21614), .B(n21270), .Y(n21271) );
  sky130_fd_sc_hd__nor2_1 U27011 ( .A(n21272), .B(n21271), .Y(n21273) );
  sky130_fd_sc_hd__a31oi_1 U27012 ( .A1(n21678), .A2(n21274), .A3(n21273), 
        .B1(n21705), .Y(n21275) );
  sky130_fd_sc_hd__o21a_1 U27013 ( .A1(n21276), .A2(n21275), .B1(n21697), .X(
        n21308) );
  sky130_fd_sc_hd__nor3_1 U27014 ( .A(n21310), .B(n21277), .C(n21308), .Y(
        n21294) );
  sky130_fd_sc_hd__nor2_1 U27015 ( .A(n21619), .B(n21279), .Y(n21280) );
  sky130_fd_sc_hd__nand2_1 U27016 ( .A(n21281), .B(n21280), .Y(n21282) );
  sky130_fd_sc_hd__nand2_1 U27017 ( .A(n21282), .B(n13275), .Y(n21313) );
  sky130_fd_sc_hd__nor4b_1 U27018 ( .D_N(n12180), .A(n21285), .B(n21284), .C(
        n21283), .Y(n21292) );
  sky130_fd_sc_hd__nand3_1 U27019 ( .A(n21628), .B(n21287), .C(n21286), .Y(
        n21290) );
  sky130_fd_sc_hd__nand2_1 U27022 ( .A(n21293), .B(n13481), .Y(n21312) );
  sky130_fd_sc_hd__nand2_1 U27023 ( .A(j202_soc_core_memory0_ram_dout0[461]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n21298) );
  sky130_fd_sc_hd__nand2_1 U27024 ( .A(j202_soc_core_memory0_ram_dout0[429]), 
        .B(n21598), .Y(n21297) );
  sky130_fd_sc_hd__nand2_1 U27025 ( .A(j202_soc_core_memory0_ram_dout0[45]), 
        .B(n21604), .Y(n21296) );
  sky130_fd_sc_hd__nand2_1 U27026 ( .A(j202_soc_core_memory0_ram_dout0[493]), 
        .B(n21771), .Y(n21315) );
  sky130_fd_sc_hd__nand4_1 U27027 ( .A(n21301), .B(n21738), .C(n21300), .D(
        n21299), .Y(n21303) );
  sky130_fd_sc_hd__nor2_1 U27028 ( .A(n21303), .B(n21302), .Y(n21306) );
  sky130_fd_sc_hd__nand4_1 U27029 ( .A(n21307), .B(n21306), .C(n21305), .D(
        n21304), .Y(n21309) );
  sky130_fd_sc_hd__nor3_1 U27030 ( .A(n21310), .B(n21309), .C(n21308), .Y(
        n21311) );
  sky130_fd_sc_hd__nand3_1 U27031 ( .A(n21315), .B(n21314), .C(n21313), .Y(
        n21339) );
  sky130_fd_sc_hd__nor2_1 U27032 ( .A(n21342), .B(n21319), .Y(n21320) );
  sky130_fd_sc_hd__xnor2_1 U27033 ( .A(n21321), .B(n21320), .Y(n25329) );
  sky130_fd_sc_hd__nand2_1 U27034 ( .A(n22596), .B(n25329), .Y(n21323) );
  sky130_fd_sc_hd__nand2_1 U27035 ( .A(n22515), .B(n27361), .Y(n21322) );
  sky130_fd_sc_hd__nand2_1 U27036 ( .A(n21334), .B(n21333), .Y(n21335) );
  sky130_fd_sc_hd__xor2_1 U27037 ( .A(n21336), .B(n21335), .X(n25316) );
  sky130_fd_sc_hd__nand2_1 U27038 ( .A(n25316), .B(n12158), .Y(n21337) );
  sky130_fd_sc_hd__nand2_1 U27039 ( .A(n21340), .B(n21339), .Y(n23694) );
  sky130_fd_sc_hd__nand2b_1 U27040 ( .A_N(n23694), .B(n22581), .Y(n21351) );
  sky130_fd_sc_hd__xnor2_1 U27041 ( .A(n21342), .B(n21341), .Y(n25291) );
  sky130_fd_sc_hd__nand2_1 U27042 ( .A(n22596), .B(n25291), .Y(n21344) );
  sky130_fd_sc_hd__nand2_1 U27043 ( .A(n22515), .B(n27365), .Y(n21343) );
  sky130_fd_sc_hd__o211a_2 U27044 ( .A1(n26708), .A2(n11143), .B1(n21344), 
        .C1(n21343), .X(n21350) );
  sky130_fd_sc_hd__nand2_1 U27045 ( .A(n21346), .B(n21345), .Y(n21348) );
  sky130_fd_sc_hd__xnor2_1 U27046 ( .A(n21348), .B(n21347), .Y(n23710) );
  sky130_fd_sc_hd__nand2_1 U27047 ( .A(n23710), .B(n12158), .Y(n21349) );
  sky130_fd_sc_hd__nand2_1 U27048 ( .A(n22321), .B(n21353), .Y(n21367) );
  sky130_fd_sc_hd__nor2_1 U27049 ( .A(n21469), .B(n21367), .Y(n21354) );
  sky130_fd_sc_hd__xnor2_1 U27050 ( .A(n19496), .B(n21354), .Y(n26390) );
  sky130_fd_sc_hd__o22a_1 U27051 ( .A1(n26426), .A2(n11143), .B1(n26413), .B2(
        n22590), .X(n21355) );
  sky130_fd_sc_hd__o21ai_1 U27052 ( .A1(n26413), .A2(n22592), .B1(n21355), .Y(
        n21356) );
  sky130_fd_sc_hd__a21oi_1 U27053 ( .A1(n26390), .A2(n22596), .B1(n21356), .Y(
        n21365) );
  sky130_fd_sc_hd__nand2_1 U27054 ( .A(n21361), .B(n21360), .Y(n21362) );
  sky130_fd_sc_hd__xor2_1 U27055 ( .A(n21363), .B(n21362), .X(n26387) );
  sky130_fd_sc_hd__nand2_1 U27056 ( .A(n26387), .B(n12158), .Y(n21364) );
  sky130_fd_sc_hd__nand2_1 U27057 ( .A(n12175), .B(n22581), .Y(n21376) );
  sky130_fd_sc_hd__xor2_1 U27058 ( .A(n21367), .B(n21469), .X(n24687) );
  sky130_fd_sc_hd__o22a_1 U27059 ( .A1(n23780), .A2(n13603), .B1(n26336), .B2(
        n11143), .X(n21368) );
  sky130_fd_sc_hd__a21oi_1 U27061 ( .A1(n27377), .A2(n22515), .B1(n21369), .Y(
        n21375) );
  sky130_fd_sc_hd__nand2_1 U27062 ( .A(n21371), .B(n21370), .Y(n21372) );
  sky130_fd_sc_hd__xor2_1 U27063 ( .A(n21373), .B(n21372), .X(n24676) );
  sky130_fd_sc_hd__nand2_1 U27064 ( .A(n24676), .B(n12158), .Y(n21374) );
  sky130_fd_sc_hd__nor2_1 U27065 ( .A(n29062), .B(n23305), .Y(n22709) );
  sky130_fd_sc_hd__nand2_1 U27066 ( .A(n22709), .B(n22668), .Y(n22677) );
  sky130_fd_sc_hd__nor2_1 U27067 ( .A(n22711), .B(n22677), .Y(n29027) );
  sky130_fd_sc_hd__nand2_1 U27068 ( .A(n11941), .B(n21813), .Y(n21377) );
  sky130_fd_sc_hd__nand3_1 U27069 ( .A(n28921), .B(n22712), .C(n22723), .Y(
        n21383) );
  sky130_fd_sc_hd__nand3_1 U27070 ( .A(n12616), .B(n21813), .C(n22723), .Y(
        n21382) );
  sky130_fd_sc_hd__nand3_1 U27071 ( .A(n12175), .B(n22715), .C(n22723), .Y(
        n21381) );
  sky130_fd_sc_hd__nand3b_1 U27072 ( .A_N(n29513), .B(n22714), .C(n22723), .Y(
        n21380) );
  sky130_fd_sc_hd__nand4_1 U27073 ( .A(n21383), .B(n21382), .C(n21381), .D(
        n21380), .Y(n26604) );
  sky130_fd_sc_hd__nand2_1 U27075 ( .A(n21387), .B(n21386), .Y(n21389) );
  sky130_fd_sc_hd__xor2_1 U27076 ( .A(n21389), .B(n21388), .X(n24128) );
  sky130_fd_sc_hd__nand2_1 U27077 ( .A(n24128), .B(n22927), .Y(n22011) );
  sky130_fd_sc_hd__mux2i_1 U27078 ( .A0(n22722), .A1(n26423), .S(n26792), .Y(
        n21403) );
  sky130_fd_sc_hd__nand2_1 U27079 ( .A(n26341), .B(n26719), .Y(n21391) );
  sky130_fd_sc_hd__nand2_1 U27080 ( .A(n26342), .B(n27425), .Y(n21390) );
  sky130_fd_sc_hd__o211ai_1 U27081 ( .A1(n26577), .A2(n26418), .B1(n21391), 
        .C1(n21390), .Y(n21402) );
  sky130_fd_sc_hd__nand2_1 U27082 ( .A(n27429), .B(n22723), .Y(n26627) );
  sky130_fd_sc_hd__nand2b_1 U27083 ( .A_N(n21972), .B(n24132), .Y(n22007) );
  sky130_fd_sc_hd__a22oi_1 U27084 ( .A1(n26329), .A2(n22009), .B1(n22723), 
        .B2(n23940), .Y(n21393) );
  sky130_fd_sc_hd__nand2_1 U27085 ( .A(n26792), .B(n26713), .Y(n26628) );
  sky130_fd_sc_hd__nand3_1 U27086 ( .A(n26628), .B(n26326), .C(n26627), .Y(
        n21392) );
  sky130_fd_sc_hd__o211ai_1 U27087 ( .A1(n26432), .A2(n26627), .B1(n21393), 
        .C1(n21392), .Y(n21395) );
  sky130_fd_sc_hd__o22ai_1 U27088 ( .A1(n25229), .A2(n26427), .B1(n27007), 
        .B2(n26424), .Y(n21394) );
  sky130_fd_sc_hd__nor2_1 U27089 ( .A(n21395), .B(n21394), .Y(n21400) );
  sky130_fd_sc_hd__nand2b_1 U27090 ( .A_N(n22925), .B(
        j202_soc_core_j22_cpu_ml_macl[3]), .Y(n22010) );
  sky130_fd_sc_hd__a22oi_1 U27091 ( .A1(n26077), .A2(n26720), .B1(n21396), 
        .B2(n26329), .Y(n21399) );
  sky130_fd_sc_hd__nand2_1 U27092 ( .A(n24483), .B(n26603), .Y(n21398) );
  sky130_fd_sc_hd__nand2_1 U27093 ( .A(n26338), .B(n27377), .Y(n21397) );
  sky130_fd_sc_hd__nand4_1 U27094 ( .A(n21400), .B(n21399), .C(n21398), .D(
        n21397), .Y(n21401) );
  sky130_fd_sc_hd__nor3_1 U27095 ( .A(n21403), .B(n21402), .C(n21401), .Y(
        n21404) );
  sky130_fd_sc_hd__o21ai_1 U27096 ( .A1(n18916), .A2(n22011), .B1(n21404), .Y(
        n21405) );
  sky130_fd_sc_hd__a21oi_1 U27097 ( .A1(n24645), .A2(n26409), .B1(n21405), .Y(
        n21409) );
  sky130_fd_sc_hd__nand2_1 U27098 ( .A(n22723), .B(n26323), .Y(n21406) );
  sky130_fd_sc_hd__nand2_1 U27099 ( .A(n21406), .B(n25159), .Y(n21407) );
  sky130_fd_sc_hd__nand2_1 U27100 ( .A(n27428), .B(n21407), .Y(n21408) );
  sky130_fd_sc_hd__nand2_1 U27101 ( .A(n21410), .B(n22873), .Y(n21417) );
  sky130_fd_sc_hd__o22ai_1 U27102 ( .A1(n21411), .A2(n22854), .B1(n20285), 
        .B2(n22860), .Y(n21412) );
  sky130_fd_sc_hd__a21oi_1 U27103 ( .A1(j202_soc_core_j22_cpu_rf_gpr[3]), .A2(
        n22866), .B1(n21412), .Y(n21416) );
  sky130_fd_sc_hd__a22oi_1 U27104 ( .A1(n21847), .A2(
        j202_soc_core_j22_cpu_rf_gbr[3]), .B1(n22864), .B2(
        j202_soc_core_j22_cpu_rf_vbr[3]), .Y(n21415) );
  sky130_fd_sc_hd__a2bb2oi_1 U27105 ( .B1(j202_soc_core_j22_cpu_rf_gpr[483]), 
        .B2(n22865), .A1_N(n21413), .A2_N(n22033), .Y(n21414) );
  sky130_fd_sc_hd__nand4_1 U27106 ( .A(n21417), .B(n21416), .C(n21415), .D(
        n21414), .Y(n22976) );
  sky130_fd_sc_hd__nand2_1 U27107 ( .A(n22976), .B(n22824), .Y(n21434) );
  sky130_fd_sc_hd__nand2_1 U27108 ( .A(n22014), .B(n21434), .Y(n21436) );
  sky130_fd_sc_hd__nand2_1 U27109 ( .A(n11139), .B(n21419), .Y(n21426) );
  sky130_fd_sc_hd__nand2_1 U27110 ( .A(n21790), .B(n21422), .Y(n21424) );
  sky130_fd_sc_hd__a21oi_1 U27111 ( .A1(n21797), .A2(n21422), .B1(n21421), .Y(
        n21423) );
  sky130_fd_sc_hd__o21ai_2 U27112 ( .A1(n21424), .A2(n22912), .B1(n21423), .Y(
        n21425) );
  sky130_fd_sc_hd__xnor2_2 U27113 ( .A(n21426), .B(n21425), .Y(n23233) );
  sky130_fd_sc_hd__nand2_1 U27114 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[3]), .Y(n24133) );
  sky130_fd_sc_hd__a21oi_1 U27115 ( .A1(n19200), .A2(n21429), .B1(n11142), .Y(
        n21433) );
  sky130_fd_sc_hd__nand2_1 U27116 ( .A(n21431), .B(n21430), .Y(n21432) );
  sky130_fd_sc_hd__xor2_1 U27117 ( .A(n21433), .B(n21432), .X(n22955) );
  sky130_fd_sc_hd__nand2_1 U27118 ( .A(n22955), .B(n24499), .Y(n24134) );
  sky130_fd_sc_hd__nand2_1 U27119 ( .A(n21439), .B(n21438), .Y(n21445) );
  sky130_fd_sc_hd__nand2_1 U27120 ( .A(n21874), .B(n21441), .Y(n21443) );
  sky130_fd_sc_hd__a21oi_1 U27121 ( .A1(n21881), .A2(n21441), .B1(n21440), .Y(
        n21442) );
  sky130_fd_sc_hd__o21ai_1 U27122 ( .A1(n21443), .A2(n22837), .B1(n21442), .Y(
        n21444) );
  sky130_fd_sc_hd__xnor2_1 U27123 ( .A(n21445), .B(n21444), .Y(n22688) );
  sky130_fd_sc_hd__nand2_1 U27124 ( .A(n22688), .B(n24499), .Y(n21457) );
  sky130_fd_sc_hd__nand2_1 U27125 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[11]), .Y(n21456) );
  sky130_fd_sc_hd__nand2_1 U27126 ( .A(n21457), .B(n21456), .Y(n24654) );
  sky130_fd_sc_hd__nand2_1 U27127 ( .A(n21447), .B(n21446), .Y(n21455) );
  sky130_fd_sc_hd__nand2_1 U27128 ( .A(n22521), .B(n21451), .Y(n21453) );
  sky130_fd_sc_hd__a21oi_1 U27129 ( .A1(n22661), .A2(n21451), .B1(n21450), .Y(
        n21452) );
  sky130_fd_sc_hd__a31oi_1 U27130 ( .A1(n21457), .A2(n26318), .A3(n21456), 
        .B1(n11713), .Y(n21458) );
  sky130_fd_sc_hd__o22a_1 U27132 ( .A1(n21972), .A2(n21459), .B1(n23972), .B2(
        n22925), .X(n24662) );
  sky130_fd_sc_hd__a21oi_1 U27133 ( .A1(n21461), .A2(n12208), .B1(n21460), .Y(
        n21464) );
  sky130_fd_sc_hd__nand2_1 U27134 ( .A(n13280), .B(n21462), .Y(n21463) );
  sky130_fd_sc_hd__xor2_1 U27135 ( .A(n21464), .B(n21463), .X(n25147) );
  sky130_fd_sc_hd__nand2_1 U27136 ( .A(n25147), .B(n22927), .Y(n24680) );
  sky130_fd_sc_hd__nand3_1 U27137 ( .A(n21465), .B(n24662), .C(n24680), .Y(
        n21466) );
  sky130_fd_sc_hd__nand2_1 U27138 ( .A(n21466), .B(n22929), .Y(n21477) );
  sky130_fd_sc_hd__nand2_1 U27139 ( .A(n21467), .B(n22873), .Y(n21475) );
  sky130_fd_sc_hd__o22ai_1 U27140 ( .A1(n21469), .A2(n22860), .B1(n22854), 
        .B2(n21468), .Y(n21470) );
  sky130_fd_sc_hd__a21oi_1 U27141 ( .A1(n22866), .A2(
        j202_soc_core_j22_cpu_rf_gpr[11]), .B1(n21470), .Y(n21474) );
  sky130_fd_sc_hd__a22oi_1 U27142 ( .A1(n21847), .A2(
        j202_soc_core_j22_cpu_rf_gbr[11]), .B1(n22864), .B2(
        j202_soc_core_j22_cpu_rf_vbr[11]), .Y(n21473) );
  sky130_fd_sc_hd__a2bb2oi_1 U27143 ( .B1(j202_soc_core_j22_cpu_rf_gpr[491]), 
        .B2(n22865), .A1_N(n21471), .A2_N(n22033), .Y(n21472) );
  sky130_fd_sc_hd__nand4_1 U27144 ( .A(n21475), .B(n21474), .C(n21473), .D(
        n21472), .Y(n22703) );
  sky130_fd_sc_hd__nand2_1 U27145 ( .A(n22703), .B(n22004), .Y(n21476) );
  sky130_fd_sc_hd__nand3_1 U27146 ( .A(n22704), .B(n21477), .C(n21476), .Y(
        n28979) );
  sky130_fd_sc_hd__nand2_1 U27147 ( .A(n12771), .B(n22581), .Y(n21488) );
  sky130_fd_sc_hd__nand2_1 U27148 ( .A(n22327), .B(n22325), .Y(n21483) );
  sky130_fd_sc_hd__xnor2_1 U27150 ( .A(n21483), .B(n22328), .Y(n24729) );
  sky130_fd_sc_hd__o22a_1 U27151 ( .A1(n25121), .A2(n22590), .B1(n25788), .B2(
        n11143), .X(n21484) );
  sky130_fd_sc_hd__o21ai_1 U27152 ( .A1(n25121), .A2(n22592), .B1(n21484), .Y(
        n21485) );
  sky130_fd_sc_hd__a21oi_1 U27153 ( .A1(n24729), .A2(n12158), .B1(n21485), .Y(
        n21487) );
  sky130_fd_sc_hd__xnor2_1 U27154 ( .A(n22861), .B(n22321), .Y(n25555) );
  sky130_fd_sc_hd__nand2_1 U27155 ( .A(n22596), .B(n25555), .Y(n21486) );
  sky130_fd_sc_hd__nand3_1 U27156 ( .A(n21488), .B(n21487), .C(n21486), .Y(
        n29032) );
  sky130_fd_sc_hd__nand2_1 U27157 ( .A(n21490), .B(n21489), .Y(n21497) );
  sky130_fd_sc_hd__nor2_1 U27158 ( .A(n21491), .B(n22617), .Y(n21493) );
  sky130_fd_sc_hd__o21ai_1 U27159 ( .A1(n21491), .A2(n22619), .B1(n21867), .Y(
        n21492) );
  sky130_fd_sc_hd__xnor2_2 U27160 ( .A(n21497), .B(n21496), .Y(n23244) );
  sky130_fd_sc_hd__nand2_1 U27161 ( .A(n23244), .B(n26863), .Y(n25325) );
  sky130_fd_sc_hd__nand2_1 U27162 ( .A(n21500), .B(n21499), .Y(n21501) );
  sky130_fd_sc_hd__xor2_1 U27163 ( .A(n22897), .B(n21501), .X(n24510) );
  sky130_fd_sc_hd__nand2_1 U27164 ( .A(n24510), .B(n24499), .Y(n25323) );
  sky130_fd_sc_hd__nand2_1 U27165 ( .A(n21502), .B(n26398), .Y(n21508) );
  sky130_fd_sc_hd__nand2_1 U27166 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[14]), .Y(n25324) );
  sky130_fd_sc_hd__nand2b_1 U27167 ( .A_N(n21972), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .Y(n25300) );
  sky130_fd_sc_hd__o21ai_1 U27168 ( .A1(n11713), .A2(n25324), .B1(n25300), .Y(
        n21503) );
  sky130_fd_sc_hd__nor2_1 U27169 ( .A(n23949), .B(n22925), .Y(n25301) );
  sky130_fd_sc_hd__nor2_1 U27170 ( .A(n21503), .B(n25301), .Y(n21507) );
  sky130_fd_sc_hd__nand2_1 U27171 ( .A(n21505), .B(n21504), .Y(n21506) );
  sky130_fd_sc_hd__xnor2_1 U27172 ( .A(n21506), .B(n18886), .Y(n24511) );
  sky130_fd_sc_hd__nand2_1 U27173 ( .A(n24511), .B(n22927), .Y(n25318) );
  sky130_fd_sc_hd__nand3_1 U27174 ( .A(n21508), .B(n21507), .C(n25318), .Y(
        n21509) );
  sky130_fd_sc_hd__nand2_1 U27175 ( .A(n21509), .B(n22929), .Y(n21581) );
  sky130_fd_sc_hd__nand2_1 U27176 ( .A(n12178), .B(n21510), .Y(n21514) );
  sky130_fd_sc_hd__o21ai_2 U27177 ( .A1(n21512), .A2(n11439), .B1(n21511), .Y(
        n21513) );
  sky130_fd_sc_hd__xnor2_2 U27178 ( .A(n21514), .B(n21513), .Y(n23234) );
  sky130_fd_sc_hd__nand2_1 U27179 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[6]), .Y(n25336) );
  sky130_fd_sc_hd__nand2_1 U27180 ( .A(n12173), .B(n21515), .Y(n21517) );
  sky130_fd_sc_hd__xnor2_1 U27181 ( .A(n21517), .B(n12599), .Y(n25345) );
  sky130_fd_sc_hd__nand2_1 U27182 ( .A(n25345), .B(n22927), .Y(n22240) );
  sky130_fd_sc_hd__nor2_1 U27183 ( .A(n18916), .B(n22240), .Y(n22243) );
  sky130_fd_sc_hd__o21a_1 U27184 ( .A1(n26802), .A2(n22243), .B1(n22768), .X(
        n22612) );
  sky130_fd_sc_hd__nand2_1 U27185 ( .A(n22613), .B(n22612), .Y(n21580) );
  sky130_fd_sc_hd__nand2_1 U27186 ( .A(n21519), .B(n21520), .Y(n23693) );
  sky130_fd_sc_hd__a21oi_1 U27187 ( .A1(n27409), .A2(n25415), .B1(n26085), .Y(
        n21525) );
  sky130_fd_sc_hd__nand2_1 U27188 ( .A(n27408), .B(n26323), .Y(n21524) );
  sky130_fd_sc_hd__nand2_1 U27189 ( .A(n21528), .B(n21527), .Y(n21533) );
  sky130_fd_sc_hd__a21oi_1 U27190 ( .A1(n21531), .A2(n21530), .B1(n21529), .Y(
        n21760) );
  sky130_fd_sc_hd__o21ai_0 U27191 ( .A1(n21756), .A2(n21760), .B1(n21757), .Y(
        n21532) );
  sky130_fd_sc_hd__xnor2_1 U27192 ( .A(n21533), .B(n21532), .Y(n25526) );
  sky130_fd_sc_hd__o22ai_1 U27193 ( .A1(n27007), .A2(n26419), .B1(n25821), 
        .B2(n26418), .Y(n21534) );
  sky130_fd_sc_hd__a21oi_1 U27194 ( .A1(n26342), .A2(n27405), .B1(n21534), .Y(
        n21546) );
  sky130_fd_sc_hd__xnor2_1 U27195 ( .A(n26600), .B(n27409), .Y(n26640) );
  sky130_fd_sc_hd__nor2_1 U27196 ( .A(n26415), .B(n26640), .Y(n21544) );
  sky130_fd_sc_hd__o22ai_1 U27197 ( .A1(n26577), .A2(n26427), .B1(n25798), 
        .B2(n26424), .Y(n21543) );
  sky130_fd_sc_hd__nand2_1 U27198 ( .A(n26338), .B(n27361), .Y(n21541) );
  sky130_fd_sc_hd__nand2b_1 U27199 ( .A_N(n21972), .B(
        j202_soc_core_j22_cpu_ml_bufa[6]), .Y(n22235) );
  sky130_fd_sc_hd__o22ai_1 U27200 ( .A1(n18916), .A2(n22235), .B1(n26423), 
        .B2(n27409), .Y(n21535) );
  sky130_fd_sc_hd__a21oi_1 U27201 ( .A1(n22731), .A2(n26508), .B1(n21535), .Y(
        n21536) );
  sky130_fd_sc_hd__o21a_1 U27202 ( .A1(n26703), .A2(n22729), .B1(n21536), .X(
        n21540) );
  sky130_fd_sc_hd__nand2_1 U27203 ( .A(n26077), .B(n26725), .Y(n21539) );
  sky130_fd_sc_hd__nor2_1 U27204 ( .A(n21537), .B(n22925), .Y(n22238) );
  sky130_fd_sc_hd__nand2_1 U27205 ( .A(n22238), .B(n26329), .Y(n21538) );
  sky130_fd_sc_hd__nand4_1 U27206 ( .A(n21541), .B(n21540), .C(n21539), .D(
        n21538), .Y(n21542) );
  sky130_fd_sc_hd__nor3_1 U27207 ( .A(n21544), .B(n21543), .C(n21542), .Y(
        n21545) );
  sky130_fd_sc_hd__o211ai_1 U27208 ( .A1(n11977), .A2(n22722), .B1(n21546), 
        .C1(n21545), .Y(n21547) );
  sky130_fd_sc_hd__a21oi_1 U27209 ( .A1(n25526), .A2(n26409), .B1(n21547), .Y(
        n21551) );
  sky130_fd_sc_hd__nand2b_1 U27210 ( .A_N(n21548), .B(n23011), .Y(n21549) );
  sky130_fd_sc_hd__nand2_1 U27211 ( .A(n24785), .B(n21549), .Y(n26351) );
  sky130_fd_sc_hd__o22ai_1 U27213 ( .A1(n21553), .A2(n22856), .B1(n21552), 
        .B2(n22854), .Y(n21557) );
  sky130_fd_sc_hd__o22ai_1 U27214 ( .A1(n21555), .A2(n22860), .B1(n21554), 
        .B2(n22858), .Y(n21556) );
  sky130_fd_sc_hd__nor2_1 U27215 ( .A(n21557), .B(n21556), .Y(n21561) );
  sky130_fd_sc_hd__a22oi_1 U27216 ( .A1(n22865), .A2(
        j202_soc_core_j22_cpu_rf_gpr[486]), .B1(n22864), .B2(
        j202_soc_core_j22_cpu_rf_vbr[6]), .Y(n21560) );
  sky130_fd_sc_hd__nand2_1 U27217 ( .A(n22866), .B(
        j202_soc_core_j22_cpu_rf_gpr[6]), .Y(n21559) );
  sky130_fd_sc_hd__nand2_1 U27218 ( .A(n22867), .B(
        j202_soc_core_j22_cpu_rf_tmp[6]), .Y(n21558) );
  sky130_fd_sc_hd__nand4_1 U27219 ( .A(n21561), .B(n21560), .C(n21559), .D(
        n21558), .Y(n21562) );
  sky130_fd_sc_hd__a21oi_1 U27220 ( .A1(n21563), .A2(n22873), .B1(n21562), .Y(
        n22352) );
  sky130_fd_sc_hd__or2_0 U27221 ( .A(n22352), .B(n23292), .X(n21564) );
  sky130_fd_sc_hd__nand2_1 U27222 ( .A(n21565), .B(n21564), .Y(n22610) );
  sky130_fd_sc_hd__o22ai_1 U27223 ( .A1(n21321), .A2(n22860), .B1(n22854), 
        .B2(n21566), .Y(n21567) );
  sky130_fd_sc_hd__a21oi_1 U27224 ( .A1(n22866), .A2(
        j202_soc_core_j22_cpu_rf_gpr[14]), .B1(n21567), .Y(n21571) );
  sky130_fd_sc_hd__a22oi_1 U27225 ( .A1(n21847), .A2(
        j202_soc_core_j22_cpu_rf_gbr[14]), .B1(n22864), .B2(
        j202_soc_core_j22_cpu_rf_vbr[14]), .Y(n21570) );
  sky130_fd_sc_hd__nand2_1 U27226 ( .A(n22865), .B(
        j202_soc_core_j22_cpu_rf_gpr[494]), .Y(n21569) );
  sky130_fd_sc_hd__nand2_1 U27227 ( .A(n22867), .B(
        j202_soc_core_j22_cpu_rf_tmp[14]), .Y(n21568) );
  sky130_fd_sc_hd__nand4_1 U27228 ( .A(n21571), .B(n21570), .C(n21569), .D(
        n21568), .Y(n21572) );
  sky130_fd_sc_hd__a21oi_1 U27229 ( .A1(n21573), .A2(n22873), .B1(n21572), .Y(
        n22611) );
  sky130_fd_sc_hd__nand2_1 U27230 ( .A(n21576), .B(n21575), .Y(n21577) );
  sky130_fd_sc_hd__xor2_1 U27231 ( .A(n22837), .B(n21577), .X(n22340) );
  sky130_fd_sc_hd__nand2_1 U27232 ( .A(n22340), .B(n24499), .Y(n23274) );
  sky130_fd_sc_hd__o22ai_1 U27233 ( .A1(n22932), .A2(n22611), .B1(n21578), 
        .B2(n23274), .Y(n21579) );
  sky130_fd_sc_hd__nand2b_1 U27234 ( .A_N(n23693), .B(n22581), .Y(n21589) );
  sky130_fd_sc_hd__nor2_1 U27235 ( .A(n21761), .B(n21762), .Y(n21582) );
  sky130_fd_sc_hd__xnor2_1 U27236 ( .A(n21555), .B(n21582), .Y(n25529) );
  sky130_fd_sc_hd__o22a_1 U27237 ( .A1(n21585), .A2(n13603), .B1(n11145), .B2(
        n11143), .X(n21583) );
  sky130_fd_sc_hd__o21ai_1 U27238 ( .A1(n21585), .A2(n21584), .B1(n21583), .Y(
        n21586) );
  sky130_fd_sc_hd__a21oi_1 U27239 ( .A1(n25526), .A2(n12158), .B1(n21586), .Y(
        n21588) );
  sky130_fd_sc_hd__nand2_1 U27240 ( .A(n22515), .B(n27409), .Y(n21587) );
  sky130_fd_sc_hd__nand3_1 U27241 ( .A(n21589), .B(n21588), .C(n21587), .Y(
        n29011) );
  sky130_fd_sc_hd__nand2_1 U27242 ( .A(j202_soc_core_memory0_ram_dout0[133]), 
        .B(n21592), .Y(n21595) );
  sky130_fd_sc_hd__nand2_1 U27243 ( .A(j202_soc_core_memory0_ram_dout0[325]), 
        .B(n21593), .Y(n21594) );
  sky130_fd_sc_hd__nand2_1 U27244 ( .A(j202_soc_core_memory0_ram_dout0[357]), 
        .B(n21596), .Y(n21602) );
  sky130_fd_sc_hd__nand2_1 U27245 ( .A(j202_soc_core_memory0_ram_dout0[389]), 
        .B(n21597), .Y(n21601) );
  sky130_fd_sc_hd__nand2_1 U27246 ( .A(j202_soc_core_memory0_ram_dout0[453]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[14]), .Y(n21600) );
  sky130_fd_sc_hd__nand2_1 U27247 ( .A(j202_soc_core_memory0_ram_dout0[421]), 
        .B(n21598), .Y(n21599) );
  sky130_fd_sc_hd__nand4_1 U27248 ( .A(n21609), .B(n21608), .C(n21607), .D(
        n21606), .Y(n21610) );
  sky130_fd_sc_hd__nor3_1 U27249 ( .A(n21612), .B(n21611), .C(n21610), .Y(
        n21623) );
  sky130_fd_sc_hd__nand2_1 U27250 ( .A(n21614), .B(n21613), .Y(n21616) );
  sky130_fd_sc_hd__nor2_1 U27251 ( .A(n21616), .B(n21615), .Y(n21712) );
  sky130_fd_sc_hd__nor3_1 U27252 ( .A(n21620), .B(n21619), .C(n21618), .Y(
        n21621) );
  sky130_fd_sc_hd__and3_1 U27253 ( .A(n21712), .B(n21683), .C(n21621), .X(
        n21622) );
  sky130_fd_sc_hd__o22ai_1 U27254 ( .A1(n21623), .A2(n21722), .B1(n21622), 
        .B2(n21705), .Y(n21640) );
  sky130_fd_sc_hd__nor4_1 U27255 ( .A(n21627), .B(n21626), .C(n21625), .D(
        n21624), .Y(n21629) );
  sky130_fd_sc_hd__a31oi_1 U27256 ( .A1(n21630), .A2(n21629), .A3(n21628), 
        .B1(n21720), .Y(n21638) );
  sky130_fd_sc_hd__nand4_1 U27257 ( .A(n21634), .B(n21633), .C(n21632), .D(
        n21631), .Y(n21635) );
  sky130_fd_sc_hd__nand2_1 U27258 ( .A(n21636), .B(n21635), .Y(n21637) );
  sky130_fd_sc_hd__nand2b_1 U27259 ( .A_N(n21638), .B(n21637), .Y(n21639) );
  sky130_fd_sc_hd__o21a_1 U27260 ( .A1(n21640), .A2(n21639), .B1(n20908), .X(
        n21747) );
  sky130_fd_sc_hd__nor3_1 U27261 ( .A(n21643), .B(n21642), .C(n21641), .Y(
        n21644) );
  sky130_fd_sc_hd__a31oi_1 U27262 ( .A1(n21683), .A2(n21645), .A3(n21644), 
        .B1(n21709), .Y(n21663) );
  sky130_fd_sc_hd__a31oi_1 U27263 ( .A1(n21710), .A2(n21647), .A3(n21646), 
        .B1(n21705), .Y(n21662) );
  sky130_fd_sc_hd__nand4_1 U27264 ( .A(n21651), .B(n21650), .C(n21649), .D(
        n21648), .Y(n21652) );
  sky130_fd_sc_hd__nor4_1 U27265 ( .A(n21654), .B(n21653), .C(n21656), .D(
        n21652), .Y(n21660) );
  sky130_fd_sc_hd__nor4_1 U27266 ( .A(n21658), .B(n21657), .C(n21656), .D(
        n21655), .Y(n21659) );
  sky130_fd_sc_hd__o22ai_1 U27267 ( .A1(n21660), .A2(n21722), .B1(n21659), 
        .B2(n21720), .Y(n21661) );
  sky130_fd_sc_hd__nor3_1 U27268 ( .A(n21663), .B(n21662), .C(n21661), .Y(
        n21665) );
  sky130_fd_sc_hd__nand2b_1 U27269 ( .A_N(n21665), .B(n13481), .Y(n21745) );
  sky130_fd_sc_hd__nand2_1 U27270 ( .A(n21666), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[69]), .Y(n21739) );
  sky130_fd_sc_hd__nand2_1 U27271 ( .A(n21667), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[13]), .Y(n21673) );
  sky130_fd_sc_hd__nand2_1 U27272 ( .A(n24376), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[21]), .Y(n21672) );
  sky130_fd_sc_hd__nand2_1 U27273 ( .A(n21668), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[5]), .Y(n21671) );
  sky130_fd_sc_hd__nand2_1 U27274 ( .A(n21669), .B(
        j202_soc_core_uart_TOP_rx_fifo_mem[29]), .Y(n21670) );
  sky130_fd_sc_hd__nand4_1 U27275 ( .A(n21673), .B(n21672), .C(n21671), .D(
        n21670), .Y(n21674) );
  sky130_fd_sc_hd__nand2_1 U27276 ( .A(n21675), .B(n21674), .Y(n21737) );
  sky130_fd_sc_hd__nand2_1 U27277 ( .A(n21676), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[5]), .Y(n21736) );
  sky130_fd_sc_hd__nand4_1 U27278 ( .A(n21739), .B(n21677), .C(n21737), .D(
        n21736), .Y(n21703) );
  sky130_fd_sc_hd__and4_1 U27279 ( .A(n21680), .B(n21679), .C(n21678), .D(
        n21681), .X(n21695) );
  sky130_fd_sc_hd__a31oi_1 U27280 ( .A1(n21683), .A2(n21682), .A3(n21681), 
        .B1(n21722), .Y(n21693) );
  sky130_fd_sc_hd__and3_1 U27281 ( .A(n21687), .B(n21686), .C(n21685), .X(
        n21691) );
  sky130_fd_sc_hd__and3_1 U27282 ( .A(n21712), .B(n21689), .C(n21688), .X(
        n21690) );
  sky130_fd_sc_hd__o22ai_1 U27283 ( .A1(n21691), .A2(n21720), .B1(n21690), 
        .B2(n21709), .Y(n21692) );
  sky130_fd_sc_hd__nor2_1 U27284 ( .A(n21693), .B(n21692), .Y(n21694) );
  sky130_fd_sc_hd__nand2_1 U27286 ( .A(n21697), .B(n21696), .Y(n21702) );
  sky130_fd_sc_hd__nand2_1 U27287 ( .A(n21698), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[101]), .Y(n21701) );
  sky130_fd_sc_hd__nand2_1 U27288 ( .A(n21699), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[37]), .Y(n21700) );
  sky130_fd_sc_hd__nand3_1 U27289 ( .A(n21702), .B(n21701), .C(n21700), .Y(
        n21740) );
  sky130_fd_sc_hd__nor2_1 U27290 ( .A(n21703), .B(n21740), .Y(n21729) );
  sky130_fd_sc_hd__a31oi_1 U27291 ( .A1(n21708), .A2(n21707), .A3(n21706), 
        .B1(n21705), .Y(n21726) );
  sky130_fd_sc_hd__a31oi_1 U27292 ( .A1(n21712), .A2(n21711), .A3(n21710), 
        .B1(n21709), .Y(n21725) );
  sky130_fd_sc_hd__nor4_1 U27293 ( .A(n21716), .B(n21715), .C(n21714), .D(
        n21713), .Y(n21723) );
  sky130_fd_sc_hd__nor3_1 U27294 ( .A(n21719), .B(n21718), .C(n21717), .Y(
        n21721) );
  sky130_fd_sc_hd__o22ai_1 U27295 ( .A1(n21723), .A2(n21722), .B1(n21721), 
        .B2(n21720), .Y(n21724) );
  sky130_fd_sc_hd__nor3_1 U27296 ( .A(n21726), .B(n21725), .C(n21724), .Y(
        n21728) );
  sky130_fd_sc_hd__nand2b_1 U27297 ( .A_N(n21728), .B(n21727), .Y(n21743) );
  sky130_fd_sc_hd__nand2_1 U27298 ( .A(n15249), .B(
        j202_soc_core_bldc_core_00_pwm_period[5]), .Y(n21742) );
  sky130_fd_sc_hd__nand4_1 U27299 ( .A(n21745), .B(n21729), .C(n21743), .D(
        n21742), .Y(n21730) );
  sky130_fd_sc_hd__nor2_1 U27300 ( .A(n21747), .B(n21730), .Y(n21731) );
  sky130_fd_sc_hd__nand2_1 U27301 ( .A(j202_soc_core_memory0_ram_dout0[485]), 
        .B(n21771), .Y(n21749) );
  sky130_fd_sc_hd__nand4_1 U27302 ( .A(n21739), .B(n21738), .C(n21737), .D(
        n21736), .Y(n21741) );
  sky130_fd_sc_hd__nor2_1 U27303 ( .A(n21741), .B(n21740), .Y(n21744) );
  sky130_fd_sc_hd__nand4_1 U27304 ( .A(n21745), .B(n21744), .C(n21743), .D(
        n21742), .Y(n21746) );
  sky130_fd_sc_hd__nor2_1 U27305 ( .A(n21747), .B(n21746), .Y(n21748) );
  sky130_fd_sc_hd__nand2_1 U27306 ( .A(n21749), .B(n21748), .Y(n21754) );
  sky130_fd_sc_hd__a22oi_1 U27307 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__5_), .B1(n21775), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__5_), .Y(n21753) );
  sky130_fd_sc_hd__nand2_1 U27308 ( .A(n21755), .B(n21754), .Y(n23695) );
  sky130_fd_sc_hd__nand2b_1 U27309 ( .A_N(n23695), .B(n22581), .Y(n21768) );
  sky130_fd_sc_hd__nand2_1 U27310 ( .A(n21758), .B(n21757), .Y(n21759) );
  sky130_fd_sc_hd__xor2_1 U27311 ( .A(n21760), .B(n21759), .X(n26889) );
  sky130_fd_sc_hd__nand2_1 U27312 ( .A(n26889), .B(n12158), .Y(n21765) );
  sky130_fd_sc_hd__xor2_1 U27313 ( .A(n21762), .B(n21761), .X(n26913) );
  sky130_fd_sc_hd__nand2_1 U27314 ( .A(n22596), .B(n26913), .Y(n21764) );
  sky130_fd_sc_hd__nand2_1 U27315 ( .A(n22510), .B(n26711), .Y(n21763) );
  sky130_fd_sc_hd__and3_1 U27316 ( .A(n21765), .B(n21764), .C(n21763), .X(
        n21767) );
  sky130_fd_sc_hd__nand2_1 U27317 ( .A(n22515), .B(n27415), .Y(n21766) );
  sky130_fd_sc_hd__nand3_1 U27318 ( .A(n21768), .B(n21767), .C(n21766), .Y(
        n29035) );
  sky130_fd_sc_hd__mux2i_1 U27319 ( .A0(n21769), .A1(n21770), .S(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n21772) );
  sky130_fd_sc_hd__nand2_1 U27320 ( .A(n21772), .B(n21771), .Y(n21774) );
  sky130_fd_sc_hd__nand2_1 U27321 ( .A(n21774), .B(n21773), .Y(n28923) );
  sky130_fd_sc_hd__nor2_1 U27322 ( .A(n21778), .B(n21777), .Y(n21779) );
  sky130_fd_sc_hd__nor2_1 U27323 ( .A(j202_soc_core_uart_BRG_sio_ce_x4_r), .B(
        n28035), .Y(n29081) );
  sky130_fd_sc_hd__nand2_1 U27324 ( .A(j202_soc_core_uart_TOP_dpll_state[0]), 
        .B(n21784), .Y(n28560) );
  sky130_fd_sc_hd__nand2_1 U27325 ( .A(n21787), .B(n21786), .Y(n21801) );
  sky130_fd_sc_hd__nor2_1 U27326 ( .A(n21794), .B(n21789), .Y(n21796) );
  sky130_fd_sc_hd__a21oi_1 U27328 ( .A1(n21797), .A2(n21796), .B1(n21795), .Y(
        n21798) );
  sky130_fd_sc_hd__xnor2_2 U27329 ( .A(n21801), .B(n21800), .Y(n23230) );
  sky130_fd_sc_hd__nor2_1 U27330 ( .A(n21805), .B(n12317), .Y(n21807) );
  sky130_fd_sc_hd__a21oi_1 U27332 ( .A1(n21807), .A2(n19200), .B1(n21806), .Y(
        n21812) );
  sky130_fd_sc_hd__nand2_1 U27333 ( .A(n21810), .B(n21809), .Y(n21811) );
  sky130_fd_sc_hd__xor2_1 U27334 ( .A(n21812), .B(n21811), .X(n22116) );
  sky130_fd_sc_hd__nand2_1 U27335 ( .A(n22116), .B(n24499), .Y(n24380) );
  sky130_fd_sc_hd__nand2_1 U27336 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[5]), .Y(n22450) );
  sky130_fd_sc_hd__nand2b_1 U27337 ( .A_N(n23694), .B(n22715), .Y(n21815) );
  sky130_fd_sc_hd__a21oi_1 U27338 ( .A1(n27415), .A2(n25415), .B1(n26085), .Y(
        n21819) );
  sky130_fd_sc_hd__nand2_1 U27339 ( .A(n12449), .B(n26323), .Y(n21818) );
  sky130_fd_sc_hd__nand2_1 U27340 ( .A(n21820), .B(n26711), .Y(n21841) );
  sky130_fd_sc_hd__nand2_1 U27341 ( .A(n21823), .B(n21822), .Y(n21825) );
  sky130_fd_sc_hd__xor2_1 U27342 ( .A(n21825), .B(n21824), .X(n24062) );
  sky130_fd_sc_hd__nand2_1 U27343 ( .A(n24062), .B(n22927), .Y(n22251) );
  sky130_fd_sc_hd__xnor2_1 U27344 ( .A(n26711), .B(n27415), .Y(n26631) );
  sky130_fd_sc_hd__o2bb2ai_1 U27345 ( .B1(n26415), .B2(n26631), .A1_N(n27365), 
        .A2_N(n26338), .Y(n21830) );
  sky130_fd_sc_hd__nand2b_1 U27346 ( .A_N(n22925), .B(
        j202_soc_core_j22_cpu_ml_macl[5]), .Y(n22250) );
  sky130_fd_sc_hd__nand2_1 U27347 ( .A(n22250), .B(n22247), .Y(n21826) );
  sky130_fd_sc_hd__nand2_1 U27348 ( .A(n21826), .B(n26329), .Y(n21828) );
  sky130_fd_sc_hd__o22a_1 U27349 ( .A1(n26713), .A2(n26419), .B1(n25798), .B2(
        n26418), .X(n21827) );
  sky130_fd_sc_hd__o211ai_1 U27350 ( .A1(n27007), .A2(n26427), .B1(n21828), 
        .C1(n21827), .Y(n21829) );
  sky130_fd_sc_hd__nor2_1 U27351 ( .A(n21830), .B(n21829), .Y(n21835) );
  sky130_fd_sc_hd__a21oi_1 U27352 ( .A1(n26341), .A2(n27183), .B1(n21831), .Y(
        n21834) );
  sky130_fd_sc_hd__mux2_2 U27353 ( .A0(n26423), .A1(n22722), .S(n27415), .X(
        n21833) );
  sky130_fd_sc_hd__nand2_1 U27354 ( .A(n26342), .B(n27412), .Y(n21832) );
  sky130_fd_sc_hd__nand4_1 U27355 ( .A(n21835), .B(n21834), .C(n21833), .D(
        n21832), .Y(n21836) );
  sky130_fd_sc_hd__a21oi_1 U27356 ( .A1(n26889), .A2(n26409), .B1(n21836), .Y(
        n21837) );
  sky130_fd_sc_hd__o21a_1 U27357 ( .A1(n18916), .A2(n22251), .B1(n21837), .X(
        n21840) );
  sky130_fd_sc_hd__o21ai_1 U27358 ( .A1(n26352), .A2(n26711), .B1(n26351), .Y(
        n21838) );
  sky130_fd_sc_hd__nand2_1 U27359 ( .A(n12449), .B(n21838), .Y(n21839) );
  sky130_fd_sc_hd__nand2_1 U27360 ( .A(n21842), .B(n24381), .Y(n21844) );
  sky130_fd_sc_hd__nand3_2 U27361 ( .A(n21844), .B(n22768), .C(n24383), .Y(
        n22257) );
  sky130_fd_sc_hd__o22ai_1 U27362 ( .A1(n21342), .A2(n22860), .B1(n22854), 
        .B2(n21845), .Y(n21846) );
  sky130_fd_sc_hd__a21oi_1 U27363 ( .A1(n22866), .A2(
        j202_soc_core_j22_cpu_rf_gpr[13]), .B1(n21846), .Y(n21851) );
  sky130_fd_sc_hd__a22oi_1 U27364 ( .A1(n21847), .A2(
        j202_soc_core_j22_cpu_rf_gbr[13]), .B1(n22864), .B2(
        j202_soc_core_j22_cpu_rf_vbr[13]), .Y(n21850) );
  sky130_fd_sc_hd__nand2_1 U27365 ( .A(n22865), .B(
        j202_soc_core_j22_cpu_rf_gpr[493]), .Y(n21849) );
  sky130_fd_sc_hd__nand2_1 U27366 ( .A(n22867), .B(
        j202_soc_core_j22_cpu_rf_tmp[13]), .Y(n21848) );
  sky130_fd_sc_hd__nand4_1 U27367 ( .A(n21851), .B(n21850), .C(n21849), .D(
        n21848), .Y(n21852) );
  sky130_fd_sc_hd__a21oi_1 U27368 ( .A1(n21853), .A2(n22873), .B1(n21852), .Y(
        n22452) );
  sky130_fd_sc_hd__nand2_1 U27369 ( .A(n21854), .B(n22873), .Y(n21866) );
  sky130_fd_sc_hd__o22ai_1 U27370 ( .A1(n21856), .A2(n22856), .B1(n21855), 
        .B2(n22854), .Y(n21859) );
  sky130_fd_sc_hd__o22ai_1 U27371 ( .A1(n21761), .A2(n22860), .B1(n21857), 
        .B2(n22858), .Y(n21858) );
  sky130_fd_sc_hd__nor2_1 U27372 ( .A(n21859), .B(n21858), .Y(n21865) );
  sky130_fd_sc_hd__o22ai_1 U27373 ( .A1(n21861), .A2(n22034), .B1(n21860), 
        .B2(n22033), .Y(n21863) );
  sky130_fd_sc_hd__a22o_1 U27374 ( .A1(j202_soc_core_j22_cpu_rf_gpr[485]), 
        .A2(n22865), .B1(n22864), .B2(j202_soc_core_j22_cpu_rf_vbr[5]), .X(
        n21862) );
  sky130_fd_sc_hd__nor2_1 U27375 ( .A(n21863), .B(n21862), .Y(n21864) );
  sky130_fd_sc_hd__nand3_1 U27376 ( .A(n21866), .B(n21865), .C(n21864), .Y(
        n22254) );
  sky130_fd_sc_hd__nand2_1 U27377 ( .A(n22254), .B(n22824), .Y(n22451) );
  sky130_fd_sc_hd__o21a_1 U27378 ( .A1(n22932), .A2(n22452), .B1(n22451), .X(
        n21901) );
  sky130_fd_sc_hd__nand2_1 U27379 ( .A(n21868), .B(n21867), .Y(n21869) );
  sky130_fd_sc_hd__nand2_1 U27380 ( .A(n21872), .B(n21871), .Y(n21885) );
  sky130_fd_sc_hd__nor2_1 U27381 ( .A(n12741), .B(n21873), .Y(n21880) );
  sky130_fd_sc_hd__nand2_1 U27382 ( .A(n21880), .B(n21874), .Y(n21883) );
  sky130_fd_sc_hd__o21ai_1 U27383 ( .A1(n12741), .A2(n21877), .B1(n21876), .Y(
        n21879) );
  sky130_fd_sc_hd__a21oi_1 U27384 ( .A1(n21881), .A2(n21880), .B1(n21879), .Y(
        n21882) );
  sky130_fd_sc_hd__o21ai_1 U27385 ( .A1(n21883), .A2(n22837), .B1(n21882), .Y(
        n21884) );
  sky130_fd_sc_hd__xnor2_1 U27386 ( .A(n21885), .B(n21884), .Y(n22437) );
  sky130_fd_sc_hd__nand2_1 U27387 ( .A(n22437), .B(n24499), .Y(n23042) );
  sky130_fd_sc_hd__nand2_1 U27388 ( .A(n25289), .B(n26398), .Y(n21898) );
  sky130_fd_sc_hd__o2bb2ai_1 U27389 ( .B1(n17585), .B2(n25338), .A1_N(
        j202_soc_core_j22_cpu_ml_mach[13]), .A2_N(n22936), .Y(n25290) );
  sky130_fd_sc_hd__nand2_1 U27390 ( .A(n22923), .B(n21887), .Y(n23049) );
  sky130_fd_sc_hd__a21oi_1 U27391 ( .A1(n25290), .A2(n26398), .B1(n21888), .Y(
        n21897) );
  sky130_fd_sc_hd__nand2_1 U27392 ( .A(n21891), .B(n21890), .Y(n21896) );
  sky130_fd_sc_hd__o21ai_1 U27393 ( .A1(n21894), .A2(n21893), .B1(n21892), .Y(
        n21895) );
  sky130_fd_sc_hd__xnor2_1 U27394 ( .A(n21896), .B(n21895), .Y(n26978) );
  sky130_fd_sc_hd__nand2_1 U27395 ( .A(n26978), .B(n22927), .Y(n23068) );
  sky130_fd_sc_hd__nand2b_1 U27396 ( .A_N(n22925), .B(
        j202_soc_core_j22_cpu_ml_macl[13]), .Y(n23050) );
  sky130_fd_sc_hd__nand4_1 U27397 ( .A(n21898), .B(n21897), .C(n23068), .D(
        n23050), .Y(n21899) );
  sky130_fd_sc_hd__nand2_1 U27398 ( .A(n21899), .B(n22929), .Y(n21900) );
  sky130_fd_sc_hd__nand2_1 U27399 ( .A(n28923), .B(n22581), .Y(n21908) );
  sky130_fd_sc_hd__o22a_1 U27400 ( .A1(n26791), .A2(n22590), .B1(n27007), .B2(
        n11143), .X(n21902) );
  sky130_fd_sc_hd__o21ai_1 U27401 ( .A1(n26791), .A2(n22592), .B1(n21902), .Y(
        n21903) );
  sky130_fd_sc_hd__a21oi_1 U27402 ( .A1(n24594), .A2(n12158), .B1(n21903), .Y(
        n21907) );
  sky130_fd_sc_hd__nand2_1 U27403 ( .A(n21904), .B(j202_soc_core_j22_cpu_pc[3]), .Y(n21905) );
  sky130_fd_sc_hd__xor2_1 U27404 ( .A(n21905), .B(n19453), .X(n25759) );
  sky130_fd_sc_hd__nand2_1 U27405 ( .A(n22596), .B(n25759), .Y(n21906) );
  sky130_fd_sc_hd__nand3_1 U27406 ( .A(n21908), .B(n21907), .C(n21906), .Y(
        n29034) );
  sky130_fd_sc_hd__nand2_1 U27407 ( .A(n22753), .B(n22751), .Y(n21913) );
  sky130_fd_sc_hd__o21ai_2 U27408 ( .A1(n21911), .A2(n22912), .B1(n21910), .Y(
        n21912) );
  sky130_fd_sc_hd__xnor2_2 U27409 ( .A(n21913), .B(n21912), .Y(n23231) );
  sky130_fd_sc_hd__nand2_1 U27410 ( .A(n28926), .B(n22712), .Y(n21917) );
  sky130_fd_sc_hd__nand2_1 U27411 ( .A(n21918), .B(n26723), .Y(n21949) );
  sky130_fd_sc_hd__nand2_1 U27412 ( .A(n21921), .B(n21920), .Y(n21922) );
  sky130_fd_sc_hd__xnor2_1 U27413 ( .A(n21923), .B(n21922), .Y(n23717) );
  sky130_fd_sc_hd__nand2_1 U27414 ( .A(n24602), .B(n22927), .Y(n22305) );
  sky130_fd_sc_hd__mux2i_1 U27415 ( .A0(n22722), .A1(n26423), .S(n23982), .Y(
        n21943) );
  sky130_fd_sc_hd__nand2_1 U27416 ( .A(n26342), .B(n27447), .Y(n21930) );
  sky130_fd_sc_hd__mux2i_1 U27417 ( .A0(n27341), .A1(n23928), .S(n27415), .Y(
        n21928) );
  sky130_fd_sc_hd__nand3_1 U27418 ( .A(n21928), .B(n23026), .C(n27435), .Y(
        n21929) );
  sky130_fd_sc_hd__nand2_1 U27419 ( .A(n21930), .B(n21929), .Y(n21942) );
  sky130_fd_sc_hd__a22oi_1 U27420 ( .A1(n26338), .A2(n27396), .B1(n26341), 
        .B2(n27045), .Y(n21940) );
  sky130_fd_sc_hd__nor2_1 U27421 ( .A(n21931), .B(n22925), .Y(n22303) );
  sky130_fd_sc_hd__a22oi_1 U27422 ( .A1(n26077), .A2(n26710), .B1(n22303), 
        .B2(n26329), .Y(n21939) );
  sky130_fd_sc_hd__nand2_1 U27423 ( .A(n27455), .B(n26723), .Y(n26746) );
  sky130_fd_sc_hd__nand2_1 U27424 ( .A(n22923), .B(n12613), .Y(n22300) );
  sky130_fd_sc_hd__nand3_1 U27425 ( .A(n21932), .B(
        j202_soc_core_j22_cpu_rfuo_sr__t_), .C(n26690), .Y(n21933) );
  sky130_fd_sc_hd__o22a_1 U27426 ( .A1(n18916), .A2(n22300), .B1(n21933), .B2(
        n24778), .X(n21935) );
  sky130_fd_sc_hd__nand2_1 U27427 ( .A(n23982), .B(n25789), .Y(n26626) );
  sky130_fd_sc_hd__nand3_1 U27428 ( .A(n26626), .B(n26326), .C(n26746), .Y(
        n21934) );
  sky130_fd_sc_hd__o211ai_1 U27429 ( .A1(n26432), .A2(n26746), .B1(n21935), 
        .C1(n21934), .Y(n21936) );
  sky130_fd_sc_hd__a21oi_1 U27430 ( .A1(n25131), .A2(n23920), .B1(n21936), .Y(
        n21938) );
  sky130_fd_sc_hd__nand2_1 U27431 ( .A(n25063), .B(n26603), .Y(n21937) );
  sky130_fd_sc_hd__nand4_1 U27432 ( .A(n21940), .B(n21939), .C(n21938), .D(
        n21937), .Y(n21941) );
  sky130_fd_sc_hd__nor3_1 U27433 ( .A(n21943), .B(n21942), .C(n21941), .Y(
        n21944) );
  sky130_fd_sc_hd__a21oi_1 U27435 ( .A1(n23717), .A2(n26409), .B1(n21945), .Y(
        n21948) );
  sky130_fd_sc_hd__o21ai_1 U27436 ( .A1(n26352), .A2(n26723), .B1(n26351), .Y(
        n21946) );
  sky130_fd_sc_hd__nand2_1 U27437 ( .A(n12417), .B(n21946), .Y(n21947) );
  sky130_fd_sc_hd__o22ai_1 U27438 ( .A1(n23928), .A2(n22856), .B1(n21950), 
        .B2(n22854), .Y(n21953) );
  sky130_fd_sc_hd__o22ai_1 U27439 ( .A1(n23720), .A2(n22860), .B1(n21951), 
        .B2(n22858), .Y(n21952) );
  sky130_fd_sc_hd__nor2_1 U27440 ( .A(n21953), .B(n21952), .Y(n21958) );
  sky130_fd_sc_hd__a22oi_1 U27441 ( .A1(n22865), .A2(
        j202_soc_core_j22_cpu_rf_gpr[480]), .B1(n22864), .B2(
        j202_soc_core_j22_cpu_rf_vbr[0]), .Y(n21957) );
  sky130_fd_sc_hd__o22a_1 U27442 ( .A1(n21955), .A2(n22034), .B1(n21954), .B2(
        n22033), .X(n21956) );
  sky130_fd_sc_hd__nand3_1 U27443 ( .A(n21958), .B(n21957), .C(n21956), .Y(
        n21959) );
  sky130_fd_sc_hd__a21oi_1 U27444 ( .A1(n21960), .A2(n22873), .B1(n21959), .Y(
        n22546) );
  sky130_fd_sc_hd__nand2_1 U27445 ( .A(n21962), .B(n22762), .Y(n21963) );
  sky130_fd_sc_hd__xor2_1 U27446 ( .A(n21961), .B(n21963), .X(n22533) );
  sky130_fd_sc_hd__nand2_1 U27447 ( .A(n22533), .B(n26862), .Y(n22298) );
  sky130_fd_sc_hd__a22oi_1 U27448 ( .A1(n12613), .A2(n27187), .B1(n22936), 
        .B2(j202_soc_core_j22_cpu_ml_mach[0]), .Y(n22299) );
  sky130_fd_sc_hd__nand2_1 U27449 ( .A(n22298), .B(n22299), .Y(n24168) );
  sky130_fd_sc_hd__nand2_1 U27450 ( .A(n24168), .B(n22459), .Y(n21964) );
  sky130_fd_sc_hd__nand2_1 U27452 ( .A(n21970), .B(n22845), .Y(n21971) );
  sky130_fd_sc_hd__xor2_1 U27453 ( .A(n22846), .B(n21971), .X(n25873) );
  sky130_fd_sc_hd__nand2_1 U27454 ( .A(n25873), .B(n22927), .Y(n25809) );
  sky130_fd_sc_hd__nand2b_1 U27455 ( .A_N(n22925), .B(
        j202_soc_core_j22_cpu_ml_macl[8]), .Y(n25792) );
  sky130_fd_sc_hd__nand2_1 U27456 ( .A(n25809), .B(n25792), .Y(n21989) );
  sky130_fd_sc_hd__nor2_1 U27457 ( .A(n25823), .B(n21972), .Y(n21985) );
  sky130_fd_sc_hd__nand2_1 U27458 ( .A(n25791), .B(n11713), .Y(n21988) );
  sky130_fd_sc_hd__nand2_1 U27459 ( .A(n21973), .B(n22906), .Y(n21979) );
  sky130_fd_sc_hd__nand2_1 U27460 ( .A(n22521), .B(n21975), .Y(n21977) );
  sky130_fd_sc_hd__o21ai_2 U27461 ( .A1(n21977), .A2(n22897), .B1(n21976), .Y(
        n21978) );
  sky130_fd_sc_hd__xnor2_2 U27462 ( .A(n21979), .B(n21978), .Y(n23235) );
  sky130_fd_sc_hd__nand2_1 U27463 ( .A(n22834), .B(n22832), .Y(n21984) );
  sky130_fd_sc_hd__xnor2_1 U27465 ( .A(n21984), .B(n21983), .Y(n22575) );
  sky130_fd_sc_hd__nand2_1 U27466 ( .A(n22575), .B(n26862), .Y(n25785) );
  sky130_fd_sc_hd__nand2_1 U27467 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[8]), .Y(n25784) );
  sky130_fd_sc_hd__nand2_1 U27468 ( .A(n25785), .B(n25784), .Y(n25787) );
  sky130_fd_sc_hd__nor2_1 U27469 ( .A(n21985), .B(n21989), .Y(n21986) );
  sky130_fd_sc_hd__nand2_1 U27470 ( .A(n25832), .B(n21986), .Y(n21987) );
  sky130_fd_sc_hd__o211ai_1 U27471 ( .A1(n21989), .A2(n21988), .B1(n22929), 
        .C1(n21987), .Y(n22006) );
  sky130_fd_sc_hd__nand2_1 U27472 ( .A(n21990), .B(n22873), .Y(n22003) );
  sky130_fd_sc_hd__o22ai_1 U27473 ( .A1(n21992), .A2(n22856), .B1(n21991), 
        .B2(n22854), .Y(n21996) );
  sky130_fd_sc_hd__o22ai_1 U27474 ( .A1(n21994), .A2(n22860), .B1(n22858), 
        .B2(n21993), .Y(n21995) );
  sky130_fd_sc_hd__nor2_1 U27475 ( .A(n21996), .B(n21995), .Y(n22002) );
  sky130_fd_sc_hd__o22ai_1 U27476 ( .A1(n21998), .A2(n22034), .B1(n21997), 
        .B2(n22033), .Y(n22000) );
  sky130_fd_sc_hd__a22o_1 U27477 ( .A1(j202_soc_core_j22_cpu_rf_gpr[488]), 
        .A2(n22865), .B1(n22864), .B2(j202_soc_core_j22_cpu_rf_vbr[8]), .X(
        n21999) );
  sky130_fd_sc_hd__nor2_1 U27478 ( .A(n22000), .B(n21999), .Y(n22001) );
  sky130_fd_sc_hd__nand3_1 U27479 ( .A(n22003), .B(n22002), .C(n22001), .Y(
        n22574) );
  sky130_fd_sc_hd__nand2_1 U27480 ( .A(n22574), .B(n22004), .Y(n22005) );
  sky130_fd_sc_hd__nand3_1 U27481 ( .A(n22580), .B(n22006), .C(n22005), .Y(
        n29007) );
  sky130_fd_sc_hd__nand3_1 U27482 ( .A(n24118), .B(n22668), .C(n29062), .Y(
        n22708) );
  sky130_fd_sc_hd__nor2_1 U27483 ( .A(n22711), .B(n22708), .Y(n29028) );
  sky130_fd_sc_hd__nand4_1 U27484 ( .A(n24135), .B(n22007), .C(n24134), .D(
        n24133), .Y(n22008) );
  sky130_fd_sc_hd__o21ai_1 U27485 ( .A1(n22009), .A2(n26398), .B1(n22008), .Y(
        n22012) );
  sky130_fd_sc_hd__nand3_1 U27486 ( .A(n22012), .B(n22011), .C(n22010), .Y(
        n22013) );
  sky130_fd_sc_hd__nand2_1 U27487 ( .A(n22013), .B(n22929), .Y(n22018) );
  sky130_fd_sc_hd__nand3_1 U27488 ( .A(n24135), .B(n11068), .C(n24134), .Y(
        n22016) );
  sky130_fd_sc_hd__inv_1 U27489 ( .A(n22014), .Y(n22015) );
  sky130_fd_sc_hd__nand2_1 U27490 ( .A(n22016), .B(n22015), .Y(n22983) );
  sky130_fd_sc_hd__nor2_1 U27491 ( .A(n23574), .B(n22039), .Y(n22318) );
  sky130_fd_sc_hd__nand2_1 U27492 ( .A(n22976), .B(n11158), .Y(n22017) );
  sky130_fd_sc_hd__nand3_1 U27493 ( .A(n22018), .B(n22983), .C(n22017), .Y(
        n29002) );
  sky130_fd_sc_hd__nand2_1 U27494 ( .A(n27773), .B(n27256), .Y(n22021) );
  sky130_fd_sc_hd__nor2_1 U27495 ( .A(n23821), .B(n22021), .Y(n22022) );
  sky130_fd_sc_hd__nand2_1 U27496 ( .A(n12728), .B(n27980), .Y(n22027) );
  sky130_fd_sc_hd__nand3_1 U27497 ( .A(n22025), .B(n22024), .C(n23195), .Y(
        n24469) );
  sky130_fd_sc_hd__nor2_1 U27498 ( .A(n26398), .B(n22978), .Y(n22654) );
  sky130_fd_sc_hd__o22ai_1 U27499 ( .A1(n25824), .A2(n17975), .B1(n22030), 
        .B2(n22952), .Y(n22031) );
  sky130_fd_sc_hd__a21oi_1 U27500 ( .A1(n22032), .A2(n26872), .B1(n22031), .Y(
        n25182) );
  sky130_fd_sc_hd__nand2_1 U27501 ( .A(n24742), .B(n22956), .Y(n25178) );
  sky130_fd_sc_hd__nand2_1 U27502 ( .A(n22864), .B(n22039), .Y(n22877) );
  sky130_fd_sc_hd__nand2_1 U27503 ( .A(n22957), .B(
        j202_soc_core_j22_cpu_rf_vbr[23]), .Y(n22038) );
  sky130_fd_sc_hd__nand2_1 U27504 ( .A(n22865), .B(n22039), .Y(n22875) );
  sky130_fd_sc_hd__nand2_1 U27505 ( .A(n22958), .B(
        j202_soc_core_j22_cpu_rf_gpr[503]), .Y(n22037) );
  sky130_fd_sc_hd__nor2_1 U27506 ( .A(n22033), .B(n23302), .Y(n22959) );
  sky130_fd_sc_hd__nand2_1 U27507 ( .A(n22959), .B(
        j202_soc_core_j22_cpu_rf_tmp[23]), .Y(n22036) );
  sky130_fd_sc_hd__nor2_1 U27508 ( .A(n22034), .B(n23302), .Y(n22960) );
  sky130_fd_sc_hd__nand2_1 U27509 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[23]), .Y(n22035) );
  sky130_fd_sc_hd__nand4_1 U27510 ( .A(n22038), .B(n22037), .C(n22036), .D(
        n22035), .Y(n22044) );
  sky130_fd_sc_hd__nand2_1 U27511 ( .A(n22040), .B(n22969), .Y(n22043) );
  sky130_fd_sc_hd__nor2_1 U27512 ( .A(n22860), .B(n23302), .Y(n22966) );
  sky130_fd_sc_hd__nand2_1 U27513 ( .A(n22965), .B(n22029), .Y(n25166) );
  sky130_fd_sc_hd__a2bb2oi_1 U27514 ( .B1(j202_soc_core_j22_cpu_pc[23]), .B2(
        n22966), .A1_N(n22978), .A2_N(n25166), .Y(n22042) );
  sky130_fd_sc_hd__nor2_1 U27515 ( .A(n22854), .B(n23302), .Y(n22968) );
  sky130_fd_sc_hd__nor2_1 U27516 ( .A(n22858), .B(n23302), .Y(n22967) );
  sky130_fd_sc_hd__a22oi_1 U27517 ( .A1(n22968), .A2(
        j202_soc_core_j22_cpu_rf_pr[23]), .B1(j202_soc_core_j22_cpu_rf_gbr[23]), .B2(n22967), .Y(n22041) );
  sky130_fd_sc_hd__nand4b_1 U27518 ( .A_N(n22044), .B(n22043), .C(n22042), .D(
        n22041), .Y(n22045) );
  sky130_fd_sc_hd__a21oi_1 U27519 ( .A1(n22226), .A2(n23574), .B1(n22045), .Y(
        n22046) );
  sky130_fd_sc_hd__o21a_1 U27520 ( .A1(n22978), .A2(n25178), .B1(n22046), .X(
        n22047) );
  sky130_fd_sc_hd__o21a_1 U27521 ( .A1(n22980), .A2(n25182), .B1(n22047), .X(
        n22111) );
  sky130_fd_sc_hd__nand2_1 U27522 ( .A(n23240), .B(n24499), .Y(n22109) );
  sky130_fd_sc_hd__nor2_1 U27523 ( .A(n12159), .B(n22048), .Y(n22074) );
  sky130_fd_sc_hd__nor2_1 U27524 ( .A(n12159), .B(n22049), .Y(n22390) );
  sky130_fd_sc_hd__nor2_1 U27525 ( .A(n22074), .B(n22050), .Y(n22555) );
  sky130_fd_sc_hd__nand2_1 U27526 ( .A(n22050), .B(n22074), .Y(n22554) );
  sky130_fd_sc_hd__nand2_1 U27527 ( .A(n22388), .B(n22554), .Y(n22108) );
  sky130_fd_sc_hd__xnor2_1 U27528 ( .A(n22052), .B(n22051), .Y(n22053) );
  sky130_fd_sc_hd__o22ai_1 U27529 ( .A1(n12159), .A2(n22056), .B1(n22055), 
        .B2(n22054), .Y(n22067) );
  sky130_fd_sc_hd__fa_1 U27530 ( .A(n22061), .B(n22060), .CIN(n22059), .COUT(
        n22076), .SUM(n17383) );
  sky130_fd_sc_hd__nor2_1 U27531 ( .A(n12135), .B(n22062), .Y(n22086) );
  sky130_fd_sc_hd__nor2_1 U27532 ( .A(n12135), .B(n22063), .Y(n22064) );
  sky130_fd_sc_hd__nor2_1 U27533 ( .A(n22079), .B(n22080), .Y(n22177) );
  sky130_fd_sc_hd__fa_1 U27534 ( .A(n22065), .B(n22068), .CIN(n22064), .COUT(
        n22080), .SUM(n22077) );
  sky130_fd_sc_hd__fa_1 U27535 ( .A(n22068), .B(n22067), .CIN(n22066), .COUT(
        n22078), .SUM(n22075) );
  sky130_fd_sc_hd__nor2_1 U27536 ( .A(n22077), .B(n22078), .Y(n22794) );
  sky130_fd_sc_hd__nor2_1 U27537 ( .A(n22177), .B(n22794), .Y(n22083) );
  sky130_fd_sc_hd__nand2_1 U27538 ( .A(n22520), .B(n22083), .Y(n22085) );
  sky130_fd_sc_hd__nor2_1 U27539 ( .A(n22085), .B(n22069), .Y(n22160) );
  sky130_fd_sc_hd__nor2_1 U27540 ( .A(n12135), .B(n22070), .Y(n22088) );
  sky130_fd_sc_hd__o21ai_1 U27541 ( .A1(n12159), .A2(n22072), .B1(n22071), .Y(
        n22094) );
  sky130_fd_sc_hd__nor2_1 U27542 ( .A(n22088), .B(n22089), .Y(n22157) );
  sky130_fd_sc_hd__nor2_1 U27543 ( .A(n22086), .B(n22087), .Y(n22937) );
  sky130_fd_sc_hd__nor2_1 U27544 ( .A(n22157), .B(n22937), .Y(n22091) );
  sky130_fd_sc_hd__nand2_1 U27545 ( .A(n22160), .B(n22091), .Y(n22093) );
  sky130_fd_sc_hd__nor2_1 U27546 ( .A(n12159), .B(n22073), .Y(n22096) );
  sky130_fd_sc_hd__nor2_1 U27547 ( .A(n22094), .B(n22095), .Y(n22361) );
  sky130_fd_sc_hd__nand2_1 U27548 ( .A(n22471), .B(n22103), .Y(n22890) );
  sky130_fd_sc_hd__nand2_1 U27549 ( .A(n22076), .B(n22075), .Y(n22519) );
  sky130_fd_sc_hd__nand2_1 U27550 ( .A(n22078), .B(n22077), .Y(n22795) );
  sky130_fd_sc_hd__nand2_1 U27551 ( .A(n22080), .B(n22079), .Y(n22178) );
  sky130_fd_sc_hd__a21oi_1 U27553 ( .A1(n22083), .A2(n22082), .B1(n22081), .Y(
        n22084) );
  sky130_fd_sc_hd__nand2_1 U27555 ( .A(n22087), .B(n22086), .Y(n22938) );
  sky130_fd_sc_hd__nand2_1 U27556 ( .A(n22089), .B(n22088), .Y(n22158) );
  sky130_fd_sc_hd__o21ai_1 U27557 ( .A1(n22938), .A2(n22157), .B1(n22158), .Y(
        n22090) );
  sky130_fd_sc_hd__a21oi_1 U27558 ( .A1(n22161), .A2(n22091), .B1(n22090), .Y(
        n22092) );
  sky130_fd_sc_hd__nand2_1 U27559 ( .A(n22095), .B(n22094), .Y(n22359) );
  sky130_fd_sc_hd__nand2_1 U27560 ( .A(n22097), .B(n22096), .Y(n22356) );
  sky130_fd_sc_hd__inv_1 U27561 ( .A(n22892), .Y(n22104) );
  sky130_fd_sc_hd__a21oi_1 U27562 ( .A1(n22944), .A2(n22105), .B1(n22104), .Y(
        n22106) );
  sky130_fd_sc_hd__nor2_1 U27563 ( .A(n11713), .B(n22978), .Y(n22950) );
  sky130_fd_sc_hd__nand2_1 U27564 ( .A(n26068), .B(n22950), .Y(n22110) );
  sky130_fd_sc_hd__nand3_1 U27565 ( .A(n22234), .B(n22111), .C(n22110), .Y(
        n28992) );
  sky130_fd_sc_hd__o22ai_1 U27566 ( .A1(n25824), .A2(n22114), .B1(n22113), 
        .B2(n22952), .Y(n22115) );
  sky130_fd_sc_hd__a21oi_1 U27567 ( .A1(n22116), .A2(n26872), .B1(n22115), .Y(
        n25398) );
  sky130_fd_sc_hd__nand2_1 U27568 ( .A(n24062), .B(n22956), .Y(n25397) );
  sky130_fd_sc_hd__nand2_1 U27569 ( .A(n22957), .B(
        j202_soc_core_j22_cpu_rf_vbr[21]), .Y(n22120) );
  sky130_fd_sc_hd__nand2_1 U27570 ( .A(n22958), .B(
        j202_soc_core_j22_cpu_rf_gpr[501]), .Y(n22119) );
  sky130_fd_sc_hd__nand2_1 U27571 ( .A(n22959), .B(
        j202_soc_core_j22_cpu_rf_tmp[21]), .Y(n22118) );
  sky130_fd_sc_hd__nand2_1 U27572 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[21]), .Y(n22117) );
  sky130_fd_sc_hd__nand4_1 U27573 ( .A(n22120), .B(n22119), .C(n22118), .D(
        n22117), .Y(n22125) );
  sky130_fd_sc_hd__nand2_1 U27574 ( .A(n22965), .B(n22112), .Y(n25393) );
  sky130_fd_sc_hd__a2bb2oi_1 U27575 ( .B1(j202_soc_core_j22_cpu_rf_pr[21]), 
        .B2(n22968), .A1_N(n22978), .A2_N(n25393), .Y(n22124) );
  sky130_fd_sc_hd__a22oi_1 U27576 ( .A1(n22966), .A2(
        j202_soc_core_j22_cpu_pc[21]), .B1(j202_soc_core_j22_cpu_rf_gbr[21]), 
        .B2(n22967), .Y(n22123) );
  sky130_fd_sc_hd__nand2_1 U27577 ( .A(n22121), .B(n22969), .Y(n22122) );
  sky130_fd_sc_hd__nand4b_1 U27578 ( .A_N(n22125), .B(n22124), .C(n22123), .D(
        n22122), .Y(n22126) );
  sky130_fd_sc_hd__a21oi_1 U27579 ( .A1(n22254), .A2(n23574), .B1(n22126), .Y(
        n22127) );
  sky130_fd_sc_hd__o21a_1 U27580 ( .A1(n22978), .A2(n25397), .B1(n22127), .X(
        n22128) );
  sky130_fd_sc_hd__o21a_1 U27581 ( .A1(n22980), .A2(n25398), .B1(n22128), .X(
        n22140) );
  sky130_fd_sc_hd__nand2_1 U27582 ( .A(n23230), .B(n26862), .Y(n25396) );
  sky130_fd_sc_hd__nand2_1 U27583 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[21]), .Y(n25394) );
  sky130_fd_sc_hd__nand2_1 U27584 ( .A(n22129), .B(n22359), .Y(n22137) );
  sky130_fd_sc_hd__nand2_1 U27585 ( .A(n22471), .B(n22131), .Y(n22358) );
  sky130_fd_sc_hd__a21oi_1 U27586 ( .A1(n22398), .A2(n22131), .B1(n22130), .Y(
        n22360) );
  sky130_fd_sc_hd__a21oi_1 U27587 ( .A1(n22944), .A2(n22133), .B1(n22132), .Y(
        n22134) );
  sky130_fd_sc_hd__o21ai_1 U27588 ( .A1(n22135), .A2(n22897), .B1(n22134), .Y(
        n22136) );
  sky130_fd_sc_hd__xnor2_1 U27589 ( .A(n22137), .B(n22136), .Y(n22138) );
  sky130_fd_sc_hd__nand2_1 U27590 ( .A(n22138), .B(n26863), .Y(n25395) );
  sky130_fd_sc_hd__nand3_1 U27591 ( .A(n25396), .B(n25394), .C(n25395), .Y(
        n27186) );
  sky130_fd_sc_hd__nand2_1 U27592 ( .A(n27186), .B(n22950), .Y(n22139) );
  sky130_fd_sc_hd__nand3_1 U27593 ( .A(n22257), .B(n22140), .C(n22139), .Y(
        n28990) );
  sky130_fd_sc_hd__o22ai_1 U27594 ( .A1(n25824), .A2(n22142), .B1(n22141), 
        .B2(n22952), .Y(n22143) );
  sky130_fd_sc_hd__a21oi_1 U27595 ( .A1(n22144), .A2(n26872), .B1(n22143), .Y(
        n24538) );
  sky130_fd_sc_hd__nand2_1 U27596 ( .A(n24586), .B(n22956), .Y(n24529) );
  sky130_fd_sc_hd__nand2_1 U27597 ( .A(n22957), .B(
        j202_soc_core_j22_cpu_rf_vbr[20]), .Y(n22148) );
  sky130_fd_sc_hd__nand2_1 U27598 ( .A(n22958), .B(
        j202_soc_core_j22_cpu_rf_gpr[500]), .Y(n22147) );
  sky130_fd_sc_hd__nand2_1 U27599 ( .A(n22959), .B(
        j202_soc_core_j22_cpu_rf_tmp[20]), .Y(n22146) );
  sky130_fd_sc_hd__nand2_1 U27600 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[20]), .Y(n22145) );
  sky130_fd_sc_hd__nand4_1 U27601 ( .A(n22148), .B(n22147), .C(n22146), .D(
        n22145), .Y(n22153) );
  sky130_fd_sc_hd__nand2_1 U27602 ( .A(n22965), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .Y(n24519) );
  sky130_fd_sc_hd__a2bb2oi_1 U27603 ( .B1(j202_soc_core_j22_cpu_rf_pr[20]), 
        .B2(n22968), .A1_N(n22978), .A2_N(n24519), .Y(n22152) );
  sky130_fd_sc_hd__a22oi_1 U27604 ( .A1(n22966), .A2(
        j202_soc_core_j22_cpu_pc[20]), .B1(j202_soc_core_j22_cpu_rf_gbr[20]), 
        .B2(n22967), .Y(n22151) );
  sky130_fd_sc_hd__nand2_1 U27605 ( .A(n22149), .B(n22969), .Y(n22150) );
  sky130_fd_sc_hd__nand4b_1 U27606 ( .A_N(n22153), .B(n22152), .C(n22151), .D(
        n22150), .Y(n22154) );
  sky130_fd_sc_hd__a21oi_1 U27607 ( .A1(n23574), .A2(n22268), .B1(n22154), .Y(
        n22155) );
  sky130_fd_sc_hd__o21a_1 U27608 ( .A1(n22978), .A2(n24529), .B1(n22155), .X(
        n22156) );
  sky130_fd_sc_hd__o21a_1 U27609 ( .A1(n22980), .A2(n24538), .B1(n22156), .X(
        n22176) );
  sky130_fd_sc_hd__nand2_1 U27610 ( .A(n23243), .B(n24499), .Y(n22174) );
  sky130_fd_sc_hd__nand2_1 U27611 ( .A(n22159), .B(n22158), .Y(n22171) );
  sky130_fd_sc_hd__nor2_1 U27612 ( .A(n22163), .B(n22180), .Y(n22165) );
  sky130_fd_sc_hd__nand2_1 U27613 ( .A(n22471), .B(n22165), .Y(n22940) );
  sky130_fd_sc_hd__nor2_1 U27614 ( .A(n22937), .B(n22940), .Y(n22167) );
  sky130_fd_sc_hd__o21ai_1 U27615 ( .A1(n22163), .A2(n22182), .B1(n22162), .Y(
        n22164) );
  sky130_fd_sc_hd__a21oi_1 U27617 ( .A1(n22944), .A2(n22167), .B1(n22166), .Y(
        n22168) );
  sky130_fd_sc_hd__o21ai_1 U27618 ( .A1(n22169), .A2(n22897), .B1(n22168), .Y(
        n22170) );
  sky130_fd_sc_hd__xnor2_1 U27619 ( .A(n22171), .B(n22170), .Y(n22172) );
  sky130_fd_sc_hd__a22oi_1 U27620 ( .A1(j202_soc_core_j22_cpu_ml_mach[20]), 
        .A2(n22936), .B1(n22172), .B2(n26863), .Y(n22173) );
  sky130_fd_sc_hd__nand2_1 U27621 ( .A(n26472), .B(n22950), .Y(n22175) );
  sky130_fd_sc_hd__nand3_1 U27622 ( .A(n12387), .B(n22176), .C(n22175), .Y(
        n28989) );
  sky130_fd_sc_hd__nand2_1 U27623 ( .A(n22179), .B(n22178), .Y(n22195) );
  sky130_fd_sc_hd__nand2_1 U27624 ( .A(n22181), .B(n22185), .Y(n22523) );
  sky130_fd_sc_hd__nor2_1 U27625 ( .A(n22187), .B(n22523), .Y(n22189) );
  sky130_fd_sc_hd__nand2_1 U27626 ( .A(n22471), .B(n22189), .Y(n22797) );
  sky130_fd_sc_hd__nor2_1 U27627 ( .A(n22794), .B(n22797), .Y(n22191) );
  sky130_fd_sc_hd__a21oi_1 U27628 ( .A1(n22186), .A2(n22185), .B1(n22184), .Y(
        n22522) );
  sky130_fd_sc_hd__o21ai_1 U27629 ( .A1(n22187), .A2(n22522), .B1(n22519), .Y(
        n22188) );
  sky130_fd_sc_hd__xnor2_1 U27631 ( .A(n22195), .B(n22194), .Y(n22196) );
  sky130_fd_sc_hd__nand2_1 U27632 ( .A(n22196), .B(n26863), .Y(n25250) );
  sky130_fd_sc_hd__nand2_1 U27633 ( .A(n22197), .B(n26872), .Y(n22201) );
  sky130_fd_sc_hd__o22ai_1 U27634 ( .A1(n25824), .A2(n22202), .B1(n22198), 
        .B2(n22952), .Y(n22199) );
  sky130_fd_sc_hd__a21oi_1 U27635 ( .A1(n24805), .A2(n26977), .B1(n22199), .Y(
        n22200) );
  sky130_fd_sc_hd__nand2_1 U27636 ( .A(n22201), .B(n22200), .Y(n25254) );
  sky130_fd_sc_hd__nand2_1 U27637 ( .A(n22968), .B(
        j202_soc_core_j22_cpu_rf_pr[18]), .Y(n22206) );
  sky130_fd_sc_hd__nand2_1 U27638 ( .A(n22966), .B(
        j202_soc_core_j22_cpu_pc[18]), .Y(n22205) );
  sky130_fd_sc_hd__nor2_1 U27639 ( .A(n22202), .B(n25338), .Y(n25247) );
  sky130_fd_sc_hd__nand2_1 U27640 ( .A(n22950), .B(n25247), .Y(n22204) );
  sky130_fd_sc_hd__nand2_1 U27641 ( .A(n22967), .B(
        j202_soc_core_j22_cpu_rf_gbr[18]), .Y(n22203) );
  sky130_fd_sc_hd__nand4_1 U27642 ( .A(n22206), .B(n22205), .C(n22204), .D(
        n22203), .Y(n22212) );
  sky130_fd_sc_hd__nand2_1 U27643 ( .A(n22957), .B(
        j202_soc_core_j22_cpu_rf_vbr[18]), .Y(n22210) );
  sky130_fd_sc_hd__nand2_1 U27644 ( .A(n22958), .B(
        j202_soc_core_j22_cpu_rf_gpr[498]), .Y(n22209) );
  sky130_fd_sc_hd__nand2_1 U27645 ( .A(n22959), .B(
        j202_soc_core_j22_cpu_rf_tmp[18]), .Y(n22208) );
  sky130_fd_sc_hd__nand2_1 U27646 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[18]), .Y(n22207) );
  sky130_fd_sc_hd__nand4_1 U27647 ( .A(n22210), .B(n22209), .C(n22208), .D(
        n22207), .Y(n22211) );
  sky130_fd_sc_hd__a211oi_1 U27648 ( .A1(n22213), .A2(n22969), .B1(n22212), 
        .C1(n22211), .Y(n22215) );
  sky130_fd_sc_hd__nand2_1 U27649 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[18]), .Y(n25249) );
  sky130_fd_sc_hd__nand2b_1 U27650 ( .A_N(n25249), .B(n22950), .Y(n22214) );
  sky130_fd_sc_hd__o211ai_1 U27651 ( .A1(n22545), .A2(n22317), .B1(n22215), 
        .C1(n22214), .Y(n22216) );
  sky130_fd_sc_hd__a21oi_1 U27652 ( .A1(n25254), .A2(n22654), .B1(n22216), .Y(
        n22217) );
  sky130_fd_sc_hd__nand2_1 U27653 ( .A(n11055), .B(n22218), .Y(n25243) );
  sky130_fd_sc_hd__nand2_1 U27654 ( .A(n25243), .B(n22219), .Y(n22319) );
  sky130_fd_sc_hd__nand2_1 U27655 ( .A(n22224), .B(n22223), .Y(n22225) );
  sky130_fd_sc_hd__a22oi_1 U27656 ( .A1(n11158), .A2(n22226), .B1(n22225), 
        .B2(n22929), .Y(n22233) );
  sky130_fd_sc_hd__nand2_1 U27658 ( .A(n25545), .B(n22230), .Y(n22231) );
  sky130_fd_sc_hd__nand2_1 U27659 ( .A(n22231), .B(n22929), .Y(n22232) );
  sky130_fd_sc_hd__nand3_1 U27660 ( .A(n22234), .B(n22233), .C(n22232), .Y(
        n29006) );
  sky130_fd_sc_hd__nand4_1 U27661 ( .A(n23275), .B(n25336), .C(n23274), .D(
        n22235), .Y(n22236) );
  sky130_fd_sc_hd__nand2_1 U27662 ( .A(n22241), .B(n22929), .Y(n22246) );
  sky130_fd_sc_hd__nand2_1 U27663 ( .A(n23278), .B(n29535), .Y(n22244) );
  sky130_fd_sc_hd__nand4_1 U27664 ( .A(n24382), .B(n22450), .C(n24380), .D(
        n22247), .Y(n22249) );
  sky130_fd_sc_hd__nand2_1 U27665 ( .A(n22247), .B(n11713), .Y(n22248) );
  sky130_fd_sc_hd__nand2_1 U27666 ( .A(n22249), .B(n22248), .Y(n22252) );
  sky130_fd_sc_hd__nand3_1 U27667 ( .A(n22252), .B(n22251), .C(n22250), .Y(
        n22253) );
  sky130_fd_sc_hd__nand2_1 U27668 ( .A(n22253), .B(n22929), .Y(n22256) );
  sky130_fd_sc_hd__nand2_1 U27669 ( .A(n22254), .B(n11158), .Y(n22255) );
  sky130_fd_sc_hd__nand4_1 U27670 ( .A(n24367), .B(n22259), .C(n22258), .D(
        n22260), .Y(n22262) );
  sky130_fd_sc_hd__nand2_1 U27671 ( .A(n22260), .B(n11713), .Y(n22261) );
  sky130_fd_sc_hd__nand2_1 U27672 ( .A(n22262), .B(n22261), .Y(n22266) );
  sky130_fd_sc_hd__nand3_1 U27673 ( .A(n22266), .B(n22265), .C(n22264), .Y(
        n22267) );
  sky130_fd_sc_hd__nand2_1 U27674 ( .A(n22267), .B(n22929), .Y(n22271) );
  sky130_fd_sc_hd__nand2_1 U27675 ( .A(n22268), .B(n11158), .Y(n22269) );
  sky130_fd_sc_hd__nand3_1 U27676 ( .A(n12387), .B(n22271), .C(n22269), .Y(
        n29003) );
  sky130_fd_sc_hd__nand3_1 U27677 ( .A(n23862), .B(n22275), .C(
        j202_soc_core_j22_cpu_opst[1]), .Y(n23597) );
  sky130_fd_sc_hd__nand2b_1 U27678 ( .A_N(n27956), .B(n22276), .Y(n27175) );
  sky130_fd_sc_hd__o21ai_1 U27679 ( .A1(j202_soc_core_j22_cpu_opst[2]), .A2(
        n27175), .B1(n27176), .Y(n22283) );
  sky130_fd_sc_hd__a31oi_1 U27680 ( .A1(n27260), .A2(n13272), .A3(n29075), 
        .B1(n22279), .Y(n22280) );
  sky130_fd_sc_hd__mux2i_1 U27681 ( .A0(n25048), .A1(n29015), .S(n11133), .Y(
        n22285) );
  sky130_fd_sc_hd__nand2_1 U27682 ( .A(n23141), .B(n12757), .Y(n22286) );
  sky130_fd_sc_hd__nand2_1 U27683 ( .A(n28926), .B(n22581), .Y(n22295) );
  sky130_fd_sc_hd__nand2_1 U27684 ( .A(n23717), .B(n12158), .Y(n22292) );
  sky130_fd_sc_hd__nand2_1 U27685 ( .A(n22596), .B(j202_soc_core_j22_cpu_pc[0]), .Y(n22291) );
  sky130_fd_sc_hd__nand2_1 U27686 ( .A(n22510), .B(n26723), .Y(n22290) );
  sky130_fd_sc_hd__and3_1 U27687 ( .A(n22292), .B(n22291), .C(n22290), .X(
        n22294) );
  sky130_fd_sc_hd__nand2_1 U27688 ( .A(n22515), .B(n27455), .Y(n22293) );
  sky130_fd_sc_hd__nor2_1 U27689 ( .A(n27622), .B(n12459), .Y(n28964) );
  sky130_fd_sc_hd__and3_1 U27690 ( .A(n22296), .B(j202_soc_core_aquc_CE__1_), 
        .C(j202_soc_core_aquc_SEL__0_), .X(n29029) );
  sky130_fd_sc_hd__nand2_1 U27691 ( .A(j202_soc_core_aquc_WE_), .B(
        j202_soc_core_aquc_CE__1_), .Y(n24572) );
  sky130_fd_sc_hd__nor2_1 U27692 ( .A(n22297), .B(n24572), .Y(n28967) );
  sky130_fd_sc_hd__nand4_1 U27693 ( .A(n24166), .B(n22299), .C(n22298), .D(
        n22300), .Y(n22302) );
  sky130_fd_sc_hd__nand2_1 U27694 ( .A(n22300), .B(n11713), .Y(n22301) );
  sky130_fd_sc_hd__nand2_1 U27695 ( .A(n22302), .B(n22301), .Y(n22306) );
  sky130_fd_sc_hd__nand2_1 U27696 ( .A(n22307), .B(n22929), .Y(n22309) );
  sky130_fd_sc_hd__nand2b_1 U27697 ( .A_N(n22546), .B(n11158), .Y(n22308) );
  sky130_fd_sc_hd__nand4_1 U27698 ( .A(n22311), .B(n22312), .C(n25230), .D(
        n22310), .Y(n22315) );
  sky130_fd_sc_hd__nand2_1 U27699 ( .A(n22312), .B(n11713), .Y(n22314) );
  sky130_fd_sc_hd__a21oi_1 U27700 ( .A1(n22315), .A2(n22314), .B1(n22313), .Y(
        n22316) );
  sky130_fd_sc_hd__nand2_1 U27701 ( .A(n28971), .B(n22581), .Y(n22336) );
  sky130_fd_sc_hd__nand2_1 U27702 ( .A(n22321), .B(j202_soc_core_j22_cpu_pc[9]), .Y(n22322) );
  sky130_fd_sc_hd__xor2_1 U27703 ( .A(n22322), .B(n19213), .X(n25053) );
  sky130_fd_sc_hd__o22a_1 U27704 ( .A1(n26325), .A2(n11143), .B1(n25057), .B2(
        n22590), .X(n22323) );
  sky130_fd_sc_hd__o21ai_1 U27705 ( .A1(n25057), .A2(n22592), .B1(n22323), .Y(
        n22324) );
  sky130_fd_sc_hd__a21oi_1 U27706 ( .A1(n25053), .A2(n22596), .B1(n22324), .Y(
        n22335) );
  sky130_fd_sc_hd__a21oi_1 U27707 ( .A1(n22328), .A2(n22327), .B1(n22326), .Y(
        n22333) );
  sky130_fd_sc_hd__nand2_1 U27708 ( .A(n22331), .B(n22330), .Y(n22332) );
  sky130_fd_sc_hd__xor2_1 U27709 ( .A(n22333), .B(n22332), .X(n25042) );
  sky130_fd_sc_hd__nand2_1 U27710 ( .A(n25042), .B(n12158), .Y(n22334) );
  sky130_fd_sc_hd__nand3_1 U27711 ( .A(n22336), .B(n22335), .C(n22334), .Y(
        n29063) );
  sky130_fd_sc_hd__o22ai_1 U27712 ( .A1(n25824), .A2(n22338), .B1(n22337), 
        .B2(n22952), .Y(n22339) );
  sky130_fd_sc_hd__a21oi_1 U27713 ( .A1(n22340), .A2(n26872), .B1(n22339), .Y(
        n26101) );
  sky130_fd_sc_hd__nand2_1 U27714 ( .A(n22957), .B(
        j202_soc_core_j22_cpu_rf_vbr[22]), .Y(n22344) );
  sky130_fd_sc_hd__nand2_1 U27715 ( .A(n22958), .B(
        j202_soc_core_j22_cpu_rf_gpr[502]), .Y(n22343) );
  sky130_fd_sc_hd__nand2_1 U27716 ( .A(n22959), .B(
        j202_soc_core_j22_cpu_rf_tmp[22]), .Y(n22342) );
  sky130_fd_sc_hd__nand2_1 U27717 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[22]), .Y(n22341) );
  sky130_fd_sc_hd__nand4_1 U27718 ( .A(n22344), .B(n22343), .C(n22342), .D(
        n22341), .Y(n22350) );
  sky130_fd_sc_hd__a22oi_1 U27719 ( .A1(n22966), .A2(
        j202_soc_core_j22_cpu_pc[22]), .B1(j202_soc_core_j22_cpu_rf_gbr[22]), 
        .B2(n22967), .Y(n22348) );
  sky130_fd_sc_hd__nand2_1 U27720 ( .A(n22345), .B(n22969), .Y(n22347) );
  sky130_fd_sc_hd__nand2_1 U27721 ( .A(n22965), .B(n12725), .Y(n26083) );
  sky130_fd_sc_hd__a2bb2oi_1 U27722 ( .B1(j202_soc_core_j22_cpu_rf_pr[22]), 
        .B2(n22968), .A1_N(n22978), .A2_N(n26083), .Y(n22346) );
  sky130_fd_sc_hd__nand3_1 U27723 ( .A(n22348), .B(n22347), .C(n22346), .Y(
        n22349) );
  sky130_fd_sc_hd__nor2_1 U27724 ( .A(n22350), .B(n22349), .Y(n22351) );
  sky130_fd_sc_hd__nand2_1 U27726 ( .A(n25345), .B(n22956), .Y(n26093) );
  sky130_fd_sc_hd__nor2_1 U27727 ( .A(n22978), .B(n26093), .Y(n22353) );
  sky130_fd_sc_hd__nor2_1 U27728 ( .A(n22354), .B(n22353), .Y(n22355) );
  sky130_fd_sc_hd__o21a_1 U27729 ( .A1(n22980), .A2(n26101), .B1(n22355), .X(
        n22370) );
  sky130_fd_sc_hd__nand2_1 U27730 ( .A(n23234), .B(n26862), .Y(n26108) );
  sky130_fd_sc_hd__nand2_1 U27731 ( .A(n22357), .B(n22356), .Y(n22367) );
  sky130_fd_sc_hd__nor2_1 U27732 ( .A(n22361), .B(n22358), .Y(n22363) );
  sky130_fd_sc_hd__a21oi_1 U27734 ( .A1(n22944), .A2(n22363), .B1(n22362), .Y(
        n22364) );
  sky130_fd_sc_hd__o21ai_1 U27735 ( .A1(n22365), .A2(n22897), .B1(n22364), .Y(
        n22366) );
  sky130_fd_sc_hd__xnor2_1 U27736 ( .A(n22367), .B(n22366), .Y(n22368) );
  sky130_fd_sc_hd__nand2_1 U27737 ( .A(n22368), .B(n26863), .Y(n26107) );
  sky130_fd_sc_hd__nand2_1 U27738 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[22]), .Y(n26106) );
  sky130_fd_sc_hd__nand2_1 U27739 ( .A(n26510), .B(n22950), .Y(n22369) );
  sky130_fd_sc_hd__nand3_1 U27740 ( .A(n22371), .B(n22370), .C(n22369), .Y(
        n28991) );
  sky130_fd_sc_hd__nand2_1 U27741 ( .A(n22957), .B(
        j202_soc_core_j22_cpu_rf_vbr[26]), .Y(n22375) );
  sky130_fd_sc_hd__nand2_1 U27742 ( .A(n22967), .B(
        j202_soc_core_j22_cpu_rf_gbr[26]), .Y(n22374) );
  sky130_fd_sc_hd__nand2_1 U27743 ( .A(n22958), .B(
        j202_soc_core_j22_cpu_rf_gpr[506]), .Y(n22373) );
  sky130_fd_sc_hd__nand2_1 U27744 ( .A(n22959), .B(
        j202_soc_core_j22_cpu_rf_tmp[26]), .Y(n22372) );
  sky130_fd_sc_hd__nand4_1 U27745 ( .A(n22375), .B(n22374), .C(n22373), .D(
        n22372), .Y(n22380) );
  sky130_fd_sc_hd__a22oi_1 U27746 ( .A1(n22968), .A2(
        j202_soc_core_j22_cpu_rf_pr[26]), .B1(j202_soc_core_j22_cpu_pc[26]), 
        .B2(n22966), .Y(n22379) );
  sky130_fd_sc_hd__nand2_1 U27747 ( .A(n22376), .B(n22969), .Y(n22378) );
  sky130_fd_sc_hd__nand2_1 U27748 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[26]), .Y(n22377) );
  sky130_fd_sc_hd__nand4b_1 U27749 ( .A_N(n22380), .B(n22379), .C(n22378), .D(
        n22377), .Y(n22381) );
  sky130_fd_sc_hd__a21oi_1 U27750 ( .A1(n22382), .A2(n22702), .B1(n22381), .Y(
        n22413) );
  sky130_fd_sc_hd__nor2_1 U27751 ( .A(n12135), .B(n22383), .Y(n22387) );
  sky130_fd_sc_hd__nor2_1 U27752 ( .A(n12135), .B(n22384), .Y(n22422) );
  sky130_fd_sc_hd__nor2_1 U27753 ( .A(n22387), .B(n22385), .Y(n22682) );
  sky130_fd_sc_hd__nand2_1 U27754 ( .A(n22385), .B(n22387), .Y(n22681) );
  sky130_fd_sc_hd__nand2_1 U27755 ( .A(n22421), .B(n22681), .Y(n22404) );
  sky130_fd_sc_hd__nor2_1 U27756 ( .A(n12159), .B(n22386), .Y(n22394) );
  sky130_fd_sc_hd__nor2_1 U27757 ( .A(n22394), .B(n22395), .Y(n22887) );
  sky130_fd_sc_hd__nand2_1 U27758 ( .A(n22388), .B(n22553), .Y(n22893) );
  sky130_fd_sc_hd__nand2_1 U27759 ( .A(n22391), .B(n22390), .Y(n22552) );
  sky130_fd_sc_hd__a21oi_1 U27760 ( .A1(n22553), .A2(n22393), .B1(n22392), .Y(
        n22891) );
  sky130_fd_sc_hd__nand2_1 U27761 ( .A(n22395), .B(n22394), .Y(n22888) );
  sky130_fd_sc_hd__o21a_1 U27762 ( .A1(n22887), .A2(n22891), .B1(n22888), .X(
        n22396) );
  sky130_fd_sc_hd__a21oi_1 U27763 ( .A1(n22944), .A2(n22400), .B1(n22399), .Y(
        n22401) );
  sky130_fd_sc_hd__xnor2_1 U27765 ( .A(n22404), .B(n22403), .Y(n22405) );
  sky130_fd_sc_hd__nand2_1 U27766 ( .A(n22405), .B(n26863), .Y(n25082) );
  sky130_fd_sc_hd__nand2_1 U27767 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[26]), .Y(n25081) );
  sky130_fd_sc_hd__a21oi_1 U27768 ( .A1(n22965), .A2(n25085), .B1(n11713), .Y(
        n22406) );
  sky130_fd_sc_hd__nand3_1 U27769 ( .A(n25083), .B(n25082), .C(n13319), .Y(
        n25075) );
  sky130_fd_sc_hd__o22ai_1 U27770 ( .A1(n25824), .A2(n22408), .B1(n22407), 
        .B2(n22952), .Y(n22409) );
  sky130_fd_sc_hd__nand2_1 U27771 ( .A(n25049), .B(n22956), .Y(n22411) );
  sky130_fd_sc_hd__nand3_1 U27772 ( .A(n23262), .B(n11713), .C(n22411), .Y(
        n25056) );
  sky130_fd_sc_hd__nand3_1 U27773 ( .A(n25075), .B(n22929), .C(n25056), .Y(
        n22412) );
  sky130_fd_sc_hd__nand2_1 U27774 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[29]), .Y(n24372) );
  sky130_fd_sc_hd__nand2_1 U27775 ( .A(n22965), .B(n18672), .Y(n22415) );
  sky130_fd_sc_hd__and3_1 U27776 ( .A(n24372), .B(n26398), .C(n22415), .X(
        n24049) );
  sky130_fd_sc_hd__nor2_1 U27777 ( .A(n12135), .B(n22416), .Y(n22420) );
  sky130_fd_sc_hd__nor2_1 U27778 ( .A(n12159), .B(n22417), .Y(n22479) );
  sky130_fd_sc_hd__nand2_1 U27779 ( .A(n22418), .B(n22420), .Y(n22472) );
  sky130_fd_sc_hd__nand2_1 U27780 ( .A(n22474), .B(n22472), .Y(n22435) );
  sky130_fd_sc_hd__nor2_1 U27781 ( .A(n12135), .B(n22419), .Y(n22426) );
  sky130_fd_sc_hd__nor2_1 U27782 ( .A(n22426), .B(n22427), .Y(n22655) );
  sky130_fd_sc_hd__nand2_1 U27783 ( .A(n22421), .B(n22679), .Y(n22659) );
  sky130_fd_sc_hd__nor2_1 U27784 ( .A(n22655), .B(n22659), .Y(n22469) );
  sky130_fd_sc_hd__nor2_1 U27785 ( .A(n22429), .B(n22680), .Y(n22431) );
  sky130_fd_sc_hd__nand2_1 U27786 ( .A(n22423), .B(n22422), .Y(n22678) );
  sky130_fd_sc_hd__a21oi_1 U27787 ( .A1(n22679), .A2(n22425), .B1(n22424), .Y(
        n22658) );
  sky130_fd_sc_hd__nand2_1 U27788 ( .A(n22427), .B(n22426), .Y(n22656) );
  sky130_fd_sc_hd__o21ai_1 U27789 ( .A1(n22655), .A2(n22658), .B1(n22656), .Y(
        n22475) );
  sky130_fd_sc_hd__a21oi_1 U27790 ( .A1(n22944), .A2(n22431), .B1(n22430), .Y(
        n22432) );
  sky130_fd_sc_hd__o21ai_1 U27791 ( .A1(n22433), .A2(n22897), .B1(n22432), .Y(
        n22434) );
  sky130_fd_sc_hd__xnor2_1 U27792 ( .A(n22435), .B(n22434), .Y(n22436) );
  sky130_fd_sc_hd__nand2_1 U27793 ( .A(n22436), .B(n26863), .Y(n24050) );
  sky130_fd_sc_hd__nand3_1 U27794 ( .A(n24051), .B(n24049), .C(n24050), .Y(
        n22440) );
  sky130_fd_sc_hd__nand2_1 U27795 ( .A(n22437), .B(n26872), .Y(n26975) );
  sky130_fd_sc_hd__nand2b_1 U27796 ( .A_N(n22952), .B(
        j202_soc_core_j22_cpu_ml_macl[29]), .Y(n26974) );
  sky130_fd_sc_hd__nand2_1 U27797 ( .A(n25344), .B(n18672), .Y(n26973) );
  sky130_fd_sc_hd__nand3_1 U27798 ( .A(n26974), .B(n11713), .C(n26973), .Y(
        n22438) );
  sky130_fd_sc_hd__a21oi_1 U27799 ( .A1(n26978), .A2(n22956), .B1(n22438), .Y(
        n22439) );
  sky130_fd_sc_hd__nand2_1 U27800 ( .A(n26975), .B(n22439), .Y(n24031) );
  sky130_fd_sc_hd__nand3_1 U27801 ( .A(n22440), .B(n22929), .C(n24031), .Y(
        n22463) );
  sky130_fd_sc_hd__a22oi_1 U27802 ( .A1(n22966), .A2(
        j202_soc_core_j22_cpu_pc[29]), .B1(j202_soc_core_j22_cpu_rf_gbr[29]), 
        .B2(n22967), .Y(n22446) );
  sky130_fd_sc_hd__a2bb2oi_1 U27803 ( .B1(j202_soc_core_j22_cpu_rf_pr[29]), 
        .B2(n22968), .A1_N(n22441), .A2_N(n22877), .Y(n22445) );
  sky130_fd_sc_hd__a2bb2oi_1 U27804 ( .B1(j202_soc_core_j22_cpu_rf_tmp[29]), 
        .B2(n22959), .A1_N(n22442), .A2_N(n22875), .Y(n22444) );
  sky130_fd_sc_hd__nand2_1 U27805 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[29]), .Y(n22443) );
  sky130_fd_sc_hd__nand4_1 U27806 ( .A(n22446), .B(n22445), .C(n22444), .D(
        n22443), .Y(n22447) );
  sky130_fd_sc_hd__a21oi_1 U27807 ( .A1(n22969), .A2(n22448), .B1(n22447), .Y(
        n22449) );
  sky130_fd_sc_hd__o21ai_1 U27808 ( .A1(n22456), .A2(n22450), .B1(n22449), .Y(
        n22454) );
  sky130_fd_sc_hd__nor2_1 U27810 ( .A(n22454), .B(n22453), .Y(n22455) );
  sky130_fd_sc_hd__a21oi_1 U27812 ( .A1(n22768), .A2(n22458), .B1(n22457), .Y(
        n22462) );
  sky130_fd_sc_hd__nand2_1 U27813 ( .A(n22460), .B(n22459), .Y(n22461) );
  sky130_fd_sc_hd__nand3_1 U27814 ( .A(n22463), .B(n22462), .C(n22461), .Y(
        n28998) );
  sky130_fd_sc_hd__nand2_1 U27815 ( .A(n26873), .B(n22927), .Y(n22492) );
  sky130_fd_sc_hd__nor2_1 U27816 ( .A(n11713), .B(n25219), .Y(n24478) );
  sky130_fd_sc_hd__nor2_1 U27817 ( .A(n12159), .B(n22464), .Y(n22466) );
  sky130_fd_sc_hd__nand2_1 U27818 ( .A(n13278), .B(n22466), .Y(n22467) );
  sky130_fd_sc_hd__nand2_1 U27819 ( .A(n22468), .B(n22467), .Y(n22486) );
  sky130_fd_sc_hd__nor2_1 U27820 ( .A(n22479), .B(n13278), .Y(n22615) );
  sky130_fd_sc_hd__nand2_1 U27821 ( .A(n22470), .B(n22477), .Y(n22620) );
  sky130_fd_sc_hd__nor2_1 U27822 ( .A(n22615), .B(n22620), .Y(n22480) );
  sky130_fd_sc_hd__a21o_1 U27823 ( .A1(n22475), .A2(n22474), .B1(n22473), .X(
        n22476) );
  sky130_fd_sc_hd__nand2_1 U27824 ( .A(n13278), .B(n22479), .Y(n22616) );
  sky130_fd_sc_hd__a21oi_1 U27825 ( .A1(n22944), .A2(n22482), .B1(n22481), .Y(
        n22483) );
  sky130_fd_sc_hd__o21ai_1 U27826 ( .A1(n22484), .A2(n22897), .B1(n22483), .Y(
        n22485) );
  sky130_fd_sc_hd__xnor2_1 U27827 ( .A(n22486), .B(n22485), .Y(n26864) );
  sky130_fd_sc_hd__nand2b_1 U27828 ( .A_N(n22952), .B(
        j202_soc_core_j22_cpu_ml_macl[31]), .Y(n26875) );
  sky130_fd_sc_hd__nand2_1 U27829 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[31]), .Y(n26867) );
  sky130_fd_sc_hd__nand2_1 U27830 ( .A(n25344), .B(n22487), .Y(n26874) );
  sky130_fd_sc_hd__a2bb2oi_1 U27831 ( .B1(n22965), .B2(n22487), .A1_N(n26398), 
        .A2_N(n26874), .Y(n22488) );
  sky130_fd_sc_hd__o21a_1 U27832 ( .A1(n11713), .A2(n26867), .B1(n22488), .X(
        n22490) );
  sky130_fd_sc_hd__nand2_1 U27833 ( .A(n26871), .B(n22956), .Y(n22489) );
  sky130_fd_sc_hd__nand2_1 U27834 ( .A(n24997), .B(n22929), .Y(n22506) );
  sky130_fd_sc_hd__a22oi_1 U27835 ( .A1(n22968), .A2(
        j202_soc_core_j22_cpu_rf_pr[31]), .B1(j202_soc_core_j22_cpu_rf_gbr[31]), .B2(n22967), .Y(n22498) );
  sky130_fd_sc_hd__a2bb2oi_1 U27836 ( .B1(j202_soc_core_j22_cpu_pc[31]), .B2(
        n22966), .A1_N(n22493), .A2_N(n22875), .Y(n22497) );
  sky130_fd_sc_hd__a2bb2oi_1 U27837 ( .B1(j202_soc_core_j22_cpu_rf_tmp[31]), 
        .B2(n22959), .A1_N(n22494), .A2_N(n22877), .Y(n22496) );
  sky130_fd_sc_hd__nand2_1 U27838 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[31]), .Y(n22495) );
  sky130_fd_sc_hd__nand4_1 U27839 ( .A(n22498), .B(n22497), .C(n22496), .D(
        n22495), .Y(n22499) );
  sky130_fd_sc_hd__a21oi_1 U27840 ( .A1(n22969), .A2(n22500), .B1(n22499), .Y(
        n22504) );
  sky130_fd_sc_hd__nand2_1 U27841 ( .A(n22501), .B(n22702), .Y(n22502) );
  sky130_fd_sc_hd__nand2_1 U27842 ( .A(n23467), .B(n26255), .Y(n25953) );
  sky130_fd_sc_hd__nor2_1 U27843 ( .A(n28243), .B(n25953), .Y(n27037) );
  sky130_fd_sc_hd__nand2_1 U27844 ( .A(j202_soc_core_qspi_wb_addr[24]), .B(
        j202_soc_core_ahb2wbqspi_00_stb_o), .Y(n23336) );
  sky130_fd_sc_hd__and3_1 U27845 ( .A(n27037), .B(n22508), .C(n29594), .X(
        n28966) );
  sky130_fd_sc_hd__nor2b_1 U27846 ( .B_N(j202_soc_core_qspi_int), .A(n28590), 
        .Y(n29057) );
  sky130_fd_sc_hd__xor2_1 U27847 ( .A(n22509), .B(n19063), .X(n25268) );
  sky130_fd_sc_hd__a22oi_1 U27848 ( .A1(n22510), .A2(n26726), .B1(n22596), 
        .B2(n25268), .Y(n22517) );
  sky130_fd_sc_hd__nand2_1 U27849 ( .A(n22512), .B(n22511), .Y(n22514) );
  sky130_fd_sc_hd__xnor2_1 U27850 ( .A(n22514), .B(n22513), .Y(n24156) );
  sky130_fd_sc_hd__a22oi_1 U27851 ( .A1(n27354), .A2(n22515), .B1(n24156), 
        .B2(n12158), .Y(n22516) );
  sky130_fd_sc_hd__nand3_1 U27852 ( .A(n22518), .B(n22517), .C(n22516), .Y(
        n29031) );
  sky130_fd_sc_hd__nand2_1 U27853 ( .A(n22520), .B(n22519), .Y(n22529) );
  sky130_fd_sc_hd__nor2_1 U27854 ( .A(n22523), .B(n22617), .Y(n22525) );
  sky130_fd_sc_hd__o21ai_1 U27855 ( .A1(n22523), .A2(n22619), .B1(n22522), .Y(
        n22524) );
  sky130_fd_sc_hd__a21oi_1 U27856 ( .A1(n22661), .A2(n22525), .B1(n22524), .Y(
        n22526) );
  sky130_fd_sc_hd__nand2_1 U27857 ( .A(n23231), .B(n24499), .Y(n23975) );
  sky130_fd_sc_hd__nand2_1 U27858 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[16]), .Y(n23977) );
  sky130_fd_sc_hd__nand3_1 U27859 ( .A(n23978), .B(n23975), .C(n23977), .Y(
        n27048) );
  sky130_fd_sc_hd__nand2_1 U27860 ( .A(n27048), .B(n22950), .Y(n22550) );
  sky130_fd_sc_hd__o22ai_1 U27861 ( .A1(n25824), .A2(n22531), .B1(n22530), 
        .B2(n22952), .Y(n22532) );
  sky130_fd_sc_hd__a21oi_1 U27862 ( .A1(n22533), .A2(n26872), .B1(n22532), .Y(
        n24171) );
  sky130_fd_sc_hd__nand2_1 U27863 ( .A(n24602), .B(n22956), .Y(n23994) );
  sky130_fd_sc_hd__nand2_1 U27864 ( .A(n22957), .B(
        j202_soc_core_j22_cpu_rf_vbr[16]), .Y(n22537) );
  sky130_fd_sc_hd__nand2_1 U27865 ( .A(n22958), .B(
        j202_soc_core_j22_cpu_rf_gpr[496]), .Y(n22536) );
  sky130_fd_sc_hd__nand2_1 U27866 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[16]), .Y(n22535) );
  sky130_fd_sc_hd__nand2_1 U27867 ( .A(n22959), .B(
        j202_soc_core_j22_cpu_rf_tmp[16]), .Y(n22534) );
  sky130_fd_sc_hd__nand4_1 U27868 ( .A(n22537), .B(n22536), .C(n22535), .D(
        n22534), .Y(n22543) );
  sky130_fd_sc_hd__a22oi_1 U27869 ( .A1(n22968), .A2(
        j202_soc_core_j22_cpu_rf_pr[16]), .B1(n22967), .B2(
        j202_soc_core_j22_cpu_rf_gbr[16]), .Y(n22541) );
  sky130_fd_sc_hd__nand2_1 U27870 ( .A(n22538), .B(n22969), .Y(n22540) );
  sky130_fd_sc_hd__nand2_1 U27871 ( .A(n22965), .B(n12577), .Y(n23985) );
  sky130_fd_sc_hd__a2bb2oi_1 U27872 ( .B1(j202_soc_core_j22_cpu_pc[16]), .B2(
        n22966), .A1_N(n22978), .A2_N(n23985), .Y(n22539) );
  sky130_fd_sc_hd__nand3_1 U27873 ( .A(n22541), .B(n22540), .C(n22539), .Y(
        n22542) );
  sky130_fd_sc_hd__nor2_1 U27874 ( .A(n22543), .B(n22542), .Y(n22544) );
  sky130_fd_sc_hd__o21a_1 U27875 ( .A1(n22546), .A2(n22545), .B1(n22544), .X(
        n22547) );
  sky130_fd_sc_hd__o21a_1 U27876 ( .A1(n22978), .A2(n23994), .B1(n22547), .X(
        n22548) );
  sky130_fd_sc_hd__o21a_1 U27877 ( .A1(n22980), .A2(n24171), .B1(n22548), .X(
        n22549) );
  sky130_fd_sc_hd__nand3_1 U27878 ( .A(n22551), .B(n22550), .C(n22549), .Y(
        n28984) );
  sky130_fd_sc_hd__nand2_1 U27879 ( .A(n23235), .B(n24499), .Y(n22563) );
  sky130_fd_sc_hd__nand2_1 U27880 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[24]), .Y(n23824) );
  sky130_fd_sc_hd__nand2_1 U27881 ( .A(n22553), .B(n22552), .Y(n22561) );
  sky130_fd_sc_hd__nor2_1 U27882 ( .A(n22555), .B(n22890), .Y(n22557) );
  sky130_fd_sc_hd__o21ai_1 U27883 ( .A1(n22555), .A2(n22892), .B1(n22554), .Y(
        n22556) );
  sky130_fd_sc_hd__a21oi_1 U27884 ( .A1(n22944), .A2(n22557), .B1(n22556), .Y(
        n22558) );
  sky130_fd_sc_hd__o21ai_1 U27885 ( .A1(n22559), .A2(n22897), .B1(n22558), .Y(
        n22560) );
  sky130_fd_sc_hd__xnor2_1 U27886 ( .A(n22561), .B(n22560), .Y(n22562) );
  sky130_fd_sc_hd__nand2_1 U27887 ( .A(n22562), .B(n26863), .Y(n23850) );
  sky130_fd_sc_hd__nand2_1 U27888 ( .A(n25873), .B(n22956), .Y(n23827) );
  sky130_fd_sc_hd__nand2_1 U27889 ( .A(n22957), .B(
        j202_soc_core_j22_cpu_rf_vbr[24]), .Y(n22567) );
  sky130_fd_sc_hd__nand2_1 U27890 ( .A(n22958), .B(
        j202_soc_core_j22_cpu_rf_gpr[504]), .Y(n22566) );
  sky130_fd_sc_hd__nand2_1 U27891 ( .A(n22959), .B(
        j202_soc_core_j22_cpu_rf_tmp[24]), .Y(n22565) );
  sky130_fd_sc_hd__nand2_1 U27892 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[24]), .Y(n22564) );
  sky130_fd_sc_hd__nand4_1 U27893 ( .A(n22567), .B(n22566), .C(n22565), .D(
        n22564), .Y(n22572) );
  sky130_fd_sc_hd__nand2_1 U27894 ( .A(n22965), .B(n24583), .Y(n23823) );
  sky130_fd_sc_hd__a2bb2oi_1 U27895 ( .B1(j202_soc_core_j22_cpu_rf_pr[24]), 
        .B2(n22968), .A1_N(n22978), .A2_N(n23823), .Y(n22571) );
  sky130_fd_sc_hd__a22oi_1 U27896 ( .A1(n22966), .A2(
        j202_soc_core_j22_cpu_pc[24]), .B1(j202_soc_core_j22_cpu_rf_gbr[24]), 
        .B2(n22967), .Y(n22570) );
  sky130_fd_sc_hd__nand2_1 U27897 ( .A(n22568), .B(n22969), .Y(n22569) );
  sky130_fd_sc_hd__nand4b_1 U27898 ( .A_N(n22572), .B(n22571), .C(n22570), .D(
        n22569), .Y(n22573) );
  sky130_fd_sc_hd__a21oi_1 U27899 ( .A1(n22574), .A2(n22702), .B1(n22573), .Y(
        n22577) );
  sky130_fd_sc_hd__nand2_1 U27900 ( .A(n22575), .B(n26872), .Y(n23829) );
  sky130_fd_sc_hd__nand2b_1 U27901 ( .A_N(n22952), .B(
        j202_soc_core_j22_cpu_ml_macl[24]), .Y(n23825) );
  sky130_fd_sc_hd__nand2_1 U27902 ( .A(n25344), .B(n24583), .Y(n23826) );
  sky130_fd_sc_hd__nand3_1 U27903 ( .A(n23829), .B(n23825), .C(n23826), .Y(
        n25874) );
  sky130_fd_sc_hd__nand2_1 U27904 ( .A(n25874), .B(n22654), .Y(n22576) );
  sky130_fd_sc_hd__o211ai_1 U27905 ( .A1(n22978), .A2(n23827), .B1(n22577), 
        .C1(n22576), .Y(n22578) );
  sky130_fd_sc_hd__a21oi_1 U27906 ( .A1(n24582), .A2(n22950), .B1(n22578), .Y(
        n22579) );
  sky130_fd_sc_hd__nand2_1 U27907 ( .A(n22580), .B(n22579), .Y(n28993) );
  sky130_fd_sc_hd__nand2_1 U27908 ( .A(n21914), .B(n22581), .Y(n22599) );
  sky130_fd_sc_hd__nand2_1 U27909 ( .A(n22584), .B(n22583), .Y(n22589) );
  sky130_fd_sc_hd__xnor2_1 U27911 ( .A(n22589), .B(n22588), .Y(n25806) );
  sky130_fd_sc_hd__o22a_1 U27912 ( .A1(n25821), .A2(n11143), .B1(n23832), .B2(
        n22590), .X(n22591) );
  sky130_fd_sc_hd__o21ai_1 U27913 ( .A1(n23832), .A2(n22592), .B1(n22591), .Y(
        n22593) );
  sky130_fd_sc_hd__a21oi_1 U27914 ( .A1(n25806), .A2(n12158), .B1(n22593), .Y(
        n22598) );
  sky130_fd_sc_hd__nand2_1 U27915 ( .A(n22594), .B(j202_soc_core_j22_cpu_pc[7]), .Y(n22595) );
  sky130_fd_sc_hd__xor2_1 U27916 ( .A(n22595), .B(n21994), .X(n25848) );
  sky130_fd_sc_hd__nand2_1 U27917 ( .A(n22596), .B(n25848), .Y(n22597) );
  sky130_fd_sc_hd__nand3_1 U27918 ( .A(n22599), .B(n22598), .C(n22597), .Y(
        n29064) );
  sky130_fd_sc_hd__nand2_1 U27919 ( .A(n22600), .B(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[1]), .Y(n24807) );
  sky130_fd_sc_hd__nor4_1 U27920 ( .A(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[2]), .B(n22601), 
        .C(n24807), .D(n25677), .Y(n29050) );
  sky130_fd_sc_hd__nor2b_1 U27921 ( .B_N(j202_soc_core_bldc_int), .A(n28590), 
        .Y(n29051) );
  sky130_fd_sc_hd__a22oi_1 U27922 ( .A1(n22968), .A2(
        j202_soc_core_j22_cpu_rf_pr[30]), .B1(j202_soc_core_j22_cpu_pc[30]), 
        .B2(n22966), .Y(n22607) );
  sky130_fd_sc_hd__a2bb2oi_1 U27923 ( .B1(j202_soc_core_j22_cpu_rf_gbr[30]), 
        .B2(n22967), .A1_N(n22602), .A2_N(n22877), .Y(n22606) );
  sky130_fd_sc_hd__a2bb2oi_1 U27924 ( .B1(j202_soc_core_j22_cpu_rf_tmp[30]), 
        .B2(n22959), .A1_N(n22603), .A2_N(n22875), .Y(n22605) );
  sky130_fd_sc_hd__nand2_1 U27925 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[30]), .Y(n22604) );
  sky130_fd_sc_hd__nand4_1 U27926 ( .A(n22607), .B(n22606), .C(n22605), .D(
        n22604), .Y(n22608) );
  sky130_fd_sc_hd__nand2_1 U27927 ( .A(n24510), .B(n22927), .Y(n26513) );
  sky130_fd_sc_hd__nand2_1 U27929 ( .A(n11147), .B(n22616), .Y(n22626) );
  sky130_fd_sc_hd__nor2_1 U27930 ( .A(n22620), .B(n22617), .Y(n22622) );
  sky130_fd_sc_hd__nand2_1 U27931 ( .A(n22521), .B(n22622), .Y(n22624) );
  sky130_fd_sc_hd__a21oi_1 U27933 ( .A1(n22944), .A2(n22622), .B1(n22621), .Y(
        n22623) );
  sky130_fd_sc_hd__o21ai_1 U27934 ( .A1(n22624), .A2(n22897), .B1(n22623), .Y(
        n22625) );
  sky130_fd_sc_hd__xnor2_1 U27935 ( .A(n22626), .B(n22625), .Y(n24500) );
  sky130_fd_sc_hd__nand2_1 U27936 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[30]), .Y(n24502) );
  sky130_fd_sc_hd__nand2_1 U27937 ( .A(n25344), .B(n24505), .Y(n24507) );
  sky130_fd_sc_hd__nor2_1 U27938 ( .A(n22628), .B(n22952), .Y(n24508) );
  sky130_fd_sc_hd__nand2_1 U27939 ( .A(n24508), .B(n11713), .Y(n22629) );
  sky130_fd_sc_hd__o211ai_1 U27940 ( .A1(n11713), .A2(n24502), .B1(n22630), 
        .C1(n22629), .Y(n22631) );
  sky130_fd_sc_hd__a21oi_1 U27941 ( .A1(n24511), .A2(n22956), .B1(n22631), .Y(
        n24492) );
  sky130_fd_sc_hd__nand2_1 U27942 ( .A(n26515), .B(n24492), .Y(n22632) );
  sky130_fd_sc_hd__nand2_1 U27943 ( .A(n22929), .B(n22632), .Y(n22633) );
  sky130_fd_sc_hd__o211a_1 U27944 ( .A1(n22978), .A2(n22635), .B1(n22634), 
        .C1(n22633), .X(n22636) );
  sky130_fd_sc_hd__nand2_1 U27945 ( .A(n12498), .B(n22636), .Y(n29000) );
  sky130_fd_sc_hd__nand2_1 U27946 ( .A(n22637), .B(n26872), .Y(n22640) );
  sky130_fd_sc_hd__o22a_1 U27947 ( .A1(n25824), .A2(n17370), .B1(n22638), .B2(
        n22952), .X(n22639) );
  sky130_fd_sc_hd__nand2_1 U27948 ( .A(n22640), .B(n22639), .Y(n24550) );
  sky130_fd_sc_hd__nand2_1 U27949 ( .A(n24551), .B(n22956), .Y(n26401) );
  sky130_fd_sc_hd__nand2_1 U27950 ( .A(n22957), .B(
        j202_soc_core_j22_cpu_rf_vbr[28]), .Y(n22644) );
  sky130_fd_sc_hd__nand2_1 U27951 ( .A(n22958), .B(
        j202_soc_core_j22_cpu_rf_gpr[508]), .Y(n22643) );
  sky130_fd_sc_hd__nand2_1 U27952 ( .A(n22959), .B(
        j202_soc_core_j22_cpu_rf_tmp[28]), .Y(n22642) );
  sky130_fd_sc_hd__nand2_1 U27953 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[28]), .Y(n22641) );
  sky130_fd_sc_hd__nand4_1 U27954 ( .A(n22644), .B(n22643), .C(n22642), .D(
        n22641), .Y(n22649) );
  sky130_fd_sc_hd__a2bb2oi_1 U27955 ( .B1(j202_soc_core_j22_cpu_rf_pr[28]), 
        .B2(n22968), .A1_N(n22978), .A2_N(n26396), .Y(n22648) );
  sky130_fd_sc_hd__a22oi_1 U27956 ( .A1(n22966), .A2(
        j202_soc_core_j22_cpu_pc[28]), .B1(j202_soc_core_j22_cpu_rf_gbr[28]), 
        .B2(n22967), .Y(n22647) );
  sky130_fd_sc_hd__nand2_1 U27957 ( .A(n22645), .B(n22969), .Y(n22646) );
  sky130_fd_sc_hd__nand4b_1 U27958 ( .A_N(n22649), .B(n22648), .C(n22647), .D(
        n22646), .Y(n22650) );
  sky130_fd_sc_hd__a21oi_1 U27959 ( .A1(n22651), .A2(n22702), .B1(n22650), .Y(
        n22652) );
  sky130_fd_sc_hd__o21ai_1 U27960 ( .A1(n22978), .A2(n26401), .B1(n22652), .Y(
        n22653) );
  sky130_fd_sc_hd__a21oi_1 U27961 ( .A1(n24550), .A2(n22654), .B1(n22653), .Y(
        n22666) );
  sky130_fd_sc_hd__nand2_1 U27962 ( .A(n26321), .B(n24499), .Y(n26400) );
  sky130_fd_sc_hd__nand2_1 U27963 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[28]), .Y(n26397) );
  sky130_fd_sc_hd__nand2_1 U27964 ( .A(n22657), .B(n22656), .Y(n22664) );
  sky130_fd_sc_hd__nor2_1 U27965 ( .A(n22659), .B(n22680), .Y(n22660) );
  sky130_fd_sc_hd__nand3_1 U27966 ( .A(n26400), .B(n26397), .C(n26399), .Y(
        n24548) );
  sky130_fd_sc_hd__nand2_1 U27967 ( .A(n24548), .B(n22950), .Y(n22665) );
  sky130_fd_sc_hd__nand3_1 U27968 ( .A(n22667), .B(n22666), .C(n22665), .Y(
        n28997) );
  sky130_fd_sc_hd__nand2_1 U27969 ( .A(j202_soc_core_qspi_wb_wdat[31]), .B(
        n29594), .Y(n27081) );
  sky130_fd_sc_hd__nand2_1 U27970 ( .A(j202_soc_core_qspi_wb_wdat[30]), .B(
        n29594), .Y(n27095) );
  sky130_fd_sc_hd__nand2_1 U27971 ( .A(j202_soc_core_qspi_wb_wdat[29]), .B(
        n29594), .Y(n26959) );
  sky130_fd_sc_hd__nand2_1 U27972 ( .A(j202_soc_core_qspi_wb_wdat[28]), .B(
        n29594), .Y(n26456) );
  sky130_fd_sc_hd__nand2_1 U27973 ( .A(j202_soc_core_qspi_wb_wdat[26]), .B(
        n29594), .Y(n25097) );
  sky130_fd_sc_hd__nand2_1 U27974 ( .A(j202_soc_core_qspi_wb_wdat[24]), .B(
        n29594), .Y(n25858) );
  sky130_fd_sc_hd__nand2_1 U27975 ( .A(j202_soc_core_qspi_wb_wdat[23]), .B(
        n29594), .Y(n27028) );
  sky130_fd_sc_hd__nand2_1 U27976 ( .A(j202_soc_core_qspi_wb_wdat[22]), .B(
        n29594), .Y(n26494) );
  sky130_fd_sc_hd__nand2_1 U27977 ( .A(j202_soc_core_qspi_wb_wdat[20]), .B(
        n29594), .Y(n28604) );
  sky130_fd_sc_hd__nand2_1 U27978 ( .A(j202_soc_core_qspi_wb_wdat[18]), .B(
        n29594), .Y(n28605) );
  sky130_fd_sc_hd__nand2_1 U27979 ( .A(j202_soc_core_qspi_wb_wdat[12]), .B(
        n29594), .Y(n28608) );
  sky130_fd_sc_hd__nand2_1 U27980 ( .A(j202_soc_core_qspi_wb_wdat[8]), .B(
        n29594), .Y(n28599) );
  sky130_fd_sc_hd__nand2_1 U27981 ( .A(j202_soc_core_qspi_wb_wdat[7]), .B(
        n29594), .Y(n28610) );
  sky130_fd_sc_hd__nand2_1 U27982 ( .A(j202_soc_core_qspi_wb_wdat[6]), .B(
        n29594), .Y(n28611) );
  sky130_fd_sc_hd__nand2_1 U27983 ( .A(j202_soc_core_qspi_wb_wdat[5]), .B(
        n29594), .Y(n28612) );
  sky130_fd_sc_hd__nand2_1 U27984 ( .A(j202_soc_core_qspi_wb_wdat[4]), .B(
        n29594), .Y(n28613) );
  sky130_fd_sc_hd__nand2_1 U27985 ( .A(j202_soc_core_qspi_wb_wdat[0]), .B(
        n29594), .Y(n28881) );
  sky130_fd_sc_hd__nor2_1 U27986 ( .A(n28946), .B(n29031), .Y(n22670) );
  sky130_fd_sc_hd__inv_2 U27987 ( .A(n28947), .Y(n22676) );
  sky130_fd_sc_hd__nand2_1 U27988 ( .A(n22676), .B(n28948), .Y(n22710) );
  sky130_fd_sc_hd__nand2_1 U27989 ( .A(n22674), .B(n22673), .Y(n22675) );
  sky130_fd_sc_hd__nand2_1 U27990 ( .A(n28947), .B(n28948), .Y(n22995) );
  sky130_fd_sc_hd__nor2_1 U27991 ( .A(n22995), .B(n22677), .Y(n29024) );
  sky130_fd_sc_hd__nor2_1 U27992 ( .A(n22710), .B(n22677), .Y(n29025) );
  sky130_fd_sc_hd__nor2_1 U27993 ( .A(n12162), .B(n22677), .Y(n29026) );
  sky130_fd_sc_hd__nand2_1 U27994 ( .A(n22679), .B(n22678), .Y(n22684) );
  sky130_fd_sc_hd__nor2_1 U27995 ( .A(n22682), .B(n22680), .Y(n22683) );
  sky130_fd_sc_hd__a21oi_1 U27996 ( .A1(n22965), .A2(n22685), .B1(n11713), .Y(
        n22686) );
  sky130_fd_sc_hd__nand2_1 U27997 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[27]), .Y(n25142) );
  sky130_fd_sc_hd__nand2_1 U27998 ( .A(n23248), .B(n24499), .Y(n25144) );
  sky130_fd_sc_hd__nand2_1 U27999 ( .A(n22687), .B(n25144), .Y(n22691) );
  sky130_fd_sc_hd__nand2_1 U28000 ( .A(n22688), .B(n26872), .Y(n23007) );
  sky130_fd_sc_hd__nand2b_1 U28001 ( .A_N(n22952), .B(
        j202_soc_core_j22_cpu_ml_macl[27]), .Y(n23003) );
  sky130_fd_sc_hd__nand2_1 U28002 ( .A(n25344), .B(n22685), .Y(n23004) );
  sky130_fd_sc_hd__nand3_1 U28003 ( .A(n23007), .B(n23003), .C(n23004), .Y(
        n25148) );
  sky130_fd_sc_hd__nand2_1 U28004 ( .A(n25147), .B(n22956), .Y(n23005) );
  sky130_fd_sc_hd__a31oi_1 U28005 ( .A1(n22689), .A2(n11713), .A3(n23005), 
        .B1(n22978), .Y(n22690) );
  sky130_fd_sc_hd__nand2_1 U28006 ( .A(n22691), .B(n22690), .Y(n22706) );
  sky130_fd_sc_hd__nand2_1 U28007 ( .A(n22957), .B(
        j202_soc_core_j22_cpu_rf_vbr[27]), .Y(n22695) );
  sky130_fd_sc_hd__nand2_1 U28008 ( .A(n22967), .B(
        j202_soc_core_j22_cpu_rf_gbr[27]), .Y(n22694) );
  sky130_fd_sc_hd__nand2_1 U28009 ( .A(n22958), .B(
        j202_soc_core_j22_cpu_rf_gpr[507]), .Y(n22693) );
  sky130_fd_sc_hd__nand2_1 U28010 ( .A(n22959), .B(
        j202_soc_core_j22_cpu_rf_tmp[27]), .Y(n22692) );
  sky130_fd_sc_hd__nand4_1 U28011 ( .A(n22695), .B(n22694), .C(n22693), .D(
        n22692), .Y(n22700) );
  sky130_fd_sc_hd__a22oi_1 U28012 ( .A1(n22968), .A2(
        j202_soc_core_j22_cpu_rf_pr[27]), .B1(j202_soc_core_j22_cpu_pc[27]), 
        .B2(n22966), .Y(n22699) );
  sky130_fd_sc_hd__nand2_1 U28013 ( .A(n22696), .B(n22969), .Y(n22698) );
  sky130_fd_sc_hd__nand2_1 U28014 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[27]), .Y(n22697) );
  sky130_fd_sc_hd__nand4b_1 U28015 ( .A_N(n22700), .B(n22699), .C(n22698), .D(
        n22697), .Y(n22701) );
  sky130_fd_sc_hd__a21oi_1 U28016 ( .A1(n22703), .A2(n22702), .B1(n22701), .Y(
        n22705) );
  sky130_fd_sc_hd__nor2b_1 U28017 ( .B_N(
        j202_soc_core_intc_core_00_rg_sint[15]), .A(n28590), .Y(n29046) );
  sky130_fd_sc_hd__nor2b_1 U28018 ( .B_N(
        j202_soc_core_intc_core_00_rg_sint[14]), .A(n28590), .Y(n29047) );
  sky130_fd_sc_hd__nor2b_1 U28019 ( .B_N(
        j202_soc_core_intc_core_00_rg_sint[13]), .A(n28590), .Y(n29049) );
  sky130_fd_sc_hd__nor2b_1 U28020 ( .B_N(
        j202_soc_core_intc_core_00_rg_sint[12]), .A(n28590), .Y(n29048) );
  sky130_fd_sc_hd__nor2b_1 U28021 ( .B_N(
        j202_soc_core_intc_core_00_rg_sint[11]), .A(n28590), .Y(n29060) );
  sky130_fd_sc_hd__nor2b_1 U28022 ( .B_N(
        j202_soc_core_intc_core_00_rg_sint[10]), .A(n28590), .Y(n29043) );
  sky130_fd_sc_hd__nor2b_1 U28023 ( .B_N(j202_soc_core_intc_core_00_rg_sint[9]), .A(n28590), .Y(n29044) );
  sky130_fd_sc_hd__nor2b_1 U28024 ( .B_N(j202_soc_core_intc_core_00_rg_sint[8]), .A(n28590), .Y(n29045) );
  sky130_fd_sc_hd__nor2b_1 U28025 ( .B_N(j202_soc_core_intc_core_00_rg_sint[7]), .A(n28590), .Y(n29042) );
  sky130_fd_sc_hd__nor2b_1 U28026 ( .B_N(j202_soc_core_intc_core_00_rg_sint[6]), .A(n28590), .Y(n29041) );
  sky130_fd_sc_hd__nor2b_1 U28027 ( .B_N(j202_soc_core_intc_core_00_rg_sint[5]), .A(n28590), .Y(n29039) );
  sky130_fd_sc_hd__nor2b_1 U28028 ( .B_N(j202_soc_core_intc_core_00_rg_sint[4]), .A(n28590), .Y(n29040) );
  sky130_fd_sc_hd__nor2b_1 U28029 ( .B_N(j202_soc_core_intc_core_00_rg_sint[3]), .A(n28590), .Y(n29037) );
  sky130_fd_sc_hd__nor2b_1 U28030 ( .B_N(j202_soc_core_intc_core_00_rg_sint[2]), .A(n28590), .Y(n29068) );
  sky130_fd_sc_hd__nor2b_1 U28031 ( .B_N(j202_soc_core_intc_core_00_rg_sint[1]), .A(n28590), .Y(n29052) );
  sky130_fd_sc_hd__nor2b_1 U28032 ( .B_N(j202_soc_core_intc_core_00_rg_sint[0]), .A(n28590), .Y(n29038) );
  sky130_fd_sc_hd__nand3_1 U28033 ( .A(n24118), .B(n29030), .C(n29062), .Y(
        n22707) );
  sky130_fd_sc_hd__nor2_1 U28034 ( .A(n22995), .B(n22707), .Y(n29074) );
  sky130_fd_sc_hd__nor2_1 U28035 ( .A(n12162), .B(n22707), .Y(n29019) );
  sky130_fd_sc_hd__nor2_1 U28036 ( .A(n22710), .B(n22707), .Y(n29020) );
  sky130_fd_sc_hd__nor2_1 U28037 ( .A(n22711), .B(n22707), .Y(n29078) );
  sky130_fd_sc_hd__nor2_1 U28038 ( .A(n22995), .B(n22708), .Y(n29023) );
  sky130_fd_sc_hd__nor2_1 U28039 ( .A(n12162), .B(n22708), .Y(n29016) );
  sky130_fd_sc_hd__nor2_1 U28040 ( .A(n22710), .B(n22708), .Y(n29073) );
  sky130_fd_sc_hd__nand2_1 U28041 ( .A(n22709), .B(n29030), .Y(n22994) );
  sky130_fd_sc_hd__nor2_1 U28042 ( .A(n12162), .B(n22994), .Y(n29017) );
  sky130_fd_sc_hd__nor2_1 U28043 ( .A(n22710), .B(n22994), .Y(n29022) );
  sky130_fd_sc_hd__nor2_1 U28044 ( .A(n22711), .B(n22994), .Y(n29021) );
  sky130_fd_sc_hd__nand2_1 U28045 ( .A(n13301), .B(n22719), .Y(n22720) );
  sky130_fd_sc_hd__xnor2_1 U28046 ( .A(n22721), .B(n22720), .Y(n24164) );
  sky130_fd_sc_hd__nand2_1 U28047 ( .A(n24164), .B(n22927), .Y(n22776) );
  sky130_fd_sc_hd__mux2i_1 U28048 ( .A0(n22722), .A1(n26423), .S(n24612), .Y(
        n22741) );
  sky130_fd_sc_hd__nand2_1 U28049 ( .A(n25131), .B(n22723), .Y(n22728) );
  sky130_fd_sc_hd__nand2_1 U28050 ( .A(n26338), .B(n27389), .Y(n22727) );
  sky130_fd_sc_hd__nand2_1 U28051 ( .A(n25743), .B(n24612), .Y(n26633) );
  sky130_fd_sc_hd__nand2_1 U28052 ( .A(n27443), .B(n26603), .Y(n26632) );
  sky130_fd_sc_hd__nand3_1 U28053 ( .A(n26633), .B(n26326), .C(n26632), .Y(
        n22726) );
  sky130_fd_sc_hd__nor2_1 U28054 ( .A(n22724), .B(n22925), .Y(n22774) );
  sky130_fd_sc_hd__nand2_1 U28055 ( .A(n22774), .B(n26329), .Y(n22725) );
  sky130_fd_sc_hd__nand4_1 U28056 ( .A(n22728), .B(n22727), .C(n22726), .D(
        n22725), .Y(n22740) );
  sky130_fd_sc_hd__nand2_1 U28057 ( .A(n26342), .B(n24613), .Y(n22738) );
  sky130_fd_sc_hd__a2bb2oi_1 U28058 ( .B1(n26077), .B2(n26721), .A1_N(n25128), 
        .A2_N(n22729), .Y(n22737) );
  sky130_fd_sc_hd__nand2_1 U28059 ( .A(n22923), .B(n22730), .Y(n22771) );
  sky130_fd_sc_hd__o21a_1 U28060 ( .A1(n26432), .A2(n26632), .B1(n22732), .X(
        n22733) );
  sky130_fd_sc_hd__o21a_1 U28061 ( .A1(n25229), .A2(n26424), .B1(n22733), .X(
        n22736) );
  sky130_fd_sc_hd__nand2_1 U28062 ( .A(n22734), .B(n26723), .Y(n22735) );
  sky130_fd_sc_hd__nand4_1 U28063 ( .A(n22738), .B(n22737), .C(n22736), .D(
        n22735), .Y(n22739) );
  sky130_fd_sc_hd__nor3_1 U28064 ( .A(n22741), .B(n22740), .C(n22739), .Y(
        n22742) );
  sky130_fd_sc_hd__o21ai_1 U28065 ( .A1(n18916), .A2(n22776), .B1(n22742), .Y(
        n22743) );
  sky130_fd_sc_hd__a21oi_1 U28066 ( .A1(n23781), .A2(n26409), .B1(n22743), .Y(
        n22746) );
  sky130_fd_sc_hd__o21ai_1 U28067 ( .A1(n24792), .A2(n26603), .B1(n25159), .Y(
        n22744) );
  sky130_fd_sc_hd__nand2_1 U28068 ( .A(n27442), .B(n22744), .Y(n22745) );
  sky130_fd_sc_hd__nand2_1 U28069 ( .A(n22749), .B(n22748), .Y(n22758) );
  sky130_fd_sc_hd__nand2_1 U28070 ( .A(n22750), .B(n22753), .Y(n22756) );
  sky130_fd_sc_hd__a21oi_1 U28071 ( .A1(n22754), .A2(n22753), .B1(n22752), .Y(
        n22755) );
  sky130_fd_sc_hd__o21ai_2 U28072 ( .A1(n22756), .A2(n22912), .B1(n22755), .Y(
        n22757) );
  sky130_fd_sc_hd__xnor2_2 U28073 ( .A(n22758), .B(n22757), .Y(n23232) );
  sky130_fd_sc_hd__nand2_1 U28075 ( .A(n22761), .B(n22760), .Y(n22765) );
  sky130_fd_sc_hd__o21ai_0 U28076 ( .A1(n22763), .A2(n21961), .B1(n22762), .Y(
        n22764) );
  sky130_fd_sc_hd__xnor2_1 U28077 ( .A(n22765), .B(n22764), .Y(n22809) );
  sky130_fd_sc_hd__nand2_1 U28078 ( .A(n22809), .B(n24499), .Y(n22769) );
  sky130_fd_sc_hd__a22oi_1 U28079 ( .A1(n22730), .A2(n27187), .B1(n22936), 
        .B2(j202_soc_core_j22_cpu_ml_mach[1]), .Y(n22770) );
  sky130_fd_sc_hd__nand4_1 U28080 ( .A(n24700), .B(n22770), .C(n22771), .D(
        n22769), .Y(n22773) );
  sky130_fd_sc_hd__nand2_1 U28081 ( .A(n22771), .B(n11713), .Y(n22772) );
  sky130_fd_sc_hd__nand2_1 U28082 ( .A(n22773), .B(n22772), .Y(n22777) );
  sky130_fd_sc_hd__nand3_1 U28083 ( .A(n22777), .B(n22776), .C(n22775), .Y(
        n22778) );
  sky130_fd_sc_hd__nand2_1 U28084 ( .A(n22778), .B(n22929), .Y(n22793) );
  sky130_fd_sc_hd__nand2_1 U28085 ( .A(n22779), .B(n22873), .Y(n22791) );
  sky130_fd_sc_hd__o22ai_1 U28086 ( .A1(n24273), .A2(n22856), .B1(n22780), 
        .B2(n22854), .Y(n22784) );
  sky130_fd_sc_hd__o22ai_1 U28087 ( .A1(n22782), .A2(n22860), .B1(n22781), 
        .B2(n22858), .Y(n22783) );
  sky130_fd_sc_hd__nor2_1 U28088 ( .A(n22784), .B(n22783), .Y(n22790) );
  sky130_fd_sc_hd__nand2_1 U28089 ( .A(n22864), .B(
        j202_soc_core_j22_cpu_rf_vbr[1]), .Y(n22788) );
  sky130_fd_sc_hd__nand2_1 U28090 ( .A(n22867), .B(
        j202_soc_core_j22_cpu_rf_tmp[1]), .Y(n22787) );
  sky130_fd_sc_hd__nand2_1 U28091 ( .A(n22865), .B(
        j202_soc_core_j22_cpu_rf_gpr[481]), .Y(n22786) );
  sky130_fd_sc_hd__nand2_1 U28092 ( .A(n22866), .B(
        j202_soc_core_j22_cpu_rf_gpr[1]), .Y(n22785) );
  sky130_fd_sc_hd__and4_1 U28093 ( .A(n22788), .B(n22787), .C(n22786), .D(
        n22785), .X(n22789) );
  sky130_fd_sc_hd__nand3_1 U28094 ( .A(n22791), .B(n22790), .C(n22789), .Y(
        n22825) );
  sky130_fd_sc_hd__nand2_1 U28095 ( .A(n22825), .B(n11158), .Y(n22792) );
  sky130_fd_sc_hd__nand3_1 U28096 ( .A(n22827), .B(n22793), .C(n22792), .Y(
        n28988) );
  sky130_fd_sc_hd__nand2_1 U28097 ( .A(j202_soc_core_qspi_wb_wdat[1]), .B(
        n29594), .Y(n28603) );
  sky130_fd_sc_hd__nand2_1 U28098 ( .A(n23232), .B(n24499), .Y(n25710) );
  sky130_fd_sc_hd__nand2_1 U28099 ( .A(n22796), .B(n22795), .Y(n22804) );
  sky130_fd_sc_hd__xnor2_1 U28100 ( .A(n22804), .B(n22803), .Y(n22805) );
  sky130_fd_sc_hd__nand2_1 U28101 ( .A(n22805), .B(n26863), .Y(n25709) );
  sky130_fd_sc_hd__nand2_1 U28102 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[17]), .Y(n25708) );
  sky130_fd_sc_hd__nand2_1 U28103 ( .A(n24634), .B(n22950), .Y(n22823) );
  sky130_fd_sc_hd__o22ai_1 U28104 ( .A1(n25824), .A2(n22807), .B1(n22806), 
        .B2(n22952), .Y(n22808) );
  sky130_fd_sc_hd__a21oi_1 U28105 ( .A1(n22809), .A2(n26872), .B1(n22808), .Y(
        n24628) );
  sky130_fd_sc_hd__nand2_1 U28106 ( .A(n24164), .B(n22956), .Y(n24624) );
  sky130_fd_sc_hd__nand2_1 U28107 ( .A(n22957), .B(
        j202_soc_core_j22_cpu_rf_vbr[17]), .Y(n22813) );
  sky130_fd_sc_hd__nand2_1 U28108 ( .A(n22958), .B(
        j202_soc_core_j22_cpu_rf_gpr[497]), .Y(n22812) );
  sky130_fd_sc_hd__nand2_1 U28109 ( .A(n22959), .B(
        j202_soc_core_j22_cpu_rf_tmp[17]), .Y(n22811) );
  sky130_fd_sc_hd__nand2_1 U28110 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[17]), .Y(n22810) );
  sky130_fd_sc_hd__nand4_1 U28111 ( .A(n22813), .B(n22812), .C(n22811), .D(
        n22810), .Y(n22818) );
  sky130_fd_sc_hd__nand2_1 U28112 ( .A(n22965), .B(n18300), .Y(n24614) );
  sky130_fd_sc_hd__a2bb2oi_1 U28113 ( .B1(j202_soc_core_j22_cpu_rf_pr[17]), 
        .B2(n22968), .A1_N(n22978), .A2_N(n24614), .Y(n22817) );
  sky130_fd_sc_hd__a22oi_1 U28114 ( .A1(n22966), .A2(
        j202_soc_core_j22_cpu_pc[17]), .B1(j202_soc_core_j22_cpu_rf_gbr[17]), 
        .B2(n22967), .Y(n22816) );
  sky130_fd_sc_hd__nand2_1 U28115 ( .A(n22814), .B(n22969), .Y(n22815) );
  sky130_fd_sc_hd__nand4b_1 U28116 ( .A_N(n22818), .B(n22817), .C(n22816), .D(
        n22815), .Y(n22819) );
  sky130_fd_sc_hd__a21oi_1 U28117 ( .A1(n22825), .A2(n23574), .B1(n22819), .Y(
        n22820) );
  sky130_fd_sc_hd__o21ba_2 U28119 ( .A1(n22980), .A2(n24628), .B1_N(n22821), 
        .X(n22822) );
  sky130_fd_sc_hd__nand3_1 U28120 ( .A(n22827), .B(n22823), .C(n22822), .Y(
        n28985) );
  sky130_fd_sc_hd__nand2_1 U28121 ( .A(j202_soc_core_qspi_wb_wdat[17]), .B(
        n29594), .Y(n28602) );
  sky130_fd_sc_hd__nand2_1 U28123 ( .A(n22830), .B(n22829), .Y(n22840) );
  sky130_fd_sc_hd__nand2_1 U28124 ( .A(n22831), .B(n22834), .Y(n22838) );
  sky130_fd_sc_hd__a21oi_1 U28125 ( .A1(n12579), .A2(n22834), .B1(n22833), .Y(
        n22836) );
  sky130_fd_sc_hd__o21ai_1 U28126 ( .A1(n22838), .A2(n22837), .B1(n22836), .Y(
        n22839) );
  sky130_fd_sc_hd__xnor2_1 U28127 ( .A(n22840), .B(n22839), .Y(n22918) );
  sky130_fd_sc_hd__o22ai_1 U28128 ( .A1(n25824), .A2(n18057), .B1(n22841), 
        .B2(n22952), .Y(n22842) );
  sky130_fd_sc_hd__a21oi_1 U28129 ( .A1(n22918), .A2(n26872), .B1(n22842), .Y(
        n23260) );
  sky130_fd_sc_hd__nand2_1 U28130 ( .A(n12364), .B(n22844), .Y(n22849) );
  sky130_fd_sc_hd__xnor2_1 U28132 ( .A(n22849), .B(n22848), .Y(n24013) );
  sky130_fd_sc_hd__nand2_1 U28133 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[25]), .Y(n25216) );
  sky130_fd_sc_hd__o22ai_1 U28134 ( .A1(n18057), .A2(n22850), .B1(n11713), 
        .B2(n25216), .Y(n22851) );
  sky130_fd_sc_hd__a21oi_1 U28135 ( .A1(n24013), .A2(n22956), .B1(n22851), .Y(
        n22852) );
  sky130_fd_sc_hd__nand2_1 U28136 ( .A(n22853), .B(n22852), .Y(n25118) );
  sky130_fd_sc_hd__o22ai_1 U28137 ( .A1(n22857), .A2(n22856), .B1(n22855), 
        .B2(n22854), .Y(n22863) );
  sky130_fd_sc_hd__o22ai_1 U28138 ( .A1(n22861), .A2(n22860), .B1(n22859), 
        .B2(n22858), .Y(n22862) );
  sky130_fd_sc_hd__nor2_1 U28139 ( .A(n22863), .B(n22862), .Y(n22871) );
  sky130_fd_sc_hd__a22oi_1 U28140 ( .A1(n22865), .A2(
        j202_soc_core_j22_cpu_rf_gpr[489]), .B1(n22864), .B2(
        j202_soc_core_j22_cpu_rf_vbr[9]), .Y(n22870) );
  sky130_fd_sc_hd__nand2_1 U28141 ( .A(n22866), .B(
        j202_soc_core_j22_cpu_rf_gpr[9]), .Y(n22869) );
  sky130_fd_sc_hd__nand2_1 U28142 ( .A(n22867), .B(
        j202_soc_core_j22_cpu_rf_tmp[9]), .Y(n22868) );
  sky130_fd_sc_hd__nand4_1 U28143 ( .A(n22871), .B(n22870), .C(n22869), .D(
        n22868), .Y(n22872) );
  sky130_fd_sc_hd__a21oi_1 U28144 ( .A1(n22874), .A2(n22873), .B1(n22872), .Y(
        n22931) );
  sky130_fd_sc_hd__a22oi_1 U28145 ( .A1(n22966), .A2(
        j202_soc_core_j22_cpu_pc[25]), .B1(j202_soc_core_j22_cpu_rf_gbr[25]), 
        .B2(n22967), .Y(n22882) );
  sky130_fd_sc_hd__a2bb2oi_1 U28146 ( .B1(j202_soc_core_j22_cpu_rf_pr[25]), 
        .B2(n22968), .A1_N(n22876), .A2_N(n22875), .Y(n22881) );
  sky130_fd_sc_hd__a2bb2oi_1 U28147 ( .B1(j202_soc_core_j22_cpu_rf_tmp[25]), 
        .B2(n22959), .A1_N(n22878), .A2_N(n22877), .Y(n22880) );
  sky130_fd_sc_hd__nand2_1 U28148 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[25]), .Y(n22879) );
  sky130_fd_sc_hd__nand4_1 U28149 ( .A(n22882), .B(n22881), .C(n22880), .D(
        n22879), .Y(n22883) );
  sky130_fd_sc_hd__a21oi_1 U28150 ( .A1(n22969), .A2(n22884), .B1(n22883), .Y(
        n22885) );
  sky130_fd_sc_hd__o21ai_1 U28151 ( .A1(n23296), .A2(n22931), .B1(n22885), .Y(
        n22886) );
  sky130_fd_sc_hd__a21oi_1 U28152 ( .A1(n25118), .A2(n22929), .B1(n22886), .Y(
        n22917) );
  sky130_fd_sc_hd__nand2_1 U28153 ( .A(n22889), .B(n22888), .Y(n22900) );
  sky130_fd_sc_hd__nor2_1 U28154 ( .A(n22893), .B(n22890), .Y(n22895) );
  sky130_fd_sc_hd__nand2_1 U28155 ( .A(n12321), .B(n22895), .Y(n22898) );
  sky130_fd_sc_hd__a21oi_1 U28157 ( .A1(n22944), .A2(n22895), .B1(n22894), .Y(
        n22896) );
  sky130_fd_sc_hd__o21ai_1 U28158 ( .A1(n22898), .A2(n22897), .B1(n22896), .Y(
        n22899) );
  sky130_fd_sc_hd__xnor2_1 U28159 ( .A(n22900), .B(n22899), .Y(n22901) );
  sky130_fd_sc_hd__nand2_1 U28160 ( .A(n22904), .B(n22903), .Y(n22915) );
  sky130_fd_sc_hd__nor2_1 U28161 ( .A(n22908), .B(n22905), .Y(n22910) );
  sky130_fd_sc_hd__nand2_1 U28162 ( .A(n22521), .B(n22910), .Y(n22913) );
  sky130_fd_sc_hd__o21ai_1 U28163 ( .A1(n22908), .A2(n22907), .B1(n22906), .Y(
        n22909) );
  sky130_fd_sc_hd__o21ai_2 U28164 ( .A1(n22913), .A2(n22897), .B1(n22911), .Y(
        n22914) );
  sky130_fd_sc_hd__xnor2_2 U28165 ( .A(n22915), .B(n22914), .Y(n23236) );
  sky130_fd_sc_hd__nand2_1 U28166 ( .A(n25117), .B(n22929), .Y(n22916) );
  sky130_fd_sc_hd__nand2_1 U28167 ( .A(n22918), .B(n24499), .Y(n22921) );
  sky130_fd_sc_hd__a22oi_1 U28168 ( .A1(n22919), .A2(n27187), .B1(n22936), 
        .B2(j202_soc_core_j22_cpu_ml_mach[9]), .Y(n22920) );
  sky130_fd_sc_hd__nand2_1 U28169 ( .A(n22921), .B(n22920), .Y(n24692) );
  sky130_fd_sc_hd__a31oi_1 U28170 ( .A1(n22921), .A2(n26318), .A3(n22920), 
        .B1(n11713), .Y(n22922) );
  sky130_fd_sc_hd__nand2_1 U28172 ( .A(n22923), .B(n22919), .Y(n22924) );
  sky130_fd_sc_hd__o21a_1 U28173 ( .A1(n22926), .A2(n22925), .B1(n22924), .X(
        n24717) );
  sky130_fd_sc_hd__nand2_1 U28174 ( .A(n24013), .B(n22927), .Y(n24732) );
  sky130_fd_sc_hd__nand3_1 U28175 ( .A(n22928), .B(n24717), .C(n24732), .Y(
        n22930) );
  sky130_fd_sc_hd__nand2_1 U28176 ( .A(n22930), .B(n22929), .Y(n22934) );
  sky130_fd_sc_hd__or2_0 U28177 ( .A(n22932), .B(n22931), .X(n22933) );
  sky130_fd_sc_hd__nand2_1 U28178 ( .A(j202_soc_core_qspi_wb_wdat[9]), .B(
        n29594), .Y(n28601) );
  sky130_fd_sc_hd__nand2_1 U28179 ( .A(j202_soc_core_qspi_wb_wdat[3]), .B(
        n29594), .Y(n28614) );
  sky130_fd_sc_hd__nand2_1 U28180 ( .A(n22936), .B(
        j202_soc_core_j22_cpu_ml_mach[19]), .Y(n25664) );
  sky130_fd_sc_hd__nand2_1 U28181 ( .A(n22939), .B(n22938), .Y(n22948) );
  sky130_fd_sc_hd__xnor2_1 U28182 ( .A(n22948), .B(n22947), .Y(n22949) );
  sky130_fd_sc_hd__nand2_1 U28183 ( .A(n25703), .B(n22950), .Y(n22982) );
  sky130_fd_sc_hd__o22ai_1 U28184 ( .A1(n25824), .A2(n17417), .B1(n22953), 
        .B2(n22952), .Y(n22954) );
  sky130_fd_sc_hd__a21oi_1 U28185 ( .A1(n22955), .A2(n26872), .B1(n22954), .Y(
        n24066) );
  sky130_fd_sc_hd__nand2_1 U28186 ( .A(n24128), .B(n22956), .Y(n24083) );
  sky130_fd_sc_hd__nand2_1 U28187 ( .A(n22957), .B(
        j202_soc_core_j22_cpu_rf_vbr[19]), .Y(n22964) );
  sky130_fd_sc_hd__nand2_1 U28188 ( .A(n22958), .B(
        j202_soc_core_j22_cpu_rf_gpr[499]), .Y(n22963) );
  sky130_fd_sc_hd__nand2_1 U28189 ( .A(n22959), .B(
        j202_soc_core_j22_cpu_rf_tmp[19]), .Y(n22962) );
  sky130_fd_sc_hd__nand2_1 U28190 ( .A(n22960), .B(
        j202_soc_core_j22_cpu_rf_gpr[19]), .Y(n22961) );
  sky130_fd_sc_hd__nand4_1 U28191 ( .A(n22964), .B(n22963), .C(n22962), .D(
        n22961), .Y(n22974) );
  sky130_fd_sc_hd__nand2_1 U28192 ( .A(n22965), .B(n22951), .Y(n24073) );
  sky130_fd_sc_hd__a2bb2oi_1 U28193 ( .B1(j202_soc_core_j22_cpu_pc[19]), .B2(
        n22966), .A1_N(n22978), .A2_N(n24073), .Y(n22973) );
  sky130_fd_sc_hd__a22oi_1 U28194 ( .A1(n22968), .A2(
        j202_soc_core_j22_cpu_rf_pr[19]), .B1(j202_soc_core_j22_cpu_rf_gbr[19]), .B2(n22967), .Y(n22972) );
  sky130_fd_sc_hd__nand2_1 U28195 ( .A(n22970), .B(n22969), .Y(n22971) );
  sky130_fd_sc_hd__nand4b_1 U28196 ( .A_N(n22974), .B(n22973), .C(n22972), .D(
        n22971), .Y(n22975) );
  sky130_fd_sc_hd__a21oi_1 U28197 ( .A1(n22976), .A2(n23574), .B1(n22975), .Y(
        n22977) );
  sky130_fd_sc_hd__o21ai_1 U28198 ( .A1(n22978), .A2(n24083), .B1(n22977), .Y(
        n22979) );
  sky130_fd_sc_hd__nand3_1 U28199 ( .A(n22983), .B(n22982), .C(n22981), .Y(
        n28987) );
  sky130_fd_sc_hd__nand2_1 U28200 ( .A(j202_soc_core_qspi_wb_wdat[19]), .B(
        n29594), .Y(n28600) );
  sky130_fd_sc_hd__nand2_1 U28201 ( .A(j202_soc_core_qspi_wb_wdat[13]), .B(
        n29594), .Y(n28598) );
  sky130_fd_sc_hd__nand2_1 U28202 ( .A(n29081), .B(n12142), .Y(n28009) );
  sky130_fd_sc_hd__nor2_1 U28203 ( .A(j202_soc_core_uart_BRG_cnt[0]), .B(
        n28009), .Y(n29082) );
  sky130_fd_sc_hd__nor2_1 U28204 ( .A(j202_soc_core_uart_BRG_cnt[1]), .B(
        j202_soc_core_uart_BRG_cnt[0]), .Y(n29090) );
  sky130_fd_sc_hd__nand2_1 U28205 ( .A(j202_soc_core_uart_sio_ce), .B(
        j202_soc_core_uart_TOP_shift_en), .Y(n24228) );
  sky130_fd_sc_hd__nor2_1 U28206 ( .A(n28590), .B(n24228), .Y(n29080) );
  sky130_fd_sc_hd__nand2_1 U28207 ( .A(j202_soc_core_qspi_wb_wdat[14]), .B(
        n29594), .Y(n28597) );
  sky130_fd_sc_hd__nand2_1 U28208 ( .A(j202_soc_core_qspi_wb_wdat[11]), .B(
        n29594), .Y(n28596) );
  sky130_fd_sc_hd__nor4_1 U28209 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[21]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[22]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[25]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[23]), .Y(n22987) );
  sky130_fd_sc_hd__nor4_1 U28210 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[26]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[27]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[29]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[30]), .Y(n22986) );
  sky130_fd_sc_hd__nor4_1 U28211 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[10]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[11]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[14]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[13]), .Y(n22985) );
  sky130_fd_sc_hd__nor4_1 U28212 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[15]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[18]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[19]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[17]), .Y(n22984) );
  sky130_fd_sc_hd__nand4_1 U28213 ( .A(n22987), .B(n22986), .C(n22985), .D(
        n22984), .Y(n22993) );
  sky130_fd_sc_hd__nor4_1 U28214 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[1]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[2]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[31]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[3]), .Y(n22991) );
  sky130_fd_sc_hd__nor4_1 U28215 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[5]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[6]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[7]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[9]), .Y(n22990) );
  sky130_fd_sc_hd__nor4_1 U28216 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[0]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[4]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[8]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[12]), .Y(n22989) );
  sky130_fd_sc_hd__nor4_1 U28217 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[16]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[20]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[24]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[28]), .Y(n22988) );
  sky130_fd_sc_hd__nand4_1 U28218 ( .A(n22991), .B(n22990), .C(n22989), .D(
        n22988), .Y(n22992) );
  sky130_fd_sc_hd__o21a_1 U28219 ( .A1(n22993), .A2(n22992), .B1(n29593), .X(
        n29058) );
  sky130_fd_sc_hd__nor2_1 U28220 ( .A(n22995), .B(n22994), .Y(n29018) );
  sky130_fd_sc_hd__nand2_1 U28221 ( .A(j202_soc_core_bldc_core_00_comm[2]), 
        .B(j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld), .Y(n28588) );
  sky130_fd_sc_hd__nor2_1 U28222 ( .A(j202_soc_core_bldc_core_00_comm[1]), .B(
        n28588), .Y(n29089) );
  sky130_fd_sc_hd__nand2_1 U28223 ( .A(n22996), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld), .Y(n28585) );
  sky130_fd_sc_hd__nor2_1 U28224 ( .A(n28583), .B(n28585), .Y(n29088) );
  sky130_fd_sc_hd__nor2_1 U28225 ( .A(n23174), .B(n23520), .Y(n22997) );
  sky130_fd_sc_hd__and4_1 U28226 ( .A(n23005), .B(n11713), .C(n23004), .D(
        n23003), .X(n23006) );
  sky130_fd_sc_hd__nand2_1 U28227 ( .A(n23007), .B(n23006), .Y(n23008) );
  sky130_fd_sc_hd__nand2_1 U28228 ( .A(n23008), .B(n26329), .Y(n23015) );
  sky130_fd_sc_hd__o21a_1 U28229 ( .A1(n23012), .A2(n25130), .B1(n23011), .X(
        n23013) );
  sky130_fd_sc_hd__nand2b_1 U28230 ( .A_N(n23016), .B(n23026), .Y(n26425) );
  sky130_fd_sc_hd__xor2_1 U28231 ( .A(n25130), .B(n24671), .X(n26621) );
  sky130_fd_sc_hd__o2bb2ai_1 U28232 ( .B1(n26336), .B2(n26425), .A1_N(n26326), 
        .A2_N(n26621), .Y(n23018) );
  sky130_fd_sc_hd__o22ai_1 U28233 ( .A1(n26702), .A2(n26418), .B1(n26706), 
        .B2(n26419), .Y(n23017) );
  sky130_fd_sc_hd__nor2_1 U28234 ( .A(n23018), .B(n23017), .Y(n23032) );
  sky130_fd_sc_hd__nand2_1 U28235 ( .A(n23019), .B(n23047), .Y(n24777) );
  sky130_fd_sc_hd__nand2_1 U28236 ( .A(n24777), .B(n24785), .Y(n26431) );
  sky130_fd_sc_hd__nand2_1 U28237 ( .A(n23021), .B(n23918), .Y(n24773) );
  sky130_fd_sc_hd__nand2_1 U28238 ( .A(n24773), .B(n24785), .Y(n26412) );
  sky130_fd_sc_hd__o22a_1 U28239 ( .A1(n27375), .A2(n26431), .B1(n24667), .B2(
        n26412), .X(n23031) );
  sky130_fd_sc_hd__a21oi_1 U28240 ( .A1(n24671), .A2(n25415), .B1(n23022), .Y(
        n23024) );
  sky130_fd_sc_hd__nand2_1 U28241 ( .A(n27375), .B(n25308), .Y(n23023) );
  sky130_fd_sc_hd__o31a_1 U28242 ( .A1(n26707), .A2(n24778), .A3(n23024), .B1(
        n23023), .X(n23025) );
  sky130_fd_sc_hd__o21ai_1 U28243 ( .A1(n26705), .A2(n26424), .B1(n23025), .Y(
        n23028) );
  sky130_fd_sc_hd__nand2_1 U28244 ( .A(n23026), .B(n27422), .Y(n26416) );
  sky130_fd_sc_hd__o22ai_1 U28245 ( .A1(n25403), .A2(n26416), .B1(n26563), 
        .B2(n26427), .Y(n23027) );
  sky130_fd_sc_hd__nor2_1 U28246 ( .A(n23028), .B(n23027), .Y(n23030) );
  sky130_fd_sc_hd__nand3_1 U28247 ( .A(n23029), .B(n27402), .C(n26603), .Y(
        n24147) );
  sky130_fd_sc_hd__nand2b_1 U28248 ( .A_N(n24147), .B(n23920), .Y(n23060) );
  sky130_fd_sc_hd__o31ai_1 U28249 ( .A1(n25743), .A2(n26566), .A3(n23919), 
        .B1(n23060), .Y(n24772) );
  sky130_fd_sc_hd__nand2_1 U28250 ( .A(n24772), .B(n24785), .Y(n26411) );
  sky130_fd_sc_hd__nand4_1 U28251 ( .A(n23032), .B(n23031), .C(n23030), .D(
        n26411), .Y(n23033) );
  sky130_fd_sc_hd__a21oi_1 U28252 ( .A1(n23786), .A2(n26409), .B1(n23033), .Y(
        n23035) );
  sky130_fd_sc_hd__nand2_1 U28253 ( .A(n23172), .B(n23036), .Y(n23038) );
  sky130_fd_sc_hd__nand2b_1 U28254 ( .A_N(n23174), .B(n12171), .Y(n23037) );
  sky130_fd_sc_hd__nand2_1 U28255 ( .A(n25158), .B(n26360), .Y(n23040) );
  sky130_fd_sc_hd__nand2_1 U28257 ( .A(n23042), .B(n23041), .Y(n23044) );
  sky130_fd_sc_hd__a31oi_1 U28258 ( .A1(n23042), .A2(n26318), .A3(n23041), 
        .B1(n29535), .Y(n23043) );
  sky130_fd_sc_hd__a21oi_1 U28259 ( .A1(n27365), .A2(n25415), .B1(n26085), .Y(
        n23046) );
  sky130_fd_sc_hd__nand2_1 U28261 ( .A(n23048), .B(n24785), .Y(n26349) );
  sky130_fd_sc_hd__nor2_1 U28262 ( .A(n26582), .B(n26349), .Y(n23055) );
  sky130_fd_sc_hd__xnor2_1 U28263 ( .A(n23070), .B(n27365), .Y(n26665) );
  sky130_fd_sc_hd__nand2_1 U28264 ( .A(n23050), .B(n23049), .Y(n23051) );
  sky130_fd_sc_hd__nand2_1 U28265 ( .A(n23051), .B(n26329), .Y(n23053) );
  sky130_fd_sc_hd__o22a_1 U28266 ( .A1(n26567), .A2(n26418), .B1(n26336), .B2(
        n26419), .X(n23052) );
  sky130_fd_sc_hd__o211ai_1 U28267 ( .A1(n26415), .A2(n26665), .B1(n23053), 
        .C1(n23052), .Y(n23054) );
  sky130_fd_sc_hd__nor2_1 U28268 ( .A(n23055), .B(n23054), .Y(n23063) );
  sky130_fd_sc_hd__a22oi_1 U28269 ( .A1(n25308), .A2(n26582), .B1(n26077), 
        .B2(n27183), .Y(n23057) );
  sky130_fd_sc_hd__nand2_1 U28270 ( .A(n26338), .B(n27415), .Y(n23056) );
  sky130_fd_sc_hd__o211ai_1 U28271 ( .A1(n26426), .A2(n26427), .B1(n23057), 
        .C1(n23056), .Y(n23058) );
  sky130_fd_sc_hd__a21oi_1 U28272 ( .A1(n26342), .A2(n24052), .B1(n23058), .Y(
        n23062) );
  sky130_fd_sc_hd__o22ai_1 U28273 ( .A1(n26577), .A2(n26416), .B1(n26565), 
        .B2(n26424), .Y(n23059) );
  sky130_fd_sc_hd__a21oi_1 U28274 ( .A1(n26341), .A2(n26971), .B1(n23059), .Y(
        n23061) );
  sky130_fd_sc_hd__nand2b_1 U28275 ( .A_N(n23060), .B(n24785), .Y(n26344) );
  sky130_fd_sc_hd__nand4_1 U28276 ( .A(n23063), .B(n23062), .C(n23061), .D(
        n26344), .Y(n23064) );
  sky130_fd_sc_hd__a21oi_1 U28277 ( .A1(n23710), .A2(n26409), .B1(n23064), .Y(
        n23067) );
  sky130_fd_sc_hd__o21ai_0 U28278 ( .A1(n26352), .A2(n23070), .B1(n26351), .Y(
        n23065) );
  sky130_fd_sc_hd__nand2_1 U28279 ( .A(n27364), .B(n23065), .Y(n23066) );
  sky130_fd_sc_hd__nand2_1 U28280 ( .A(n12355), .B(n26360), .Y(n23075) );
  sky130_fd_sc_hd__nand2_1 U28281 ( .A(n11611), .B(n23073), .Y(n23074) );
  sky130_fd_sc_hd__nand2_1 U28282 ( .A(n23075), .B(n23074), .Y(
        j202_soc_core_j22_cpu_rf_N2729) );
  sky130_fd_sc_hd__nand2_1 U28283 ( .A(n23172), .B(n23080), .Y(n23078) );
  sky130_fd_sc_hd__nand2b_1 U28284 ( .A_N(n23174), .B(n23076), .Y(n23077) );
  sky130_fd_sc_hd__nand2_1 U28285 ( .A(n12355), .B(n26379), .Y(n23084) );
  sky130_fd_sc_hd__nand2_1 U28286 ( .A(n11611), .B(n23082), .Y(n23083) );
  sky130_fd_sc_hd__nand2_1 U28287 ( .A(n23084), .B(n23083), .Y(
        j202_soc_core_j22_cpu_rf_N3136) );
  sky130_fd_sc_hd__nand2_1 U28288 ( .A(n23172), .B(n23088), .Y(n23087) );
  sky130_fd_sc_hd__nand2b_1 U28289 ( .A_N(n23174), .B(n29568), .Y(n23086) );
  sky130_fd_sc_hd__nand3_2 U28290 ( .A(n23177), .B(n23087), .C(n23086), .Y(
        n27465) );
  sky130_fd_sc_hd__nand2_1 U28291 ( .A(n12355), .B(n25818), .Y(n23093) );
  sky130_fd_sc_hd__nand2_1 U28292 ( .A(n11611), .B(n23091), .Y(n23092) );
  sky130_fd_sc_hd__nand2_1 U28293 ( .A(n23093), .B(n23092), .Y(
        j202_soc_core_j22_cpu_rf_N2766) );
  sky130_fd_sc_hd__nand2_1 U28294 ( .A(n23172), .B(n23097), .Y(n23096) );
  sky130_fd_sc_hd__nand2b_1 U28295 ( .A_N(n23174), .B(n23094), .Y(n23095) );
  sky130_fd_sc_hd__nand2_1 U28296 ( .A(n12355), .B(n26374), .Y(n23101) );
  sky130_fd_sc_hd__nand2_1 U28297 ( .A(n11611), .B(n11136), .Y(n23100) );
  sky130_fd_sc_hd__nand2_1 U28298 ( .A(n23101), .B(n23100), .Y(
        j202_soc_core_j22_cpu_rf_N2877) );
  sky130_fd_sc_hd__nand2_1 U28299 ( .A(n23172), .B(n23104), .Y(n23103) );
  sky130_fd_sc_hd__nand2b_1 U28300 ( .A_N(n23174), .B(n12172), .Y(n23102) );
  sky130_fd_sc_hd__nand3_2 U28301 ( .A(n23177), .B(n23103), .C(n23102), .Y(
        n27212) );
  sky130_fd_sc_hd__nand2_1 U28302 ( .A(n12355), .B(n26362), .Y(n23108) );
  sky130_fd_sc_hd__nand2_1 U28303 ( .A(n11611), .B(n23106), .Y(n23107) );
  sky130_fd_sc_hd__nand2_1 U28304 ( .A(n23108), .B(n23107), .Y(
        j202_soc_core_j22_cpu_rf_N2803) );
  sky130_fd_sc_hd__nand2_1 U28305 ( .A(n23172), .B(n23112), .Y(n23111) );
  sky130_fd_sc_hd__nand2b_1 U28306 ( .A_N(n23174), .B(n23109), .Y(n23110) );
  sky130_fd_sc_hd__nand2_1 U28307 ( .A(n12355), .B(n25819), .Y(n23117) );
  sky130_fd_sc_hd__nand2_1 U28308 ( .A(n11611), .B(n23115), .Y(n23116) );
  sky130_fd_sc_hd__nand2_1 U28309 ( .A(n23117), .B(n23116), .Y(
        j202_soc_core_j22_cpu_rf_N2840) );
  sky130_fd_sc_hd__nand2_1 U28310 ( .A(n23172), .B(n23121), .Y(n23120) );
  sky130_fd_sc_hd__nand2b_1 U28311 ( .A_N(n23174), .B(n23118), .Y(n23119) );
  sky130_fd_sc_hd__nand2_1 U28312 ( .A(n12355), .B(n11109), .Y(n23125) );
  sky130_fd_sc_hd__o2bb2ai_1 U28313 ( .B1(n11115), .B2(n23172), .A1_N(n23121), 
        .A2_N(n23174), .Y(n23123) );
  sky130_fd_sc_hd__nand2_1 U28314 ( .A(n11611), .B(n11108), .Y(n23124) );
  sky130_fd_sc_hd__nand2_1 U28315 ( .A(n23125), .B(n23124), .Y(
        j202_soc_core_j22_cpu_rf_N3099) );
  sky130_fd_sc_hd__nand2_1 U28316 ( .A(n23172), .B(n23129), .Y(n23128) );
  sky130_fd_sc_hd__nand2b_1 U28317 ( .A_N(n23174), .B(n23126), .Y(n23127) );
  sky130_fd_sc_hd__nand2_1 U28318 ( .A(n12355), .B(n26369), .Y(n23134) );
  sky130_fd_sc_hd__nand2_1 U28319 ( .A(n11611), .B(n23132), .Y(n23133) );
  sky130_fd_sc_hd__nand2_1 U28320 ( .A(n23134), .B(n23133), .Y(
        j202_soc_core_j22_cpu_rf_N2988) );
  sky130_fd_sc_hd__nand2_1 U28321 ( .A(n12641), .B(n24257), .Y(n23135) );
  sky130_fd_sc_hd__inv_1 U28322 ( .A(n23211), .Y(n24399) );
  sky130_fd_sc_hd__nand2_1 U28323 ( .A(n23135), .B(n12665), .Y(n23136) );
  sky130_fd_sc_hd__inv_1 U28324 ( .A(n23606), .Y(n24400) );
  sky130_fd_sc_hd__nand4_1 U28326 ( .A(n27964), .B(n27947), .C(n24436), .D(
        n24456), .Y(n23137) );
  sky130_fd_sc_hd__nand2_1 U28327 ( .A(n12475), .B(n27898), .Y(n23138) );
  sky130_fd_sc_hd__inv_1 U28328 ( .A(n24705), .Y(n23142) );
  sky130_fd_sc_hd__nand2_1 U28329 ( .A(n27298), .B(n29071), .Y(n23162) );
  sky130_fd_sc_hd__nor2_1 U28330 ( .A(n23606), .B(n12362), .Y(n23202) );
  sky130_fd_sc_hd__nand2_1 U28331 ( .A(n24360), .B(n27230), .Y(n27789) );
  sky130_fd_sc_hd__nand2_1 U28332 ( .A(n23202), .B(n24386), .Y(n23187) );
  sky130_fd_sc_hd__inv_1 U28333 ( .A(n23148), .Y(n23149) );
  sky130_fd_sc_hd__o21a_1 U28335 ( .A1(n23150), .A2(n24353), .B1(n23802), .X(
        n23153) );
  sky130_fd_sc_hd__nand2_1 U28336 ( .A(n12462), .B(n29075), .Y(n27891) );
  sky130_fd_sc_hd__nand2_1 U28337 ( .A(n24265), .B(n13271), .Y(n23203) );
  sky130_fd_sc_hd__o22ai_1 U28338 ( .A1(n27891), .A2(n23606), .B1(n23203), 
        .B2(n29548), .Y(n23151) );
  sky130_fd_sc_hd__nor2_1 U28339 ( .A(n29071), .B(n23586), .Y(n23156) );
  sky130_fd_sc_hd__nand2_1 U28340 ( .A(n23211), .B(n27298), .Y(n23155) );
  sky130_fd_sc_hd__and2_1 U28341 ( .A(n12150), .B(n24335), .X(n27691) );
  sky130_fd_sc_hd__nand2_1 U28342 ( .A(n23164), .B(n24350), .Y(n24253) );
  sky130_fd_sc_hd__nand2_1 U28343 ( .A(n27947), .B(n27928), .Y(n27949) );
  sky130_fd_sc_hd__o2bb2ai_1 U28344 ( .B1(n23168), .B2(n23172), .A1_N(n23171), 
        .A2_N(n23174), .Y(n23170) );
  sky130_fd_sc_hd__nand2_1 U28345 ( .A(n23172), .B(n23171), .Y(n23176) );
  sky130_fd_sc_hd__nand2b_1 U28346 ( .A_N(n23174), .B(n23173), .Y(n23175) );
  sky130_fd_sc_hd__nand2_1 U28347 ( .A(n29009), .B(n29015), .Y(n23599) );
  sky130_fd_sc_hd__o21ai_1 U28348 ( .A1(n24094), .A2(n11646), .B1(n12436), .Y(
        n23181) );
  sky130_fd_sc_hd__nand4_1 U28349 ( .A(n12665), .B(n27892), .C(n23182), .D(
        n23181), .Y(n23183) );
  sky130_fd_sc_hd__nand2_1 U28350 ( .A(n29077), .B(n29015), .Y(n23186) );
  sky130_fd_sc_hd__nand2b_1 U28351 ( .A_N(n27817), .B(n23195), .Y(n23190) );
  sky130_fd_sc_hd__nand2b_1 U28352 ( .A_N(n23197), .B(n27904), .Y(n27164) );
  sky130_fd_sc_hd__nand2_1 U28353 ( .A(n23190), .B(n27164), .Y(n23858) );
  sky130_fd_sc_hd__nor2_1 U28354 ( .A(n23191), .B(n27956), .Y(n24407) );
  sky130_fd_sc_hd__nor2_1 U28355 ( .A(n27978), .B(n27947), .Y(n27900) );
  sky130_fd_sc_hd__or3_1 U28356 ( .A(n27919), .B(n24407), .C(n27900), .X(
        n23201) );
  sky130_fd_sc_hd__nand2b_1 U28357 ( .A_N(n27175), .B(
        j202_soc_core_j22_cpu_opst[2]), .Y(n23193) );
  sky130_fd_sc_hd__nand3_1 U28358 ( .A(n23196), .B(n27904), .C(n23195), .Y(
        n23596) );
  sky130_fd_sc_hd__nand2b_1 U28359 ( .A_N(n27956), .B(n23192), .Y(n24364) );
  sky130_fd_sc_hd__nand2_1 U28360 ( .A(n23193), .B(n24364), .Y(n27264) );
  sky130_fd_sc_hd__nand2_1 U28361 ( .A(n27905), .B(
        j202_soc_core_j22_cpu_opst[2]), .Y(n24343) );
  sky130_fd_sc_hd__nand2_1 U28362 ( .A(n27166), .B(n24343), .Y(n23598) );
  sky130_fd_sc_hd__nand2_1 U28363 ( .A(n27932), .B(n23598), .Y(n23199) );
  sky130_fd_sc_hd__and3_1 U28364 ( .A(n23863), .B(n23196), .C(n23195), .X(
        n24103) );
  sky130_fd_sc_hd__nand2_1 U28365 ( .A(j202_soc_core_j22_cpu_opst[2]), .B(
        j202_soc_core_j22_cpu_opst[0]), .Y(n23595) );
  sky130_fd_sc_hd__nor2_1 U28366 ( .A(n23595), .B(n23197), .Y(n24393) );
  sky130_fd_sc_hd__nor2_1 U28367 ( .A(n24103), .B(n24393), .Y(n23957) );
  sky130_fd_sc_hd__nand2b_1 U28368 ( .A_N(n27956), .B(n23198), .Y(n27942) );
  sky130_fd_sc_hd__o211a_2 U28369 ( .A1(j202_soc_core_j22_cpu_opst[0]), .A2(
        n27947), .B1(n23199), .C1(n27942), .X(n23200) );
  sky130_fd_sc_hd__nand2b_1 U28370 ( .A_N(n27264), .B(n23200), .Y(n24404) );
  sky130_fd_sc_hd__inv_1 U28371 ( .A(n23202), .Y(n23205) );
  sky130_fd_sc_hd__nand2_1 U28372 ( .A(n24262), .B(n23204), .Y(n24389) );
  sky130_fd_sc_hd__nand2_1 U28373 ( .A(n23205), .B(n24389), .Y(n24325) );
  sky130_fd_sc_hd__nand2_1 U28375 ( .A(n23208), .B(n27928), .Y(n23209) );
  sky130_fd_sc_hd__nand2_1 U28376 ( .A(n23954), .B(n11792), .Y(n24324) );
  sky130_fd_sc_hd__nand2_1 U28377 ( .A(n27957), .B(n24324), .Y(n23212) );
  sky130_fd_sc_hd__nor2_1 U28378 ( .A(n23232), .B(n23233), .Y(n23217) );
  sky130_fd_sc_hd__nor2_1 U28379 ( .A(n23236), .B(n23235), .Y(n23216) );
  sky130_fd_sc_hd__nor2_1 U28380 ( .A(n23231), .B(n23230), .Y(n23215) );
  sky130_fd_sc_hd__nor2_1 U28381 ( .A(n23237), .B(n23234), .Y(n23214) );
  sky130_fd_sc_hd__nand4_1 U28382 ( .A(n23216), .B(n23217), .C(n23215), .D(
        n23214), .Y(n23218) );
  sky130_fd_sc_hd__inv_2 U28383 ( .A(n23218), .Y(n23229) );
  sky130_fd_sc_hd__nor2_1 U28384 ( .A(n23242), .B(n23244), .Y(n23221) );
  sky130_fd_sc_hd__nor2_1 U28385 ( .A(n23243), .B(n26873), .Y(n23220) );
  sky130_fd_sc_hd__nor2_1 U28386 ( .A(n23248), .B(n23241), .Y(n23219) );
  sky130_fd_sc_hd__nand3_1 U28387 ( .A(n23221), .B(n23219), .C(n23220), .Y(
        n23222) );
  sky130_fd_sc_hd__inv_2 U28388 ( .A(n23222), .Y(n23228) );
  sky130_fd_sc_hd__inv_2 U28389 ( .A(n23247), .Y(n23268) );
  sky130_fd_sc_hd__nand4_1 U28390 ( .A(n23225), .B(n23268), .C(n23224), .D(
        n23223), .Y(n23226) );
  sky130_fd_sc_hd__inv_2 U28391 ( .A(n23226), .Y(n23227) );
  sky130_fd_sc_hd__nand4_1 U28392 ( .A(n23233), .B(n23232), .C(n23231), .D(
        n23230), .Y(n23239) );
  sky130_fd_sc_hd__nand4_1 U28393 ( .A(n23237), .B(n23236), .C(n23235), .D(
        n23234), .Y(n23238) );
  sky130_fd_sc_hd__nand2_1 U28394 ( .A(n23241), .B(n23240), .Y(n23246) );
  sky130_fd_sc_hd__nand4_1 U28395 ( .A(n23244), .B(n23243), .C(n26873), .D(
        n23242), .Y(n23245) );
  sky130_fd_sc_hd__nor2_1 U28396 ( .A(n23246), .B(n23245), .Y(n23251) );
  sky130_fd_sc_hd__and4_1 U28397 ( .A(n11128), .B(n23249), .C(n23248), .D(
        n23247), .X(n23250) );
  sky130_fd_sc_hd__nand2_1 U28398 ( .A(n11614), .B(n23255), .Y(n23254) );
  sky130_fd_sc_hd__inv_2 U28399 ( .A(n12917), .Y(n24169) );
  sky130_fd_sc_hd__nand2_1 U28400 ( .A(n24169), .B(n25345), .Y(n23258) );
  sky130_fd_sc_hd__nand2_1 U28401 ( .A(n13286), .B(n23258), .Y(
        j202_soc_core_j22_cpu_ml_maclj[22]) );
  sky130_fd_sc_hd__nand2_1 U28402 ( .A(n24169), .B(n24062), .Y(n23259) );
  sky130_fd_sc_hd__nand2_1 U28403 ( .A(n13285), .B(n23259), .Y(
        j202_soc_core_j22_cpu_ml_maclj[21]) );
  sky130_fd_sc_hd__nand2_1 U28404 ( .A(n24169), .B(n24013), .Y(n23261) );
  sky130_fd_sc_hd__nand2_1 U28405 ( .A(n13299), .B(n23261), .Y(
        j202_soc_core_j22_cpu_ml_maclj[25]) );
  sky130_fd_sc_hd__nand2_1 U28406 ( .A(n24169), .B(n25049), .Y(n23263) );
  sky130_fd_sc_hd__nand2_1 U28407 ( .A(n13284), .B(n23263), .Y(
        j202_soc_core_j22_cpu_ml_maclj[26]) );
  sky130_fd_sc_hd__nand2_1 U28408 ( .A(n24169), .B(n24586), .Y(n23264) );
  sky130_fd_sc_hd__nand2_1 U28409 ( .A(n13283), .B(n23264), .Y(
        j202_soc_core_j22_cpu_ml_maclj[20]) );
  sky130_fd_sc_hd__nand2_1 U28410 ( .A(n24169), .B(n24742), .Y(n23265) );
  sky130_fd_sc_hd__nand2_1 U28411 ( .A(n13282), .B(n23265), .Y(
        j202_soc_core_j22_cpu_ml_maclj[23]) );
  sky130_fd_sc_hd__nand2_1 U28412 ( .A(n24169), .B(n24128), .Y(n23266) );
  sky130_fd_sc_hd__nand2_1 U28413 ( .A(n13281), .B(n23266), .Y(
        j202_soc_core_j22_cpu_ml_maclj[19]) );
  sky130_fd_sc_hd__nand2_4 U28414 ( .A(n12487), .B(n26865), .Y(n27273) );
  sky130_fd_sc_hd__inv_2 U28415 ( .A(n27273), .Y(n25829) );
  sky130_fd_sc_hd__a21oi_1 U28416 ( .A1(j202_soc_core_j22_cpu_ml_bufa[12]), 
        .A2(n27187), .B1(n25829), .Y(n23273) );
  sky130_fd_sc_hd__nand2_1 U28417 ( .A(n23273), .B(n23272), .Y(
        j202_soc_core_j22_cpu_ml_machj[12]) );
  sky130_fd_sc_hd__nand2_1 U28418 ( .A(n26802), .B(n23276), .Y(n23277) );
  sky130_fd_sc_hd__nor2_1 U28419 ( .A(j202_soc_core_j22_cpu_regop_We__1_), .B(
        n12366), .Y(n23529) );
  sky130_fd_sc_hd__nand3_1 U28420 ( .A(n23529), .B(
        j202_soc_core_j22_cpu_regop_We__3_), .C(n23279), .Y(n26805) );
  sky130_fd_sc_hd__nand2b_1 U28421 ( .A_N(n14849), .B(n26801), .Y(n27334) );
  sky130_fd_sc_hd__nor2_1 U28422 ( .A(j202_soc_core_j22_cpu_intack), .B(n27334), .Y(n25756) );
  sky130_fd_sc_hd__nand2_1 U28423 ( .A(n23280), .B(n25756), .Y(n23287) );
  sky130_fd_sc_hd__nand2b_1 U28424 ( .A_N(n14849), .B(
        j202_soc_core_j22_cpu_intack), .Y(n25451) );
  sky130_fd_sc_hd__nand2_1 U28425 ( .A(n27334), .B(n25451), .Y(n25539) );
  sky130_fd_sc_hd__nand2b_1 U28426 ( .A_N(n24113), .B(n23282), .Y(n23531) );
  sky130_fd_sc_hd__nor2_1 U28427 ( .A(n23283), .B(n23531), .Y(n23547) );
  sky130_fd_sc_hd__o22ai_1 U28428 ( .A1(n23284), .A2(n25451), .B1(n23547), 
        .B2(n25539), .Y(n26906) );
  sky130_fd_sc_hd__a21oi_1 U28429 ( .A1(j202_soc_core_intr_level__2_), .A2(
        n26907), .B1(n26906), .Y(n23285) );
  sky130_fd_sc_hd__o21a_1 U28430 ( .A1(n25539), .A2(n26556), .B1(n23285), .X(
        n23286) );
  sky130_fd_sc_hd__nand2_1 U28431 ( .A(n23287), .B(n23286), .Y(
        j202_soc_core_j22_cpu_rf_N3390) );
  sky130_fd_sc_hd__nand2_1 U28432 ( .A(n28964), .B(n29559), .Y(n23307) );
  sky130_fd_sc_hd__nor2_1 U28433 ( .A(j202_soc_core_j22_cpu_memop_MEM__2_), 
        .B(n27721), .Y(n23290) );
  sky130_fd_sc_hd__nand2b_1 U28434 ( .A_N(n23573), .B(n23289), .Y(n23294) );
  sky130_fd_sc_hd__nand2_1 U28435 ( .A(n23290), .B(
        j202_soc_core_j22_cpu_memop_MEM__1_), .Y(n23291) );
  sky130_fd_sc_hd__nand3_1 U28436 ( .A(n23293), .B(n23292), .C(n23291), .Y(
        n23575) );
  sky130_fd_sc_hd__a21oi_1 U28437 ( .A1(n29033), .A2(n23294), .B1(n23575), .Y(
        n23563) );
  sky130_fd_sc_hd__nand2_1 U28438 ( .A(n29033), .B(n27914), .Y(n23295) );
  sky130_fd_sc_hd__o211ai_1 U28439 ( .A1(n23298), .A2(n23297), .B1(n23296), 
        .C1(n23295), .Y(n27621) );
  sky130_fd_sc_hd__nand2b_1 U28440 ( .A_N(n29033), .B(n23299), .Y(n23303) );
  sky130_fd_sc_hd__nand2_1 U28441 ( .A(n23300), .B(n24280), .Y(n23301) );
  sky130_fd_sc_hd__nand3_1 U28442 ( .A(n23303), .B(n23302), .C(n23301), .Y(
        n27620) );
  sky130_fd_sc_hd__a21oi_1 U28443 ( .A1(n29559), .A2(n27621), .B1(n27620), .Y(
        n23304) );
  sky130_fd_sc_hd__nand2_1 U28445 ( .A(n23307), .B(n13335), .Y(
        j202_soc_core_ahb2aqu_00_N163) );
  sky130_fd_sc_hd__clkbuf_1 U28446 ( .A(la_data_out[16]), .X(io_out[36]) );
  sky130_fd_sc_hd__and3_1 U28447 ( .A(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[0]), .C(n23455), .X(io_oeb[12]) );
  sky130_fd_sc_hd__clkbuf_1 U28448 ( .A(la_data_out[15]), .X(io_out[35]) );
  sky130_fd_sc_hd__clkbuf_1 U28449 ( .A(io_oeb[12]), .X(io_oeb[10]) );
  sky130_fd_sc_hd__clkbuf_1 U28450 ( .A(la_data_out[14]), .X(io_out[34]) );
  sky130_fd_sc_hd__clkbuf_1 U28451 ( .A(la_data_out[13]), .X(io_out[33]) );
  sky130_fd_sc_hd__clkbuf_1 U28452 ( .A(la_data_out[12]), .X(io_out[32]) );
  sky130_fd_sc_hd__clkbuf_1 U28453 ( .A(la_data_out[0]), .X(io_out[0]) );
  sky130_fd_sc_hd__clkbuf_1 U28454 ( .A(la_data_out[10]), .X(io_out[30]) );
  sky130_fd_sc_hd__clkbuf_1 U28455 ( .A(la_data_out[1]), .X(io_out[1]) );
  sky130_fd_sc_hd__clkbuf_1 U28456 ( .A(la_data_out[9]), .X(io_out[29]) );
  sky130_fd_sc_hd__clkbuf_1 U28457 ( .A(la_data_out[8]), .X(io_out[28]) );
  sky130_fd_sc_hd__clkbuf_1 U28458 ( .A(la_data_out[7]), .X(io_out[27]) );
  sky130_fd_sc_hd__clkbuf_1 U28459 ( .A(la_data_out[6]), .X(io_out[26]) );
  sky130_fd_sc_hd__clkbuf_1 U28460 ( .A(la_data_out[3]), .X(io_out[3]) );
  sky130_fd_sc_hd__clkbuf_1 U28461 ( .A(la_data_out[5]), .X(io_out[7]) );
  sky130_fd_sc_hd__clkbuf_1 U28462 ( .A(la_data_out[4]), .X(io_out[4]) );
  sky130_fd_sc_hd__nand2_1 U28463 ( .A(j202_soc_core_uart_TOP_rx_go), .B(
        j202_soc_core_uart_TOP_rx_sio_ce), .Y(n28000) );
  sky130_fd_sc_hd__o21ai_1 U28464 ( .A1(n23309), .A2(n23308), .B1(
        j202_soc_core_uart_TOP_rx_valid), .Y(n23310) );
  sky130_fd_sc_hd__nor2_1 U28465 ( .A(j202_soc_core_uart_TOP_rx_valid_r), .B(
        n23310), .Y(n27138) );
  sky130_fd_sc_hd__nand2_1 U28466 ( .A(n27138), .B(
        j202_soc_core_uart_TOP_rx_fifo_wp[0]), .Y(n27133) );
  sky130_fd_sc_hd__nor2_1 U28467 ( .A(n27134), .B(n27133), .Y(n29355) );
  sky130_fd_sc_hd__clkinv_1 U28468 ( .A(gpio_en_o[12]), .Y(io_oeb[32]) );
  sky130_fd_sc_hd__nand2_1 U28469 ( .A(n23453), .B(
        j202_soc_core_gpio_core_00_reg_addr[3]), .Y(n27652) );
  sky130_fd_sc_hd__and4_1 U28470 ( .A(j202_soc_core_pstrb[1]), .B(
        j202_soc_core_pstrb[0]), .C(j202_soc_core_pstrb[3]), .D(
        j202_soc_core_pstrb[2]), .X(n23311) );
  sky130_fd_sc_hd__nand2_1 U28471 ( .A(j202_soc_core_pwrite[2]), .B(n23311), 
        .Y(n23313) );
  sky130_fd_sc_hd__nand3_1 U28472 ( .A(n24316), .B(n23312), .C(
        j202_soc_core_ahb2apb_02_state[1]), .Y(n27648) );
  sky130_fd_sc_hd__nor2_1 U28473 ( .A(n23313), .B(n27648), .Y(n24173) );
  sky130_fd_sc_hd__nor2_1 U28474 ( .A(j202_soc_core_gpio_core_00_reg_addr[7]), 
        .B(j202_soc_core_gpio_core_00_reg_addr[1]), .Y(n23315) );
  sky130_fd_sc_hd__nor2_1 U28475 ( .A(j202_soc_core_gpio_core_00_reg_addr[5]), 
        .B(j202_soc_core_gpio_core_00_reg_addr[6]), .Y(n23314) );
  sky130_fd_sc_hd__nand3_1 U28476 ( .A(n23315), .B(n23314), .C(n27633), .Y(
        n27651) );
  sky130_fd_sc_hd__nand3_1 U28477 ( .A(n24173), .B(n23316), .C(n23452), .Y(
        n27640) );
  sky130_fd_sc_hd__o21ai_2 U28478 ( .A1(n27652), .A2(n27640), .B1(n12142), .Y(
        n10675) );
  sky130_fd_sc_hd__nor2_1 U28479 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[0]), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[1]), .Y(n28749) );
  sky130_fd_sc_hd__nand3_1 U28480 ( .A(n28749), .B(n25023), .C(n23317), .Y(
        n28056) );
  sky130_fd_sc_hd__nand2b_1 U28481 ( .A_N(
        j202_soc_core_wbqspiflash_00_reset_counter[4]), .B(n23318), .Y(n28059)
         );
  sky130_fd_sc_hd__nor2_1 U28482 ( .A(n28059), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[5]), .Y(n28061) );
  sky130_fd_sc_hd__nand2b_1 U28483 ( .A_N(
        j202_soc_core_wbqspiflash_00_reset_counter[6]), .B(n28061), .Y(n28064)
         );
  sky130_fd_sc_hd__nor2_1 U28484 ( .A(n28064), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[7]), .Y(n25014) );
  sky130_fd_sc_hd__nand2_1 U28485 ( .A(n25014), .B(n23319), .Y(n25016) );
  sky130_fd_sc_hd__nand2b_1 U28486 ( .A_N(n25016), .B(n25022), .Y(n26183) );
  sky130_fd_sc_hd__nand2_1 U28487 ( .A(n23320), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n25024) );
  sky130_fd_sc_hd__nand2_1 U28488 ( .A(n26035), .B(n25916), .Y(n28063) );
  sky130_fd_sc_hd__nand2_1 U28489 ( .A(n23324), .B(n23329), .Y(n24053) );
  sky130_fd_sc_hd__nor2_1 U28490 ( .A(n27456), .B(n27438), .Y(n27454) );
  sky130_fd_sc_hd__o31ai_1 U28491 ( .A1(j202_soc_core_j22_cpu_macop_MAC_[4]), 
        .A2(n23332), .A3(n24278), .B1(n27454), .Y(n23325) );
  sky130_fd_sc_hd__nand2_1 U28492 ( .A(n23331), .B(n23330), .Y(n24023) );
  sky130_fd_sc_hd__nand2_1 U28493 ( .A(n26255), .B(
        j202_soc_core_wbqspiflash_00_state[2]), .Y(n26008) );
  sky130_fd_sc_hd__nand2_1 U28494 ( .A(n25954), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n26007) );
  sky130_fd_sc_hd__nor2_1 U28495 ( .A(n26008), .B(n26007), .Y(n25982) );
  sky130_fd_sc_hd__nand2b_1 U28496 ( .A_N(n26007), .B(n26035), .Y(n26242) );
  sky130_fd_sc_hd__nand2_1 U28497 ( .A(n28268), .B(
        j202_soc_core_wbqspiflash_00_spi_valid), .Y(n26244) );
  sky130_fd_sc_hd__nand3_1 U28498 ( .A(j202_soc_core_wbqspiflash_00_spi_valid), 
        .B(n23333), .C(n26226), .Y(n23334) );
  sky130_fd_sc_hd__nor2_1 U28499 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(n26008), .Y(n28228) );
  sky130_fd_sc_hd__nand2_1 U28500 ( .A(n25954), .B(n28228), .Y(n25929) );
  sky130_fd_sc_hd__o22ai_1 U28501 ( .A1(n26242), .A2(n26244), .B1(n23334), 
        .B2(n25929), .Y(n23335) );
  sky130_fd_sc_hd__a21oi_1 U28502 ( .A1(j202_soc_core_wbqspiflash_00_spi_valid), .A2(n25982), .B1(n23335), .Y(n26142) );
  sky130_fd_sc_hd__nand2_1 U28503 ( .A(n27037), .B(n28058), .Y(n25993) );
  sky130_fd_sc_hd__nor2_1 U28504 ( .A(n10958), .B(n23336), .Y(n26032) );
  sky130_fd_sc_hd__nand2_1 U28505 ( .A(n28106), .B(n28116), .Y(n26148) );
  sky130_fd_sc_hd__nor2_1 U28506 ( .A(
        j202_soc_core_wbqspiflash_00_write_in_progress), .B(n26148), .Y(n25972) );
  sky130_fd_sc_hd__nand2_1 U28507 ( .A(j202_soc_core_wbqspiflash_00_state[1]), 
        .B(j202_soc_core_wbqspiflash_00_state[3]), .Y(n26046) );
  sky130_fd_sc_hd__nand2_1 U28508 ( .A(n28228), .B(n25926), .Y(n26115) );
  sky130_fd_sc_hd__nor2_1 U28509 ( .A(n26476), .B(n26115), .Y(n24995) );
  sky130_fd_sc_hd__a31oi_1 U28510 ( .A1(n26155), .A2(n26032), .A3(n25972), 
        .B1(n24995), .Y(n23337) );
  sky130_fd_sc_hd__a21o_1 U28511 ( .A1(n26142), .A2(n23337), .B1(n28590), .X(
        n23338) );
  sky130_fd_sc_hd__nand4_1 U28512 ( .A(n28966), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .C(n25949), .D(n10959), .Y(
        n26159) );
  sky130_fd_sc_hd__nor2_1 U28513 ( .A(n25880), .B(n26244), .Y(n26127) );
  sky130_fd_sc_hd__nor2_1 U28514 ( .A(j202_soc_core_wbqspiflash_00_state[4]), 
        .B(n28243), .Y(n28230) );
  sky130_fd_sc_hd__nor2_1 U28515 ( .A(j202_soc_core_qspi_wb_addr[24]), .B(
        n26131), .Y(n26149) );
  sky130_fd_sc_hd__nand2_1 U28516 ( .A(n10958), .B(n26149), .Y(n23339) );
  sky130_fd_sc_hd__nor2_1 U28517 ( .A(n23339), .B(n12292), .Y(n23439) );
  sky130_fd_sc_hd__nor2_1 U28518 ( .A(j202_soc_core_qspi_wb_addr[23]), .B(
        n23340), .Y(n23438) );
  sky130_fd_sc_hd__xor2_1 U28519 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .B(
        j202_soc_core_qspi_wb_addr[22]), .X(n23342) );
  sky130_fd_sc_hd__xnor2_1 U28520 ( .A(n23343), .B(n23342), .Y(n23431) );
  sky130_fd_sc_hd__xnor2_1 U28521 ( .A(n23345), .B(n13311), .Y(n23424) );
  sky130_fd_sc_hd__xor2_1 U28522 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .B(
        j202_soc_core_qspi_wb_addr[18]), .X(n23347) );
  sky130_fd_sc_hd__xnor2_1 U28523 ( .A(n23348), .B(n23347), .Y(n23417) );
  sky130_fd_sc_hd__xor2_1 U28524 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]), .B(
        j202_soc_core_qspi_wb_addr[16]), .X(n23350) );
  sky130_fd_sc_hd__xnor2_1 U28525 ( .A(n23351), .B(n23350), .Y(n23410) );
  sky130_fd_sc_hd__xor2_1 U28526 ( .A(j202_soc_core_qspi_wb_addr[9]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[9]), .X(n23353) );
  sky130_fd_sc_hd__xnor2_1 U28527 ( .A(n23354), .B(n23353), .Y(n23357) );
  sky130_fd_sc_hd__xnor2_1 U28528 ( .A(n23355), .B(n12292), .Y(n23356) );
  sky130_fd_sc_hd__nor2_1 U28529 ( .A(n23357), .B(n23356), .Y(n23367) );
  sky130_fd_sc_hd__xnor2_1 U28530 ( .A(j202_soc_core_qspi_wb_addr[7]), .B(
        n23358), .Y(n23359) );
  sky130_fd_sc_hd__xnor2_1 U28531 ( .A(n23360), .B(n23359), .Y(n23365) );
  sky130_fd_sc_hd__xnor2_1 U28532 ( .A(j202_soc_core_qspi_wb_addr[6]), .B(
        n23361), .Y(n23362) );
  sky130_fd_sc_hd__xnor2_1 U28533 ( .A(n23363), .B(n23362), .Y(n23364) );
  sky130_fd_sc_hd__nor2_1 U28534 ( .A(n23365), .B(n23364), .Y(n23366) );
  sky130_fd_sc_hd__nand2_1 U28535 ( .A(n23367), .B(n23366), .Y(n23382) );
  sky130_fd_sc_hd__xnor2_1 U28536 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .B(
        j202_soc_core_qspi_wb_addr[2]), .Y(n23370) );
  sky130_fd_sc_hd__xnor2_1 U28537 ( .A(j202_soc_core_qspi_wb_addr[3]), .B(
        n23470), .Y(n23368) );
  sky130_fd_sc_hd__xnor2_1 U28538 ( .A(n23469), .B(n23368), .Y(n23369) );
  sky130_fd_sc_hd__nor2_1 U28539 ( .A(n23370), .B(n23369), .Y(n23380) );
  sky130_fd_sc_hd__xnor2_1 U28540 ( .A(j202_soc_core_qspi_wb_addr[5]), .B(
        n23371), .Y(n23372) );
  sky130_fd_sc_hd__xnor2_1 U28541 ( .A(n23373), .B(n23372), .Y(n23378) );
  sky130_fd_sc_hd__xnor2_1 U28542 ( .A(j202_soc_core_qspi_wb_addr[4]), .B(
        n23374), .Y(n23375) );
  sky130_fd_sc_hd__xnor2_1 U28543 ( .A(n23376), .B(n23375), .Y(n23377) );
  sky130_fd_sc_hd__nor2_1 U28544 ( .A(n23378), .B(n23377), .Y(n23379) );
  sky130_fd_sc_hd__nand2_1 U28545 ( .A(n23380), .B(n23379), .Y(n23381) );
  sky130_fd_sc_hd__nor2_1 U28546 ( .A(n23382), .B(n23381), .Y(n23408) );
  sky130_fd_sc_hd__xor2_1 U28547 ( .A(n23384), .B(n13313), .X(n23389) );
  sky130_fd_sc_hd__xor2_1 U28548 ( .A(j202_soc_core_qspi_wb_addr[15]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[15]), .X(n23386) );
  sky130_fd_sc_hd__xor2_1 U28549 ( .A(n23387), .B(n23386), .X(n23388) );
  sky130_fd_sc_hd__nand2_1 U28550 ( .A(n23389), .B(n23388), .Y(n23406) );
  sky130_fd_sc_hd__xnor2_1 U28551 ( .A(n23391), .B(n13297), .Y(n23395) );
  sky130_fd_sc_hd__xnor2_1 U28552 ( .A(n23393), .B(n13298), .Y(n23394) );
  sky130_fd_sc_hd__nor2_1 U28553 ( .A(n23395), .B(n23394), .Y(n23404) );
  sky130_fd_sc_hd__xnor2_1 U28554 ( .A(n23397), .B(n13312), .Y(n23402) );
  sky130_fd_sc_hd__xor2_1 U28555 ( .A(j202_soc_core_qspi_wb_addr[12]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[12]), .X(n23399) );
  sky130_fd_sc_hd__xnor2_1 U28556 ( .A(n23400), .B(n23399), .Y(n23401) );
  sky130_fd_sc_hd__nor2_1 U28557 ( .A(n23402), .B(n23401), .Y(n23403) );
  sky130_fd_sc_hd__nand2_1 U28558 ( .A(n23404), .B(n23403), .Y(n23405) );
  sky130_fd_sc_hd__nor2_1 U28559 ( .A(n23406), .B(n23405), .Y(n23407) );
  sky130_fd_sc_hd__nand2_1 U28560 ( .A(n23408), .B(n23407), .Y(n23409) );
  sky130_fd_sc_hd__nor2_1 U28561 ( .A(n23410), .B(n23409), .Y(n23415) );
  sky130_fd_sc_hd__xor2_1 U28562 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]), .B(
        j202_soc_core_qspi_wb_addr[17]), .X(n23412) );
  sky130_fd_sc_hd__xor2_1 U28563 ( .A(n23413), .B(n23412), .X(n23414) );
  sky130_fd_sc_hd__nand2_1 U28564 ( .A(n23415), .B(n23414), .Y(n23416) );
  sky130_fd_sc_hd__nor2_1 U28565 ( .A(n23417), .B(n23416), .Y(n23422) );
  sky130_fd_sc_hd__xor2_1 U28566 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .B(
        j202_soc_core_qspi_wb_addr[19]), .X(n23419) );
  sky130_fd_sc_hd__xor2_1 U28567 ( .A(n23420), .B(n23419), .X(n23421) );
  sky130_fd_sc_hd__nand2_1 U28568 ( .A(n23422), .B(n23421), .Y(n23423) );
  sky130_fd_sc_hd__nor2_1 U28569 ( .A(n23424), .B(n23423), .Y(n23429) );
  sky130_fd_sc_hd__xor2_1 U28570 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]), .B(
        j202_soc_core_qspi_wb_addr[21]), .X(n23426) );
  sky130_fd_sc_hd__xor2_1 U28571 ( .A(n23427), .B(n23426), .X(n23428) );
  sky130_fd_sc_hd__nand2_1 U28572 ( .A(n23429), .B(n23428), .Y(n23430) );
  sky130_fd_sc_hd__nor2_1 U28573 ( .A(n23431), .B(n23430), .Y(n23436) );
  sky130_fd_sc_hd__xor2_1 U28574 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]), .B(
        j202_soc_core_qspi_wb_addr[23]), .X(n23433) );
  sky130_fd_sc_hd__xor2_1 U28575 ( .A(n23434), .B(n23433), .X(n23435) );
  sky130_fd_sc_hd__nand2_1 U28576 ( .A(n23436), .B(n23435), .Y(n23437) );
  sky130_fd_sc_hd__nor2_1 U28577 ( .A(n23438), .B(n23437), .Y(n26181) );
  sky130_fd_sc_hd__nand2_1 U28578 ( .A(n23439), .B(n26181), .Y(n25882) );
  sky130_fd_sc_hd__nor2_1 U28579 ( .A(j202_soc_core_wbqspiflash_00_spi_wr), 
        .B(n25882), .Y(n26000) );
  sky130_fd_sc_hd__nor2_1 U28580 ( .A(n28058), .B(n28243), .Y(n26009) );
  sky130_fd_sc_hd__and3_1 U28581 ( .A(n26000), .B(j202_soc_core_qspi_wb_cyc), 
        .C(n26009), .X(n23440) );
  sky130_fd_sc_hd__nor2_1 U28582 ( .A(j202_soc_core_wbqspiflash_00_state[2]), 
        .B(n26255), .Y(n26188) );
  sky130_fd_sc_hd__nor2_1 U28583 ( .A(n26188), .B(n28080), .Y(n28067) );
  sky130_fd_sc_hd__nand2_1 U28585 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__1_), 
        .B(j202_soc_core_j22_cpu_regop_M_Rn__0_), .Y(n23541) );
  sky130_fd_sc_hd__nand4_1 U28586 ( .A(n24291), .B(n23493), .C(
        j202_soc_core_j22_cpu_regop_M_Rn__3_), .D(
        j202_soc_core_j22_cpu_regop_M_Rn__2_), .Y(n23537) );
  sky130_fd_sc_hd__nand2_1 U28587 ( .A(n23444), .B(n23443), .Y(n23451) );
  sky130_fd_sc_hd__nand2_1 U28588 ( .A(n23445), .B(n12365), .Y(n23447) );
  sky130_fd_sc_hd__nand3_1 U28589 ( .A(n23447), .B(
        j202_soc_core_j22_cpu_regop_We__1_), .C(n23446), .Y(n23450) );
  sky130_fd_sc_hd__nand2_1 U28590 ( .A(n23520), .B(n29566), .Y(n23449) );
  sky130_fd_sc_hd__nor2_1 U28591 ( .A(n23452), .B(n27651), .Y(n27657) );
  sky130_fd_sc_hd__nand2_1 U28592 ( .A(n27657), .B(n23453), .Y(n27658) );
  sky130_fd_sc_hd__nand2_1 U28593 ( .A(n23455), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_cs_n), .Y(n23457) );
  sky130_fd_sc_hd__nand2_1 U28594 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .B(
        j202_soc_core_wbqspiflash_00_alt_cmd), .Y(n23456) );
  sky130_fd_sc_hd__nor2_1 U28595 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(j202_soc_core_wbqspiflash_00_state[2]), .Y(n26187) );
  sky130_fd_sc_hd__nand2_1 U28596 ( .A(n26187), .B(n25984), .Y(n26049) );
  sky130_fd_sc_hd__nand2_1 U28597 ( .A(n23467), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n25980) );
  sky130_fd_sc_hd__a21oi_1 U28598 ( .A1(n26049), .A2(n25980), .B1(n26042), .Y(
        n23458) );
  sky130_fd_sc_hd__nor2_1 U28599 ( .A(n28080), .B(n26007), .Y(n26053) );
  sky130_fd_sc_hd__nor2_1 U28600 ( .A(n23458), .B(n26053), .Y(n25885) );
  sky130_fd_sc_hd__nand2_1 U28601 ( .A(n26135), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .Y(n28210) );
  sky130_fd_sc_hd__nand2_1 U28602 ( .A(n28210), .B(
        j202_soc_core_wbqspiflash_00_spif_ctrl), .Y(n26141) );
  sky130_fd_sc_hd__nor2_1 U28603 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(n28243), .Y(n25004) );
  sky130_fd_sc_hd__nor2_1 U28604 ( .A(j202_soc_core_wbqspiflash_00_spi_busy), 
        .B(n26255), .Y(n26138) );
  sky130_fd_sc_hd__nand3_1 U28605 ( .A(n25004), .B(n26138), .C(io_out[8]), .Y(
        n25897) );
  sky130_fd_sc_hd__nor2_1 U28606 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(n23467), .Y(n25955) );
  sky130_fd_sc_hd__nand2_1 U28607 ( .A(n28079), .B(n25955), .Y(n26050) );
  sky130_fd_sc_hd__nand2_1 U28608 ( .A(n28230), .B(n28058), .Y(n26013) );
  sky130_fd_sc_hd__nand3_1 U28609 ( .A(n23459), .B(n26131), .C(
        j202_soc_core_wbqspiflash_00_write_in_progress), .Y(n25971) );
  sky130_fd_sc_hd__nor2_1 U28610 ( .A(n25988), .B(n26032), .Y(n26012) );
  sky130_fd_sc_hd__nand2_1 U28611 ( .A(n10958), .B(
        j202_soc_core_ahb2wbqspi_00_stb_o), .Y(n25991) );
  sky130_fd_sc_hd__nor2_1 U28612 ( .A(n26153), .B(n25991), .Y(n26147) );
  sky130_fd_sc_hd__nand2_1 U28613 ( .A(j202_soc_core_qspi_wb_addr[3]), .B(
        j202_soc_core_qspi_wb_addr[2]), .Y(n28222) );
  sky130_fd_sc_hd__nand3_1 U28614 ( .A(n26147), .B(n26148), .C(n28222), .Y(
        n25886) );
  sky130_fd_sc_hd__nand2_1 U28616 ( .A(n26149), .B(n10959), .Y(n28231) );
  sky130_fd_sc_hd__nand2_1 U28617 ( .A(n26147), .B(
        j202_soc_core_qspi_wb_wdat[31]), .Y(n26029) );
  sky130_fd_sc_hd__nand2_1 U28619 ( .A(n26467), .B(n23460), .Y(n23461) );
  sky130_fd_sc_hd__nand3b_1 U28620 ( .A_N(n23462), .B(n28231), .C(n23461), .Y(
        n25938) );
  sky130_fd_sc_hd__a21oi_1 U28621 ( .A1(
        j202_soc_core_wbqspiflash_00_write_in_progress), .A2(n23464), .B1(
        n23463), .Y(n23636) );
  sky130_fd_sc_hd__nand2b_1 U28622 ( .A_N(n26013), .B(n23636), .Y(n23465) );
  sky130_fd_sc_hd__o211ai_1 U28623 ( .A1(n23466), .A2(n25897), .B1(n26050), 
        .C1(n23465), .Y(n26170) );
  sky130_fd_sc_hd__nand2_1 U28624 ( .A(n25880), .B(n25944), .Y(n25921) );
  sky130_fd_sc_hd__nand2_1 U28625 ( .A(io_out[8]), .B(n26116), .Y(n26167) );
  sky130_fd_sc_hd__nor2_1 U28626 ( .A(n23467), .B(n26167), .Y(n23472) );
  sky130_fd_sc_hd__nor2_1 U28627 ( .A(j202_soc_core_wbqspiflash_00_spif_ctrl), 
        .B(n26135), .Y(n26017) );
  sky130_fd_sc_hd__nand2_1 U28628 ( .A(j202_soc_core_wbqspiflash_00_spif_ctrl), 
        .B(j202_soc_core_wbqspiflash_00_spif_cmd), .Y(n25951) );
  sky130_fd_sc_hd__o211ai_1 U28629 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[31]), .B1(n23470), .C1(n23471), 
        .Y(n25891) );
  sky130_fd_sc_hd__a31oi_1 U28630 ( .A1(n26017), .A2(n26171), .A3(n26467), 
        .B1(n23468), .Y(n26041) );
  sky130_fd_sc_hd__nand2_1 U28631 ( .A(n23470), .B(n23469), .Y(n27040) );
  sky130_fd_sc_hd__nand2_1 U28632 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .Y(n28236) );
  sky130_fd_sc_hd__nand3_1 U28633 ( .A(n27040), .B(n23471), .C(n28236), .Y(
        n25958) );
  sky130_fd_sc_hd__nor2_1 U28634 ( .A(j202_soc_core_wbqspiflash_00_spif_cmd), 
        .B(n26134), .Y(n28237) );
  sky130_fd_sc_hd__nand2_1 U28635 ( .A(n28237), .B(n27040), .Y(n25890) );
  sky130_fd_sc_hd__nand3_1 U28636 ( .A(n26041), .B(n25958), .C(n25890), .Y(
        n26164) );
  sky130_fd_sc_hd__a21oi_1 U28637 ( .A1(n23472), .A2(n26164), .B1(n26138), .Y(
        n23474) );
  sky130_fd_sc_hd__a21oi_1 U28638 ( .A1(n23474), .A2(n25024), .B1(n23473), .Y(
        n23478) );
  sky130_fd_sc_hd__nand2_1 U28639 ( .A(n25916), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n25961) );
  sky130_fd_sc_hd__nor2_1 U28640 ( .A(n26035), .B(n25961), .Y(n26194) );
  sky130_fd_sc_hd__nand3_1 U28641 ( .A(n25949), .B(
        j202_soc_core_qspi_wb_addr[24]), .C(n10959), .Y(n23475) );
  sky130_fd_sc_hd__nand3_1 U28642 ( .A(n27037), .B(n23476), .C(n23475), .Y(
        n25924) );
  sky130_fd_sc_hd__nand2_1 U28643 ( .A(n26009), .B(n28080), .Y(n25884) );
  sky130_fd_sc_hd__nand2_1 U28644 ( .A(n25924), .B(n25884), .Y(n26169) );
  sky130_fd_sc_hd__nor2_1 U28645 ( .A(n26194), .B(n26169), .Y(n23477) );
  sky130_fd_sc_hd__nand2b_1 U28646 ( .A_N(n23478), .B(n23477), .Y(n23640) );
  sky130_fd_sc_hd__nor4_1 U28647 ( .A(n26185), .B(n23479), .C(n26170), .D(
        n23640), .Y(n23480) );
  sky130_fd_sc_hd__nor2_2 U28648 ( .A(n28590), .B(n23480), .Y(n29361) );
  sky130_fd_sc_hd__nor2_1 U28649 ( .A(n28590), .B(n23485), .Y(n23699) );
  sky130_fd_sc_hd__nor2_1 U28650 ( .A(j202_soc_core_j22_cpu_regop_We__2_), .B(
        n14849), .Y(n23508) );
  sky130_fd_sc_hd__nand2b_1 U28651 ( .A_N(n23558), .B(
        j202_soc_core_j22_cpu_regop_We__1_), .Y(n23482) );
  sky130_fd_sc_hd__nand3_1 U28652 ( .A(n26812), .B(
        j202_soc_core_j22_cpu_regop_We__2_), .C(n23481), .Y(n23556) );
  sky130_fd_sc_hd__nand2b_1 U28653 ( .A_N(n23556), .B(
        j202_soc_core_j22_cpu_regop_We__3_), .Y(n24643) );
  sky130_fd_sc_hd__nand2_1 U28654 ( .A(n23482), .B(n24643), .Y(n23703) );
  sky130_fd_sc_hd__o22ai_1 U28655 ( .A1(n24291), .A2(n26897), .B1(n23483), 
        .B2(n23703), .Y(n23492) );
  sky130_fd_sc_hd__nor2_1 U28656 ( .A(j202_soc_core_j22_cpu_rte4), .B(n23485), 
        .Y(n23486) );
  sky130_fd_sc_hd__nand2_1 U28657 ( .A(n23487), .B(n23486), .Y(n23489) );
  sky130_fd_sc_hd__nor2_1 U28658 ( .A(n23489), .B(n23488), .Y(n23491) );
  sky130_fd_sc_hd__nand3_1 U28659 ( .A(n24471), .B(n23491), .C(n24468), .Y(
        n23704) );
  sky130_fd_sc_hd__nand4_1 U28660 ( .A(n24291), .B(n23493), .C(
        j202_soc_core_j22_cpu_regop_M_Rn__3_), .D(n23534), .Y(n23543) );
  sky130_fd_sc_hd__nand2_1 U28661 ( .A(n23494), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__0_), .Y(n23540) );
  sky130_fd_sc_hd__nand2_1 U28662 ( .A(n23174), .B(n23496), .Y(n23498) );
  sky130_fd_sc_hd__nand2_1 U28663 ( .A(n23520), .B(n11160), .Y(n23497) );
  sky130_fd_sc_hd__a21o_2 U28664 ( .A1(n23498), .A2(n23497), .B1(n14849), .X(
        n27222) );
  sky130_fd_sc_hd__nand2_1 U28665 ( .A(n23499), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__1_), .Y(n23539) );
  sky130_fd_sc_hd__nand2_1 U28666 ( .A(n23174), .B(n23501), .Y(n23504) );
  sky130_fd_sc_hd__nand2_1 U28667 ( .A(n23520), .B(n23502), .Y(n23503) );
  sky130_fd_sc_hd__a21o_2 U28668 ( .A1(n23504), .A2(n23503), .B1(n14849), .X(
        n27210) );
  sky130_fd_sc_hd__nor2_1 U28669 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__1_), 
        .B(j202_soc_core_j22_cpu_regop_M_Wm__2_), .Y(n24428) );
  sky130_fd_sc_hd__nand2_1 U28670 ( .A(n24428), .B(n23505), .Y(n23506) );
  sky130_fd_sc_hd__nor3_1 U28671 ( .A(n23507), .B(n23506), .C(n24113), .Y(
        n23943) );
  sky130_fd_sc_hd__nand3_1 U28672 ( .A(n23508), .B(
        j202_soc_core_j22_cpu_regop_We__3_), .C(
        j202_soc_core_j22_cpu_regop_We__1_), .Y(n23856) );
  sky130_fd_sc_hd__nand2_1 U28673 ( .A(n23174), .B(n23510), .Y(n23512) );
  sky130_fd_sc_hd__nand2_1 U28674 ( .A(n23520), .B(n15983), .Y(n23511) );
  sky130_fd_sc_hd__nand3_1 U28675 ( .A(n24291), .B(n23535), .C(
        j202_soc_core_j22_cpu_regop_M_Rn__2_), .Y(n23542) );
  sky130_fd_sc_hd__nand2_1 U28676 ( .A(n23174), .B(n23514), .Y(n23517) );
  sky130_fd_sc_hd__nand2_1 U28677 ( .A(n23520), .B(n23515), .Y(n23516) );
  sky130_fd_sc_hd__o21ai_2 U28678 ( .A1(n23539), .A2(n23542), .B1(n27214), .Y(
        j202_soc_core_j22_cpu_rf_N2931) );
  sky130_fd_sc_hd__nand2_1 U28679 ( .A(n23174), .B(n23519), .Y(n23522) );
  sky130_fd_sc_hd__nand2_1 U28680 ( .A(n23520), .B(n16493), .Y(n23521) );
  sky130_fd_sc_hd__o21ai_2 U28681 ( .A1(n23541), .A2(n23542), .B1(n27224), .Y(
        j202_soc_core_j22_cpu_rf_N2968) );
  sky130_fd_sc_hd__nand2b_1 U28682 ( .A_N(n23558), .B(n23529), .Y(n23530) );
  sky130_fd_sc_hd__nand3_1 U28683 ( .A(n24291), .B(n23535), .C(n23534), .Y(
        n23538) );
  sky130_fd_sc_hd__o21ai_2 U28684 ( .A1(n23542), .A2(n23540), .B1(n27220), .Y(
        j202_soc_core_j22_cpu_rf_N2894) );
  sky130_fd_sc_hd__o21ai_2 U28685 ( .A1(n23544), .A2(n23542), .B1(n27216), .Y(
        j202_soc_core_j22_cpu_rf_N2857) );
  sky130_fd_sc_hd__o21ai_2 U28686 ( .A1(n23544), .A2(n23543), .B1(n27218), .Y(
        j202_soc_core_j22_cpu_rf_N3005) );
  sky130_fd_sc_hd__nand3_1 U28687 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[2]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_sck), .C(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .Y(n23545) );
  sky130_fd_sc_hd__nand2_1 U28688 ( .A(n26202), .B(n25010), .Y(n28646) );
  sky130_fd_sc_hd__nor2_1 U28689 ( .A(j202_soc_core_wbqspiflash_00_w_qspi_sck), 
        .B(n28646), .Y(n28640) );
  sky130_fd_sc_hd__nor2_1 U28690 ( .A(j202_soc_core_wbqspiflash_00_w_qspi_sck), 
        .B(n26202), .Y(n26199) );
  sky130_fd_sc_hd__nand2_1 U28691 ( .A(n26225), .B(n24575), .Y(n26200) );
  sky130_fd_sc_hd__nor2_1 U28692 ( .A(n29033), .B(n29061), .Y(n25106) );
  sky130_fd_sc_hd__o21a_1 U28693 ( .A1(n23563), .A2(n25106), .B1(n11936), .X(
        n23561) );
  sky130_fd_sc_hd__nor2b_1 U28694 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[29]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N32) );
  sky130_fd_sc_hd__nor2b_1 U28695 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[16]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N19) );
  sky130_fd_sc_hd__nor2b_1 U28696 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[24]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N27) );
  sky130_fd_sc_hd__nor2b_1 U28697 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[17]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N20) );
  sky130_fd_sc_hd__nor2b_1 U28698 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[3]), .A(n28590), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N6) );
  sky130_fd_sc_hd__nor2b_1 U28699 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[28]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N31) );
  sky130_fd_sc_hd__nand3_1 U28700 ( .A(n28281), .B(
        j202_soc_core_uart_TOP_tx_fifo_wp[0]), .C(j202_soc_core_uart_WRTXD1), 
        .Y(n24695) );
  sky130_fd_sc_hd__nor2_1 U28701 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[1]), 
        .B(n24695), .Y(n29352) );
  sky130_fd_sc_hd__nand2_1 U28702 ( .A(n28229), .B(
        j202_soc_core_wbqspiflash_00_state[3]), .Y(n25901) );
  sky130_fd_sc_hd__nor2_1 U28703 ( .A(n25984), .B(n25901), .Y(n26191) );
  sky130_fd_sc_hd__nand2_1 U28704 ( .A(n26191), .B(
        j202_soc_core_wbqspiflash_00_state[4]), .Y(n28187) );
  sky130_fd_sc_hd__nand2_1 U28705 ( .A(n28187), .B(n29594), .Y(
        j202_soc_core_wbqspiflash_00_N710) );
  sky130_fd_sc_hd__nand2_1 U28706 ( .A(n27334), .B(n23548), .Y(
        j202_soc_core_j22_cpu_rf_N2627) );
  sky130_fd_sc_hd__nand2_1 U28707 ( .A(n28969), .B(n29594), .Y(n23549) );
  sky130_fd_sc_hd__nor2b_1 U28708 ( .B_N(j202_soc_core_prdata[2]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N130) );
  sky130_fd_sc_hd__nor2b_1 U28709 ( .B_N(j202_soc_core_prdata[11]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N139) );
  sky130_fd_sc_hd__nor2b_1 U28710 ( .B_N(j202_soc_core_prdata[13]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N141) );
  sky130_fd_sc_hd__nor2b_1 U28711 ( .B_N(j202_soc_core_prdata[3]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N131) );
  sky130_fd_sc_hd__nor2b_1 U28712 ( .B_N(j202_soc_core_prdata[5]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N133) );
  sky130_fd_sc_hd__nor2b_1 U28713 ( .B_N(j202_soc_core_prdata[4]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N132) );
  sky130_fd_sc_hd__nor2b_1 U28714 ( .B_N(j202_soc_core_prdata[8]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N136) );
  sky130_fd_sc_hd__nor2b_1 U28715 ( .B_N(j202_soc_core_prdata[15]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N143) );
  sky130_fd_sc_hd__nor2b_1 U28716 ( .B_N(j202_soc_core_prdata[1]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N129) );
  sky130_fd_sc_hd__nor2b_1 U28717 ( .B_N(j202_soc_core_prdata[9]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N137) );
  sky130_fd_sc_hd__nor2b_1 U28718 ( .B_N(j202_soc_core_prdata[6]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N134) );
  sky130_fd_sc_hd__nor2b_1 U28719 ( .B_N(j202_soc_core_prdata[14]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N142) );
  sky130_fd_sc_hd__nor2b_1 U28720 ( .B_N(j202_soc_core_prdata[12]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N140) );
  sky130_fd_sc_hd__nor2b_1 U28721 ( .B_N(j202_soc_core_prdata[7]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N135) );
  sky130_fd_sc_hd__nor2b_1 U28722 ( .B_N(j202_soc_core_prdata[0]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N128) );
  sky130_fd_sc_hd__nor2b_1 U28723 ( .B_N(j202_soc_core_prdata[10]), .A(n23549), 
        .Y(j202_soc_core_ahb2apb_00_N138) );
  sky130_fd_sc_hd__nand2_1 U28724 ( .A(n12200), .B(n29594), .Y(n10562) );
  sky130_fd_sc_hd__nand2_1 U28725 ( .A(n23555), .B(n12366), .Y(n23557) );
  sky130_fd_sc_hd__nand2_1 U28726 ( .A(n12365), .B(
        j202_soc_core_j22_cpu_regop_We__1_), .Y(n23559) );
  sky130_fd_sc_hd__nor2_1 U28727 ( .A(n29033), .B(n27622), .Y(n23562) );
  sky130_fd_sc_hd__inv_1 U28728 ( .A(n23565), .Y(n23567) );
  sky130_fd_sc_hd__nor2_1 U28729 ( .A(n23567), .B(n23566), .Y(n24460) );
  sky130_fd_sc_hd__nand2_1 U28730 ( .A(n23821), .B(n29036), .Y(n23568) );
  sky130_fd_sc_hd__nand2_1 U28731 ( .A(n24294), .B(n23568), .Y(n23569) );
  sky130_fd_sc_hd__nand2_1 U28732 ( .A(n23603), .B(n12595), .Y(n23570) );
  sky130_fd_sc_hd__nor2_1 U28733 ( .A(n23820), .B(n27924), .Y(n23571) );
  sky130_fd_sc_hd__nand2_1 U28734 ( .A(n12729), .B(n12731), .Y(n24309) );
  sky130_fd_sc_hd__nand4_1 U28735 ( .A(n24460), .B(n27788), .C(n23571), .D(
        n24309), .Y(n23572) );
  sky130_fd_sc_hd__o2bb2ai_1 U28736 ( .B1(n23859), .B2(n27956), .A1_N(n27980), 
        .A2_N(n23572), .Y(n10504) );
  sky130_fd_sc_hd__nor2_1 U28738 ( .A(n23574), .B(n23573), .Y(n23577) );
  sky130_fd_sc_hd__o21a_1 U28739 ( .A1(n23577), .A2(n29033), .B1(n23576), .X(
        n24117) );
  sky130_fd_sc_hd__a21o_1 U28740 ( .A1(n29033), .A2(n29061), .B1(n24117), .X(
        n23578) );
  sky130_fd_sc_hd__nor2_1 U28741 ( .A(n29061), .B(n29559), .Y(n23580) );
  sky130_fd_sc_hd__nand2_1 U28742 ( .A(n11798), .B(n23586), .Y(n23587) );
  sky130_fd_sc_hd__nor2_1 U28743 ( .A(n23587), .B(n12658), .Y(n23588) );
  sky130_fd_sc_hd__nor2_1 U28744 ( .A(n23588), .B(n27561), .Y(n24345) );
  sky130_fd_sc_hd__a21oi_1 U28745 ( .A1(n24257), .A2(n12475), .B1(n27688), .Y(
        n23593) );
  sky130_fd_sc_hd__nand2_1 U28746 ( .A(n27550), .B(n27892), .Y(n23591) );
  sky130_fd_sc_hd__nor3_1 U28747 ( .A(n23589), .B(n12060), .C(n24357), .Y(
        n23590) );
  sky130_fd_sc_hd__nor2_1 U28748 ( .A(n23591), .B(n23590), .Y(n23592) );
  sky130_fd_sc_hd__nand4_1 U28749 ( .A(n11048), .B(n24345), .C(n23593), .D(
        n23592), .Y(n23594) );
  sky130_fd_sc_hd__o2bb2ai_1 U28750 ( .B1(n27175), .B2(n23595), .A1_N(n27980), 
        .A2_N(n23594), .Y(n10598) );
  sky130_fd_sc_hd__nand4b_1 U28751 ( .A_N(n23598), .B(n23957), .C(n23597), .D(
        n23596), .Y(n23857) );
  sky130_fd_sc_hd__nand2_1 U28752 ( .A(n11873), .B(n23599), .Y(n23600) );
  sky130_fd_sc_hd__nand2_1 U28753 ( .A(n12436), .B(n23600), .Y(n23601) );
  sky130_fd_sc_hd__nand2_1 U28754 ( .A(n12436), .B(n24094), .Y(n24336) );
  sky130_fd_sc_hd__nand2_1 U28755 ( .A(n23604), .B(n24265), .Y(n27786) );
  sky130_fd_sc_hd__nand2_1 U28756 ( .A(n23604), .B(n12150), .Y(n27781) );
  sky130_fd_sc_hd__nand2_1 U28757 ( .A(n27786), .B(n27781), .Y(n23610) );
  sky130_fd_sc_hd__nand2b_1 U28758 ( .A_N(n24353), .B(n29569), .Y(n27787) );
  sky130_fd_sc_hd__nand4_1 U28759 ( .A(n27782), .B(n27772), .C(n27787), .D(
        n23605), .Y(n23609) );
  sky130_fd_sc_hd__nor3_1 U28760 ( .A(n23610), .B(n23609), .C(n27875), .Y(
        n23612) );
  sky130_fd_sc_hd__nand3_1 U28761 ( .A(n23612), .B(n27794), .C(n27785), .Y(
        n23613) );
  sky130_fd_sc_hd__o2bb2ai_1 U28762 ( .B1(n23614), .B2(n27956), .A1_N(n27980), 
        .A2_N(n23613), .Y(n10592) );
  sky130_fd_sc_hd__nand2_1 U28763 ( .A(j202_soc_core_uart_TOP_load), .B(
        j202_soc_core_uart_sio_ce), .Y(n28776) );
  sky130_fd_sc_hd__nor2b_1 U28764 ( .B_N(j202_soc_core_uart_TOP_hold_reg[1]), 
        .A(n28003), .Y(j202_soc_core_uart_TOP_N25) );
  sky130_fd_sc_hd__nor2b_1 U28765 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[1]), .A(n28590), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N4) );
  sky130_fd_sc_hd__nor2b_1 U28766 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[0]), .A(n28590), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N3) );
  sky130_fd_sc_hd__nor2b_1 U28767 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[5]), .A(n28590), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N8) );
  sky130_fd_sc_hd__nor2b_1 U28768 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[2]), .A(n28590), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N5) );
  sky130_fd_sc_hd__nor2b_1 U28769 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[23]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N26) );
  sky130_fd_sc_hd__nor2b_1 U28770 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[6]), .A(n28590), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N9) );
  sky130_fd_sc_hd__nor2b_1 U28771 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[12]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N15) );
  sky130_fd_sc_hd__nor2b_1 U28772 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[30]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N33) );
  sky130_fd_sc_hd__nor2b_1 U28773 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[7]), .A(n28590), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N10) );
  sky130_fd_sc_hd__nor2b_1 U28774 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[20]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N23) );
  sky130_fd_sc_hd__nor2b_1 U28775 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[21]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N24) );
  sky130_fd_sc_hd__nor2b_1 U28776 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[8]), .A(n28590), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N11) );
  sky130_fd_sc_hd__nor2b_1 U28777 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[9]), .A(n28590), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N12) );
  sky130_fd_sc_hd__nor2b_1 U28778 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[10]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N13) );
  sky130_fd_sc_hd__nor2b_1 U28779 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[14]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N17) );
  sky130_fd_sc_hd__nor2b_1 U28780 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[18]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N21) );
  sky130_fd_sc_hd__nor2b_1 U28781 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[15]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N18) );
  sky130_fd_sc_hd__nor2b_1 U28782 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[19]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N22) );
  sky130_fd_sc_hd__nor2b_1 U28783 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[26]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N29) );
  sky130_fd_sc_hd__nor2b_1 U28784 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[13]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N16) );
  sky130_fd_sc_hd__nor2b_1 U28785 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[25]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N28) );
  sky130_fd_sc_hd__nor2b_1 U28786 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[4]), .A(n28590), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N7) );
  sky130_fd_sc_hd__nor2b_1 U28787 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[22]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N25) );
  sky130_fd_sc_hd__nor2b_1 U28788 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[27]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N30) );
  sky130_fd_sc_hd__nor2b_1 U28789 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[31]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N34) );
  sky130_fd_sc_hd__nor2b_1 U28790 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[11]), .A(n28590), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N14) );
  sky130_fd_sc_hd__nor2_1 U28791 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[28]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n23616) );
  sky130_fd_sc_hd__nor2_1 U28792 ( .A(n28901), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[25]), .Y(n23615) );
  sky130_fd_sc_hd__nor2_1 U28793 ( .A(n23616), .B(n23615), .Y(n23882) );
  sky130_fd_sc_hd__a2bb2oi_1 U28794 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23617), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[27]), .Y(n23883) );
  sky130_fd_sc_hd__a2bb2oi_1 U28795 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23618), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[26]), .Y(n23884) );
  sky130_fd_sc_hd__a2bb2oi_1 U28796 ( .B1(n28901), .B2(n23618), .A1_N(n28901), 
        .A2_N(j202_soc_core_wbqspiflash_00_lldriver_r_input[20]), .Y(n23900)
         );
  sky130_fd_sc_hd__a2bb2oi_1 U28797 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23630), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[22]), .Y(n23887) );
  sky130_fd_sc_hd__a2bb2oi_1 U28798 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23619), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[3]), .Y(n23899) );
  sky130_fd_sc_hd__a2bb2oi_1 U28799 ( .B1(n28901), .B2(n23622), .A1_N(n28901), 
        .A2_N(j202_soc_core_wbqspiflash_00_lldriver_r_input[18]), .Y(n23901)
         );
  sky130_fd_sc_hd__nor2_1 U28800 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[29]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n23621) );
  sky130_fd_sc_hd__nor2_1 U28801 ( .A(n28901), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[26]), .Y(n23620) );
  sky130_fd_sc_hd__nor2_1 U28802 ( .A(n23621), .B(n23620), .Y(n23881) );
  sky130_fd_sc_hd__a2bb2oi_1 U28803 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23622), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[24]), .Y(n23886) );
  sky130_fd_sc_hd__a2bb2oi_1 U28804 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23623), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[10]), .Y(n23894) );
  sky130_fd_sc_hd__a2bb2oi_1 U28805 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23629), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[18]), .Y(n23889) );
  sky130_fd_sc_hd__a2bb2oi_1 U28806 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23624), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[11]), .Y(n23893) );
  sky130_fd_sc_hd__a2bb2oi_1 U28807 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23625), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[4]), .Y(n23898) );
  sky130_fd_sc_hd__a2bb2oi_1 U28808 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23626), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[20]), .Y(n23888) );
  sky130_fd_sc_hd__a2bb2oi_1 U28809 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23635), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[17]), .Y(n23890) );
  sky130_fd_sc_hd__a2bb2oi_1 U28810 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23632), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[16]), .Y(n23891) );
  sky130_fd_sc_hd__a2bb2oi_1 U28811 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23627), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[25]), .Y(n23885) );
  sky130_fd_sc_hd__a2bb2oi_1 U28812 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23628), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[7]), .Y(n23897) );
  sky130_fd_sc_hd__a2bb2oi_1 U28813 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23631), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[8]), .Y(n23896) );
  sky130_fd_sc_hd__a2bb2oi_1 U28814 ( .B1(n28901), .B2(n23629), .A1_N(n28901), 
        .A2_N(j202_soc_core_wbqspiflash_00_lldriver_r_input[12]), .Y(n23903)
         );
  sky130_fd_sc_hd__a2bb2oi_1 U28815 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23633), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[9]), .Y(n23895) );
  sky130_fd_sc_hd__a2bb2oi_1 U28816 ( .B1(n28901), .B2(n23630), .A1_N(n28901), 
        .A2_N(j202_soc_core_wbqspiflash_00_lldriver_r_input[16]), .Y(n23902)
         );
  sky130_fd_sc_hd__a2bb2oi_1 U28817 ( .B1(n28901), .B2(n23631), .A1_N(n28901), 
        .A2_N(j202_soc_core_wbqspiflash_00_lldriver_r_input[2]), .Y(n23908) );
  sky130_fd_sc_hd__a2bb2oi_1 U28818 ( .B1(n28901), .B2(n23632), .A1_N(n28901), 
        .A2_N(j202_soc_core_wbqspiflash_00_lldriver_r_input[10]), .Y(n23905)
         );
  sky130_fd_sc_hd__a2bb2oi_1 U28819 ( .B1(n28901), .B2(n23633), .A1_N(n28901), 
        .A2_N(j202_soc_core_wbqspiflash_00_lldriver_r_input[3]), .Y(n23906) );
  sky130_fd_sc_hd__a2bb2oi_1 U28820 ( .B1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B2(n23634), .A1_N(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2_N(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[12]), .Y(n23892) );
  sky130_fd_sc_hd__a2bb2oi_1 U28821 ( .B1(n28901), .B2(n23635), .A1_N(n28901), 
        .A2_N(j202_soc_core_wbqspiflash_00_lldriver_r_input[11]), .Y(n23904)
         );
  sky130_fd_sc_hd__nand2_1 U28822 ( .A(n26161), .B(n28058), .Y(n26254) );
  sky130_fd_sc_hd__nand2_1 U28823 ( .A(n26254), .B(n25954), .Y(n23638) );
  sky130_fd_sc_hd__a21oi_1 U28825 ( .A1(n23638), .A2(n23637), .B1(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n23642) );
  sky130_fd_sc_hd__nor2_1 U28826 ( .A(n28080), .B(n23638), .Y(n23639) );
  sky130_fd_sc_hd__nand2_1 U28827 ( .A(n26119), .B(n25926), .Y(n28096) );
  sky130_fd_sc_hd__or4_1 U28828 ( .A(n28968), .B(n23639), .C(n26191), .D(
        n26192), .X(n23641) );
  sky130_fd_sc_hd__or3_1 U28829 ( .A(n23642), .B(n23641), .C(n23640), .X(
        j202_soc_core_wbqspiflash_00_N735) );
  sky130_fd_sc_hd__o2bb2ai_1 U28830 ( .B1(n28730), .B2(n28723), .A1_N(n28733), 
        .A2_N(j202_soc_core_wbqspiflash_00_lldriver_r_word[29]), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N317) );
  sky130_fd_sc_hd__nor2_1 U28831 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[1]), 
        .B(n28623), .Y(n27996) );
  sky130_fd_sc_hd__nor2b_1 U28832 ( .B_N(j202_soc_core_uart_TOP_rx_bit_cnt[3]), 
        .A(j202_soc_core_uart_TOP_rx_bit_cnt[2]), .Y(n28624) );
  sky130_fd_sc_hd__nand2_1 U28833 ( .A(j202_soc_core_cmt_core_00_str0), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[0]), .Y(n24823) );
  sky130_fd_sc_hd__nor2_1 U28834 ( .A(n24824), .B(n24823), .Y(n24825) );
  sky130_fd_sc_hd__nand2_1 U28835 ( .A(n24825), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[2]), .Y(n24828) );
  sky130_fd_sc_hd__nand2b_1 U28836 ( .A_N(n24828), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[3]), .Y(n24831) );
  sky130_fd_sc_hd__nor2_1 U28837 ( .A(n24832), .B(n24831), .Y(n24830) );
  sky130_fd_sc_hd__nand3_1 U28838 ( .A(n23643), .B(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[1]), .C(
        j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_2), .Y(n23669) );
  sky130_fd_sc_hd__nand3_1 U28839 ( .A(n23646), .B(n23645), .C(n23644), .Y(
        n23668) );
  sky130_fd_sc_hd__nor2_1 U28840 ( .A(j202_soc_core_cmt_core_00_reg_addr[4]), 
        .B(j202_soc_core_cmt_core_00_reg_addr[5]), .Y(n23647) );
  sky130_fd_sc_hd__nand3_1 U28841 ( .A(n23648), .B(n23647), .C(n23666), .Y(
        n24951) );
  sky130_fd_sc_hd__nor2_1 U28842 ( .A(n23669), .B(n24951), .Y(n24843) );
  sky130_fd_sc_hd__nand2_1 U28843 ( .A(j202_soc_core_cmt_core_00_reg_addr[3]), 
        .B(j202_soc_core_cmt_core_00_reg_addr[2]), .Y(n24960) );
  sky130_fd_sc_hd__nand2_1 U28844 ( .A(n24843), .B(n23649), .Y(n27473) );
  sky130_fd_sc_hd__a22oi_1 U28845 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[3]), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[7]), .B1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[5]), .B2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[9]), .Y(n23655) );
  sky130_fd_sc_hd__o21ai_1 U28846 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[7]), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[3]), .B1(
        j202_soc_core_cmt_core_00_cks0[0]), .Y(n23654) );
  sky130_fd_sc_hd__nand3_1 U28847 ( .A(n23651), .B(n23650), .C(
        j202_soc_core_cmt_core_00_cks0[1]), .Y(n23653) );
  sky130_fd_sc_hd__and4_1 U28849 ( .A(n23655), .B(n23654), .C(n23653), .D(
        n23652), .X(n23662) );
  sky130_fd_sc_hd__nand2_1 U28850 ( .A(n23656), .B(n24832), .Y(n23657) );
  sky130_fd_sc_hd__nor3_1 U28851 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[0]), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[1]), .C(n23657), .Y(
        n23661) );
  sky130_fd_sc_hd__nor2_1 U28852 ( .A(j202_soc_core_cmt_core_00_cks0[1]), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[5]), .Y(n23659) );
  sky130_fd_sc_hd__nand2_1 U28853 ( .A(n24833), .B(n24839), .Y(n23658) );
  sky130_fd_sc_hd__a21oi_1 U28854 ( .A1(n23659), .A2(n24829), .B1(n23658), .Y(
        n23660) );
  sky130_fd_sc_hd__nand3_1 U28855 ( .A(n23662), .B(n23661), .C(n23660), .Y(
        n24874) );
  sky130_fd_sc_hd__nand2_1 U28856 ( .A(n27473), .B(n24874), .Y(n26284) );
  sky130_fd_sc_hd__nand2_1 U28857 ( .A(n24830), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[5]), .Y(n24834) );
  sky130_fd_sc_hd__o211a_2 U28858 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[5]), .A2(n24830), .B1(
        n28619), .C1(n24834), .X(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[5]) );
  sky130_fd_sc_hd__nor2_1 U28859 ( .A(n24833), .B(n24834), .Y(n24836) );
  sky130_fd_sc_hd__nand2_1 U28860 ( .A(n24836), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[7]), .Y(n24838) );
  sky130_fd_sc_hd__o211a_2 U28861 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[7]), .A2(n24836), .B1(
        n28619), .C1(n24838), .X(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[7]) );
  sky130_fd_sc_hd__nand2_1 U28862 ( .A(n27138), .B(n27135), .Y(n27132) );
  sky130_fd_sc_hd__nor2_1 U28863 ( .A(j202_soc_core_uart_TOP_rx_fifo_wp[1]), 
        .B(n27132), .Y(n29350) );
  sky130_fd_sc_hd__nor2_1 U28864 ( .A(n27134), .B(n27132), .Y(n29349) );
  sky130_fd_sc_hd__nor2_1 U28865 ( .A(j202_soc_core_uart_TOP_rx_fifo_wp[1]), 
        .B(n27133), .Y(n29351) );
  sky130_fd_sc_hd__nand3_1 U28866 ( .A(n28281), .B(j202_soc_core_uart_WRTXD1), 
        .C(n24694), .Y(n23663) );
  sky130_fd_sc_hd__nor2_1 U28867 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[1]), 
        .B(n23663), .Y(n29345) );
  sky130_fd_sc_hd__nor2_1 U28868 ( .A(n23664), .B(n23663), .Y(n29344) );
  sky130_fd_sc_hd__nor2_1 U28869 ( .A(n23664), .B(n24695), .Y(n29346) );
  sky130_fd_sc_hd__nand2_1 U28870 ( .A(j202_soc_core_cmt_core_00_str1), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[0]), .Y(n24885) );
  sky130_fd_sc_hd__nor2_1 U28871 ( .A(n24886), .B(n24885), .Y(n24887) );
  sky130_fd_sc_hd__nand2_1 U28872 ( .A(n24887), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[2]), .Y(n24890) );
  sky130_fd_sc_hd__nor2_1 U28873 ( .A(n24891), .B(n24890), .Y(n24889) );
  sky130_fd_sc_hd__nand2_1 U28874 ( .A(n24889), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[4]), .Y(n24893) );
  sky130_fd_sc_hd__nor2_1 U28875 ( .A(n24894), .B(n24893), .Y(n24892) );
  sky130_fd_sc_hd__nand2_1 U28876 ( .A(n24892), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[6]), .Y(n24899) );
  sky130_fd_sc_hd__nor2_1 U28877 ( .A(n24900), .B(n24899), .Y(n24898) );
  sky130_fd_sc_hd__nand3_1 U28878 ( .A(n23666), .B(n23665), .C(
        j202_soc_core_cmt_core_00_reg_addr[4]), .Y(n23667) );
  sky130_fd_sc_hd__nor2_1 U28879 ( .A(n23668), .B(n23667), .Y(n24955) );
  sky130_fd_sc_hd__nor2_1 U28880 ( .A(j202_soc_core_cmt_core_00_reg_addr[3]), 
        .B(j202_soc_core_cmt_core_00_reg_addr[2]), .Y(n24954) );
  sky130_fd_sc_hd__nand3_1 U28881 ( .A(n24955), .B(n24896), .C(n24954), .Y(
        n27491) );
  sky130_fd_sc_hd__nand2_1 U28882 ( .A(n24902), .B(
        j202_soc_core_cmt_core_00_cks1[0]), .Y(n23670) );
  sky130_fd_sc_hd__nand2_1 U28883 ( .A(n23670), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[5]), .Y(n23674) );
  sky130_fd_sc_hd__nand2_1 U28884 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[3]), .B(
        j202_soc_core_cmt_core_00_cks1[0]), .Y(n23673) );
  sky130_fd_sc_hd__nand2_1 U28885 ( .A(n23671), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[9]), .Y(n23672) );
  sky130_fd_sc_hd__and3_1 U28886 ( .A(n23674), .B(n23673), .C(n23672), .X(
        n23684) );
  sky130_fd_sc_hd__nor2_1 U28888 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[2]), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[6]), .Y(n23677) );
  sky130_fd_sc_hd__nor2_1 U28889 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[0]), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[1]), .Y(n23676) );
  sky130_fd_sc_hd__nor2_1 U28890 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[4]), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[8]), .Y(n23675) );
  sky130_fd_sc_hd__and4_1 U28891 ( .A(n23678), .B(n23677), .C(n23676), .D(
        n23675), .X(n23683) );
  sky130_fd_sc_hd__nand3_1 U28892 ( .A(n23679), .B(n24894), .C(n24891), .Y(
        n23681) );
  sky130_fd_sc_hd__nand3_1 U28893 ( .A(n24900), .B(n24902), .C(
        j202_soc_core_cmt_core_00_cks1[1]), .Y(n23680) );
  sky130_fd_sc_hd__nand3_1 U28894 ( .A(n23684), .B(n23683), .C(n23682), .Y(
        n24905) );
  sky130_fd_sc_hd__nand2_1 U28895 ( .A(n27491), .B(n24905), .Y(n26300) );
  sky130_fd_sc_hd__nand2_1 U28896 ( .A(n24898), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[8]), .Y(n24901) );
  sky130_fd_sc_hd__o211a_2 U28897 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[8]), .A2(n24898), .B1(
        n28622), .C1(n24901), .X(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[8]) );
  sky130_fd_sc_hd__nor2_1 U28898 ( .A(n28623), .B(n23685), .Y(n23686) );
  sky130_fd_sc_hd__nor2_1 U28899 ( .A(n28590), .B(n28000), .Y(n23911) );
  sky130_fd_sc_hd__nand2_1 U28900 ( .A(n23686), .B(
        j202_soc_core_uart_TOP_rx_bit_cnt[2]), .Y(n27998) );
  sky130_fd_sc_hd__o211a_2 U28901 ( .A1(j202_soc_core_uart_TOP_rx_bit_cnt[2]), 
        .A2(n23686), .B1(n23911), .C1(n27998), .X(j202_soc_core_uart_TOP_N88)
         );
  sky130_fd_sc_hd__nand2_1 U28902 ( .A(n25954), .B(n26188), .Y(n26022) );
  sky130_fd_sc_hd__nor2_1 U28903 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(n26022), .Y(n28199) );
  sky130_fd_sc_hd__nand2_1 U28904 ( .A(n25916), .B(
        j202_soc_core_wbqspiflash_00_state[4]), .Y(n26174) );
  sky130_fd_sc_hd__nor3_1 U28905 ( .A(j202_soc_core_wbqspiflash_00_spi_out[0]), 
        .B(n26476), .C(n25980), .Y(n23687) );
  sky130_fd_sc_hd__nand2b_1 U28906 ( .A_N(n26174), .B(n23687), .Y(n26248) );
  sky130_fd_sc_hd__a21oi_1 U28908 ( .A1(n26116), .A2(n28199), .B1(n23688), .Y(
        n25941) );
  sky130_fd_sc_hd__nand2_1 U28909 ( .A(n25982), .B(
        j202_soc_core_wbqspiflash_00_spi_valid), .Y(n23689) );
  sky130_fd_sc_hd__a21oi_1 U28910 ( .A1(n25941), .A2(n23689), .B1(n28590), .Y(
        n29358) );
  sky130_fd_sc_hd__nand2_1 U28911 ( .A(n23691), .B(n29594), .Y(
        j202_soc_core_ahb2apb_00_N127) );
  sky130_fd_sc_hd__nand2_1 U28912 ( .A(n14849), .B(n29594), .Y(n10565) );
  sky130_fd_sc_hd__nand2_1 U28913 ( .A(n23692), .B(n27176), .Y(n10563) );
  sky130_fd_sc_hd__nand2_1 U28914 ( .A(n27360), .B(n11157), .Y(n23709) );
  sky130_fd_sc_hd__o22a_1 U28915 ( .A1(n23704), .A2(n23703), .B1(n23702), .B2(
        n23705), .X(n23784) );
  sky130_fd_sc_hd__a22oi_1 U28916 ( .A1(n23794), .A2(n27361), .B1(n26895), 
        .B2(n25329), .Y(n23708) );
  sky130_fd_sc_hd__nand2_1 U28917 ( .A(n25316), .B(n24593), .Y(n23707) );
  sky130_fd_sc_hd__nand3_1 U28918 ( .A(n23709), .B(n23708), .C(n23707), .Y(
        j202_soc_core_j22_cpu_rf_N312) );
  sky130_fd_sc_hd__nand2_1 U28919 ( .A(n11611), .B(n11157), .Y(n23713) );
  sky130_fd_sc_hd__a22oi_1 U28920 ( .A1(n23794), .A2(n27365), .B1(n26895), 
        .B2(n25291), .Y(n23712) );
  sky130_fd_sc_hd__nand2_1 U28921 ( .A(n23710), .B(n24593), .Y(n23711) );
  sky130_fd_sc_hd__nand3_1 U28922 ( .A(n23713), .B(n23712), .C(n23711), .Y(
        j202_soc_core_j22_cpu_rf_N311) );
  sky130_fd_sc_hd__a22oi_1 U28923 ( .A1(n23731), .A2(n23762), .B1(n21914), 
        .B2(n23777), .Y(n26553) );
  sky130_fd_sc_hd__nand2_1 U28924 ( .A(n27395), .B(n11157), .Y(n23716) );
  sky130_fd_sc_hd__a22oi_1 U28925 ( .A1(n23794), .A2(n27396), .B1(n25806), 
        .B2(n24593), .Y(n23715) );
  sky130_fd_sc_hd__nand2_1 U28926 ( .A(n26895), .B(n25848), .Y(n23714) );
  sky130_fd_sc_hd__nand3_1 U28927 ( .A(n23716), .B(n23715), .C(n23714), .Y(
        j202_soc_core_j22_cpu_rf_N306) );
  sky130_fd_sc_hd__a22oi_1 U28928 ( .A1(n23794), .A2(n27455), .B1(n23717), 
        .B2(n24593), .Y(n23719) );
  sky130_fd_sc_hd__nand2_1 U28929 ( .A(n12417), .B(n11157), .Y(n23718) );
  sky130_fd_sc_hd__o211ai_1 U28930 ( .A1(n23784), .A2(n23720), .B1(n23719), 
        .C1(n23718), .Y(j202_soc_core_j22_cpu_rf_N298) );
  sky130_fd_sc_hd__nand2_1 U28931 ( .A(n12389), .B(n11157), .Y(n23723) );
  sky130_fd_sc_hd__a22oi_1 U28932 ( .A1(n23794), .A2(n27389), .B1(n24729), 
        .B2(n24593), .Y(n23722) );
  sky130_fd_sc_hd__nand2_1 U28933 ( .A(n26895), .B(n25555), .Y(n23721) );
  sky130_fd_sc_hd__nand3_1 U28934 ( .A(n23723), .B(n23722), .C(n23721), .Y(
        j202_soc_core_j22_cpu_rf_N307) );
  sky130_fd_sc_hd__nand2_1 U28935 ( .A(n11764), .B(n11157), .Y(n23726) );
  sky130_fd_sc_hd__a22oi_1 U28936 ( .A1(n23794), .A2(n27447), .B1(n26895), 
        .B2(n25261), .Y(n23725) );
  sky130_fd_sc_hd__nand2_1 U28937 ( .A(n23996), .B(n24593), .Y(n23724) );
  sky130_fd_sc_hd__nand3_1 U28938 ( .A(n23726), .B(n23725), .C(n23724), .Y(
        j202_soc_core_j22_cpu_rf_N314) );
  sky130_fd_sc_hd__nand2_1 U28939 ( .A(n26557), .B(n11157), .Y(n23730) );
  sky130_fd_sc_hd__a22oi_1 U28940 ( .A1(n23794), .A2(n27368), .B1(n26895), 
        .B2(n26446), .Y(n23729) );
  sky130_fd_sc_hd__nand2_1 U28941 ( .A(n26410), .B(n24593), .Y(n23728) );
  sky130_fd_sc_hd__nand3_1 U28942 ( .A(n23730), .B(n23729), .C(n23728), .Y(
        j202_soc_core_j22_cpu_rf_N326) );
  sky130_fd_sc_hd__nand2_1 U28943 ( .A(n12647), .B(n11157), .Y(n23734) );
  sky130_fd_sc_hd__a22oi_1 U28944 ( .A1(n23794), .A2(n27392), .B1(n26895), 
        .B2(n25851), .Y(n23733) );
  sky130_fd_sc_hd__nand2_1 U28945 ( .A(n23831), .B(n24593), .Y(n23732) );
  sky130_fd_sc_hd__nand3_1 U28946 ( .A(n23734), .B(n23733), .C(n23732), .Y(
        j202_soc_core_j22_cpu_rf_N322) );
  sky130_fd_sc_hd__nor2_1 U28947 ( .A(n27928), .B(n27895), .Y(
        j202_soc_core_j22_cpu_id_idec_N900) );
  sky130_fd_sc_hd__nand2_1 U28948 ( .A(n11612), .B(n11157), .Y(n23738) );
  sky130_fd_sc_hd__a22oi_1 U28949 ( .A1(n23794), .A2(n24052), .B1(n26895), 
        .B2(n26949), .Y(n23737) );
  sky130_fd_sc_hd__nand2_1 U28950 ( .A(n24044), .B(n24593), .Y(n23736) );
  sky130_fd_sc_hd__nand3_1 U28951 ( .A(n23738), .B(n23737), .C(n23736), .Y(
        j202_soc_core_j22_cpu_rf_N327) );
  sky130_fd_sc_hd__nand2_1 U28952 ( .A(n11770), .B(n11157), .Y(n23741) );
  sky130_fd_sc_hd__a22oi_1 U28953 ( .A1(n23794), .A2(n27425), .B1(n26895), 
        .B2(n25669), .Y(n23740) );
  sky130_fd_sc_hd__nand2_1 U28954 ( .A(n24085), .B(n24593), .Y(n23739) );
  sky130_fd_sc_hd__nand3_1 U28955 ( .A(n23741), .B(n23740), .C(n23739), .Y(
        j202_soc_core_j22_cpu_rf_N317) );
  sky130_fd_sc_hd__nand2_1 U28956 ( .A(n11771), .B(n11157), .Y(n23745) );
  sky130_fd_sc_hd__a22oi_1 U28957 ( .A1(n23794), .A2(n27357), .B1(n26895), 
        .B2(n26520), .Y(n23744) );
  sky130_fd_sc_hd__nand2_1 U28958 ( .A(n24490), .B(n24593), .Y(n23743) );
  sky130_fd_sc_hd__nand3_1 U28959 ( .A(n23745), .B(n23744), .C(n23743), .Y(
        j202_soc_core_j22_cpu_rf_N328) );
  sky130_fd_sc_hd__nor2_1 U28960 ( .A(n26548), .B(n10967), .Y(n25417) );
  sky130_fd_sc_hd__nand2_1 U28961 ( .A(n29549), .B(n11157), .Y(n23749) );
  sky130_fd_sc_hd__a22oi_1 U28962 ( .A1(n23794), .A2(n27412), .B1(n26895), 
        .B2(n25423), .Y(n23748) );
  sky130_fd_sc_hd__nand2_1 U28963 ( .A(n25412), .B(n24593), .Y(n23747) );
  sky130_fd_sc_hd__nand3_1 U28964 ( .A(n23749), .B(n23748), .C(n23747), .Y(
        j202_soc_core_j22_cpu_rf_N319) );
  sky130_fd_sc_hd__nand2_1 U28965 ( .A(n25259), .B(n11157), .Y(n23752) );
  sky130_fd_sc_hd__inv_2 U28966 ( .A(n23794), .Y(n26892) );
  sky130_fd_sc_hd__a22oi_1 U28967 ( .A1(n23794), .A2(n27432), .B1(n26895), 
        .B2(n24799), .Y(n23751) );
  sky130_fd_sc_hd__nand2_1 U28968 ( .A(n24766), .B(n24593), .Y(n23750) );
  sky130_fd_sc_hd__nand3_1 U28969 ( .A(n23752), .B(n23751), .C(n23750), .Y(
        j202_soc_core_j22_cpu_rf_N316) );
  sky130_fd_sc_hd__nand2_1 U28970 ( .A(n11589), .B(n11157), .Y(n23756) );
  sky130_fd_sc_hd__a22oi_1 U28971 ( .A1(n23794), .A2(n27399), .B1(n26895), 
        .B2(n26069), .Y(n23755) );
  sky130_fd_sc_hd__nand2_1 U28972 ( .A(n25176), .B(n24593), .Y(n23754) );
  sky130_fd_sc_hd__nand3_1 U28973 ( .A(n23756), .B(n23755), .C(n23754), .Y(
        j202_soc_core_j22_cpu_rf_N321) );
  sky130_fd_sc_hd__nand2_1 U28974 ( .A(n26507), .B(n11157), .Y(n23761) );
  sky130_fd_sc_hd__a22oi_1 U28975 ( .A1(n23794), .A2(n27405), .B1(n26895), 
        .B2(n26111), .Y(n23760) );
  sky130_fd_sc_hd__nand2_1 U28976 ( .A(n26096), .B(n24593), .Y(n23759) );
  sky130_fd_sc_hd__nand3_1 U28977 ( .A(n23761), .B(n23760), .C(n23759), .Y(
        j202_soc_core_j22_cpu_rf_N320) );
  sky130_fd_sc_hd__nand2_1 U28978 ( .A(n23763), .B(n23762), .Y(n23765) );
  sky130_fd_sc_hd__nand2_1 U28979 ( .A(n28971), .B(n23777), .Y(n23764) );
  sky130_fd_sc_hd__nand2_1 U28980 ( .A(n12645), .B(n11157), .Y(n23768) );
  sky130_fd_sc_hd__a22oi_1 U28981 ( .A1(n23794), .A2(n27383), .B1(n25042), 
        .B2(n24593), .Y(n23767) );
  sky130_fd_sc_hd__nand2_1 U28982 ( .A(n26895), .B(n25053), .Y(n23766) );
  sky130_fd_sc_hd__nand3_1 U28983 ( .A(n23768), .B(n23767), .C(n23766), .Y(
        j202_soc_core_j22_cpu_rf_N308) );
  sky130_fd_sc_hd__a22oi_1 U28984 ( .A1(n23794), .A2(n27419), .B1(n26895), 
        .B2(n24542), .Y(n23772) );
  sky130_fd_sc_hd__nand2_1 U28985 ( .A(n24531), .B(n24593), .Y(n23771) );
  sky130_fd_sc_hd__o211ai_1 U28986 ( .A1(n26897), .A2(n24546), .B1(n23772), 
        .C1(n23771), .Y(j202_soc_core_j22_cpu_rf_N318) );
  sky130_fd_sc_hd__a22oi_1 U28987 ( .A1(n23794), .A2(n27402), .B1(n23773), 
        .B2(n24593), .Y(n23775) );
  sky130_fd_sc_hd__nand2_1 U28988 ( .A(n12455), .B(n11157), .Y(n23774) );
  sky130_fd_sc_hd__o211ai_1 U28989 ( .A1(n23784), .A2(n23776), .B1(n23775), 
        .C1(n23774), .Y(j202_soc_core_j22_cpu_rf_N305) );
  sky130_fd_sc_hd__a22oi_1 U28990 ( .A1(n23794), .A2(n27377), .B1(n24676), 
        .B2(n24593), .Y(n23779) );
  sky130_fd_sc_hd__nand2_1 U28991 ( .A(n11766), .B(n11157), .Y(n23778) );
  sky130_fd_sc_hd__o211ai_1 U28992 ( .A1(n23784), .A2(n23780), .B1(n23779), 
        .C1(n23778), .Y(j202_soc_core_j22_cpu_rf_N309) );
  sky130_fd_sc_hd__a22oi_1 U28993 ( .A1(n23794), .A2(n27443), .B1(n23781), 
        .B2(n24593), .Y(n23783) );
  sky130_fd_sc_hd__nand2_1 U28994 ( .A(n27442), .B(n11157), .Y(n23782) );
  sky130_fd_sc_hd__o211ai_1 U28995 ( .A1(j202_soc_core_j22_cpu_pc[1]), .A2(
        n23784), .B1(n23783), .C1(n23782), .Y(j202_soc_core_j22_cpu_rf_N299)
         );
  sky130_fd_sc_hd__a22oi_1 U28996 ( .A1(n23794), .A2(n24671), .B1(n26895), 
        .B2(n23785), .Y(n23788) );
  sky130_fd_sc_hd__nand2_1 U28997 ( .A(n23786), .B(n24593), .Y(n23787) );
  sky130_fd_sc_hd__o211ai_1 U28998 ( .A1(n26897), .A2(n25157), .B1(n23788), 
        .C1(n23787), .Y(j202_soc_core_j22_cpu_rf_N325) );
  sky130_fd_sc_hd__a22oi_1 U28999 ( .A1(n23794), .A2(n25122), .B1(n26895), 
        .B2(n25188), .Y(n23791) );
  sky130_fd_sc_hd__nand2_1 U29000 ( .A(n25136), .B(n24593), .Y(n23790) );
  sky130_fd_sc_hd__a22oi_1 U29001 ( .A1(n23794), .A2(n27354), .B1(n24156), 
        .B2(n24593), .Y(n23793) );
  sky130_fd_sc_hd__nand2_1 U29002 ( .A(n26895), .B(n25268), .Y(n23792) );
  sky130_fd_sc_hd__o211ai_1 U29003 ( .A1(n26897), .A2(n25276), .B1(n23793), 
        .C1(n23792), .Y(j202_soc_core_j22_cpu_rf_N313) );
  sky130_fd_sc_hd__a22oi_1 U29004 ( .A1(n23794), .A2(n24613), .B1(n26895), 
        .B2(n25715), .Y(n23796) );
  sky130_fd_sc_hd__nand2_1 U29005 ( .A(n24626), .B(n24593), .Y(n23795) );
  sky130_fd_sc_hd__o211ai_1 U29006 ( .A1(n26897), .A2(n11103), .B1(n23796), 
        .C1(n23795), .Y(j202_soc_core_j22_cpu_rf_N315) );
  sky130_fd_sc_hd__a22oi_1 U29007 ( .A1(n23794), .A2(n25061), .B1(n26895), 
        .B2(n25077), .Y(n23799) );
  sky130_fd_sc_hd__nand2_1 U29008 ( .A(n25070), .B(n24593), .Y(n23798) );
  sky130_fd_sc_hd__o211ai_1 U29009 ( .A1(n26897), .A2(n11102), .B1(n23799), 
        .C1(n23798), .Y(j202_soc_core_j22_cpu_rf_N324) );
  sky130_fd_sc_hd__nor2_1 U29010 ( .A(n28590), .B(
        j202_soc_core_ahb2aqu_00_aqu_st_0_), .Y(n24562) );
  sky130_fd_sc_hd__nand2_1 U29011 ( .A(n12456), .B(n24562), .Y(
        j202_soc_core_ahb2aqu_00_N95) );
  sky130_fd_sc_hd__nand2_1 U29012 ( .A(n11798), .B(n24350), .Y(n27685) );
  sky130_fd_sc_hd__o21ai_1 U29013 ( .A1(n23800), .A2(n27685), .B1(n27877), .Y(
        n23806) );
  sky130_fd_sc_hd__nand2_1 U29014 ( .A(n11132), .B(n11792), .Y(n27170) );
  sky130_fd_sc_hd__nand3_1 U29015 ( .A(n23801), .B(n27686), .C(n27170), .Y(
        n23804) );
  sky130_fd_sc_hd__nor2_1 U29016 ( .A(n12595), .B(n24704), .Y(n23805) );
  sky130_fd_sc_hd__o21a_1 U29017 ( .A1(n23806), .A2(n23805), .B1(n27980), .X(
        j202_soc_core_j22_cpu_id_idec_N917) );
  sky130_fd_sc_hd__nand3_1 U29018 ( .A(n24091), .B(n24455), .C(n27256), .Y(
        n27883) );
  sky130_fd_sc_hd__nand2_1 U29019 ( .A(n23818), .B(n24266), .Y(n23822) );
  sky130_fd_sc_hd__nor2_1 U29020 ( .A(n24446), .B(n24448), .Y(n24256) );
  sky130_fd_sc_hd__o21a_1 U29021 ( .A1(n12757), .A2(n27772), .B1(n24353), .X(
        n23819) );
  sky130_fd_sc_hd__nand2_1 U29022 ( .A(n24575), .B(n29594), .Y(n29113) );
  sky130_fd_sc_hd__nand3_1 U29023 ( .A(n23824), .B(n26398), .C(n23823), .Y(
        n23830) );
  sky130_fd_sc_hd__and4_1 U29024 ( .A(n23827), .B(n11713), .C(n23826), .D(
        n23825), .X(n23828) );
  sky130_fd_sc_hd__nand2_1 U29025 ( .A(n23830), .B(n23852), .Y(n23846) );
  sky130_fd_sc_hd__nand2_1 U29026 ( .A(n23831), .B(n26409), .Y(n23844) );
  sky130_fd_sc_hd__o22ai_1 U29027 ( .A1(n23834), .A2(n26431), .B1(n23832), 
        .B2(n26412), .Y(n23842) );
  sky130_fd_sc_hd__o22ai_1 U29028 ( .A1(n26581), .A2(n26416), .B1(n26706), 
        .B2(n26424), .Y(n23833) );
  sky130_fd_sc_hd__a21oi_1 U29029 ( .A1(n25131), .A2(n26718), .B1(n23833), .Y(
        n23840) );
  sky130_fd_sc_hd__o22a_1 U29030 ( .A1(n26704), .A2(n26427), .B1(n25821), .B2(
        n26425), .X(n23839) );
  sky130_fd_sc_hd__nand2_1 U29031 ( .A(n27392), .B(n25871), .Y(n26613) );
  sky130_fd_sc_hd__nand2_1 U29032 ( .A(n23834), .B(n26701), .Y(n26614) );
  sky130_fd_sc_hd__nand3_1 U29033 ( .A(n26614), .B(n26326), .C(n26613), .Y(
        n23835) );
  sky130_fd_sc_hd__o211ai_1 U29034 ( .A1(n26432), .A2(n26613), .B1(n23836), 
        .C1(n23835), .Y(n23837) );
  sky130_fd_sc_hd__a21oi_1 U29035 ( .A1(n24483), .A2(n26508), .B1(n23837), .Y(
        n23838) );
  sky130_fd_sc_hd__nand4_1 U29036 ( .A(n23840), .B(n26411), .C(n23839), .D(
        n23838), .Y(n23841) );
  sky130_fd_sc_hd__nor2_1 U29037 ( .A(n23842), .B(n23841), .Y(n23843) );
  sky130_fd_sc_hd__nand2_1 U29038 ( .A(n23844), .B(n23843), .Y(n23845) );
  sky130_fd_sc_hd__nand2_1 U29039 ( .A(n23847), .B(n24785), .Y(n23848) );
  sky130_fd_sc_hd__nand2_1 U29040 ( .A(n23848), .B(n26407), .Y(n23849) );
  sky130_fd_sc_hd__nand2_1 U29041 ( .A(n23851), .B(n23852), .Y(n23854) );
  sky130_fd_sc_hd__nand3_1 U29042 ( .A(n23235), .B(n26862), .C(n23852), .Y(
        n23853) );
  sky130_fd_sc_hd__nor2_1 U29044 ( .A(n23858), .B(n23857), .Y(n24332) );
  sky130_fd_sc_hd__nand3_1 U29045 ( .A(n24332), .B(n23859), .C(n24469), .Y(
        n27771) );
  sky130_fd_sc_hd__nand2_1 U29046 ( .A(n23860), .B(
        j202_soc_core_j22_cpu_opst[0]), .Y(n25779) );
  sky130_fd_sc_hd__a31oi_1 U29047 ( .A1(n23863), .A2(
        j202_soc_core_j22_cpu_opst[1]), .A3(n23862), .B1(n23861), .Y(n23864)
         );
  sky130_fd_sc_hd__nand2_1 U29048 ( .A(n25779), .B(n23864), .Y(n23865) );
  sky130_fd_sc_hd__o31a_1 U29049 ( .A1(n27919), .A2(n27771), .A3(n23865), .B1(
        n10607), .X(n29117) );
  sky130_fd_sc_hd__and3_1 U29050 ( .A(n23866), .B(la_data_in[31]), .C(n29594), 
        .X(n29121) );
  sky130_fd_sc_hd__and3_1 U29051 ( .A(n23867), .B(la_data_in[30]), .C(n29594), 
        .X(n29122) );
  sky130_fd_sc_hd__and3_1 U29052 ( .A(n23868), .B(la_data_in[29]), .C(n29595), 
        .X(n29123) );
  sky130_fd_sc_hd__and3_1 U29053 ( .A(n23869), .B(la_data_in[28]), .C(n29594), 
        .X(n29124) );
  sky130_fd_sc_hd__and3_1 U29054 ( .A(n23870), .B(la_data_in[27]), .C(n29594), 
        .X(n29125) );
  sky130_fd_sc_hd__and3_1 U29055 ( .A(n23871), .B(la_data_in[26]), .C(n29595), 
        .X(n29126) );
  sky130_fd_sc_hd__and3_1 U29056 ( .A(n23872), .B(la_data_in[25]), .C(n29594), 
        .X(n29127) );
  sky130_fd_sc_hd__and3_1 U29057 ( .A(n23873), .B(la_data_in[24]), .C(n29594), 
        .X(n29128) );
  sky130_fd_sc_hd__and3_1 U29058 ( .A(n23874), .B(la_data_in[23]), .C(n29595), 
        .X(n29129) );
  sky130_fd_sc_hd__and3_1 U29059 ( .A(n23875), .B(la_data_in[22]), .C(n29595), 
        .X(n29130) );
  sky130_fd_sc_hd__and3_1 U29060 ( .A(n23876), .B(la_data_in[21]), .C(n29595), 
        .X(n29131) );
  sky130_fd_sc_hd__and3_1 U29061 ( .A(n23877), .B(la_data_in[20]), .C(n12142), 
        .X(n29132) );
  sky130_fd_sc_hd__and3_1 U29062 ( .A(n23878), .B(la_data_in[19]), .C(n29594), 
        .X(n29133) );
  sky130_fd_sc_hd__and3_1 U29063 ( .A(n23879), .B(la_data_in[18]), .C(n29595), 
        .X(n29134) );
  sky130_fd_sc_hd__and3_1 U29064 ( .A(n23880), .B(la_data_in[17]), .C(n29594), 
        .X(n29135) );
  sky130_fd_sc_hd__o211a_2 U29065 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[6]), .A2(n24892), .B1(
        n28622), .C1(n24899), .X(n29153) );
  sky130_fd_sc_hd__o211a_2 U29066 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[4]), .A2(n24889), .B1(
        n28622), .C1(n24893), .X(n29154) );
  sky130_fd_sc_hd__nand2_1 U29067 ( .A(n26242), .B(n25929), .Y(n27719) );
  sky130_fd_sc_hd__nand2b_1 U29068 ( .A_N(n25961), .B(n26035), .Y(n28751) );
  sky130_fd_sc_hd__and4_1 U29069 ( .A(n24814), .B(n29595), .C(
        j202_soc_core_ahb2apb_00_state[0]), .D(
        j202_soc_core_ahb2apb_00_state[1]), .X(n29221) );
  sky130_fd_sc_hd__and3_1 U29070 ( .A(n23910), .B(n23909), .C(
        j202_soc_core_aquc_WE_), .X(n29231) );
  sky130_fd_sc_hd__nand2_1 U29071 ( .A(n28743), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[1]), .Y(n26204) );
  sky130_fd_sc_hd__nand2_1 U29072 ( .A(n28743), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[0]), .Y(n26196) );
  sky130_fd_sc_hd__nand2_1 U29073 ( .A(n29056), .B(n28110), .Y(n23913) );
  sky130_fd_sc_hd__nor2_1 U29074 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd), .B(n26260), .Y(n26233)
         );
  sky130_fd_sc_hd__o211ai_1 U29075 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd), .A2(n26202), .B1(n23913), 
        .C1(n23912), .Y(n26197) );
  sky130_fd_sc_hd__nand2_1 U29076 ( .A(n26196), .B(n26197), .Y(n26205) );
  sky130_fd_sc_hd__nand2_1 U29077 ( .A(n26204), .B(n23914), .Y(
        DP_OP_1508J1_126_2326_n4) );
  sky130_fd_sc_hd__nand2_1 U29078 ( .A(n23922), .B(n18916), .Y(n23916) );
  sky130_fd_sc_hd__o211ai_1 U29079 ( .A1(n26859), .A2(n23916), .B1(n26407), 
        .C1(n23915), .Y(n23917) );
  sky130_fd_sc_hd__nand2_1 U29081 ( .A(n23921), .B(n27354), .Y(n23923) );
  sky130_fd_sc_hd__nand2_1 U29082 ( .A(n23923), .B(n23922), .Y(n23926) );
  sky130_fd_sc_hd__nand2_1 U29083 ( .A(n26883), .B(n26409), .Y(n23924) );
  sky130_fd_sc_hd__nand2_1 U29084 ( .A(n23924), .B(n24778), .Y(n23925) );
  sky130_fd_sc_hd__nor2_1 U29086 ( .A(n23927), .B(n26746), .Y(n23930) );
  sky130_fd_sc_hd__nor2_1 U29087 ( .A(n23928), .B(n26424), .Y(n23929) );
  sky130_fd_sc_hd__mux2_2 U29088 ( .A0(n23930), .A1(n23929), .S(n27415), .X(
        n23936) );
  sky130_fd_sc_hd__xnor2_1 U29089 ( .A(n26859), .B(n27347), .Y(n26700) );
  sky130_fd_sc_hd__o22a_1 U29090 ( .A1(n26415), .A2(n26700), .B1(n26702), .B2(
        n26419), .X(n23934) );
  sky130_fd_sc_hd__o22ai_1 U29091 ( .A1(n26423), .A2(n27347), .B1(n26704), 
        .B2(n26416), .Y(n23932) );
  sky130_fd_sc_hd__o22ai_1 U29092 ( .A1(n26578), .A2(n26427), .B1(n26567), 
        .B2(n26425), .Y(n23931) );
  sky130_fd_sc_hd__nor2_1 U29093 ( .A(n23932), .B(n23931), .Y(n23933) );
  sky130_fd_sc_hd__o211ai_1 U29094 ( .A1(n26885), .A2(n26431), .B1(n23934), 
        .C1(n23933), .Y(n23935) );
  sky130_fd_sc_hd__a21oi_1 U29095 ( .A1(n27435), .A2(n23936), .B1(n23935), .Y(
        n23937) );
  sky130_fd_sc_hd__nand2_1 U29096 ( .A(n23938), .B(n23937), .Y(n23939) );
  sky130_fd_sc_hd__a21oi_1 U29097 ( .A1(n27347), .A2(n25415), .B1(n23940), .Y(
        n23942) );
  sky130_fd_sc_hd__nand3_1 U29098 ( .A(n25063), .B(n25237), .C(n27415), .Y(
        n23941) );
  sky130_fd_sc_hd__o22ai_1 U29099 ( .A1(n27466), .A2(n27349), .B1(n27465), 
        .B2(n23944), .Y(j202_soc_core_j22_cpu_rf_N2787) );
  sky130_fd_sc_hd__o22ai_1 U29100 ( .A1(n27209), .A2(n27349), .B1(n23039), 
        .B2(n23944), .Y(j202_soc_core_j22_cpu_rf_N2750) );
  sky130_fd_sc_hd__o22ai_1 U29101 ( .A1(n27213), .A2(n27349), .B1(n27212), 
        .B2(n23944), .Y(j202_soc_core_j22_cpu_rf_N2824) );
  sky130_fd_sc_hd__o22ai_1 U29102 ( .A1(n27226), .A2(n27349), .B1(n23079), 
        .B2(n12478), .Y(j202_soc_core_j22_cpu_rf_N3157) );
  sky130_fd_sc_hd__o22ai_1 U29103 ( .A1(n27221), .A2(n27349), .B1(n27220), 
        .B2(n23944), .Y(j202_soc_core_j22_cpu_rf_N2898) );
  sky130_fd_sc_hd__o22ai_1 U29104 ( .A1(n27217), .A2(n27349), .B1(n27216), 
        .B2(n23944), .Y(j202_soc_core_j22_cpu_rf_N2861) );
  sky130_fd_sc_hd__o22ai_1 U29105 ( .A1(n27219), .A2(n27349), .B1(n27218), 
        .B2(n23944), .Y(j202_soc_core_j22_cpu_rf_N3009) );
  sky130_fd_sc_hd__o22ai_1 U29106 ( .A1(n27575), .A2(n27349), .B1(n27574), 
        .B2(n23944), .Y(j202_soc_core_j22_cpu_rf_N3120) );
  sky130_fd_sc_hd__o22ai_1 U29107 ( .A1(n27333), .A2(n27349), .B1(n23178), 
        .B2(n23944), .Y(j202_soc_core_j22_cpu_rf_N3083) );
  sky130_fd_sc_hd__o22ai_1 U29108 ( .A1(n26378), .A2(n27349), .B1(n26449), 
        .B2(n12478), .Y(j202_soc_core_j22_cpu_rf_N3268) );
  sky130_fd_sc_hd__o22ai_1 U29109 ( .A1(n11141), .A2(n27349), .B1(n27124), 
        .B2(n12478), .Y(j202_soc_core_j22_cpu_rf_N2713) );
  sky130_fd_sc_hd__o22ai_1 U29110 ( .A1(n27211), .A2(n27349), .B1(n27210), 
        .B2(n12478), .Y(j202_soc_core_j22_cpu_rf_N3231) );
  sky130_fd_sc_hd__o22ai_1 U29111 ( .A1(n27223), .A2(n27349), .B1(n27222), 
        .B2(n12478), .Y(j202_soc_core_j22_cpu_rf_N3046) );
  sky130_fd_sc_hd__o22ai_1 U29112 ( .A1(n27215), .A2(n27349), .B1(n27214), 
        .B2(n12478), .Y(j202_soc_core_j22_cpu_rf_N2935) );
  sky130_fd_sc_hd__o22ai_1 U29113 ( .A1(n27225), .A2(n27349), .B1(n27224), 
        .B2(n12478), .Y(j202_soc_core_j22_cpu_rf_N2972) );
  sky130_fd_sc_hd__nand2_1 U29114 ( .A(n26898), .B(n23943), .Y(n26899) );
  sky130_fd_sc_hd__o22ai_1 U29115 ( .A1(n27349), .A2(n26899), .B1(n26898), 
        .B2(n12478), .Y(j202_soc_core_j22_cpu_rf_N3343) );
  sky130_fd_sc_hd__o22ai_1 U29116 ( .A1(n27228), .A2(n27349), .B1(n27227), 
        .B2(n12478), .Y(j202_soc_core_j22_cpu_rf_N3194) );
  sky130_fd_sc_hd__inv_4 U29117 ( .A(n25822), .Y(n26976) );
  sky130_fd_sc_hd__a21oi_1 U29118 ( .A1(n25344), .A2(
        j202_soc_core_j22_cpu_ml_bufa[12]), .B1(n26976), .Y(n23946) );
  sky130_fd_sc_hd__nand3_1 U29119 ( .A(n12356), .B(n24551), .C(n26872), .Y(
        n23945) );
  sky130_fd_sc_hd__nand3_1 U29120 ( .A(n25875), .B(n24511), .C(n26872), .Y(
        n23948) );
  sky130_fd_sc_hd__nor2_1 U29121 ( .A(n29015), .B(n29077), .Y(n23955) );
  sky130_fd_sc_hd__nand2_1 U29122 ( .A(n12757), .B(n11873), .Y(n23952) );
  sky130_fd_sc_hd__a21o_1 U29123 ( .A1(n23957), .A2(n27166), .B1(n27956), .X(
        n23958) );
  sky130_fd_sc_hd__nand2_1 U29124 ( .A(n12515), .B(n27980), .Y(n23960) );
  sky130_fd_sc_hd__nand2b_1 U29125 ( .A_N(n23967), .B(n23966), .Y(n23968) );
  sky130_fd_sc_hd__a21oi_1 U29126 ( .A1(n25344), .A2(n18147), .B1(n26976), .Y(
        n23971) );
  sky130_fd_sc_hd__nand3_1 U29127 ( .A(n12357), .B(n25147), .C(n26872), .Y(
        n23970) );
  sky130_fd_sc_hd__buf_6 U29129 ( .A(n23974), .X(n29312) );
  sky130_fd_sc_hd__buf_6 U29130 ( .A(n23974), .X(n29313) );
  sky130_fd_sc_hd__nand2_1 U29131 ( .A(n23976), .B(n26802), .Y(n24003) );
  sky130_fd_sc_hd__nand2_1 U29132 ( .A(n23978), .B(n23977), .Y(n23979) );
  sky130_fd_sc_hd__nand2_1 U29133 ( .A(n23979), .B(n26802), .Y(n24002) );
  sky130_fd_sc_hd__a21oi_1 U29134 ( .A1(n27447), .A2(n25415), .B1(n26085), .Y(
        n23980) );
  sky130_fd_sc_hd__nand2_1 U29135 ( .A(n26329), .B(n11713), .Y(n26102) );
  sky130_fd_sc_hd__o22ai_1 U29136 ( .A1(n26580), .A2(n26431), .B1(n23982), 
        .B2(n26412), .Y(n23992) );
  sky130_fd_sc_hd__o22ai_1 U29137 ( .A1(n26567), .A2(n26427), .B1(n25821), 
        .B2(n26416), .Y(n23984) );
  sky130_fd_sc_hd__o22ai_1 U29138 ( .A1(n25128), .A2(n26424), .B1(n25789), 
        .B2(n26425), .Y(n23983) );
  sky130_fd_sc_hd__nor2_1 U29139 ( .A(n23984), .B(n23983), .Y(n23990) );
  sky130_fd_sc_hd__xor2_1 U29140 ( .A(n27045), .B(n27447), .X(n26645) );
  sky130_fd_sc_hd__o22ai_1 U29141 ( .A1(n18916), .A2(n23985), .B1(n26423), 
        .B2(n27447), .Y(n23986) );
  sky130_fd_sc_hd__a21o_1 U29142 ( .A1(n26077), .A2(n25871), .B1(n23986), .X(
        n23987) );
  sky130_fd_sc_hd__a21oi_1 U29143 ( .A1(n26326), .A2(n26645), .B1(n23987), .Y(
        n23989) );
  sky130_fd_sc_hd__o22a_1 U29144 ( .A1(n26571), .A2(n26418), .B1(n26565), .B2(
        n26419), .X(n23988) );
  sky130_fd_sc_hd__nand4_1 U29145 ( .A(n23990), .B(n26411), .C(n23989), .D(
        n23988), .Y(n23991) );
  sky130_fd_sc_hd__nor2_1 U29146 ( .A(n23992), .B(n23991), .Y(n23993) );
  sky130_fd_sc_hd__o21ai_1 U29147 ( .A1(n18916), .A2(n23994), .B1(n23993), .Y(
        n23995) );
  sky130_fd_sc_hd__a21oi_1 U29148 ( .A1(n23996), .A2(n26409), .B1(n23995), .Y(
        n23999) );
  sky130_fd_sc_hd__o21ai_1 U29149 ( .A1(n26352), .A2(n27045), .B1(n26351), .Y(
        n23997) );
  sky130_fd_sc_hd__nand2_1 U29150 ( .A(n27044), .B(n23997), .Y(n23998) );
  sky130_fd_sc_hd__o211ai_1 U29151 ( .A1(n26102), .A2(n24171), .B1(n23999), 
        .C1(n23998), .Y(n24000) );
  sky130_fd_sc_hd__o22ai_1 U29152 ( .A1(n27209), .A2(n27451), .B1(n23039), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N2733) );
  sky130_fd_sc_hd__o22ai_1 U29153 ( .A1(n27333), .A2(n27451), .B1(n23178), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N3066) );
  sky130_fd_sc_hd__o22ai_1 U29154 ( .A1(n27466), .A2(n27451), .B1(n27465), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N2770) );
  sky130_fd_sc_hd__o22ai_1 U29155 ( .A1(n27213), .A2(n27451), .B1(n27212), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N2807) );
  sky130_fd_sc_hd__o22ai_1 U29156 ( .A1(n27221), .A2(n27451), .B1(n27220), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N2881) );
  sky130_fd_sc_hd__o22ai_1 U29157 ( .A1(n27217), .A2(n27451), .B1(n27216), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N2844) );
  sky130_fd_sc_hd__o22ai_1 U29158 ( .A1(n27219), .A2(n27451), .B1(n27218), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N2992) );
  sky130_fd_sc_hd__o22ai_1 U29159 ( .A1(n27575), .A2(n27451), .B1(n27574), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N3103) );
  sky130_fd_sc_hd__o22ai_1 U29160 ( .A1(n26378), .A2(n27451), .B1(n26449), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N3251) );
  sky130_fd_sc_hd__o22ai_1 U29161 ( .A1(n27211), .A2(n27451), .B1(n27210), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N3214) );
  sky130_fd_sc_hd__o22ai_1 U29162 ( .A1(n27223), .A2(n27451), .B1(n27222), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N3029) );
  sky130_fd_sc_hd__o22ai_1 U29163 ( .A1(n27215), .A2(n27451), .B1(n27214), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N2918) );
  sky130_fd_sc_hd__o22ai_1 U29164 ( .A1(n27451), .A2(n26899), .B1(n26898), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N3327) );
  sky130_fd_sc_hd__o22ai_1 U29165 ( .A1(n11141), .A2(n27451), .B1(n27124), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N2696) );
  sky130_fd_sc_hd__o22ai_1 U29166 ( .A1(n27225), .A2(n27451), .B1(n27224), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N2955) );
  sky130_fd_sc_hd__o22ai_1 U29167 ( .A1(n27228), .A2(n27451), .B1(n27227), 
        .B2(n12383), .Y(j202_soc_core_j22_cpu_rf_N3177) );
  sky130_fd_sc_hd__nor2_1 U29168 ( .A(j202_soc_core_intc_core_00_bs_addr[1]), 
        .B(j202_soc_core_intc_core_00_bs_addr[0]), .Y(n27066) );
  sky130_fd_sc_hd__nand2_1 U29169 ( .A(n27066), .B(n28890), .Y(n24969) );
  sky130_fd_sc_hd__nand3_1 U29170 ( .A(n24319), .B(n24005), .C(
        j202_soc_core_ahb2apb_01_state[1]), .Y(n24172) );
  sky130_fd_sc_hd__nor2_1 U29171 ( .A(j202_soc_core_intc_core_00_bs_addr[10]), 
        .B(j202_soc_core_intc_core_00_bs_addr[11]), .Y(n24008) );
  sky130_fd_sc_hd__nand4_1 U29172 ( .A(j202_soc_core_pstrb[5]), .B(
        j202_soc_core_pstrb[4]), .C(j202_soc_core_pstrb[6]), .D(
        j202_soc_core_pstrb[7]), .Y(n24006) );
  sky130_fd_sc_hd__nand2_1 U29173 ( .A(j202_soc_core_pwrite[1]), .B(n24006), 
        .Y(n24007) );
  sky130_fd_sc_hd__nand2_1 U29174 ( .A(n24008), .B(n24007), .Y(n24009) );
  sky130_fd_sc_hd__nor2_1 U29175 ( .A(n24172), .B(n24009), .Y(n24972) );
  sky130_fd_sc_hd__and4_1 U29176 ( .A(n28884), .B(n24751), .C(n28892), .D(
        j202_soc_core_intc_core_00_bs_addr[9]), .X(n24010) );
  sky130_fd_sc_hd__nand3_1 U29177 ( .A(n24011), .B(n24972), .C(n24010), .Y(
        n24607) );
  sky130_fd_sc_hd__nor2_1 U29178 ( .A(j202_soc_core_intc_core_00_bs_addr[3]), 
        .B(j202_soc_core_intc_core_00_bs_addr[2]), .Y(n28888) );
  sky130_fd_sc_hd__nand3_1 U29179 ( .A(n24755), .B(n28888), .C(n24756), .Y(
        n24753) );
  sky130_fd_sc_hd__o22ai_1 U29180 ( .A1(n28615), .A2(n25534), .B1(n24987), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U29182 ( .A1(n27226), .A2(n27394), .B1(n23079), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N3149) );
  sky130_fd_sc_hd__o22ai_1 U29183 ( .A1(n27209), .A2(n27394), .B1(n23039), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N2742) );
  sky130_fd_sc_hd__o22ai_1 U29184 ( .A1(n27333), .A2(n27394), .B1(n23178), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N3075) );
  sky130_fd_sc_hd__o22ai_1 U29185 ( .A1(n27217), .A2(n27394), .B1(n27216), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N2853) );
  sky130_fd_sc_hd__o22ai_1 U29186 ( .A1(n27213), .A2(n27394), .B1(n27212), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N2816) );
  sky130_fd_sc_hd__o22ai_1 U29187 ( .A1(n27221), .A2(n27394), .B1(n27220), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N2890) );
  sky130_fd_sc_hd__o22ai_1 U29188 ( .A1(n27466), .A2(n27394), .B1(n27465), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N2779) );
  sky130_fd_sc_hd__o22ai_1 U29189 ( .A1(n27219), .A2(n27394), .B1(n27218), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N3001) );
  sky130_fd_sc_hd__o22ai_1 U29190 ( .A1(n27575), .A2(n27394), .B1(n27574), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N3112) );
  sky130_fd_sc_hd__o22ai_1 U29191 ( .A1(n26378), .A2(n27394), .B1(n26449), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N3260) );
  sky130_fd_sc_hd__o22ai_1 U29192 ( .A1(n11141), .A2(n27394), .B1(n27124), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N2705) );
  sky130_fd_sc_hd__o22ai_1 U29193 ( .A1(n27223), .A2(n27394), .B1(n27222), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N3038) );
  sky130_fd_sc_hd__o22ai_1 U29194 ( .A1(n27215), .A2(n27394), .B1(n27214), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N2927) );
  sky130_fd_sc_hd__o22ai_1 U29195 ( .A1(n27211), .A2(n27394), .B1(n27210), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N3223) );
  sky130_fd_sc_hd__o22ai_1 U29196 ( .A1(n27225), .A2(n27394), .B1(n27224), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N2964) );
  sky130_fd_sc_hd__o22ai_1 U29197 ( .A1(n27394), .A2(n26899), .B1(n26898), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N3336) );
  sky130_fd_sc_hd__o22ai_1 U29198 ( .A1(n27228), .A2(n27394), .B1(n27227), 
        .B2(n25853), .Y(j202_soc_core_j22_cpu_rf_N3186) );
  sky130_fd_sc_hd__a21oi_1 U29199 ( .A1(n25344), .A2(n22919), .B1(n26976), .Y(
        n24016) );
  sky130_fd_sc_hd__nand3_1 U29200 ( .A(n12356), .B(n24013), .C(n26872), .Y(
        n24015) );
  sky130_fd_sc_hd__nand3_1 U29201 ( .A(n12916), .B(
        j202_soc_core_j22_cpu_ml_macl[9]), .C(n25826), .Y(n24014) );
  sky130_fd_sc_hd__nand3_1 U29202 ( .A(n24016), .B(n24015), .C(n24014), .Y(
        j202_soc_core_j22_cpu_ml_maclj[9]) );
  sky130_fd_sc_hd__nand3_1 U29203 ( .A(n27338), .B(
        j202_soc_core_j22_cpu_macop_MAC_[1]), .C(
        j202_soc_core_j22_cpu_macop_MAC_[3]), .Y(n24021) );
  sky130_fd_sc_hd__nand2_1 U29204 ( .A(n24017), .B(n11713), .Y(n27342) );
  sky130_fd_sc_hd__o21ai_1 U29205 ( .A1(n24019), .A2(n24018), .B1(n27342), .Y(
        n24020) );
  sky130_fd_sc_hd__nand2_1 U29206 ( .A(n27006), .B(n24020), .Y(n25215) );
  sky130_fd_sc_hd__nand2_1 U29207 ( .A(n11104), .B(n27339), .Y(n24025) );
  sky130_fd_sc_hd__nor2_1 U29208 ( .A(n11713), .B(n24021), .Y(n27351) );
  sky130_fd_sc_hd__nor2_1 U29209 ( .A(n24022), .B(n27343), .Y(n24024) );
  sky130_fd_sc_hd__inv_2 U29210 ( .A(n24163), .Y(n27356) );
  sky130_fd_sc_hd__o2bb2a_2 U29211 ( .A1_N(n24024), .A2_N(n26726), .B1(n24023), 
        .B2(n27356), .X(n27346) );
  sky130_fd_sc_hd__o211ai_1 U29212 ( .A1(n26707), .A2(n25215), .B1(n24025), 
        .C1(n27346), .Y(j202_soc_core_j22_cpu_ml_N331) );
  sky130_fd_sc_hd__nor2_1 U29213 ( .A(n24026), .B(n24607), .Y(n24760) );
  sky130_fd_sc_hd__nand3_1 U29214 ( .A(n24760), .B(n28886), .C(n24756), .Y(
        n24754) );
  sky130_fd_sc_hd__nor2_1 U29215 ( .A(n28882), .B(n24754), .Y(n25482) );
  sky130_fd_sc_hd__nor2_1 U29216 ( .A(n28590), .B(n25482), .Y(n25481) );
  sky130_fd_sc_hd__o22ai_1 U29217 ( .A1(n28601), .A2(n27021), .B1(n24027), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__nand2_1 U29218 ( .A(n24629), .B(n27339), .Y(n24028) );
  sky130_fd_sc_hd__o211ai_1 U29219 ( .A1(n25128), .A2(n25215), .B1(n24028), 
        .C1(n27346), .Y(j202_soc_core_j22_cpu_ml_N320) );
  sky130_fd_sc_hd__o22ai_1 U29220 ( .A1(n26456), .A2(n25534), .B1(n24029), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U29221 ( .A1(n28601), .A2(n25534), .B1(n24030), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U29222 ( .A1(n26556), .A2(n27209), .B1(n23039), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N2721) );
  sky130_fd_sc_hd__o22ai_1 U29223 ( .A1(n26556), .A2(n27226), .B1(n23079), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N3128) );
  sky130_fd_sc_hd__o22ai_1 U29224 ( .A1(n26556), .A2(n27211), .B1(n27210), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N3202) );
  sky130_fd_sc_hd__o22ai_1 U29225 ( .A1(n26556), .A2(n27215), .B1(n27214), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N2906) );
  sky130_fd_sc_hd__o22ai_1 U29226 ( .A1(n26556), .A2(n27225), .B1(n27224), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N2943) );
  sky130_fd_sc_hd__o22ai_1 U29227 ( .A1(n26556), .A2(n27228), .B1(n27227), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N3165) );
  sky130_fd_sc_hd__o22ai_1 U29228 ( .A1(n26556), .A2(n27333), .B1(n23178), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N3054) );
  sky130_fd_sc_hd__o22ai_1 U29229 ( .A1(n26556), .A2(n26378), .B1(n26449), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N3239) );
  sky130_fd_sc_hd__o22ai_1 U29230 ( .A1(n26556), .A2(n11141), .B1(n27124), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N2684) );
  sky130_fd_sc_hd__o22ai_1 U29231 ( .A1(n28611), .A2(n25534), .B1(n27544), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__xnor2_1 U29232 ( .A(n26971), .B(n26970), .Y(n24048) );
  sky130_fd_sc_hd__a21oi_1 U29233 ( .A1(n26971), .A2(n26323), .B1(n24067), .Y(
        n24046) );
  sky130_fd_sc_hd__o22ai_1 U29234 ( .A1(n26570), .A2(n26416), .B1(n26708), 
        .B2(n26425), .Y(n24037) );
  sky130_fd_sc_hd__nand2_1 U29235 ( .A(n24052), .B(n26971), .Y(n26615) );
  sky130_fd_sc_hd__o22ai_1 U29236 ( .A1(n26423), .A2(n24052), .B1(n26422), 
        .B2(n26702), .Y(n24032) );
  sky130_fd_sc_hd__a21oi_1 U29237 ( .A1(n24033), .A2(n25415), .B1(n24032), .Y(
        n24035) );
  sky130_fd_sc_hd__nand2_1 U29238 ( .A(n24038), .B(n26702), .Y(n26616) );
  sky130_fd_sc_hd__nand3_1 U29239 ( .A(n26616), .B(n26326), .C(n26615), .Y(
        n24034) );
  sky130_fd_sc_hd__o211ai_1 U29240 ( .A1(n26707), .A2(n26419), .B1(n24035), 
        .C1(n24034), .Y(n24036) );
  sky130_fd_sc_hd__nor2_1 U29241 ( .A(n24037), .B(n24036), .Y(n24042) );
  sky130_fd_sc_hd__o22a_1 U29242 ( .A1(n24038), .A2(n26431), .B1(n26582), .B2(
        n26412), .X(n24041) );
  sky130_fd_sc_hd__o22ai_1 U29243 ( .A1(n26705), .A2(n26427), .B1(n26578), 
        .B2(n26424), .Y(n24039) );
  sky130_fd_sc_hd__a21oi_1 U29244 ( .A1(n25131), .A2(n26859), .B1(n24039), .Y(
        n24040) );
  sky130_fd_sc_hd__nand4_1 U29245 ( .A(n24042), .B(n24041), .C(n24040), .D(
        n26411), .Y(n24043) );
  sky130_fd_sc_hd__a21oi_1 U29246 ( .A1(n24044), .A2(n26409), .B1(n24043), .Y(
        n24045) );
  sky130_fd_sc_hd__o22ai_1 U29247 ( .A1(n27575), .A2(n24055), .B1(n27574), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N3118) );
  sky130_fd_sc_hd__o22ai_1 U29248 ( .A1(n27219), .A2(n24055), .B1(n27218), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N3007) );
  sky130_fd_sc_hd__o22ai_1 U29249 ( .A1(n27217), .A2(n24055), .B1(n27216), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N2859) );
  sky130_fd_sc_hd__o22ai_1 U29250 ( .A1(n27466), .A2(n24055), .B1(n27465), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N2785) );
  sky130_fd_sc_hd__o22ai_1 U29251 ( .A1(n27213), .A2(n24055), .B1(n27212), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N2822) );
  sky130_fd_sc_hd__o22ai_1 U29252 ( .A1(n27221), .A2(n24055), .B1(n27220), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N2896) );
  sky130_fd_sc_hd__o22ai_1 U29253 ( .A1(n27209), .A2(n24055), .B1(n23039), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N2748) );
  sky130_fd_sc_hd__o22ai_1 U29254 ( .A1(n26378), .A2(n24055), .B1(n26449), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N3266) );
  sky130_fd_sc_hd__o22ai_1 U29255 ( .A1(n27225), .A2(n24055), .B1(n27224), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N2970) );
  sky130_fd_sc_hd__o22ai_1 U29256 ( .A1(n27215), .A2(n24055), .B1(n27214), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N2933) );
  sky130_fd_sc_hd__o22ai_1 U29257 ( .A1(n27223), .A2(n24055), .B1(n27222), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N3044) );
  sky130_fd_sc_hd__o22ai_1 U29258 ( .A1(n27211), .A2(n24055), .B1(n27210), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N3229) );
  sky130_fd_sc_hd__o22ai_1 U29259 ( .A1(n27228), .A2(n24055), .B1(n27227), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N3192) );
  sky130_fd_sc_hd__o22ai_1 U29260 ( .A1(n11141), .A2(n24055), .B1(n27124), 
        .B2(n11047), .Y(j202_soc_core_j22_cpu_rf_N2711) );
  sky130_fd_sc_hd__nand2_1 U29261 ( .A(n24052), .B(n27446), .Y(n24054) );
  sky130_fd_sc_hd__o211ai_1 U29263 ( .A1(n24055), .A2(n27450), .B1(n24054), 
        .C1(n27448), .Y(j202_soc_core_j22_cpu_ml_N368) );
  sky130_fd_sc_hd__o22ai_1 U29264 ( .A1(n28612), .A2(n25534), .B1(n24056), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U29265 ( .A1(n25858), .A2(n25534), .B1(n25863), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__a21oi_1 U29266 ( .A1(n25344), .A2(n22730), .B1(n26976), .Y(
        n24059) );
  sky130_fd_sc_hd__nand3_1 U29267 ( .A(n12356), .B(n24164), .C(n26872), .Y(
        n24057) );
  sky130_fd_sc_hd__nand3_1 U29268 ( .A(n12357), .B(n24062), .C(n26872), .Y(
        n24064) );
  sky130_fd_sc_hd__nand2b_1 U29269 ( .A_N(n24066), .B(n25181), .Y(n24090) );
  sky130_fd_sc_hd__a21oi_1 U29270 ( .A1(n26719), .A2(n26323), .B1(n24067), .Y(
        n24088) );
  sky130_fd_sc_hd__nand2_1 U29271 ( .A(n24072), .B(n25403), .Y(n26658) );
  sky130_fd_sc_hd__nand2_1 U29272 ( .A(n27425), .B(n26719), .Y(n26657) );
  sky130_fd_sc_hd__nand3_1 U29273 ( .A(n26658), .B(n26326), .C(n26657), .Y(
        n24069) );
  sky130_fd_sc_hd__nand2_1 U29274 ( .A(n26077), .B(n25130), .Y(n24068) );
  sky130_fd_sc_hd__o211ai_1 U29275 ( .A1(n26336), .A2(n26416), .B1(n24069), 
        .C1(n24068), .Y(n24071) );
  sky130_fd_sc_hd__o22ai_1 U29276 ( .A1(n25128), .A2(n26419), .B1(n26570), 
        .B2(n26418), .Y(n24070) );
  sky130_fd_sc_hd__nor2_1 U29277 ( .A(n24071), .B(n24070), .Y(n24081) );
  sky130_fd_sc_hd__o22a_1 U29278 ( .A1(n24072), .A2(n26431), .B1(n26792), .B2(
        n26412), .X(n24080) );
  sky130_fd_sc_hd__o22ai_1 U29279 ( .A1(n18916), .A2(n24073), .B1(n26423), 
        .B2(n27425), .Y(n24074) );
  sky130_fd_sc_hd__a21oi_1 U29280 ( .A1(n26085), .A2(n26719), .B1(n24074), .Y(
        n24075) );
  sky130_fd_sc_hd__o21ai_0 U29281 ( .A1(n26432), .A2(n26657), .B1(n24075), .Y(
        n24078) );
  sky130_fd_sc_hd__nor2_1 U29282 ( .A(n26417), .B(n26424), .Y(n24077) );
  sky130_fd_sc_hd__o22ai_1 U29283 ( .A1(n26571), .A2(n26427), .B1(n26713), 
        .B2(n26425), .Y(n24076) );
  sky130_fd_sc_hd__nor3_1 U29284 ( .A(n24078), .B(n24077), .C(n24076), .Y(
        n24079) );
  sky130_fd_sc_hd__nand4_1 U29285 ( .A(n24081), .B(n24080), .C(n26411), .D(
        n24079), .Y(n24082) );
  sky130_fd_sc_hd__o21bai_1 U29286 ( .A1(n18916), .A2(n24083), .B1_N(n24082), 
        .Y(n24084) );
  sky130_fd_sc_hd__a21oi_1 U29287 ( .A1(n24085), .A2(n26409), .B1(n24084), .Y(
        n24086) );
  sky130_fd_sc_hd__nor2_1 U29288 ( .A(n26946), .B(n12474), .Y(
        j202_soc_core_j22_cpu_rf_N2663) );
  sky130_fd_sc_hd__o22ai_1 U29289 ( .A1(n27221), .A2(n27427), .B1(n27220), 
        .B2(n12473), .Y(j202_soc_core_j22_cpu_rf_N2884) );
  sky130_fd_sc_hd__o22ai_1 U29290 ( .A1(n27427), .A2(n26899), .B1(n26898), 
        .B2(n12474), .Y(j202_soc_core_j22_cpu_rf_N3330) );
  sky130_fd_sc_hd__o22ai_1 U29291 ( .A1(n11141), .A2(n27427), .B1(n27124), 
        .B2(n12474), .Y(j202_soc_core_j22_cpu_rf_N2699) );
  sky130_fd_sc_hd__o22ai_1 U29292 ( .A1(n27209), .A2(n27427), .B1(n23039), 
        .B2(n12473), .Y(j202_soc_core_j22_cpu_rf_N2736) );
  sky130_fd_sc_hd__o22ai_1 U29293 ( .A1(n27213), .A2(n27427), .B1(n27212), 
        .B2(n12473), .Y(j202_soc_core_j22_cpu_rf_N2810) );
  sky130_fd_sc_hd__o22ai_1 U29294 ( .A1(n27211), .A2(n27427), .B1(n27210), 
        .B2(n12474), .Y(j202_soc_core_j22_cpu_rf_N3217) );
  sky130_fd_sc_hd__o22ai_1 U29295 ( .A1(n27223), .A2(n27427), .B1(n27222), 
        .B2(n12474), .Y(j202_soc_core_j22_cpu_rf_N3032) );
  sky130_fd_sc_hd__o22ai_1 U29296 ( .A1(n27215), .A2(n27427), .B1(n27214), 
        .B2(n12474), .Y(j202_soc_core_j22_cpu_rf_N2921) );
  sky130_fd_sc_hd__o22ai_1 U29297 ( .A1(n27466), .A2(n27427), .B1(n27465), 
        .B2(n12474), .Y(j202_soc_core_j22_cpu_rf_N2773) );
  sky130_fd_sc_hd__o22ai_1 U29298 ( .A1(n27225), .A2(n27427), .B1(n27224), 
        .B2(n12474), .Y(j202_soc_core_j22_cpu_rf_N2958) );
  sky130_fd_sc_hd__o22ai_1 U29299 ( .A1(n27228), .A2(n27427), .B1(n27227), 
        .B2(n12474), .Y(j202_soc_core_j22_cpu_rf_N3180) );
  sky130_fd_sc_hd__o22ai_1 U29300 ( .A1(n27217), .A2(n27427), .B1(n27216), 
        .B2(n12473), .Y(j202_soc_core_j22_cpu_rf_N2847) );
  sky130_fd_sc_hd__o22ai_1 U29301 ( .A1(n27219), .A2(n27427), .B1(n27218), 
        .B2(n12473), .Y(j202_soc_core_j22_cpu_rf_N2995) );
  sky130_fd_sc_hd__o22ai_1 U29302 ( .A1(n27333), .A2(n27427), .B1(n23178), 
        .B2(n12473), .Y(j202_soc_core_j22_cpu_rf_N3069) );
  sky130_fd_sc_hd__o22ai_1 U29303 ( .A1(n27575), .A2(n27427), .B1(n27574), 
        .B2(n12473), .Y(j202_soc_core_j22_cpu_rf_N3106) );
  sky130_fd_sc_hd__o22ai_1 U29304 ( .A1(n26378), .A2(n27427), .B1(n26449), 
        .B2(n12474), .Y(j202_soc_core_j22_cpu_rf_N3254) );
  sky130_fd_sc_hd__nand2_1 U29305 ( .A(n27947), .B(n27176), .Y(n24658) );
  sky130_fd_sc_hd__nand2b_1 U29306 ( .A_N(n27175), .B(n27904), .Y(n27967) );
  sky130_fd_sc_hd__nand2_1 U29307 ( .A(n27232), .B(n29071), .Y(n24098) );
  sky130_fd_sc_hd__nand2_1 U29308 ( .A(n23185), .B(n24095), .Y(n24639) );
  sky130_fd_sc_hd__nand3_1 U29309 ( .A(n27787), .B(n27942), .C(n27967), .Y(
        n24096) );
  sky130_fd_sc_hd__a211oi_1 U29310 ( .A1(n29036), .A2(n24639), .B1(n24096), 
        .C1(n27934), .Y(n24097) );
  sky130_fd_sc_hd__nand3_1 U29311 ( .A(n24098), .B(n24460), .C(n24097), .Y(
        n24099) );
  sky130_fd_sc_hd__inv_1 U29312 ( .A(n24704), .Y(n24101) );
  sky130_fd_sc_hd__nand3_1 U29313 ( .A(n24101), .B(n27980), .C(n13180), .Y(
        n24102) );
  sky130_fd_sc_hd__nand2_1 U29314 ( .A(n27934), .B(n27980), .Y(n27961) );
  sky130_fd_sc_hd__nand2b_1 U29315 ( .A_N(n27956), .B(n24103), .Y(n27969) );
  sky130_fd_sc_hd__nor2_1 U29316 ( .A(n23589), .B(n24357), .Y(n24104) );
  sky130_fd_sc_hd__nor2_1 U29317 ( .A(n24104), .B(n24327), .Y(n27168) );
  sky130_fd_sc_hd__nand3_1 U29318 ( .A(n27168), .B(n24106), .C(n24105), .Y(
        n24107) );
  sky130_fd_sc_hd__nor2_1 U29319 ( .A(n24108), .B(n24659), .Y(n24109) );
  sky130_fd_sc_hd__nand2_1 U29320 ( .A(n12472), .B(n27980), .Y(n24660) );
  sky130_fd_sc_hd__nand2_1 U29321 ( .A(n27882), .B(n25815), .Y(n24110) );
  sky130_fd_sc_hd__nand2_1 U29322 ( .A(n24112), .B(n24290), .Y(n24114) );
  sky130_fd_sc_hd__nor2_1 U29323 ( .A(n24114), .B(n24113), .Y(n27269) );
  sky130_fd_sc_hd__nand2_1 U29324 ( .A(n26812), .B(n24275), .Y(n27272) );
  sky130_fd_sc_hd__o22ai_1 U29325 ( .A1(n24116), .A2(n24115), .B1(n24278), 
        .B2(n27272), .Y(j202_soc_core_j22_cpu_ml_N155) );
  sky130_fd_sc_hd__nor2_1 U29326 ( .A(n27635), .B(n12458), .Y(
        j202_soc_core_ahb2aqu_00_N132) );
  sky130_fd_sc_hd__nor2_1 U29327 ( .A(n27634), .B(n12458), .Y(
        j202_soc_core_ahb2aqu_00_N133) );
  sky130_fd_sc_hd__nor2_1 U29328 ( .A(n27637), .B(n12458), .Y(
        j202_soc_core_ahb2aqu_00_N136) );
  sky130_fd_sc_hd__nor2_1 U29329 ( .A(n27638), .B(n12458), .Y(
        j202_soc_core_ahb2aqu_00_N135) );
  sky130_fd_sc_hd__nor2_1 U29330 ( .A(n27639), .B(n12458), .Y(
        j202_soc_core_ahb2aqu_00_N134) );
  sky130_fd_sc_hd__nor2_1 U29331 ( .A(n27636), .B(n12458), .Y(
        j202_soc_core_ahb2aqu_00_N131) );
  sky130_fd_sc_hd__a21oi_1 U29332 ( .A1(n29033), .A2(n27621), .B1(n27620), .Y(
        n24122) );
  sky130_fd_sc_hd__o21ai_1 U29333 ( .A1(n24119), .A2(n24118), .B1(n24117), .Y(
        n24121) );
  sky130_fd_sc_hd__nand2_1 U29334 ( .A(n28976), .B(n29061), .Y(n24120) );
  sky130_fd_sc_hd__nand4_1 U29335 ( .A(n25225), .B(n29347), .C(n12400), .D(
        n24123), .Y(n24126) );
  sky130_fd_sc_hd__nor3_1 U29336 ( .A(n12456), .B(n24126), .C(n24125), .Y(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_N487) );
  sky130_fd_sc_hd__a21oi_1 U29337 ( .A1(n25344), .A2(n24132), .B1(n26976), .Y(
        n24131) );
  sky130_fd_sc_hd__nand3_1 U29338 ( .A(n12916), .B(
        j202_soc_core_j22_cpu_ml_macl[3]), .C(n25826), .Y(n24130) );
  sky130_fd_sc_hd__nand3_1 U29339 ( .A(n12357), .B(n24128), .C(n26872), .Y(
        n24129) );
  sky130_fd_sc_hd__nand3_1 U29340 ( .A(n24131), .B(n24130), .C(n24129), .Y(
        j202_soc_core_j22_cpu_ml_maclj[3]) );
  sky130_fd_sc_hd__o211ai_1 U29341 ( .A1(n24137), .A2(n25338), .B1(n27273), 
        .C1(n24136), .Y(j202_soc_core_j22_cpu_ml_machj[3]) );
  sky130_fd_sc_hd__nor2_2 U29342 ( .A(n24139), .B(n24138), .Y(n25270) );
  sky130_fd_sc_hd__xnor2_1 U29343 ( .A(n26726), .B(n27354), .Y(n26669) );
  sky130_fd_sc_hd__o22a_1 U29344 ( .A1(n26415), .A2(n26669), .B1(n25128), .B2(
        n26418), .X(n24140) );
  sky130_fd_sc_hd__o211ai_1 U29345 ( .A1(n26708), .A2(n26419), .B1(n24141), 
        .C1(n24140), .Y(n24149) );
  sky130_fd_sc_hd__nand2_1 U29346 ( .A(n26338), .B(n27402), .Y(n24146) );
  sky130_fd_sc_hd__nand2_1 U29347 ( .A(n24143), .B(n24142), .Y(n24144) );
  sky130_fd_sc_hd__nand2_1 U29348 ( .A(n24144), .B(n26329), .Y(n24145) );
  sky130_fd_sc_hd__o211ai_1 U29349 ( .A1(n24778), .A2(n24147), .B1(n24146), 
        .C1(n24145), .Y(n24148) );
  sky130_fd_sc_hd__nor2_1 U29350 ( .A(n24149), .B(n24148), .Y(n24154) );
  sky130_fd_sc_hd__o22ai_1 U29351 ( .A1(n25798), .A2(n26416), .B1(n26565), 
        .B2(n26427), .Y(n24150) );
  sky130_fd_sc_hd__a21oi_1 U29352 ( .A1(n26341), .A2(n26859), .B1(n24150), .Y(
        n24153) );
  sky130_fd_sc_hd__mux2_2 U29353 ( .A0(n26423), .A1(n26349), .S(n27354), .X(
        n24152) );
  sky130_fd_sc_hd__nand2_1 U29354 ( .A(n26342), .B(n27347), .Y(n24151) );
  sky130_fd_sc_hd__nand4_1 U29355 ( .A(n24154), .B(n24153), .C(n24152), .D(
        n24151), .Y(n24155) );
  sky130_fd_sc_hd__a21oi_1 U29356 ( .A1(n24156), .A2(n26409), .B1(n24155), .Y(
        n24158) );
  sky130_fd_sc_hd__nand2_1 U29358 ( .A(n27354), .B(n25415), .Y(n24160) );
  sky130_fd_sc_hd__nand2_1 U29359 ( .A(n24160), .B(n26422), .Y(n24162) );
  sky130_fd_sc_hd__nor2_1 U29360 ( .A(n26946), .B(n12161), .Y(
        j202_soc_core_j22_cpu_rf_N2658) );
  sky130_fd_sc_hd__o22ai_1 U29361 ( .A1(n27219), .A2(n25276), .B1(n27218), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N2991) );
  sky130_fd_sc_hd__o22ai_1 U29362 ( .A1(n27226), .A2(n25276), .B1(n23079), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N3139) );
  sky130_fd_sc_hd__o22ai_1 U29363 ( .A1(n26378), .A2(n25276), .B1(n26449), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N3250) );
  sky130_fd_sc_hd__o22ai_1 U29364 ( .A1(n27217), .A2(n25276), .B1(n27216), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N2843) );
  sky130_fd_sc_hd__o22ai_1 U29365 ( .A1(n27466), .A2(n25276), .B1(n27465), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N2769) );
  sky130_fd_sc_hd__o22ai_1 U29366 ( .A1(n27213), .A2(n25276), .B1(n27212), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N2806) );
  sky130_fd_sc_hd__o22ai_1 U29367 ( .A1(n27221), .A2(n25276), .B1(n27220), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N2880) );
  sky130_fd_sc_hd__o22ai_1 U29368 ( .A1(n27209), .A2(n25276), .B1(n23039), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N2732) );
  sky130_fd_sc_hd__o22ai_1 U29369 ( .A1(n27333), .A2(n25276), .B1(n23178), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N3065) );
  sky130_fd_sc_hd__o22ai_1 U29370 ( .A1(n25276), .A2(n26899), .B1(n26898), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N3326) );
  sky130_fd_sc_hd__o22ai_1 U29371 ( .A1(n11141), .A2(n27356), .B1(n27124), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N2695) );
  sky130_fd_sc_hd__o22ai_1 U29372 ( .A1(n27223), .A2(n25276), .B1(n27222), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N3028) );
  sky130_fd_sc_hd__o22ai_1 U29373 ( .A1(n27215), .A2(n27356), .B1(n27214), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N2917) );
  sky130_fd_sc_hd__o22ai_1 U29374 ( .A1(n27211), .A2(n25276), .B1(n27210), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N3213) );
  sky130_fd_sc_hd__o22ai_1 U29375 ( .A1(n27228), .A2(n27356), .B1(n27227), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N3176) );
  sky130_fd_sc_hd__o22ai_1 U29376 ( .A1(n27225), .A2(n25276), .B1(n27224), 
        .B2(n12161), .Y(j202_soc_core_j22_cpu_rf_N2954) );
  sky130_fd_sc_hd__nand2b_1 U29377 ( .A_N(n12917), .B(n24164), .Y(n24165) );
  sky130_fd_sc_hd__o211ai_1 U29378 ( .A1(n24628), .A2(n26981), .B1(n25822), 
        .C1(n24165), .Y(j202_soc_core_j22_cpu_ml_maclj[17]) );
  sky130_fd_sc_hd__nor2_1 U29379 ( .A(n24168), .B(n24167), .Y(n26807) );
  sky130_fd_sc_hd__o211ai_1 U29380 ( .A1(n26807), .A2(n27274), .B1(n27273), 
        .C1(n12356), .Y(j202_soc_core_j22_cpu_ml_machj[0]) );
  sky130_fd_sc_hd__nand2_1 U29381 ( .A(n12999), .B(n24602), .Y(n24170) );
  sky130_fd_sc_hd__o211ai_1 U29382 ( .A1(n26981), .A2(n24171), .B1(n25822), 
        .C1(n24170), .Y(j202_soc_core_j22_cpu_ml_maclj[16]) );
  sky130_fd_sc_hd__nand2_1 U29383 ( .A(n27648), .B(n29594), .Y(n29234) );
  sky130_fd_sc_hd__nand3_1 U29384 ( .A(n26946), .B(n29593), .C(n24643), .Y(
        n29235) );
  sky130_fd_sc_hd__nand2_1 U29385 ( .A(n24172), .B(n29594), .Y(n29238) );
  sky130_fd_sc_hd__nand2_1 U29386 ( .A(n27659), .B(
        j202_soc_core_gpio_core_00_reg_addr[4]), .Y(n27654) );
  sky130_fd_sc_hd__buf_6 U29387 ( .A(n13276), .X(n29251) );
  sky130_fd_sc_hd__buf_6 U29388 ( .A(n13276), .X(n29252) );
  sky130_fd_sc_hd__nand2_1 U29389 ( .A(n28978), .B(n27824), .Y(n24174) );
  sky130_fd_sc_hd__buf_6 U29390 ( .A(n24175), .X(n29253) );
  sky130_fd_sc_hd__nand2_1 U29391 ( .A(n28979), .B(n24225), .Y(n24176) );
  sky130_fd_sc_hd__buf_6 U29392 ( .A(n24177), .X(n29255) );
  sky130_fd_sc_hd__buf_6 U29393 ( .A(n24177), .X(n29256) );
  sky130_fd_sc_hd__buf_6 U29394 ( .A(n24179), .X(n29257) );
  sky130_fd_sc_hd__buf_6 U29395 ( .A(n24179), .X(n29258) );
  sky130_fd_sc_hd__nand2_1 U29396 ( .A(n28982), .B(n24225), .Y(n24182) );
  sky130_fd_sc_hd__buf_6 U29397 ( .A(n24183), .X(n29261) );
  sky130_fd_sc_hd__buf_6 U29398 ( .A(n24183), .X(n29262) );
  sky130_fd_sc_hd__nand2_1 U29399 ( .A(n28983), .B(n27824), .Y(n24184) );
  sky130_fd_sc_hd__inv_2 U29400 ( .A(n24184), .Y(n24185) );
  sky130_fd_sc_hd__buf_6 U29401 ( .A(n24185), .X(n29263) );
  sky130_fd_sc_hd__buf_6 U29402 ( .A(n24185), .X(n29264) );
  sky130_fd_sc_hd__nand2_1 U29403 ( .A(n28984), .B(n24225), .Y(n24186) );
  sky130_fd_sc_hd__buf_6 U29404 ( .A(n24187), .X(n29265) );
  sky130_fd_sc_hd__buf_6 U29405 ( .A(n24187), .X(n29266) );
  sky130_fd_sc_hd__buf_4 U29406 ( .A(n24190), .X(n29269) );
  sky130_fd_sc_hd__buf_4 U29407 ( .A(n24190), .X(n29270) );
  sky130_fd_sc_hd__buf_6 U29409 ( .A(n29571), .X(n29271) );
  sky130_fd_sc_hd__buf_6 U29410 ( .A(n29571), .X(n29272) );
  sky130_fd_sc_hd__nand2_1 U29411 ( .A(n28988), .B(n24225), .Y(n24193) );
  sky130_fd_sc_hd__buf_6 U29412 ( .A(n24194), .X(n29273) );
  sky130_fd_sc_hd__buf_6 U29413 ( .A(n24194), .X(n29274) );
  sky130_fd_sc_hd__nand2_1 U29414 ( .A(n28989), .B(n24225), .Y(n24195) );
  sky130_fd_sc_hd__buf_6 U29415 ( .A(n24196), .X(n29275) );
  sky130_fd_sc_hd__buf_6 U29416 ( .A(n24196), .X(n29276) );
  sky130_fd_sc_hd__nand2_1 U29417 ( .A(n28990), .B(n24225), .Y(n24197) );
  sky130_fd_sc_hd__buf_6 U29418 ( .A(n24198), .X(n29277) );
  sky130_fd_sc_hd__nand2_1 U29419 ( .A(n28991), .B(n24225), .Y(n24199) );
  sky130_fd_sc_hd__buf_6 U29420 ( .A(n24200), .X(n29279) );
  sky130_fd_sc_hd__buf_6 U29421 ( .A(n24200), .X(n29280) );
  sky130_fd_sc_hd__nand2_1 U29422 ( .A(n28992), .B(n24225), .Y(n24201) );
  sky130_fd_sc_hd__buf_4 U29423 ( .A(n24202), .X(n29281) );
  sky130_fd_sc_hd__buf_4 U29424 ( .A(n24202), .X(n29282) );
  sky130_fd_sc_hd__buf_6 U29427 ( .A(n24203), .X(n29285) );
  sky130_fd_sc_hd__buf_6 U29428 ( .A(n24203), .X(n29286) );
  sky130_fd_sc_hd__buf_6 U29429 ( .A(n24204), .X(n29287) );
  sky130_fd_sc_hd__buf_6 U29430 ( .A(n24204), .X(n29288) );
  sky130_fd_sc_hd__buf_6 U29431 ( .A(n24205), .X(n29289) );
  sky130_fd_sc_hd__buf_6 U29432 ( .A(n24205), .X(n29290) );
  sky130_fd_sc_hd__nand2_1 U29433 ( .A(n28997), .B(n27824), .Y(n24206) );
  sky130_fd_sc_hd__buf_6 U29434 ( .A(n24207), .X(n29291) );
  sky130_fd_sc_hd__buf_6 U29435 ( .A(n24207), .X(n29292) );
  sky130_fd_sc_hd__buf_4 U29436 ( .A(n11080), .X(n29293) );
  sky130_fd_sc_hd__buf_4 U29437 ( .A(n11080), .X(n29294) );
  sky130_fd_sc_hd__buf_6 U29438 ( .A(n24209), .X(n29295) );
  sky130_fd_sc_hd__buf_6 U29439 ( .A(n24209), .X(n29296) );
  sky130_fd_sc_hd__nand2_1 U29440 ( .A(n29000), .B(n27824), .Y(n24211) );
  sky130_fd_sc_hd__buf_6 U29441 ( .A(n24212), .X(n29297) );
  sky130_fd_sc_hd__buf_6 U29442 ( .A(n24212), .X(n29298) );
  sky130_fd_sc_hd__nand2_1 U29443 ( .A(n29001), .B(n11127), .Y(n24213) );
  sky130_fd_sc_hd__buf_6 U29444 ( .A(n24214), .X(n29299) );
  sky130_fd_sc_hd__buf_6 U29445 ( .A(n24214), .X(n29300) );
  sky130_fd_sc_hd__nand2_1 U29446 ( .A(n29002), .B(n27824), .Y(n24215) );
  sky130_fd_sc_hd__buf_6 U29447 ( .A(n24216), .X(n29301) );
  sky130_fd_sc_hd__nand2_1 U29448 ( .A(n29003), .B(n24225), .Y(n24217) );
  sky130_fd_sc_hd__buf_6 U29449 ( .A(n24218), .X(n29302) );
  sky130_fd_sc_hd__buf_6 U29450 ( .A(n24218), .X(n29303) );
  sky130_fd_sc_hd__nand2_1 U29451 ( .A(n29004), .B(n24225), .Y(n24219) );
  sky130_fd_sc_hd__buf_6 U29452 ( .A(n24220), .X(n29304) );
  sky130_fd_sc_hd__buf_6 U29453 ( .A(n24222), .X(n29306) );
  sky130_fd_sc_hd__buf_6 U29456 ( .A(n29570), .X(n29308) );
  sky130_fd_sc_hd__buf_6 U29457 ( .A(n29570), .X(n29309) );
  sky130_fd_sc_hd__nand2_1 U29458 ( .A(n29007), .B(n24225), .Y(n24226) );
  sky130_fd_sc_hd__buf_6 U29459 ( .A(n24227), .X(n29310) );
  sky130_fd_sc_hd__buf_6 U29460 ( .A(n24227), .X(n29311) );
  sky130_fd_sc_hd__nand2_1 U29461 ( .A(n24228), .B(n28776), .Y(
        j202_soc_core_uart_TOP_N24) );
  sky130_fd_sc_hd__xnor2_1 U29462 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .Y(n24229) );
  sky130_fd_sc_hd__nor2_1 U29463 ( .A(n24229), .B(n24233), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[1]) );
  sky130_fd_sc_hd__and3_1 U29464 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[2]), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .C(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .X(n24232) );
  sky130_fd_sc_hd__a2bb2oi_1 U29465 ( .B1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[2]), .B2(n28581), .A1_N(
        n24230), .A2_N(n29008), .Y(n24231) );
  sky130_fd_sc_hd__nor2_1 U29466 ( .A(n24232), .B(n24231), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[2]) );
  sky130_fd_sc_hd__nand2_1 U29467 ( .A(n24232), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[3]), .Y(n24236) );
  sky130_fd_sc_hd__nor2_1 U29469 ( .A(n24234), .B(n24233), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[3]) );
  sky130_fd_sc_hd__nor2_1 U29470 ( .A(n24237), .B(n24236), .Y(n24241) );
  sky130_fd_sc_hd__nand2_1 U29471 ( .A(n24235), .B(n28581), .Y(n24239) );
  sky130_fd_sc_hd__a21oi_1 U29472 ( .A1(n24237), .A2(n24236), .B1(n24239), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[4]) );
  sky130_fd_sc_hd__nand3_1 U29473 ( .A(n28581), .B(n24241), .C(n24240), .Y(
        n24238) );
  sky130_fd_sc_hd__o21ai_1 U29474 ( .A1(n24240), .A2(n24239), .B1(n24238), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[5]) );
  sky130_fd_sc_hd__nand3_1 U29475 ( .A(n28581), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]), .C(n24241), .Y(
        n24244) );
  sky130_fd_sc_hd__nand3_1 U29476 ( .A(n24244), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .C(n28581), .Y(
        n24242) );
  sky130_fd_sc_hd__o21ai_1 U29477 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .A2(n24244), .B1(
        n24242), .Y(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[6]) );
  sky130_fd_sc_hd__nand2_1 U29478 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .Y(n24243) );
  sky130_fd_sc_hd__nor2_1 U29479 ( .A(n24243), .B(n24244), .Y(n24249) );
  sky130_fd_sc_hd__a22oi_1 U29480 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]), .A2(n28581), .B1(
        n24245), .B2(j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .Y(
        n24246) );
  sky130_fd_sc_hd__nor2_1 U29481 ( .A(n24249), .B(n24246), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[7]) );
  sky130_fd_sc_hd__nand3_1 U29482 ( .A(n24248), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .C(n28581), .Y(
        n24247) );
  sky130_fd_sc_hd__o21ai_1 U29483 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .A2(n24248), .B1(
        n24247), .Y(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[8]) );
  sky130_fd_sc_hd__a22oi_1 U29484 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]), .A2(n28581), .B1(
        n24249), .B2(j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .Y(
        n24250) );
  sky130_fd_sc_hd__and3_1 U29485 ( .A(n24249), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .C(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]), .X(n27985) );
  sky130_fd_sc_hd__nor2_1 U29486 ( .A(n24250), .B(n27985), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[9]) );
  sky130_fd_sc_hd__nand3_1 U29487 ( .A(n24252), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .C(n28581), .Y(
        n24251) );
  sky130_fd_sc_hd__o21ai_1 U29488 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .A2(n24252), .B1(
        n24251), .Y(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[10]) );
  sky130_fd_sc_hd__nand2_1 U29489 ( .A(n24253), .B(n24266), .Y(n24255) );
  sky130_fd_sc_hd__a21oi_1 U29490 ( .A1(n24255), .A2(n27980), .B1(n24254), .Y(
        n24259) );
  sky130_fd_sc_hd__o211ai_1 U29492 ( .A1(n29569), .A2(n24257), .B1(n27980), 
        .C1(n12641), .Y(n24258) );
  sky130_fd_sc_hd__nand2_1 U29493 ( .A(n24259), .B(n24258), .Y(n10588) );
  sky130_fd_sc_hd__nor2_1 U29494 ( .A(n24260), .B(n27175), .Y(n24703) );
  sky130_fd_sc_hd__o21ai_0 U29495 ( .A1(n27928), .A2(n24455), .B1(n24270), .Y(
        n10590) );
  sky130_fd_sc_hd__nand2_1 U29496 ( .A(n11798), .B(n12482), .Y(n27565) );
  sky130_fd_sc_hd__nand3_1 U29497 ( .A(n13236), .B(n24262), .C(n24261), .Y(
        n24263) );
  sky130_fd_sc_hd__nand3_1 U29498 ( .A(n12732), .B(n24265), .C(n29532), .Y(
        n24267) );
  sky130_fd_sc_hd__o211ai_1 U29499 ( .A1(n27230), .A2(n11833), .B1(n24267), 
        .C1(n24266), .Y(n24268) );
  sky130_fd_sc_hd__o21ai_1 U29500 ( .A1(n24269), .A2(n24268), .B1(n27980), .Y(
        n24271) );
  sky130_fd_sc_hd__nand2_1 U29501 ( .A(n24271), .B(n24270), .Y(n10586) );
  sky130_fd_sc_hd__nor3_1 U29502 ( .A(n26398), .B(n24273), .C(n24272), .Y(
        n24281) );
  sky130_fd_sc_hd__or4_1 U29503 ( .A(n24275), .B(n24281), .C(n12200), .D(
        n24274), .X(n27337) );
  sky130_fd_sc_hd__and3_1 U29504 ( .A(n24276), .B(
        j202_soc_core_j22_cpu_rfuo_sr__s_), .C(n26398), .X(n24277) );
  sky130_fd_sc_hd__nand4b_1 U29505 ( .A_N(n12200), .B(
        j202_soc_core_j22_cpu_macop_MAC_[3]), .C(
        j202_soc_core_j22_cpu_macop_MAC_[2]), .D(n24277), .Y(n27336) );
  sky130_fd_sc_hd__nand2_1 U29507 ( .A(n27720), .B(n29347), .Y(n27267) );
  sky130_fd_sc_hd__nor2_1 U29508 ( .A(n24279), .B(n27267), .Y(
        j202_soc_core_j22_cpu_ma_N55) );
  sky130_fd_sc_hd__nor2_1 U29509 ( .A(n24280), .B(n27267), .Y(
        j202_soc_core_j22_cpu_ma_N56) );
  sky130_fd_sc_hd__nand2_1 U29510 ( .A(j202_soc_core_ahbcs_6__HREADY_), .B(
        n24281), .Y(n24289) );
  sky130_fd_sc_hd__o211ai_1 U29511 ( .A1(n24288), .A2(n27337), .B1(n27336), 
        .C1(n24289), .Y(j202_soc_core_j22_cpu_ml_N192) );
  sky130_fd_sc_hd__o21ai_1 U29512 ( .A1(n26398), .A2(n27337), .B1(n27336), .Y(
        j202_soc_core_j22_cpu_ml_N191) );
  sky130_fd_sc_hd__a21oi_1 U29514 ( .A1(n27269), .A2(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]), .B1(n24283), .Y(n24284) );
  sky130_fd_sc_hd__a21oi_1 U29517 ( .A1(n27269), .A2(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .B1(n24286), .Y(n24287) );
  sky130_fd_sc_hd__a31oi_1 U29520 ( .A1(n24291), .A2(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[4]), .A3(n24290), .B1(n27456), 
        .Y(n24292) );
  sky130_fd_sc_hd__o21ai_1 U29521 ( .A1(n24293), .A2(n27272), .B1(n24292), .Y(
        j202_soc_core_j22_cpu_ml_N156) );
  sky130_fd_sc_hd__nand2_1 U29522 ( .A(n24294), .B(n27957), .Y(n24295) );
  sky130_fd_sc_hd__nand3_1 U29523 ( .A(n12598), .B(n24386), .C(n11626), .Y(
        n24299) );
  sky130_fd_sc_hd__o21a_1 U29524 ( .A1(n11675), .A2(n24307), .B1(n24299), .X(
        n24301) );
  sky130_fd_sc_hd__nand2_1 U29525 ( .A(n24302), .B(n27176), .Y(n10578) );
  sky130_fd_sc_hd__nand2_1 U29526 ( .A(n24303), .B(n27956), .Y(n10574) );
  sky130_fd_sc_hd__nand2_1 U29527 ( .A(n12376), .B(n27980), .Y(n24304) );
  sky130_fd_sc_hd__nand2_1 U29528 ( .A(n24304), .B(n27956), .Y(n10575) );
  sky130_fd_sc_hd__nand2_1 U29529 ( .A(n29077), .B(n27980), .Y(n24305) );
  sky130_fd_sc_hd__nand2_1 U29530 ( .A(n24305), .B(n27956), .Y(n10576) );
  sky130_fd_sc_hd__nand2_1 U29531 ( .A(n29009), .B(n27980), .Y(n24306) );
  sky130_fd_sc_hd__nand2_1 U29532 ( .A(n24306), .B(n27956), .Y(n10577) );
  sky130_fd_sc_hd__inv_1 U29533 ( .A(n27783), .Y(n27938) );
  sky130_fd_sc_hd__a21oi_1 U29534 ( .A1(n24310), .A2(n12729), .B1(n12511), .Y(
        n24311) );
  sky130_fd_sc_hd__nand2_1 U29535 ( .A(n27938), .B(n24311), .Y(n24313) );
  sky130_fd_sc_hd__nand2_1 U29536 ( .A(n27947), .B(n27969), .Y(n24312) );
  sky130_fd_sc_hd__a21oi_1 U29537 ( .A1(n24313), .A2(n27980), .B1(n24312), .Y(
        n24314) );
  sky130_fd_sc_hd__nand2_1 U29539 ( .A(n24316), .B(
        j202_soc_core_ahb2apb_02_state[0]), .Y(n24318) );
  sky130_fd_sc_hd__nor3_1 U29540 ( .A(n28590), .B(n24315), .C(n24318), .Y(
        j202_soc_core_ahb2apb_02_N91) );
  sky130_fd_sc_hd__nor3_1 U29541 ( .A(j202_soc_core_ahb2apb_02_state[1]), .B(
        n28590), .C(n24318), .Y(j202_soc_core_ahb2apb_02_N90) );
  sky130_fd_sc_hd__nand2_1 U29542 ( .A(n24319), .B(
        j202_soc_core_ahb2apb_01_state[0]), .Y(n24323) );
  sky130_fd_sc_hd__nor3_1 U29543 ( .A(n28590), .B(n24320), .C(n24323), .Y(
        j202_soc_core_ahb2apb_01_N91) );
  sky130_fd_sc_hd__nor2_1 U29544 ( .A(j202_soc_core_ahb2apb_01_state[2]), .B(
        n24321), .Y(n24322) );
  sky130_fd_sc_hd__nor3_1 U29545 ( .A(j202_soc_core_ahb2apb_01_state[1]), .B(
        n28590), .C(n24323), .Y(j202_soc_core_ahb2apb_01_N90) );
  sky130_fd_sc_hd__nand2_1 U29546 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[0]), 
        .B(j202_soc_core_ahb2apb_01_hsize_buf[1]), .Y(
        j202_soc_core_ahb2apb_01_N123) );
  sky130_fd_sc_hd__nand3_1 U29547 ( .A(n12665), .B(n27957), .C(n24324), .Y(
        n24326) );
  sky130_fd_sc_hd__nor2_1 U29548 ( .A(n24328), .B(n24327), .Y(n24348) );
  sky130_fd_sc_hd__inv_1 U29549 ( .A(n12511), .Y(n24329) );
  sky130_fd_sc_hd__nand4_1 U29550 ( .A(n24330), .B(n24348), .C(n24402), .D(
        n24329), .Y(n24331) );
  sky130_fd_sc_hd__mux2i_1 U29551 ( .A0(n27064), .A1(n25789), .S(n27006), .Y(
        j202_soc_core_j22_cpu_ml_N303) );
  sky130_fd_sc_hd__nand2_1 U29552 ( .A(n24340), .B(n12060), .Y(n24334) );
  sky130_fd_sc_hd__nand3_1 U29553 ( .A(n12475), .B(n12482), .C(n29036), .Y(
        n24333) );
  sky130_fd_sc_hd__o211ai_1 U29554 ( .A1(n12376), .A2(n27892), .B1(n27564), 
        .C1(n27171), .Y(n24339) );
  sky130_fd_sc_hd__nand2_1 U29556 ( .A(n24340), .B(n23589), .Y(n27563) );
  sky130_fd_sc_hd__nand2_1 U29557 ( .A(n24342), .B(n27980), .Y(n24344) );
  sky130_fd_sc_hd__nand2_1 U29558 ( .A(n27264), .B(n27978), .Y(n27695) );
  sky130_fd_sc_hd__nor2_1 U29559 ( .A(n24343), .B(n27956), .Y(n27979) );
  sky130_fd_sc_hd__nand3_1 U29560 ( .A(n24344), .B(n27695), .C(n27599), .Y(
        n10596) );
  sky130_fd_sc_hd__nand2_1 U29561 ( .A(n11048), .B(n24345), .Y(n24346) );
  sky130_fd_sc_hd__nand2_1 U29562 ( .A(n24346), .B(n27980), .Y(n24366) );
  sky130_fd_sc_hd__nand2_1 U29563 ( .A(n24348), .B(n24347), .Y(n27571) );
  sky130_fd_sc_hd__nand2_1 U29564 ( .A(n12475), .B(n12731), .Y(n24349) );
  sky130_fd_sc_hd__o211ai_1 U29565 ( .A1(n25048), .A2(n27892), .B1(n27564), 
        .C1(n24349), .Y(n24359) );
  sky130_fd_sc_hd__nand2_1 U29566 ( .A(n12060), .B(n12376), .Y(n27889) );
  sky130_fd_sc_hd__nor2_1 U29567 ( .A(n13317), .B(n24351), .Y(n24352) );
  sky130_fd_sc_hd__nand2_1 U29568 ( .A(n24352), .B(n13274), .Y(n24355) );
  sky130_fd_sc_hd__o211ai_1 U29569 ( .A1(n27889), .A2(n24357), .B1(n27877), 
        .C1(n24356), .Y(n24358) );
  sky130_fd_sc_hd__nor2_1 U29570 ( .A(n24359), .B(n24358), .Y(n24362) );
  sky130_fd_sc_hd__nand3_1 U29571 ( .A(n13236), .B(n12461), .C(n12598), .Y(
        n27690) );
  sky130_fd_sc_hd__nor2_1 U29572 ( .A(n27565), .B(n27690), .Y(n27595) );
  sky130_fd_sc_hd__nand2_1 U29573 ( .A(n27595), .B(n27230), .Y(n24361) );
  sky130_fd_sc_hd__nand3b_1 U29574 ( .A_N(n27571), .B(n24362), .C(n24361), .Y(
        n24363) );
  sky130_fd_sc_hd__nand2_1 U29575 ( .A(n24363), .B(n27980), .Y(n24365) );
  sky130_fd_sc_hd__nand2_1 U29576 ( .A(n27979), .B(
        j202_soc_core_j22_cpu_opst[0]), .Y(n27265) );
  sky130_fd_sc_hd__nand3_1 U29577 ( .A(n24365), .B(n24366), .C(n27177), .Y(
        n10595) );
  sky130_fd_sc_hd__nand2_1 U29578 ( .A(n24370), .B(n27273), .Y(
        j202_soc_core_j22_cpu_ml_machj[4]) );
  sky130_fd_sc_hd__a21oi_1 U29579 ( .A1(n24373), .A2(n24372), .B1(n26865), .Y(
        n24374) );
  sky130_fd_sc_hd__a21oi_1 U29580 ( .A1(n18672), .A2(n27187), .B1(n24374), .Y(
        n24375) );
  sky130_fd_sc_hd__nand2_1 U29581 ( .A(n27189), .B(n24375), .Y(
        j202_soc_core_j22_cpu_ml_machj[29]) );
  sky130_fd_sc_hd__nand2_1 U29582 ( .A(n24377), .B(j202_soc_core_uart_RDRXD1), 
        .Y(n27141) );
  sky130_fd_sc_hd__nor2_1 U29583 ( .A(n27137), .B(n27141), .Y(n27131) );
  sky130_fd_sc_hd__o22ai_1 U29584 ( .A1(n24379), .A2(n27141), .B1(n24378), 
        .B2(n27131), .Y(n93) );
  sky130_fd_sc_hd__mux2i_1 U29585 ( .A0(n27417), .A1(n26577), .S(n27006), .Y(
        j202_soc_core_j22_cpu_ml_N308) );
  sky130_fd_sc_hd__nand2_4 U29586 ( .A(n24384), .B(n24383), .Y(n26915) );
  sky130_fd_sc_hd__nor2_1 U29587 ( .A(n26946), .B(n26915), .Y(
        j202_soc_core_j22_cpu_rf_N2647) );
  sky130_fd_sc_hd__nand2_1 U29588 ( .A(n24387), .B(n24386), .Y(n24390) );
  sky130_fd_sc_hd__nand4_1 U29589 ( .A(n11867), .B(n24390), .C(n24389), .D(
        n24388), .Y(n24392) );
  sky130_fd_sc_hd__nand2_1 U29590 ( .A(n24392), .B(n27980), .Y(n24398) );
  sky130_fd_sc_hd__nand2b_1 U29591 ( .A_N(n27956), .B(n24394), .Y(n27954) );
  sky130_fd_sc_hd__nand2b_1 U29593 ( .A_N(n27264), .B(n27599), .Y(n27820) );
  sky130_fd_sc_hd__nor2_1 U29594 ( .A(n24396), .B(n27820), .Y(n24397) );
  sky130_fd_sc_hd__nand2_1 U29595 ( .A(n24398), .B(n24397), .Y(n10489) );
  sky130_fd_sc_hd__nand2_1 U29596 ( .A(n29534), .B(n11626), .Y(n27894) );
  sky130_fd_sc_hd__nand3_1 U29597 ( .A(n24400), .B(n12598), .C(n24399), .Y(
        n24401) );
  sky130_fd_sc_hd__nand3_1 U29598 ( .A(n27894), .B(n24402), .C(n24401), .Y(
        n24403) );
  sky130_fd_sc_hd__nand2_1 U29599 ( .A(n24403), .B(n27980), .Y(n24406) );
  sky130_fd_sc_hd__nand3_1 U29600 ( .A(n27961), .B(n24406), .C(n24405), .Y(
        n10488) );
  sky130_fd_sc_hd__nor3_1 U29601 ( .A(n24408), .B(n24407), .C(n27820), .Y(
        n24413) );
  sky130_fd_sc_hd__nand2_1 U29602 ( .A(n12377), .B(n24411), .Y(n24702) );
  sky130_fd_sc_hd__o211ai_1 U29603 ( .A1(n24414), .A2(n27928), .B1(n24413), 
        .C1(n24412), .Y(n10490) );
  sky130_fd_sc_hd__nand2_1 U29604 ( .A(n24415), .B(n27947), .Y(n10605) );
  sky130_fd_sc_hd__mux2i_1 U29605 ( .A0(n26915), .A1(n27417), .S(n27460), .Y(
        j202_soc_core_j22_cpu_rf_N3275) );
  sky130_fd_sc_hd__nand2_1 U29606 ( .A(n12729), .B(n29569), .Y(n24435) );
  sky130_fd_sc_hd__nand2_1 U29607 ( .A(n24418), .B(n27980), .Y(n24419) );
  sky130_fd_sc_hd__nand2_1 U29608 ( .A(n24419), .B(n27942), .Y(n10600) );
  sky130_fd_sc_hd__inv_1 U29609 ( .A(n29514), .Y(n24422) );
  sky130_fd_sc_hd__nand4_1 U29610 ( .A(n27782), .B(n24422), .C(n24421), .D(
        n27261), .Y(n24426) );
  sky130_fd_sc_hd__inv_1 U29611 ( .A(n24423), .Y(n27822) );
  sky130_fd_sc_hd__nand2_1 U29613 ( .A(n24427), .B(n27942), .Y(n10602) );
  sky130_fd_sc_hd__nor2_1 U29614 ( .A(n28590), .B(n27919), .Y(n27951) );
  sky130_fd_sc_hd__nand3_1 U29615 ( .A(n14849), .B(n24429), .C(n24428), .Y(
        n24431) );
  sky130_fd_sc_hd__nand2_1 U29616 ( .A(n24431), .B(n24430), .Y(n24434) );
  sky130_fd_sc_hd__nor2_1 U29617 ( .A(n24432), .B(n24434), .Y(n29362) );
  sky130_fd_sc_hd__nand2_1 U29618 ( .A(n29362), .B(n26812), .Y(n24443) );
  sky130_fd_sc_hd__nor2_1 U29619 ( .A(n24433), .B(n24443), .Y(
        j202_soc_core_j22_cpu_id_idec_N958) );
  sky130_fd_sc_hd__nand2_1 U29620 ( .A(n24434), .B(n27951), .Y(n10561) );
  sky130_fd_sc_hd__o21ai_1 U29622 ( .A1(n24439), .A2(n24438), .B1(n27980), .Y(
        n24440) );
  sky130_fd_sc_hd__nand3_1 U29623 ( .A(n24440), .B(n13303), .C(n27954), .Y(
        n10601) );
  sky130_fd_sc_hd__nor2_1 U29624 ( .A(n24441), .B(n24443), .Y(
        j202_soc_core_j22_cpu_id_idec_N957) );
  sky130_fd_sc_hd__nor2_1 U29625 ( .A(n24442), .B(n24443), .Y(
        j202_soc_core_j22_cpu_id_idec_N959) );
  sky130_fd_sc_hd__nor2_1 U29626 ( .A(n24444), .B(n24443), .Y(
        j202_soc_core_j22_cpu_id_idec_N956) );
  sky130_fd_sc_hd__o22ai_1 U29627 ( .A1(n27417), .A2(n26378), .B1(n26449), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N3238) );
  sky130_fd_sc_hd__nor2_1 U29628 ( .A(n24446), .B(n24445), .Y(n24450) );
  sky130_fd_sc_hd__nor2_1 U29629 ( .A(n24448), .B(n12485), .Y(n24449) );
  sky130_fd_sc_hd__nor2_1 U29630 ( .A(n24453), .B(n27925), .Y(n24454) );
  sky130_fd_sc_hd__nor3_1 U29631 ( .A(n24457), .B(n27568), .C(n12679), .Y(
        n24459) );
  sky130_fd_sc_hd__nand4_1 U29632 ( .A(n24461), .B(n24460), .C(n24459), .D(
        n24458), .Y(n24462) );
  sky130_fd_sc_hd__nand2_1 U29633 ( .A(n24462), .B(n27980), .Y(n24463) );
  sky130_fd_sc_hd__nand2_1 U29634 ( .A(n24463), .B(n27947), .Y(n10606) );
  sky130_fd_sc_hd__nor2_1 U29635 ( .A(n26946), .B(n27063), .Y(
        j202_soc_core_j22_cpu_rf_N2642) );
  sky130_fd_sc_hd__o22ai_1 U29636 ( .A1(n27064), .A2(n26378), .B1(n26449), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N3233) );
  sky130_fd_sc_hd__nand3_1 U29637 ( .A(n24468), .B(n29493), .C(n24466), .Y(
        n24473) );
  sky130_fd_sc_hd__a21oi_1 U29638 ( .A1(n24470), .A2(n24469), .B1(n27906), .Y(
        n24472) );
  sky130_fd_sc_hd__o31ai_1 U29639 ( .A1(n24473), .A2(n24472), .A3(n24471), 
        .B1(n12142), .Y(n10559) );
  sky130_fd_sc_hd__nand2_1 U29640 ( .A(n27601), .B(n24474), .Y(n10608) );
  sky130_fd_sc_hd__nand2_1 U29641 ( .A(n29347), .B(n24475), .Y(n24476) );
  sky130_fd_sc_hd__nor2_1 U29642 ( .A(n24476), .B(n14849), .Y(
        j202_soc_core_j22_cpu_N8) );
  sky130_fd_sc_hd__o22ai_1 U29643 ( .A1(n27064), .A2(n26899), .B1(n26898), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N3307) );
  sky130_fd_sc_hd__o22ai_1 U29644 ( .A1(n27064), .A2(n11141), .B1(n27124), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N2678) );
  sky130_fd_sc_hd__nand2_1 U29645 ( .A(n26515), .B(n26513), .Y(n24477) );
  sky130_fd_sc_hd__nand2_1 U29646 ( .A(n24477), .B(n26329), .Y(n24495) );
  sky130_fd_sc_hd__nand2_1 U29647 ( .A(n26519), .B(n26716), .Y(n24479) );
  sky130_fd_sc_hd__nand2_1 U29648 ( .A(n24479), .B(n24785), .Y(n24480) );
  sky130_fd_sc_hd__o22a_1 U29649 ( .A1(n26579), .A2(n26431), .B1(n26564), .B2(
        n26412), .X(n24488) );
  sky130_fd_sc_hd__o22ai_1 U29650 ( .A1(n26423), .A2(n27357), .B1(n27341), 
        .B2(n26424), .Y(n24482) );
  sky130_fd_sc_hd__a21oi_1 U29651 ( .A1(n24483), .A2(n26414), .B1(n24482), .Y(
        n24487) );
  sky130_fd_sc_hd__xor2_1 U29652 ( .A(n26716), .B(n27357), .X(n26620) );
  sky130_fd_sc_hd__o2bb2ai_1 U29653 ( .B1(n26565), .B2(n26425), .A1_N(n26326), 
        .A2_N(n26620), .Y(n24485) );
  sky130_fd_sc_hd__o22ai_1 U29654 ( .A1(n26703), .A2(n26416), .B1(n26702), 
        .B2(n26427), .Y(n24484) );
  sky130_fd_sc_hd__nor2_1 U29655 ( .A(n24485), .B(n24484), .Y(n24486) );
  sky130_fd_sc_hd__nand4_1 U29656 ( .A(n24488), .B(n24487), .C(n24486), .D(
        n26411), .Y(n24489) );
  sky130_fd_sc_hd__a21oi_1 U29657 ( .A1(n24490), .A2(n26409), .B1(n24489), .Y(
        n24491) );
  sky130_fd_sc_hd__nand2_1 U29659 ( .A(n24497), .B(n27192), .Y(n24496) );
  sky130_fd_sc_hd__o21ai_1 U29660 ( .A1(n27192), .A2(n27359), .B1(n24496), .Y(
        j202_soc_core_j22_cpu_rf_N3304) );
  sky130_fd_sc_hd__o22ai_1 U29661 ( .A1(n27359), .A2(n26899), .B1(n26898), 
        .B2(n26523), .Y(j202_soc_core_j22_cpu_rf_N3342) );
  sky130_fd_sc_hd__o22ai_1 U29662 ( .A1(n26378), .A2(n27359), .B1(n26449), 
        .B2(n26523), .Y(j202_soc_core_j22_cpu_rf_N3267) );
  sky130_fd_sc_hd__o22ai_1 U29663 ( .A1(n11141), .A2(n27359), .B1(n27124), 
        .B2(n26523), .Y(j202_soc_core_j22_cpu_rf_N2712) );
  sky130_fd_sc_hd__a22oi_1 U29664 ( .A1(n27184), .A2(n26716), .B1(n11771), 
        .B2(n27339), .Y(n24498) );
  sky130_fd_sc_hd__nand2_1 U29665 ( .A(n27346), .B(n24498), .Y(
        j202_soc_core_j22_cpu_ml_N334) );
  sky130_fd_sc_hd__nand2_1 U29666 ( .A(n23244), .B(n24499), .Y(n24503) );
  sky130_fd_sc_hd__nand2_1 U29667 ( .A(n24500), .B(n26863), .Y(n24501) );
  sky130_fd_sc_hd__a31oi_1 U29668 ( .A1(n24503), .A2(n24502), .A3(n24501), 
        .B1(n26865), .Y(n24504) );
  sky130_fd_sc_hd__a21oi_1 U29669 ( .A1(n24505), .A2(n27187), .B1(n24504), .Y(
        n24506) );
  sky130_fd_sc_hd__nand2_1 U29670 ( .A(n27189), .B(n24506), .Y(
        j202_soc_core_j22_cpu_ml_machj[30]) );
  sky130_fd_sc_hd__a211oi_1 U29671 ( .A1(n24510), .A2(n26872), .B1(n24509), 
        .C1(n24508), .Y(n24513) );
  sky130_fd_sc_hd__nand2_1 U29673 ( .A(n26472), .B(n26802), .Y(n24540) );
  sky130_fd_sc_hd__nand2_1 U29674 ( .A(n26077), .B(n26414), .Y(n24515) );
  sky130_fd_sc_hd__nand2_1 U29675 ( .A(n24518), .B(n26417), .Y(n26649) );
  sky130_fd_sc_hd__nand2_1 U29676 ( .A(n27419), .B(n26717), .Y(n26648) );
  sky130_fd_sc_hd__nand3_1 U29677 ( .A(n26649), .B(n26326), .C(n26648), .Y(
        n24514) );
  sky130_fd_sc_hd__o211ai_1 U29678 ( .A1(n27007), .A2(n26425), .B1(n24515), 
        .C1(n24514), .Y(n24517) );
  sky130_fd_sc_hd__o22ai_1 U29679 ( .A1(n26571), .A2(n26419), .B1(n26703), 
        .B2(n26418), .Y(n24516) );
  sky130_fd_sc_hd__nor2_1 U29680 ( .A(n24517), .B(n24516), .Y(n24527) );
  sky130_fd_sc_hd__o22a_1 U29681 ( .A1(n24518), .A2(n26431), .B1(n26791), .B2(
        n26412), .X(n24526) );
  sky130_fd_sc_hd__o22ai_1 U29682 ( .A1(n18916), .A2(n24519), .B1(n26423), 
        .B2(n27419), .Y(n24520) );
  sky130_fd_sc_hd__a21oi_1 U29683 ( .A1(n26085), .A2(n26717), .B1(n24520), .Y(
        n24521) );
  sky130_fd_sc_hd__o21ai_0 U29684 ( .A1(n26432), .A2(n26648), .B1(n24521), .Y(
        n24524) );
  sky130_fd_sc_hd__nor2_1 U29685 ( .A(n26570), .B(n26424), .Y(n24523) );
  sky130_fd_sc_hd__o22ai_1 U29686 ( .A1(n25403), .A2(n26427), .B1(n26426), 
        .B2(n26416), .Y(n24522) );
  sky130_fd_sc_hd__nor3_1 U29687 ( .A(n24524), .B(n24523), .C(n24522), .Y(
        n24525) );
  sky130_fd_sc_hd__nand4_1 U29688 ( .A(n24527), .B(n24526), .C(n26411), .D(
        n24525), .Y(n24528) );
  sky130_fd_sc_hd__o21bai_1 U29689 ( .A1(n18916), .A2(n24529), .B1_N(n24528), 
        .Y(n24530) );
  sky130_fd_sc_hd__a21oi_1 U29690 ( .A1(n24531), .A2(n26409), .B1(n24530), .Y(
        n24536) );
  sky130_fd_sc_hd__nand2_1 U29691 ( .A(n26717), .B(n26323), .Y(n24532) );
  sky130_fd_sc_hd__o211ai_1 U29692 ( .A1(n26352), .A2(n26717), .B1(n26351), 
        .C1(n24532), .Y(n24533) );
  sky130_fd_sc_hd__nand2_1 U29693 ( .A(n24534), .B(n24533), .Y(n24535) );
  sky130_fd_sc_hd__nand2b_1 U29694 ( .A_N(n24538), .B(n25181), .Y(n24539) );
  sky130_fd_sc_hd__nand2_1 U29695 ( .A(n12435), .B(n27192), .Y(n24541) );
  sky130_fd_sc_hd__o21ai_0 U29696 ( .A1(n27192), .A2(n24546), .B1(n24541), .Y(
        j202_soc_core_j22_cpu_rf_N3292) );
  sky130_fd_sc_hd__o22ai_1 U29697 ( .A1(n24546), .A2(n26899), .B1(n26898), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N3331) );
  sky130_fd_sc_hd__o22ai_1 U29698 ( .A1(n26378), .A2(n24546), .B1(n26449), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N3255) );
  sky130_fd_sc_hd__o22ai_1 U29699 ( .A1(n11141), .A2(n24546), .B1(n27124), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N2700) );
  sky130_fd_sc_hd__nand2_1 U29700 ( .A(n12435), .B(n26516), .Y(n24545) );
  sky130_fd_sc_hd__o22a_1 U29701 ( .A1(n24543), .A2(n26070), .B1(n25714), .B2(
        n24546), .X(n24544) );
  sky130_fd_sc_hd__nand2_1 U29702 ( .A(n24545), .B(n24544), .Y(
        j202_soc_core_j22_cpu_rf_N3367) );
  sky130_fd_sc_hd__o22ai_1 U29703 ( .A1(n27219), .A2(n24546), .B1(n27218), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N2996) );
  sky130_fd_sc_hd__o22ai_1 U29704 ( .A1(n27217), .A2(n24546), .B1(n27216), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N2848) );
  sky130_fd_sc_hd__o22ai_1 U29705 ( .A1(n27228), .A2(n24546), .B1(n27227), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N3181) );
  sky130_fd_sc_hd__o22ai_1 U29706 ( .A1(n27225), .A2(n24546), .B1(n27224), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N2959) );
  sky130_fd_sc_hd__o22ai_1 U29707 ( .A1(n27215), .A2(n24546), .B1(n27214), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N2922) );
  sky130_fd_sc_hd__o22ai_1 U29708 ( .A1(n27223), .A2(n24546), .B1(n27222), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N3033) );
  sky130_fd_sc_hd__o22ai_1 U29709 ( .A1(n27211), .A2(n24546), .B1(n27210), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N3218) );
  sky130_fd_sc_hd__o22ai_1 U29710 ( .A1(n27221), .A2(n24546), .B1(n27220), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N2885) );
  sky130_fd_sc_hd__o22ai_1 U29711 ( .A1(n27226), .A2(n24546), .B1(n23079), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N3144) );
  sky130_fd_sc_hd__o22ai_1 U29712 ( .A1(n27213), .A2(n24546), .B1(n27212), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N2811) );
  sky130_fd_sc_hd__o22ai_1 U29713 ( .A1(n27209), .A2(n24546), .B1(n23039), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N2737) );
  sky130_fd_sc_hd__a22oi_1 U29714 ( .A1(n27184), .A2(n26414), .B1(n26557), 
        .B2(n27339), .Y(n24547) );
  sky130_fd_sc_hd__nand2_1 U29715 ( .A(n27346), .B(n24547), .Y(
        j202_soc_core_j22_cpu_ml_N332) );
  sky130_fd_sc_hd__nand2_1 U29716 ( .A(n27189), .B(n24549), .Y(
        j202_soc_core_j22_cpu_ml_machj[28]) );
  sky130_fd_sc_hd__o21ai_1 U29717 ( .A1(n26981), .A2(n26402), .B1(n24552), .Y(
        j202_soc_core_j22_cpu_ml_maclj[28]) );
  sky130_fd_sc_hd__nand2_1 U29718 ( .A(n12355), .B(n26371), .Y(n24553) );
  sky130_fd_sc_hd__nand2_1 U29719 ( .A(n12355), .B(n27211), .Y(n24554) );
  sky130_fd_sc_hd__o21ai_1 U29720 ( .A1(n27211), .A2(n27461), .B1(n24554), .Y(
        j202_soc_core_j22_cpu_rf_N3210) );
  sky130_fd_sc_hd__nand2_1 U29722 ( .A(n27459), .B(n27223), .Y(n24556) );
  sky130_fd_sc_hd__nand2_1 U29723 ( .A(n27459), .B(n27225), .Y(n24557) );
  sky130_fd_sc_hd__nand2_1 U29724 ( .A(n27459), .B(n26378), .Y(n24558) );
  sky130_fd_sc_hd__nand2_1 U29725 ( .A(n12355), .B(n11141), .Y(n24559) );
  sky130_fd_sc_hd__nand2_1 U29726 ( .A(n27459), .B(n27228), .Y(n24560) );
  sky130_fd_sc_hd__nor3_1 U29728 ( .A(n29063), .B(n29032), .C(n29030), .Y(
        n24566) );
  sky130_fd_sc_hd__nor2_1 U29729 ( .A(n29062), .B(n29031), .Y(n24564) );
  sky130_fd_sc_hd__nand3_1 U29730 ( .A(n24566), .B(n24565), .C(n24564), .Y(
        n27128) );
  sky130_fd_sc_hd__nor2_1 U29731 ( .A(n29064), .B(n27128), .Y(n24567) );
  sky130_fd_sc_hd__nand2_1 U29733 ( .A(n24808), .B(n27603), .Y(n24569) );
  sky130_fd_sc_hd__nand2_1 U29734 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[23]), .Y(n24570) );
  sky130_fd_sc_hd__o21ai_1 U29735 ( .A1(n24571), .A2(n27983), .B1(n24570), .Y(
        n49) );
  sky130_fd_sc_hd__nand2_1 U29736 ( .A(n27593), .B(j202_soc_core_uart_div1[7]), 
        .Y(n24573) );
  sky130_fd_sc_hd__o21ai_1 U29737 ( .A1(n24574), .A2(n27593), .B1(n24573), .Y(
        n111) );
  sky130_fd_sc_hd__o22ai_1 U29738 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(io_in[11]), .B1(
        n28901), .B2(io_in[10]), .Y(n24576) );
  sky130_fd_sc_hd__nor2_1 U29739 ( .A(n24575), .B(n24576), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N323) );
  sky130_fd_sc_hd__o22ai_1 U29740 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[0]), .B1(n28901), .B2(
        io_in[11]), .Y(n24993) );
  sky130_fd_sc_hd__nor2_1 U29741 ( .A(n24575), .B(n24993), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N324) );
  sky130_fd_sc_hd__o22ai_1 U29742 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[1]), .B1(n28901), .B2(
        io_in[12]), .Y(n24992) );
  sky130_fd_sc_hd__nor2_1 U29743 ( .A(n24575), .B(n24992), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N325) );
  sky130_fd_sc_hd__o22ai_1 U29744 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[2]), .B1(n28901), .B2(
        io_in[13]), .Y(n27873) );
  sky130_fd_sc_hd__nor2_1 U29745 ( .A(n24575), .B(n27873), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N326) );
  sky130_fd_sc_hd__nor2_1 U29746 ( .A(n26211), .B(n24576), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N358) );
  sky130_fd_sc_hd__nand2_1 U29747 ( .A(n27039), .B(n28096), .Y(n24580) );
  sky130_fd_sc_hd__nand2_1 U29748 ( .A(n26009), .B(n26161), .Y(n26251) );
  sky130_fd_sc_hd__nand2b_1 U29749 ( .A_N(n26049), .B(
        j202_soc_core_wbqspiflash_00_state[3]), .Y(n28217) );
  sky130_fd_sc_hd__a21oi_1 U29750 ( .A1(n28217), .A2(n25901), .B1(n26255), .Y(
        n24577) );
  sky130_fd_sc_hd__a211oi_1 U29751 ( .A1(n24580), .A2(
        j202_soc_core_wbqspiflash_00_spi_out[0]), .B1(n24579), .C1(n24577), 
        .Y(n24578) );
  sky130_fd_sc_hd__nor2_1 U29752 ( .A(n28590), .B(n24578), .Y(
        j202_soc_core_wbqspiflash_00_N709) );
  sky130_fd_sc_hd__nor2_1 U29753 ( .A(n25921), .B(n26022), .Y(n26175) );
  sky130_fd_sc_hd__nor2_1 U29754 ( .A(n26175), .B(n24579), .Y(n24581) );
  sky130_fd_sc_hd__nand2_1 U29755 ( .A(n24580), .B(
        j202_soc_core_wbqspiflash_00_spi_valid), .Y(n26474) );
  sky130_fd_sc_hd__nand4_1 U29756 ( .A(n27123), .B(n24581), .C(n26248), .D(
        n26474), .Y(j202_soc_core_wbqspiflash_00_N708) );
  sky130_fd_sc_hd__a22oi_1 U29757 ( .A1(n27187), .A2(n24583), .B1(n27273), 
        .B2(n24582), .Y(n24584) );
  sky130_fd_sc_hd__nand2_1 U29758 ( .A(n27189), .B(n24584), .Y(
        j202_soc_core_j22_cpu_ml_machj[24]) );
  sky130_fd_sc_hd__a21oi_1 U29759 ( .A1(n25344), .A2(n10968), .B1(n26976), .Y(
        n24589) );
  sky130_fd_sc_hd__nand3_1 U29760 ( .A(n12356), .B(n24586), .C(n26872), .Y(
        n24588) );
  sky130_fd_sc_hd__o21ai_0 U29761 ( .A1(n26946), .A2(n27208), .B1(n24643), .Y(
        j202_soc_core_j22_cpu_rf_N2646) );
  sky130_fd_sc_hd__mux2i_1 U29762 ( .A0(n27208), .A1(n27234), .S(n27460), .Y(
        j202_soc_core_j22_cpu_rf_N3274) );
  sky130_fd_sc_hd__o22ai_1 U29763 ( .A1(n27234), .A2(n26378), .B1(n26449), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N3237) );
  sky130_fd_sc_hd__nand2_1 U29764 ( .A(n11704), .B(n11157), .Y(n24598) );
  sky130_fd_sc_hd__o22ai_1 U29765 ( .A1(n26791), .A2(n26892), .B1(n26891), 
        .B2(n24595), .Y(n24596) );
  sky130_fd_sc_hd__a21oi_1 U29766 ( .A1(n25759), .A2(n26895), .B1(n24596), .Y(
        n24597) );
  sky130_fd_sc_hd__nand2_1 U29767 ( .A(n24598), .B(n24597), .Y(
        j202_soc_core_j22_cpu_rf_N302) );
  sky130_fd_sc_hd__o22ai_1 U29768 ( .A1(n27234), .A2(n26899), .B1(n26898), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N3314) );
  sky130_fd_sc_hd__o22ai_1 U29769 ( .A1(n27234), .A2(n11141), .B1(n27124), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N2682) );
  sky130_fd_sc_hd__nor2_1 U29770 ( .A(j202_soc_core_intc_core_00_bs_addr[2]), 
        .B(n28886), .Y(n28885) );
  sky130_fd_sc_hd__nand3_1 U29771 ( .A(n24755), .B(n28885), .C(n24756), .Y(
        n24761) );
  sky130_fd_sc_hd__nor2_1 U29772 ( .A(n28882), .B(n24761), .Y(n27752) );
  sky130_fd_sc_hd__nor2_1 U29773 ( .A(n28590), .B(n27752), .Y(n27751) );
  sky130_fd_sc_hd__o22ai_1 U29774 ( .A1(n28613), .A2(n27990), .B1(n24599), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U29775 ( .A1(n28606), .A2(n27990), .B1(n24600), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U29776 ( .A1(n28613), .A2(n25534), .B1(n24601), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__a21oi_1 U29777 ( .A1(n25344), .A2(n12613), .B1(n26976), .Y(
        n24605) );
  sky130_fd_sc_hd__nand3_1 U29778 ( .A(n12357), .B(n24602), .C(n26872), .Y(
        n24603) );
  sky130_fd_sc_hd__o22ai_1 U29779 ( .A1(n28881), .A2(n25534), .B1(n24606), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__nand2b_1 U29780 ( .A_N(n24607), .B(n24749), .Y(n24762) );
  sky130_fd_sc_hd__nor2_1 U29781 ( .A(n28882), .B(n24762), .Y(n27154) );
  sky130_fd_sc_hd__nor2_1 U29782 ( .A(n28590), .B(
        j202_soc_core_qspi_wb_wdat[4]), .Y(n28300) );
  sky130_fd_sc_hd__o22ai_1 U29783 ( .A1(n27154), .A2(n26997), .B1(n28300), 
        .B2(n27152), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__nand2_1 U29784 ( .A(n24634), .B(n26802), .Y(n24632) );
  sky130_fd_sc_hd__nand2_1 U29785 ( .A(n27439), .B(n25128), .Y(n26651) );
  sky130_fd_sc_hd__nand2_1 U29786 ( .A(n24613), .B(n26724), .Y(n26650) );
  sky130_fd_sc_hd__nand3_1 U29787 ( .A(n26651), .B(n26326), .C(n26650), .Y(
        n24609) );
  sky130_fd_sc_hd__nand2_1 U29788 ( .A(n26077), .B(n25137), .Y(n24608) );
  sky130_fd_sc_hd__o211ai_1 U29789 ( .A1(n26581), .A2(n26427), .B1(n24609), 
        .C1(n24608), .Y(n24611) );
  sky130_fd_sc_hd__o22ai_1 U29790 ( .A1(n26567), .A2(n26419), .B1(n25403), 
        .B2(n26418), .Y(n24610) );
  sky130_fd_sc_hd__nor2_1 U29791 ( .A(n24611), .B(n24610), .Y(n24622) );
  sky130_fd_sc_hd__o22a_1 U29792 ( .A1(n27439), .A2(n26431), .B1(n24612), .B2(
        n26412), .X(n24621) );
  sky130_fd_sc_hd__o22ai_1 U29793 ( .A1(n18916), .A2(n24614), .B1(n26423), 
        .B2(n24613), .Y(n24615) );
  sky130_fd_sc_hd__a21oi_1 U29794 ( .A1(n26085), .A2(n26724), .B1(n24615), .Y(
        n24616) );
  sky130_fd_sc_hd__o21ai_0 U29795 ( .A1(n26432), .A2(n26650), .B1(n24616), .Y(
        n24619) );
  sky130_fd_sc_hd__nor2_1 U29796 ( .A(n26571), .B(n26424), .Y(n24618) );
  sky130_fd_sc_hd__o22ai_1 U29797 ( .A1(n25788), .A2(n26416), .B1(n25743), 
        .B2(n26425), .Y(n24617) );
  sky130_fd_sc_hd__nor3_1 U29798 ( .A(n24619), .B(n24618), .C(n24617), .Y(
        n24620) );
  sky130_fd_sc_hd__nand4_1 U29799 ( .A(n24622), .B(n24621), .C(n26411), .D(
        n24620), .Y(n24623) );
  sky130_fd_sc_hd__o21bai_1 U29800 ( .A1(n18916), .A2(n24624), .B1_N(n24623), 
        .Y(n24625) );
  sky130_fd_sc_hd__a21oi_1 U29801 ( .A1(n24626), .A2(n26409), .B1(n24625), .Y(
        n24627) );
  sky130_fd_sc_hd__o21a_1 U29802 ( .A1(n26102), .A2(n24628), .B1(n24627), .X(
        n24631) );
  sky130_fd_sc_hd__nand2_1 U29803 ( .A(n26724), .B(n26323), .Y(n24630) );
  sky130_fd_sc_hd__o22ai_1 U29804 ( .A1(n27209), .A2(n11103), .B1(n23039), 
        .B2(n25707), .Y(j202_soc_core_j22_cpu_rf_N2734) );
  sky130_fd_sc_hd__o22ai_1 U29805 ( .A1(n27215), .A2(n11103), .B1(n27214), 
        .B2(n12468), .Y(j202_soc_core_j22_cpu_rf_N2919) );
  sky130_fd_sc_hd__o22ai_1 U29806 ( .A1(n27225), .A2(n11103), .B1(n27224), 
        .B2(n12468), .Y(j202_soc_core_j22_cpu_rf_N2956) );
  sky130_fd_sc_hd__o22ai_1 U29807 ( .A1(n26378), .A2(n11103), .B1(n26449), 
        .B2(n25707), .Y(j202_soc_core_j22_cpu_rf_N3252) );
  sky130_fd_sc_hd__o22ai_1 U29808 ( .A1(n27219), .A2(n11103), .B1(n27218), 
        .B2(n25707), .Y(j202_soc_core_j22_cpu_rf_N2993) );
  sky130_fd_sc_hd__o22ai_1 U29809 ( .A1(n27228), .A2(n11103), .B1(n27227), 
        .B2(n12468), .Y(j202_soc_core_j22_cpu_rf_N3178) );
  sky130_fd_sc_hd__o22ai_1 U29810 ( .A1(n11141), .A2(n11103), .B1(n27124), 
        .B2(n12468), .Y(j202_soc_core_j22_cpu_rf_N2697) );
  sky130_fd_sc_hd__o22ai_1 U29811 ( .A1(n27466), .A2(n11103), .B1(n27465), 
        .B2(n25707), .Y(j202_soc_core_j22_cpu_rf_N2771) );
  sky130_fd_sc_hd__o22ai_1 U29812 ( .A1(n27211), .A2(n11103), .B1(n27210), 
        .B2(n12468), .Y(j202_soc_core_j22_cpu_rf_N3215) );
  sky130_fd_sc_hd__o22ai_1 U29813 ( .A1(n27223), .A2(n11103), .B1(n27222), 
        .B2(n12468), .Y(j202_soc_core_j22_cpu_rf_N3030) );
  sky130_fd_sc_hd__o22ai_1 U29814 ( .A1(n27217), .A2(n11103), .B1(n27216), 
        .B2(n25707), .Y(j202_soc_core_j22_cpu_rf_N2845) );
  sky130_fd_sc_hd__o22ai_1 U29815 ( .A1(n27575), .A2(n11103), .B1(n27574), 
        .B2(n25707), .Y(j202_soc_core_j22_cpu_rf_N3104) );
  sky130_fd_sc_hd__o22ai_1 U29816 ( .A1(n27226), .A2(n11103), .B1(n23079), 
        .B2(n12468), .Y(j202_soc_core_j22_cpu_rf_N3141) );
  sky130_fd_sc_hd__a22oi_1 U29817 ( .A1(n27187), .A2(n18300), .B1(n24634), 
        .B2(n27047), .Y(n24635) );
  sky130_fd_sc_hd__nand2_1 U29818 ( .A(n27189), .B(n24635), .Y(
        j202_soc_core_j22_cpu_ml_machj[17]) );
  sky130_fd_sc_hd__mux2i_1 U29819 ( .A0(n27576), .A1(n26713), .S(n27006), .Y(
        j202_soc_core_j22_cpu_ml_N306) );
  sky130_fd_sc_hd__o22ai_1 U29820 ( .A1(n27576), .A2(n27209), .B1(n23039), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N2718) );
  sky130_fd_sc_hd__o22ai_1 U29821 ( .A1(n27576), .A2(n27215), .B1(n27214), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N2903) );
  sky130_fd_sc_hd__o22ai_1 U29822 ( .A1(n27576), .A2(n27225), .B1(n27224), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N2940) );
  sky130_fd_sc_hd__o22ai_1 U29823 ( .A1(n27576), .A2(n11141), .B1(n27124), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N2681) );
  sky130_fd_sc_hd__o22ai_1 U29824 ( .A1(n27576), .A2(n27226), .B1(n23079), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N3125) );
  sky130_fd_sc_hd__o22ai_1 U29825 ( .A1(n27576), .A2(n27219), .B1(n27218), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N2977) );
  sky130_fd_sc_hd__o22ai_1 U29826 ( .A1(n27576), .A2(n27228), .B1(n27227), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N3162) );
  sky130_fd_sc_hd__o22ai_1 U29827 ( .A1(n11793), .A2(n27297), .B1(n27298), 
        .B2(n24704), .Y(n24641) );
  sky130_fd_sc_hd__nor2_1 U29828 ( .A(n13271), .B(n11130), .Y(n24640) );
  sky130_fd_sc_hd__o21ai_1 U29829 ( .A1(n24641), .A2(n24640), .B1(n27980), .Y(
        n24642) );
  sky130_fd_sc_hd__nand2_1 U29830 ( .A(n24642), .B(n27300), .Y(n10500) );
  sky130_fd_sc_hd__o22ai_1 U29831 ( .A1(n12366), .A2(n24643), .B1(n26946), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N2645) );
  sky130_fd_sc_hd__o22ai_1 U29832 ( .A1(n27576), .A2(n27333), .B1(n23178), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N3051) );
  sky130_fd_sc_hd__o22ai_1 U29833 ( .A1(n27576), .A2(n27466), .B1(n27465), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N2755) );
  sky130_fd_sc_hd__o22ai_1 U29834 ( .A1(n27576), .A2(n27221), .B1(n27220), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N2866) );
  sky130_fd_sc_hd__o22ai_1 U29835 ( .A1(n27576), .A2(n27211), .B1(n27210), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N3199) );
  sky130_fd_sc_hd__o22ai_1 U29836 ( .A1(n27576), .A2(n27213), .B1(n27212), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N2792) );
  sky130_fd_sc_hd__o22ai_1 U29837 ( .A1(n27576), .A2(n27223), .B1(n27222), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N3014) );
  sky130_fd_sc_hd__o22ai_1 U29838 ( .A1(n27576), .A2(n27217), .B1(n27216), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N2829) );
  sky130_fd_sc_hd__o22ai_1 U29839 ( .A1(n27576), .A2(n26378), .B1(n26449), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N3236) );
  sky130_fd_sc_hd__mux2i_1 U29840 ( .A0(n24644), .A1(n27576), .S(n27460), .Y(
        j202_soc_core_j22_cpu_rf_N3273) );
  sky130_fd_sc_hd__nand2_1 U29841 ( .A(n12120), .B(n11157), .Y(n24649) );
  sky130_fd_sc_hd__o22ai_1 U29842 ( .A1(n26792), .A2(n26892), .B1(n26891), 
        .B2(n24646), .Y(n24647) );
  sky130_fd_sc_hd__a21oi_1 U29843 ( .A1(n24651), .A2(n26895), .B1(n24647), .Y(
        n24648) );
  sky130_fd_sc_hd__nand2_1 U29844 ( .A(n24649), .B(n24648), .Y(
        j202_soc_core_j22_cpu_rf_N301) );
  sky130_fd_sc_hd__o22ai_1 U29845 ( .A1(n27576), .A2(n26899), .B1(n26898), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N3313) );
  sky130_fd_sc_hd__a22oi_1 U29846 ( .A1(n24651), .A2(n26948), .B1(n12120), 
        .B2(n24650), .Y(n24652) );
  sky130_fd_sc_hd__o21ai_1 U29847 ( .A1(n26951), .A2(n24644), .B1(n24652), .Y(
        j202_soc_core_j22_cpu_rf_N3348) );
  sky130_fd_sc_hd__nand2_1 U29848 ( .A(n11766), .B(n27343), .Y(n24653) );
  sky130_fd_sc_hd__o21ai_1 U29849 ( .A1(n26336), .A2(n27343), .B1(n24653), .Y(
        j202_soc_core_j22_cpu_ml_N314) );
  sky130_fd_sc_hd__a21oi_1 U29850 ( .A1(n18147), .A2(n27187), .B1(n25829), .Y(
        n24655) );
  sky130_fd_sc_hd__o21ai_1 U29851 ( .A1(n27274), .A2(n24691), .B1(n24655), .Y(
        j202_soc_core_j22_cpu_ml_machj[11]) );
  sky130_fd_sc_hd__inv_1 U29852 ( .A(n29516), .Y(n24657) );
  sky130_fd_sc_hd__nand2_1 U29853 ( .A(n24657), .B(n27980), .Y(n25816) );
  sky130_fd_sc_hd__a21oi_1 U29854 ( .A1(n27377), .A2(n25415), .B1(n26085), .Y(
        n24661) );
  sky130_fd_sc_hd__xnor2_1 U29855 ( .A(n26720), .B(n27377), .Y(n26675) );
  sky130_fd_sc_hd__o22ai_1 U29856 ( .A1(n26415), .A2(n26675), .B1(n18916), 
        .B2(n24662), .Y(n24664) );
  sky130_fd_sc_hd__o22ai_1 U29857 ( .A1(n26708), .A2(n26418), .B1(n25788), 
        .B2(n26419), .Y(n24663) );
  sky130_fd_sc_hd__a211oi_1 U29858 ( .A1(n24665), .A2(n27377), .B1(n24664), 
        .C1(n24663), .Y(n24674) );
  sky130_fd_sc_hd__o22ai_1 U29859 ( .A1(n26713), .A2(n26416), .B1(n26426), 
        .B2(n26424), .Y(n24666) );
  sky130_fd_sc_hd__a21oi_1 U29860 ( .A1(n26341), .A2(n25130), .B1(n24666), .Y(
        n24673) );
  sky130_fd_sc_hd__a22oi_1 U29861 ( .A1(n25308), .A2(n24667), .B1(n26077), 
        .B2(n26719), .Y(n24669) );
  sky130_fd_sc_hd__nand2_1 U29862 ( .A(n26338), .B(n27429), .Y(n24668) );
  sky130_fd_sc_hd__o211ai_1 U29863 ( .A1(n26325), .A2(n26427), .B1(n24669), 
        .C1(n24668), .Y(n24670) );
  sky130_fd_sc_hd__a21oi_1 U29864 ( .A1(n26342), .A2(n24671), .B1(n24670), .Y(
        n24672) );
  sky130_fd_sc_hd__nand4_1 U29865 ( .A(n24674), .B(n24673), .C(n24672), .D(
        n26344), .Y(n24675) );
  sky130_fd_sc_hd__a21oi_1 U29866 ( .A1(n24676), .A2(n26409), .B1(n24675), .Y(
        n24679) );
  sky130_fd_sc_hd__o21ai_1 U29867 ( .A1(n26352), .A2(n26720), .B1(n26351), .Y(
        n24677) );
  sky130_fd_sc_hd__nand2_1 U29868 ( .A(n12374), .B(n24677), .Y(n24678) );
  sky130_fd_sc_hd__nand2_1 U29870 ( .A(n24686), .B(n27192), .Y(n24685) );
  sky130_fd_sc_hd__nand2_1 U29871 ( .A(n11766), .B(n27460), .Y(n24684) );
  sky130_fd_sc_hd__nand2_1 U29872 ( .A(n24685), .B(n24684), .Y(
        j202_soc_core_j22_cpu_rf_N3282) );
  sky130_fd_sc_hd__o22ai_1 U29873 ( .A1(n27464), .A2(n26899), .B1(n26898), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N3322) );
  sky130_fd_sc_hd__o22ai_1 U29874 ( .A1(n26378), .A2(n27464), .B1(n26449), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N3245) );
  sky130_fd_sc_hd__o22ai_1 U29875 ( .A1(n11141), .A2(n27464), .B1(n27124), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N2690) );
  sky130_fd_sc_hd__nand2_1 U29876 ( .A(n26516), .B(n26802), .Y(n25335) );
  sky130_fd_sc_hd__a22oi_1 U29877 ( .A1(n26948), .A2(n24687), .B1(n11766), 
        .B2(n24650), .Y(n24688) );
  sky130_fd_sc_hd__o21ai_1 U29879 ( .A1(n25547), .A2(n27274), .B1(n27273), .Y(
        j202_soc_core_j22_cpu_ml_machj[9]) );
  sky130_fd_sc_hd__nor2_1 U29880 ( .A(n28776), .B(n28753), .Y(n24696) );
  sky130_fd_sc_hd__a21oi_1 U29881 ( .A1(n28776), .A2(n28753), .B1(n24696), .Y(
        n23) );
  sky130_fd_sc_hd__nand2_1 U29882 ( .A(n28281), .B(j202_soc_core_uart_WRTXD1), 
        .Y(n24697) );
  sky130_fd_sc_hd__a21oi_1 U29883 ( .A1(n24694), .A2(n24697), .B1(n24693), .Y(
        n87) );
  sky130_fd_sc_hd__a21o_1 U29884 ( .A1(j202_soc_core_uart_TOP_tx_fifo_wp[1]), 
        .A2(n24695), .B1(n29352), .X(n86) );
  sky130_fd_sc_hd__xor2_1 U29885 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[1]), 
        .B(n24696), .X(n22) );
  sky130_fd_sc_hd__a211o_1 U29886 ( .A1(n24698), .A2(n27991), .B1(n24697), 
        .C1(n27993), .X(n24699) );
  sky130_fd_sc_hd__nor2_1 U29887 ( .A(n28590), .B(n24699), .Y(
        j202_soc_core_uart_TOP_tx_fifo_N42) );
  sky130_fd_sc_hd__nand3_1 U29888 ( .A(n24699), .B(n28776), .C(n29593), .Y(
        j202_soc_core_uart_TOP_tx_fifo_N41) );
  sky130_fd_sc_hd__nand2_1 U29889 ( .A(n24700), .B(n13318), .Y(n25744) );
  sky130_fd_sc_hd__nor2_1 U29890 ( .A(n26946), .B(n29565), .Y(
        j202_soc_core_j22_cpu_rf_N2643) );
  sky130_fd_sc_hd__mux2i_1 U29891 ( .A0(n29565), .A1(n27335), .S(n27460), .Y(
        j202_soc_core_j22_cpu_rf_N3271) );
  sky130_fd_sc_hd__o22ai_1 U29892 ( .A1(n27335), .A2(n26378), .B1(n26449), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N3234) );
  sky130_fd_sc_hd__o22ai_1 U29893 ( .A1(n27335), .A2(n27575), .B1(n27574), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N3086) );
  sky130_fd_sc_hd__o22ai_1 U29894 ( .A1(n27335), .A2(n27219), .B1(n27218), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N2975) );
  sky130_fd_sc_hd__o22ai_1 U29895 ( .A1(n27335), .A2(n27217), .B1(n27216), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N2827) );
  sky130_fd_sc_hd__o22ai_1 U29896 ( .A1(n27335), .A2(n27228), .B1(n27227), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N3160) );
  sky130_fd_sc_hd__o22ai_1 U29897 ( .A1(n27335), .A2(n27225), .B1(n27224), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N2938) );
  sky130_fd_sc_hd__o22ai_1 U29898 ( .A1(n27335), .A2(n27466), .B1(n27465), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N2753) );
  sky130_fd_sc_hd__o22ai_1 U29899 ( .A1(n27335), .A2(n27215), .B1(n27214), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N2901) );
  sky130_fd_sc_hd__o22ai_1 U29900 ( .A1(n27335), .A2(n27223), .B1(n27222), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N3012) );
  sky130_fd_sc_hd__o22ai_1 U29901 ( .A1(n27335), .A2(n27211), .B1(n27210), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N3197) );
  sky130_fd_sc_hd__o22ai_1 U29902 ( .A1(n27335), .A2(n27221), .B1(n27220), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N2864) );
  sky130_fd_sc_hd__o22ai_1 U29903 ( .A1(n27335), .A2(n27226), .B1(n23079), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N3123) );
  sky130_fd_sc_hd__o22ai_1 U29904 ( .A1(n27335), .A2(n27213), .B1(n27212), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N2790) );
  sky130_fd_sc_hd__o22ai_1 U29905 ( .A1(n27335), .A2(n27209), .B1(n23039), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N2716) );
  sky130_fd_sc_hd__o22ai_1 U29906 ( .A1(n27335), .A2(n11141), .B1(n27124), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N2679) );
  sky130_fd_sc_hd__nor2_1 U29907 ( .A(n24703), .B(n24702), .Y(n24709) );
  sky130_fd_sc_hd__nand2_1 U29908 ( .A(n27232), .B(n29036), .Y(n24706) );
  sky130_fd_sc_hd__o22ai_1 U29911 ( .A1(n27335), .A2(n26899), .B1(n26898), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N3309) );
  sky130_fd_sc_hd__nand2_1 U29912 ( .A(n25744), .B(n26067), .Y(n24714) );
  sky130_fd_sc_hd__nand2_1 U29913 ( .A(n27442), .B(n24650), .Y(n24710) );
  sky130_fd_sc_hd__o21ai_1 U29914 ( .A1(j202_soc_core_j22_cpu_pc[1]), .A2(
        n26070), .B1(n24710), .Y(n24711) );
  sky130_fd_sc_hd__a21oi_1 U29915 ( .A1(n26516), .A2(n12591), .B1(n24711), .Y(
        n24713) );
  sky130_fd_sc_hd__nand2_1 U29916 ( .A(n24714), .B(n24713), .Y(
        j202_soc_core_j22_cpu_rf_N3346) );
  sky130_fd_sc_hd__inv_2 U29917 ( .A(n12389), .Y(n25640) );
  sky130_fd_sc_hd__o22ai_1 U29918 ( .A1(n25798), .A2(n26419), .B1(n26336), 
        .B2(n26418), .Y(n24719) );
  sky130_fd_sc_hd__nand2_1 U29919 ( .A(n25121), .B(n25788), .Y(n26674) );
  sky130_fd_sc_hd__nand2_1 U29920 ( .A(n27389), .B(n26721), .Y(n26673) );
  sky130_fd_sc_hd__nand3_1 U29921 ( .A(n26674), .B(n26326), .C(n26673), .Y(
        n24715) );
  sky130_fd_sc_hd__o21ai_0 U29922 ( .A1(n18916), .A2(n24717), .B1(n24716), .Y(
        n24718) );
  sky130_fd_sc_hd__nor2_1 U29923 ( .A(n24719), .B(n24718), .Y(n24727) );
  sky130_fd_sc_hd__o22ai_1 U29924 ( .A1(n25743), .A2(n26416), .B1(n25821), 
        .B2(n26427), .Y(n24720) );
  sky130_fd_sc_hd__a21oi_1 U29925 ( .A1(n26338), .A2(n27443), .B1(n24720), .Y(
        n24725) );
  sky130_fd_sc_hd__o22a_1 U29926 ( .A1(n26423), .A2(n27389), .B1(n26432), .B2(
        n26673), .X(n24721) );
  sky130_fd_sc_hd__o21ai_0 U29927 ( .A1(n26325), .A2(n26424), .B1(n24721), .Y(
        n24722) );
  sky130_fd_sc_hd__a21oi_1 U29928 ( .A1(n26341), .A2(n25137), .B1(n24722), .Y(
        n24724) );
  sky130_fd_sc_hd__nand2_1 U29929 ( .A(n26342), .B(n25122), .Y(n24723) );
  sky130_fd_sc_hd__and4_1 U29930 ( .A(n24725), .B(n24724), .C(n26344), .D(
        n24723), .X(n24726) );
  sky130_fd_sc_hd__o211ai_1 U29931 ( .A1(n25121), .A2(n26349), .B1(n24727), 
        .C1(n24726), .Y(n24728) );
  sky130_fd_sc_hd__a21oi_1 U29932 ( .A1(n24729), .A2(n26409), .B1(n24728), .Y(
        n24731) );
  sky130_fd_sc_hd__o21ai_1 U29933 ( .A1(n26352), .A2(n26721), .B1(n26351), .Y(
        n24730) );
  sky130_fd_sc_hd__o22ai_1 U29934 ( .A1(n27575), .A2(n25640), .B1(n27574), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N3095) );
  sky130_fd_sc_hd__o22ai_1 U29935 ( .A1(n27219), .A2(n25640), .B1(n27218), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N2984) );
  sky130_fd_sc_hd__o22ai_1 U29936 ( .A1(n27217), .A2(n25640), .B1(n27216), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N2836) );
  sky130_fd_sc_hd__o22ai_1 U29937 ( .A1(n27228), .A2(n25640), .B1(n27227), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N3169) );
  sky130_fd_sc_hd__o22ai_1 U29938 ( .A1(n27225), .A2(n25640), .B1(n27224), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N2947) );
  sky130_fd_sc_hd__o22ai_1 U29939 ( .A1(n27466), .A2(n25640), .B1(n27465), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N2762) );
  sky130_fd_sc_hd__o22ai_1 U29940 ( .A1(n27215), .A2(n25640), .B1(n27214), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N2910) );
  sky130_fd_sc_hd__o22ai_1 U29941 ( .A1(n27223), .A2(n25640), .B1(n27222), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N3021) );
  sky130_fd_sc_hd__o22ai_1 U29942 ( .A1(n27211), .A2(n25640), .B1(n27210), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N3206) );
  sky130_fd_sc_hd__o22ai_1 U29943 ( .A1(n27221), .A2(n25640), .B1(n27220), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N2873) );
  sky130_fd_sc_hd__o22ai_1 U29944 ( .A1(n27226), .A2(n25640), .B1(n23079), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N3132) );
  sky130_fd_sc_hd__o22ai_1 U29945 ( .A1(n27213), .A2(n25640), .B1(n27212), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N2799) );
  sky130_fd_sc_hd__o22ai_1 U29946 ( .A1(n26378), .A2(n25640), .B1(n26449), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N3243) );
  sky130_fd_sc_hd__o22ai_1 U29947 ( .A1(n27209), .A2(n25640), .B1(n23039), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N2725) );
  sky130_fd_sc_hd__o22ai_1 U29948 ( .A1(n11141), .A2(n25640), .B1(n27124), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N2688) );
  sky130_fd_sc_hd__nand2_1 U29949 ( .A(n24733), .B(n27192), .Y(n24734) );
  sky130_fd_sc_hd__o22ai_1 U29951 ( .A1(n25640), .A2(n26899), .B1(n26898), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N3319) );
  sky130_fd_sc_hd__mux2i_1 U29952 ( .A0(n27467), .A1(n25798), .S(n27006), .Y(
        j202_soc_core_j22_cpu_ml_N310) );
  sky130_fd_sc_hd__o21ai_0 U29953 ( .A1(n26318), .A2(n23223), .B1(n12177), .Y(
        n24736) );
  sky130_fd_sc_hd__mux2i_1 U29954 ( .A0(n11120), .A1(n27467), .S(n27460), .Y(
        j202_soc_core_j22_cpu_rf_N3278) );
  sky130_fd_sc_hd__o22ai_1 U29955 ( .A1(n27467), .A2(n26899), .B1(n26898), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N3317) );
  sky130_fd_sc_hd__o22ai_1 U29956 ( .A1(n27467), .A2(n26378), .B1(n26449), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N3241) );
  sky130_fd_sc_hd__nor2_1 U29957 ( .A(n26946), .B(n11120), .Y(
        j202_soc_core_j22_cpu_rf_N2649) );
  sky130_fd_sc_hd__a22oi_1 U29958 ( .A1(n24738), .A2(n26948), .B1(n12455), 
        .B2(n24650), .Y(n24739) );
  sky130_fd_sc_hd__o21ai_1 U29959 ( .A1(n26951), .A2(n11120), .B1(n24739), .Y(
        j202_soc_core_j22_cpu_rf_N3352) );
  sky130_fd_sc_hd__o22ai_1 U29960 ( .A1(n27467), .A2(n27575), .B1(n27574), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N3093) );
  sky130_fd_sc_hd__o22ai_1 U29962 ( .A1(n27467), .A2(n27333), .B1(n23178), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N3056) );
  sky130_fd_sc_hd__o22ai_1 U29963 ( .A1(n27467), .A2(n27219), .B1(n27218), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N2982) );
  sky130_fd_sc_hd__o22ai_1 U29964 ( .A1(n27467), .A2(n27217), .B1(n27216), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N2834) );
  sky130_fd_sc_hd__o22ai_1 U29965 ( .A1(n27467), .A2(n27228), .B1(n27227), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N3167) );
  sky130_fd_sc_hd__o22ai_1 U29966 ( .A1(n27467), .A2(n27225), .B1(n27224), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N2945) );
  sky130_fd_sc_hd__o22ai_1 U29967 ( .A1(n27467), .A2(n27215), .B1(n27214), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N2908) );
  sky130_fd_sc_hd__o22ai_1 U29968 ( .A1(n27467), .A2(n27223), .B1(n27222), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N3019) );
  sky130_fd_sc_hd__o22ai_1 U29969 ( .A1(n27467), .A2(n27211), .B1(n27210), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N3204) );
  sky130_fd_sc_hd__o22ai_1 U29970 ( .A1(n27467), .A2(n27221), .B1(n27220), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N2871) );
  sky130_fd_sc_hd__o22ai_1 U29971 ( .A1(n27467), .A2(n27226), .B1(n23079), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N3130) );
  sky130_fd_sc_hd__o22ai_1 U29972 ( .A1(n27467), .A2(n27213), .B1(n27212), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N2797) );
  sky130_fd_sc_hd__o22ai_1 U29973 ( .A1(n27467), .A2(n27209), .B1(n23039), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N2723) );
  sky130_fd_sc_hd__o21ai_0 U29974 ( .A1(n25824), .A2(n17718), .B1(n25822), .Y(
        n24741) );
  sky130_fd_sc_hd__nand3_1 U29975 ( .A(n12357), .B(n24742), .C(n26872), .Y(
        n24743) );
  sky130_fd_sc_hd__nand2_1 U29976 ( .A(n24744), .B(n24743), .Y(
        j202_soc_core_j22_cpu_ml_maclj[7]) );
  sky130_fd_sc_hd__o22ai_1 U29977 ( .A1(n28610), .A2(n25534), .B1(n24745), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U29978 ( .A1(n28614), .A2(n25534), .B1(n24746), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__mux2i_1 U29979 ( .A0(n12161), .A1(n25276), .S(n27460), .Y(
        j202_soc_core_j22_cpu_rf_N3287) );
  sky130_fd_sc_hd__nand2_1 U29980 ( .A(n12644), .B(n27192), .Y(n24747) );
  sky130_fd_sc_hd__nand2_1 U29982 ( .A(n29594), .B(
        j202_soc_core_intc_core_00_bs_addr[6]), .Y(n24750) );
  sky130_fd_sc_hd__nor2_1 U29983 ( .A(j202_soc_core_intc_core_00_bs_addr[5]), 
        .B(j202_soc_core_intc_core_00_bs_addr[4]), .Y(n28894) );
  sky130_fd_sc_hd__and3_1 U29984 ( .A(n27066), .B(n28894), .C(n24970), .X(
        n24748) );
  sky130_fd_sc_hd__nand3_1 U29985 ( .A(n24749), .B(n24972), .C(n24748), .Y(
        n25094) );
  sky130_fd_sc_hd__nand3_1 U29986 ( .A(n29594), .B(n28884), .C(n24751), .Y(
        n24752) );
  sky130_fd_sc_hd__a222oi_1 U29987 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[18]), .B1(n27851), .B2(
        j202_soc_core_intc_core_00_rg_ipr[18]), .C1(n27862), .C2(
        j202_soc_core_intc_core_00_rg_ipr[50]), .Y(n24758) );
  sky130_fd_sc_hd__nand3_1 U29988 ( .A(n24755), .B(
        j202_soc_core_intc_core_00_bs_addr[8]), .C(n28885), .Y(n24977) );
  sky130_fd_sc_hd__nand3_1 U29989 ( .A(n24760), .B(
        j202_soc_core_intc_core_00_bs_addr[3]), .C(n24756), .Y(n24979) );
  sky130_fd_sc_hd__a22oi_1 U29990 ( .A1(n27856), .A2(
        j202_soc_core_intc_core_00_rg_itgt[84]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[114]), .Y(n24757) );
  sky130_fd_sc_hd__nand2_1 U29991 ( .A(n24758), .B(n24757), .Y(n24759) );
  sky130_fd_sc_hd__a21oi_1 U29992 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[18]), .B1(n24759), .Y(n24765) );
  sky130_fd_sc_hd__nand3_1 U29993 ( .A(n24760), .B(
        j202_soc_core_intc_core_00_bs_addr[8]), .C(
        j202_soc_core_intc_core_00_bs_addr[3]), .Y(n24975) );
  sky130_fd_sc_hd__a22oi_1 U29994 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[92]), .B1(n27869), .B2(
        j202_soc_core_intc_core_00_rg_itgt[76]), .Y(n24764) );
  sky130_fd_sc_hd__a22oi_1 U29995 ( .A1(j202_soc_core_intc_core_00_rg_ipr[82]), 
        .A2(n27852), .B1(n27850), .B2(j202_soc_core_intc_core_00_rg_itgt[68]), 
        .Y(n24763) );
  sky130_fd_sc_hd__nand2_1 U29996 ( .A(n27864), .B(
        j202_soc_core_intc_core_00_bs_addr[7]), .Y(n27865) );
  sky130_fd_sc_hd__nand4_1 U29997 ( .A(n24765), .B(n24764), .C(n24763), .D(
        n27865), .Y(j202_soc_core_ahb2apb_01_N146) );
  sky130_fd_sc_hd__nor2_1 U29998 ( .A(n11713), .B(n25247), .Y(n24767) );
  sky130_fd_sc_hd__nand2_1 U29999 ( .A(n24766), .B(n26409), .Y(n24768) );
  sky130_fd_sc_hd__nand2_1 U30000 ( .A(n24768), .B(n11713), .Y(n24769) );
  sky130_fd_sc_hd__o22ai_1 U30001 ( .A1(n26329), .A2(n24770), .B1(n24769), 
        .B2(n25254), .Y(n24798) );
  sky130_fd_sc_hd__a21oi_1 U30002 ( .A1(n27435), .A2(n24773), .B1(n24772), .Y(
        n24780) );
  sky130_fd_sc_hd__xnor2_1 U30003 ( .A(n26728), .B(n27432), .Y(n26659) );
  sky130_fd_sc_hd__o22ai_1 U30004 ( .A1(n24775), .A2(n27432), .B1(n27908), 
        .B2(n26659), .Y(n24776) );
  sky130_fd_sc_hd__a21oi_1 U30005 ( .A1(n27432), .A2(n24777), .B1(n24776), .Y(
        n24779) );
  sky130_fd_sc_hd__a21oi_1 U30006 ( .A1(n24780), .A2(n24779), .B1(n24778), .Y(
        n24797) );
  sky130_fd_sc_hd__o211ai_1 U30007 ( .A1(n26572), .A2(n24784), .B1(n24783), 
        .C1(n24782), .Y(n24786) );
  sky130_fd_sc_hd__nand3_1 U30008 ( .A(n24786), .B(n24785), .C(n26728), .Y(
        n24796) );
  sky130_fd_sc_hd__o22ai_1 U30009 ( .A1(n26325), .A2(n26416), .B1(n25229), 
        .B2(n26425), .Y(n24790) );
  sky130_fd_sc_hd__o22ai_1 U30010 ( .A1(n25128), .A2(n26427), .B1(n26417), 
        .B2(n26418), .Y(n24789) );
  sky130_fd_sc_hd__o21ai_1 U30011 ( .A1(n26581), .A2(n26419), .B1(n24787), .Y(
        n24788) );
  sky130_fd_sc_hd__nor3_1 U30012 ( .A(n24790), .B(n24789), .C(n24788), .Y(
        n24795) );
  sky130_fd_sc_hd__nand2_1 U30013 ( .A(n26728), .B(n26323), .Y(n24791) );
  sky130_fd_sc_hd__o211ai_1 U30014 ( .A1(n24792), .A2(n26728), .B1(n25159), 
        .C1(n24791), .Y(n24793) );
  sky130_fd_sc_hd__o22ai_1 U30015 ( .A1(n26378), .A2(n27434), .B1(n26449), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N3253) );
  sky130_fd_sc_hd__o22ai_1 U30016 ( .A1(n27434), .A2(n26899), .B1(n26898), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N3329) );
  sky130_fd_sc_hd__a22oi_1 U30017 ( .A1(n24799), .A2(n26948), .B1(n25259), 
        .B2(n24650), .Y(n24800) );
  sky130_fd_sc_hd__o21ai_1 U30018 ( .A1(n26951), .A2(n12433), .B1(n24800), .Y(
        j202_soc_core_j22_cpu_rf_N3365) );
  sky130_fd_sc_hd__nor2_1 U30019 ( .A(n26946), .B(n12433), .Y(
        j202_soc_core_j22_cpu_rf_N2662) );
  sky130_fd_sc_hd__a22oi_1 U30020 ( .A1(n27184), .A2(n26728), .B1(n25259), 
        .B2(n27339), .Y(n24801) );
  sky130_fd_sc_hd__nand2_1 U30021 ( .A(n27346), .B(n24801), .Y(
        j202_soc_core_j22_cpu_ml_N321) );
  sky130_fd_sc_hd__o22ai_1 U30022 ( .A1(n11141), .A2(n27434), .B1(n27124), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N2698) );
  sky130_fd_sc_hd__o22ai_1 U30023 ( .A1(n27575), .A2(n27434), .B1(n27574), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N3105) );
  sky130_fd_sc_hd__o22ai_1 U30024 ( .A1(n27219), .A2(n27434), .B1(n27218), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N2994) );
  sky130_fd_sc_hd__o22ai_1 U30025 ( .A1(n27217), .A2(n27434), .B1(n27216), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N2846) );
  sky130_fd_sc_hd__o22ai_1 U30026 ( .A1(n27228), .A2(n27434), .B1(n27227), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N3179) );
  sky130_fd_sc_hd__o22ai_1 U30027 ( .A1(n27225), .A2(n27434), .B1(n27224), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N2957) );
  sky130_fd_sc_hd__o22ai_1 U30028 ( .A1(n27466), .A2(n27434), .B1(n27465), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N2772) );
  sky130_fd_sc_hd__o22ai_1 U30029 ( .A1(n27215), .A2(n27434), .B1(n27214), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N2920) );
  sky130_fd_sc_hd__o22ai_1 U30030 ( .A1(n27223), .A2(n27434), .B1(n27222), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N3031) );
  sky130_fd_sc_hd__o22ai_1 U30031 ( .A1(n27211), .A2(n27434), .B1(n27210), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N3216) );
  sky130_fd_sc_hd__o22ai_1 U30032 ( .A1(n27221), .A2(n27434), .B1(n27220), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N2883) );
  sky130_fd_sc_hd__o22ai_1 U30033 ( .A1(n27226), .A2(n27434), .B1(n23079), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N3142) );
  sky130_fd_sc_hd__o22ai_1 U30034 ( .A1(n27213), .A2(n27434), .B1(n27212), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N2809) );
  sky130_fd_sc_hd__o22ai_1 U30035 ( .A1(n27209), .A2(n27434), .B1(n23039), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N2735) );
  sky130_fd_sc_hd__nand2_1 U30036 ( .A(n24802), .B(
        j202_soc_core_bldc_core_00_hall_value[2]), .Y(n24804) );
  sky130_fd_sc_hd__nand2_1 U30037 ( .A(n24804), .B(n24803), .Y(n138) );
  sky130_fd_sc_hd__nor2_1 U30038 ( .A(n24808), .B(n24807), .Y(n27604) );
  sky130_fd_sc_hd__nand2_1 U30039 ( .A(n24809), .B(n27604), .Y(n27728) );
  sky130_fd_sc_hd__mux2_2 U30040 ( .A0(j202_soc_core_bldc_core_00_wdata[2]), 
        .A1(j202_soc_core_bldc_core_00_comm[2]), .S(n27728), .X(n46) );
  sky130_fd_sc_hd__nor2_1 U30041 ( .A(n27635), .B(n11894), .Y(
        j202_soc_core_ahb2apb_00_N26) );
  sky130_fd_sc_hd__nor2_1 U30042 ( .A(n27636), .B(n11894), .Y(
        j202_soc_core_ahb2apb_00_N25) );
  sky130_fd_sc_hd__nor2_1 U30043 ( .A(n27622), .B(n11894), .Y(
        j202_soc_core_ahb2apb_00_N23) );
  sky130_fd_sc_hd__nor2_1 U30044 ( .A(n27634), .B(n11894), .Y(
        j202_soc_core_ahb2apb_00_N27) );
  sky130_fd_sc_hd__nor2_1 U30045 ( .A(n27639), .B(n11894), .Y(
        j202_soc_core_ahb2apb_00_N28) );
  sky130_fd_sc_hd__nor2_1 U30046 ( .A(n27638), .B(n11894), .Y(
        j202_soc_core_ahb2apb_00_N29) );
  sky130_fd_sc_hd__nor2_1 U30047 ( .A(n29559), .B(n11894), .Y(
        j202_soc_core_ahb2apb_00_N24) );
  sky130_fd_sc_hd__nor2_1 U30048 ( .A(n27637), .B(n11894), .Y(
        j202_soc_core_ahb2apb_00_N30) );
  sky130_fd_sc_hd__nand2_1 U30049 ( .A(n24811), .B(n24810), .Y(n24813) );
  sky130_fd_sc_hd__nand3_1 U30050 ( .A(n24814), .B(n24812), .C(
        j202_soc_core_ahb2apb_00_state[0]), .Y(n24949) );
  sky130_fd_sc_hd__a21oi_1 U30051 ( .A1(n24813), .A2(n24949), .B1(n28590), .Y(
        j202_soc_core_ahb2apb_00_N90) );
  sky130_fd_sc_hd__nand2_1 U30052 ( .A(n24815), .B(n24814), .Y(n24816) );
  sky130_fd_sc_hd__nor2_1 U30053 ( .A(n24816), .B(n11894), .Y(
        j202_soc_core_ahb2apb_00_N89) );
  sky130_fd_sc_hd__nand3_1 U30054 ( .A(n24818), .B(n24817), .C(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[0]), .Y(n24819) );
  sky130_fd_sc_hd__o21ai_1 U30055 ( .A1(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[0]), .A2(n24949), .B1(
        n24819), .Y(j202_soc_core_cmt_core_00_cmt_apb_00_nxt_state_0_) );
  sky130_fd_sc_hd__nor2_1 U30057 ( .A(n27619), .B(n11894), .Y(
        j202_soc_core_ahb2apb_00_N55) );
  sky130_fd_sc_hd__nor2_1 U30058 ( .A(n24820), .B(n24949), .Y(
        j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen) );
  sky130_fd_sc_hd__nand2_1 U30059 ( .A(n24896), .B(n27732), .Y(n24883) );
  sky130_fd_sc_hd__nand2_1 U30060 ( .A(n24883), .B(
        j202_soc_core_cmt_core_00_str0), .Y(n24821) );
  sky130_fd_sc_hd__o21ai_1 U30062 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[0]), .A2(
        j202_soc_core_cmt_core_00_str0), .B1(n24823), .Y(n24822) );
  sky130_fd_sc_hd__nand2_1 U30063 ( .A(n28619), .B(n24822), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[0]) );
  sky130_fd_sc_hd__a211oi_1 U30064 ( .A1(n24824), .A2(n24823), .B1(n24825), 
        .C1(n26284), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[1])
         );
  sky130_fd_sc_hd__nor2_1 U30066 ( .A(n24826), .B(n26284), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[2]) );
  sky130_fd_sc_hd__a211oi_1 U30067 ( .A1(n24829), .A2(n24828), .B1(n24827), 
        .C1(n26284), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[3])
         );
  sky130_fd_sc_hd__a211oi_1 U30068 ( .A1(n24832), .A2(n24831), .B1(n26284), 
        .C1(n24830), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[4])
         );
  sky130_fd_sc_hd__nand2_1 U30069 ( .A(n24834), .B(n24833), .Y(n24835) );
  sky130_fd_sc_hd__nand2_1 U30070 ( .A(n24835), .B(n28619), .Y(n24837) );
  sky130_fd_sc_hd__nor2_1 U30071 ( .A(n24837), .B(n24836), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[6]) );
  sky130_fd_sc_hd__nor2_1 U30072 ( .A(n24839), .B(n24838), .Y(n24840) );
  sky130_fd_sc_hd__a211oi_1 U30073 ( .A1(n24839), .A2(n24838), .B1(n26284), 
        .C1(n24840), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[8])
         );
  sky130_fd_sc_hd__xnor2_1 U30074 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[9]), .B(n24840), .Y(
        n24841) );
  sky130_fd_sc_hd__nor2_1 U30075 ( .A(n26284), .B(n24841), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[9]) );
  sky130_fd_sc_hd__nor2_1 U30076 ( .A(j202_soc_core_cmt_core_00_reg_addr[3]), 
        .B(n24842), .Y(n24956) );
  sky130_fd_sc_hd__nand2_1 U30077 ( .A(n24843), .B(n24956), .Y(n27829) );
  sky130_fd_sc_hd__nand2_1 U30078 ( .A(n24845), .B(
        j202_soc_core_cmt_core_00_wdata_cnt0[0]), .Y(n24844) );
  sky130_fd_sc_hd__o21ai_1 U30079 ( .A1(n24846), .A2(n24845), .B1(n24844), .Y(
        n81) );
  sky130_fd_sc_hd__nand2_1 U30080 ( .A(n27829), .B(
        j202_soc_core_cmt_core_00_cks0[1]), .Y(n24847) );
  sky130_fd_sc_hd__xnor2_1 U30082 ( .A(j202_soc_core_cmt_core_00_const0[1]), 
        .B(j202_soc_core_cmt_core_00_cnt0[1]), .Y(n24849) );
  sky130_fd_sc_hd__xnor2_1 U30083 ( .A(j202_soc_core_cmt_core_00_const0[3]), 
        .B(j202_soc_core_cmt_core_00_cnt0[3]), .Y(n24848) );
  sky130_fd_sc_hd__xnor2_1 U30084 ( .A(j202_soc_core_cmt_core_00_const0[8]), 
        .B(j202_soc_core_cmt_core_00_cnt0[8]), .Y(n24851) );
  sky130_fd_sc_hd__xnor2_1 U30085 ( .A(j202_soc_core_cmt_core_00_const0[2]), 
        .B(j202_soc_core_cmt_core_00_cnt0[2]), .Y(n24850) );
  sky130_fd_sc_hd__xor2_1 U30086 ( .A(j202_soc_core_cmt_core_00_const0[9]), 
        .B(j202_soc_core_cmt_core_00_cnt0[9]), .X(n24853) );
  sky130_fd_sc_hd__xor2_1 U30087 ( .A(j202_soc_core_cmt_core_00_const0[0]), 
        .B(j202_soc_core_cmt_core_00_cnt0[0]), .X(n24852) );
  sky130_fd_sc_hd__nor2_1 U30088 ( .A(n24853), .B(n24852), .Y(n24857) );
  sky130_fd_sc_hd__xnor2_1 U30089 ( .A(j202_soc_core_cmt_core_00_const0[6]), 
        .B(j202_soc_core_cmt_core_00_cnt0[6]), .Y(n24855) );
  sky130_fd_sc_hd__xnor2_1 U30090 ( .A(j202_soc_core_cmt_core_00_const0[5]), 
        .B(j202_soc_core_cmt_core_00_cnt0[5]), .Y(n24854) );
  sky130_fd_sc_hd__nand4_1 U30091 ( .A(n24859), .B(n24858), .C(n24857), .D(
        n24856), .Y(n28618) );
  sky130_fd_sc_hd__xnor2_1 U30092 ( .A(j202_soc_core_cmt_core_00_const0[10]), 
        .B(j202_soc_core_cmt_core_00_cnt0[10]), .Y(n24861) );
  sky130_fd_sc_hd__xnor2_1 U30093 ( .A(j202_soc_core_cmt_core_00_const0[12]), 
        .B(j202_soc_core_cmt_core_00_cnt0[12]), .Y(n24860) );
  sky130_fd_sc_hd__xnor2_1 U30094 ( .A(j202_soc_core_cmt_core_00_const0[4]), 
        .B(j202_soc_core_cmt_core_00_cnt0[4]), .Y(n24863) );
  sky130_fd_sc_hd__xnor2_1 U30095 ( .A(j202_soc_core_cmt_core_00_const0[7]), 
        .B(j202_soc_core_cmt_core_00_cnt0[7]), .Y(n24862) );
  sky130_fd_sc_hd__xnor2_1 U30096 ( .A(j202_soc_core_cmt_core_00_const0[14]), 
        .B(j202_soc_core_cmt_core_00_cnt0[14]), .Y(n24865) );
  sky130_fd_sc_hd__xnor2_1 U30097 ( .A(j202_soc_core_cmt_core_00_const0[13]), 
        .B(j202_soc_core_cmt_core_00_cnt0[13]), .Y(n24864) );
  sky130_fd_sc_hd__xnor2_1 U30098 ( .A(j202_soc_core_cmt_core_00_const0[15]), 
        .B(j202_soc_core_cmt_core_00_cnt0[15]), .Y(n24867) );
  sky130_fd_sc_hd__xnor2_1 U30099 ( .A(j202_soc_core_cmt_core_00_const0[11]), 
        .B(j202_soc_core_cmt_core_00_cnt0[11]), .Y(n24866) );
  sky130_fd_sc_hd__nand4_1 U30100 ( .A(n24871), .B(n24870), .C(n24869), .D(
        n24868), .Y(n28617) );
  sky130_fd_sc_hd__nor2_1 U30101 ( .A(n28618), .B(n28617), .Y(n24872) );
  sky130_fd_sc_hd__nor2_1 U30102 ( .A(n27482), .B(n24872), .Y(n27471) );
  sky130_fd_sc_hd__nand2_1 U30103 ( .A(n27471), .B(n24873), .Y(n26288) );
  sky130_fd_sc_hd__nor2_1 U30104 ( .A(j202_soc_core_cmt_core_00_cnt0[0]), .B(
        n24874), .Y(n24875) );
  sky130_fd_sc_hd__a21oi_1 U30105 ( .A1(n26288), .A2(
        j202_soc_core_cmt_core_00_cnt0[0]), .B1(n24875), .Y(n24877) );
  sky130_fd_sc_hd__nand2_1 U30106 ( .A(n27482), .B(
        j202_soc_core_cmt_core_00_wdata_cnt0[0]), .Y(n24876) );
  sky130_fd_sc_hd__o21ai_1 U30107 ( .A1(n27482), .A2(n24877), .B1(n24876), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[0]) );
  sky130_fd_sc_hd__a21oi_1 U30108 ( .A1(n26281), .A2(
        j202_soc_core_cmt_core_00_cnt0[0]), .B1(
        j202_soc_core_cmt_core_00_cnt0[1]), .Y(n24878) );
  sky130_fd_sc_hd__nand2_1 U30109 ( .A(j202_soc_core_cmt_core_00_cnt0[0]), .B(
        j202_soc_core_cmt_core_00_cnt0[1]), .Y(n25568) );
  sky130_fd_sc_hd__nor2_1 U30110 ( .A(n28619), .B(n27471), .Y(n26283) );
  sky130_fd_sc_hd__o22ai_1 U30112 ( .A1(n27473), .A2(n27611), .B1(n24878), 
        .B2(n25560), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[1])
         );
  sky130_fd_sc_hd__nor2_1 U30113 ( .A(n25568), .B(n26288), .Y(n25563) );
  sky130_fd_sc_hd__a22oi_1 U30114 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[2]), .A2(n27482), .B1(n25563), 
        .B2(n25562), .Y(n24879) );
  sky130_fd_sc_hd__nand3_1 U30116 ( .A(n24896), .B(n24955), .C(n24956), .Y(
        n27827) );
  sky130_fd_sc_hd__nand2_1 U30117 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[2]), .Y(n24880) );
  sky130_fd_sc_hd__o21ai_1 U30118 ( .A1(n24948), .A2(n27827), .B1(n24880), .Y(
        n77) );
  sky130_fd_sc_hd__nand2_1 U30119 ( .A(n27829), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[2]), .Y(n24881) );
  sky130_fd_sc_hd__nand2_1 U30121 ( .A(n24883), .B(
        j202_soc_core_cmt_core_00_str1), .Y(n24882) );
  sky130_fd_sc_hd__o21ai_1 U30122 ( .A1(n27611), .A2(n24883), .B1(n24882), .Y(
        n32) );
  sky130_fd_sc_hd__o21ai_1 U30123 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[0]), .A2(
        j202_soc_core_cmt_core_00_str1), .B1(n24885), .Y(n24884) );
  sky130_fd_sc_hd__nand2_1 U30124 ( .A(n28622), .B(n24884), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[0]) );
  sky130_fd_sc_hd__a211oi_1 U30125 ( .A1(n24886), .A2(n24885), .B1(n24887), 
        .C1(n26300), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[1])
         );
  sky130_fd_sc_hd__nor2_1 U30127 ( .A(n24888), .B(n26300), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[2]) );
  sky130_fd_sc_hd__a211oi_1 U30128 ( .A1(n24891), .A2(n24890), .B1(n24889), 
        .C1(n26300), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[3])
         );
  sky130_fd_sc_hd__a211oi_1 U30129 ( .A1(n24894), .A2(n24893), .B1(n26300), 
        .C1(n24892), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[5])
         );
  sky130_fd_sc_hd__nor2_1 U30130 ( .A(j202_soc_core_cmt_core_00_reg_addr[2]), 
        .B(n24895), .Y(n24950) );
  sky130_fd_sc_hd__nand2_1 U30131 ( .A(n24946), .B(n24957), .Y(n27831) );
  sky130_fd_sc_hd__nand2_1 U30132 ( .A(n27831), .B(
        j202_soc_core_cmt_core_00_cks1[0]), .Y(n24897) );
  sky130_fd_sc_hd__o21ai_1 U30133 ( .A1(n27731), .A2(n27831), .B1(n24897), .Y(
        n82) );
  sky130_fd_sc_hd__a211oi_1 U30134 ( .A1(n24900), .A2(n24899), .B1(n26300), 
        .C1(n24898), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[7])
         );
  sky130_fd_sc_hd__xnor2_1 U30135 ( .A(n24902), .B(n24901), .Y(n24903) );
  sky130_fd_sc_hd__nor2_1 U30136 ( .A(n26300), .B(n24903), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[9]) );
  sky130_fd_sc_hd__nand2_1 U30137 ( .A(n27831), .B(
        j202_soc_core_cmt_core_00_cks1[1]), .Y(n24904) );
  sky130_fd_sc_hd__o21ai_1 U30138 ( .A1(n27611), .A2(n27831), .B1(n24904), .Y(
        n34) );
  sky130_fd_sc_hd__nand2_1 U30139 ( .A(n24906), .B(n27491), .Y(n24935) );
  sky130_fd_sc_hd__xnor2_1 U30140 ( .A(j202_soc_core_cmt_core_00_const1[6]), 
        .B(j202_soc_core_cmt_core_00_cnt1[6]), .Y(n24908) );
  sky130_fd_sc_hd__xnor2_1 U30141 ( .A(j202_soc_core_cmt_core_00_const1[10]), 
        .B(j202_soc_core_cmt_core_00_cnt1[10]), .Y(n24907) );
  sky130_fd_sc_hd__xnor2_1 U30142 ( .A(j202_soc_core_cmt_core_00_const1[14]), 
        .B(j202_soc_core_cmt_core_00_cnt1[14]), .Y(n24910) );
  sky130_fd_sc_hd__xnor2_1 U30143 ( .A(j202_soc_core_cmt_core_00_const1[1]), 
        .B(j202_soc_core_cmt_core_00_cnt1[1]), .Y(n24909) );
  sky130_fd_sc_hd__xor2_1 U30144 ( .A(j202_soc_core_cmt_core_00_const1[9]), 
        .B(j202_soc_core_cmt_core_00_cnt1[9]), .X(n24912) );
  sky130_fd_sc_hd__xor2_1 U30145 ( .A(j202_soc_core_cmt_core_00_const1[0]), 
        .B(j202_soc_core_cmt_core_00_cnt1[0]), .X(n24911) );
  sky130_fd_sc_hd__nor2_1 U30146 ( .A(n24912), .B(n24911), .Y(n24916) );
  sky130_fd_sc_hd__xnor2_1 U30147 ( .A(j202_soc_core_cmt_core_00_const1[7]), 
        .B(j202_soc_core_cmt_core_00_cnt1[7]), .Y(n24914) );
  sky130_fd_sc_hd__xnor2_1 U30148 ( .A(j202_soc_core_cmt_core_00_const1[13]), 
        .B(j202_soc_core_cmt_core_00_cnt1[13]), .Y(n24913) );
  sky130_fd_sc_hd__nand4_1 U30149 ( .A(n24918), .B(n24917), .C(n24916), .D(
        n24915), .Y(n24932) );
  sky130_fd_sc_hd__xnor2_1 U30150 ( .A(j202_soc_core_cmt_core_00_const1[11]), 
        .B(j202_soc_core_cmt_core_00_cnt1[11]), .Y(n24920) );
  sky130_fd_sc_hd__xnor2_1 U30151 ( .A(j202_soc_core_cmt_core_00_const1[4]), 
        .B(j202_soc_core_cmt_core_00_cnt1[4]), .Y(n24919) );
  sky130_fd_sc_hd__xnor2_1 U30152 ( .A(j202_soc_core_cmt_core_00_const1[12]), 
        .B(j202_soc_core_cmt_core_00_cnt1[12]), .Y(n24922) );
  sky130_fd_sc_hd__xnor2_1 U30153 ( .A(j202_soc_core_cmt_core_00_const1[2]), 
        .B(j202_soc_core_cmt_core_00_cnt1[2]), .Y(n24921) );
  sky130_fd_sc_hd__xnor2_1 U30154 ( .A(j202_soc_core_cmt_core_00_const1[3]), 
        .B(j202_soc_core_cmt_core_00_cnt1[3]), .Y(n24924) );
  sky130_fd_sc_hd__xnor2_1 U30155 ( .A(j202_soc_core_cmt_core_00_const1[15]), 
        .B(j202_soc_core_cmt_core_00_cnt1[15]), .Y(n24923) );
  sky130_fd_sc_hd__xnor2_1 U30156 ( .A(j202_soc_core_cmt_core_00_const1[8]), 
        .B(j202_soc_core_cmt_core_00_cnt1[8]), .Y(n24926) );
  sky130_fd_sc_hd__xnor2_1 U30157 ( .A(j202_soc_core_cmt_core_00_const1[5]), 
        .B(j202_soc_core_cmt_core_00_cnt1[5]), .Y(n24925) );
  sky130_fd_sc_hd__nand4_1 U30158 ( .A(n24930), .B(n24929), .C(n24928), .D(
        n24927), .Y(n24931) );
  sky130_fd_sc_hd__nor2_1 U30159 ( .A(n24932), .B(n24931), .Y(n28620) );
  sky130_fd_sc_hd__nor2_1 U30160 ( .A(n24939), .B(n28620), .Y(n24934) );
  sky130_fd_sc_hd__a22oi_1 U30161 ( .A1(n27498), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[0]), .B1(n28622), .B2(
        j202_soc_core_cmt_core_00_cnt1[0]), .Y(n24933) );
  sky130_fd_sc_hd__o21ai_1 U30162 ( .A1(n24935), .A2(n24934), .B1(n24933), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[0]) );
  sky130_fd_sc_hd__nor2_1 U30163 ( .A(n28620), .B(n24935), .Y(n27489) );
  sky130_fd_sc_hd__a21oi_1 U30164 ( .A1(n27489), .A2(n24939), .B1(n28622), .Y(
        n24943) );
  sky130_fd_sc_hd__nor3_1 U30165 ( .A(j202_soc_core_cmt_core_00_cnt1[1]), .B(
        n26301), .C(n24939), .Y(n24936) );
  sky130_fd_sc_hd__a21oi_1 U30166 ( .A1(n27498), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[1]), .B1(n24936), .Y(n24937) );
  sky130_fd_sc_hd__nand2_1 U30168 ( .A(n27498), .B(
        j202_soc_core_cmt_core_00_wdata_cnt0[2]), .Y(n24942) );
  sky130_fd_sc_hd__o211ai_1 U30170 ( .A1(j202_soc_core_cmt_core_00_cnt1[2]), 
        .A2(j202_soc_core_cmt_core_00_cnt1[1]), .B1(n27489), .C1(n24940), .Y(
        n24941) );
  sky130_fd_sc_hd__o211ai_1 U30171 ( .A1(n24944), .A2(n24943), .B1(n24942), 
        .C1(n24941), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[2])
         );
  sky130_fd_sc_hd__nand2_1 U30172 ( .A(n27831), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[2]), .Y(n24945) );
  sky130_fd_sc_hd__o21ai_1 U30173 ( .A1(n24948), .A2(n27831), .B1(n24945), .Y(
        n76) );
  sky130_fd_sc_hd__nand2_1 U30174 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[2]), .Y(n24947) );
  sky130_fd_sc_hd__o21ai_1 U30175 ( .A1(n24948), .A2(n27833), .B1(n24947), .Y(
        n78) );
  sky130_fd_sc_hd__nor2_1 U30176 ( .A(j202_soc_core_pwrite[0]), .B(n24949), 
        .Y(n27733) );
  sky130_fd_sc_hd__nand2_1 U30177 ( .A(n27733), .B(n24950), .Y(n24952) );
  sky130_fd_sc_hd__nor2_1 U30178 ( .A(n24951), .B(n24952), .Y(n27836) );
  sky130_fd_sc_hd__a22oi_1 U30179 ( .A1(n27836), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[2]), .B1(n27835), .B2(
        j202_soc_core_cmt_core_00_const1[2]), .Y(n24964) );
  sky130_fd_sc_hd__and3_1 U30180 ( .A(n24955), .B(n27733), .C(n24956), .X(
        n27838) );
  sky130_fd_sc_hd__and3_1 U30181 ( .A(n24955), .B(n27733), .C(n24954), .X(
        n27837) );
  sky130_fd_sc_hd__a22oi_1 U30182 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[2]), .B1(n27837), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[2]), .Y(
        n24963) );
  sky130_fd_sc_hd__nand2_1 U30183 ( .A(n24957), .B(n27733), .Y(n24959) );
  sky130_fd_sc_hd__nor2_1 U30184 ( .A(n24958), .B(n24959), .Y(n27839) );
  sky130_fd_sc_hd__nand2_1 U30185 ( .A(n27839), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[2]), .Y(n24962) );
  sky130_fd_sc_hd__nor2_1 U30186 ( .A(n24960), .B(n24959), .Y(n27840) );
  sky130_fd_sc_hd__nand2_1 U30187 ( .A(n27840), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[2]), .Y(
        n24961) );
  sky130_fd_sc_hd__nand4_1 U30188 ( .A(n24964), .B(n24963), .C(n24962), .D(
        n24961), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[2]) );
  sky130_fd_sc_hd__nand2_1 U30189 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[2]), .Y(n24965) );
  sky130_fd_sc_hd__o21ai_1 U30190 ( .A1(n24966), .A2(n27983), .B1(n24965), .Y(
        n51) );
  sky130_fd_sc_hd__o22ai_1 U30191 ( .A1(n28615), .A2(n27021), .B1(n24967), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U30192 ( .A1(n28615), .A2(n27990), .B1(n24968), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U30193 ( .A1(n28615), .A2(n28535), .B1(n24983), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__nand4b_1 U30194 ( .A_N(n24969), .B(n28888), .C(
        j202_soc_core_intc_core_00_bs_addr[5]), .D(n28884), .Y(n24973) );
  sky130_fd_sc_hd__nor2_1 U30195 ( .A(j202_soc_core_intc_core_00_bs_addr[8]), 
        .B(j202_soc_core_intc_core_00_bs_addr[7]), .Y(n24971) );
  sky130_fd_sc_hd__nand3_1 U30196 ( .A(n24972), .B(n24971), .C(n24970), .Y(
        n28883) );
  sky130_fd_sc_hd__nor2_1 U30197 ( .A(n24973), .B(n28883), .Y(n27308) );
  sky130_fd_sc_hd__nand2_1 U30198 ( .A(n27308), .B(j202_soc_core_pwrite[1]), 
        .Y(n28526) );
  sky130_fd_sc_hd__o22ai_1 U30199 ( .A1(n28615), .A2(n28526), .B1(n24974), 
        .B2(n28524), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__nor2_1 U30200 ( .A(n28882), .B(n24975), .Y(n27757) );
  sky130_fd_sc_hd__o22ai_1 U30201 ( .A1(n28615), .A2(n28547), .B1(n24976), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__nor2_1 U30202 ( .A(n28882), .B(n24977), .Y(n27583) );
  sky130_fd_sc_hd__o22ai_1 U30203 ( .A1(n28615), .A2(n28538), .B1(n24978), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__nor2_1 U30204 ( .A(n28882), .B(n24979), .Y(n28520) );
  sky130_fd_sc_hd__nor2_1 U30205 ( .A(n28590), .B(n28520), .Y(n28519) );
  sky130_fd_sc_hd__o22ai_1 U30206 ( .A1(n28615), .A2(n28541), .B1(n24980), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__nor2_1 U30207 ( .A(n28882), .B(n27306), .Y(n27010) );
  sky130_fd_sc_hd__o22ai_1 U30208 ( .A1(n28544), .A2(n28615), .B1(n24981), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__a21oi_1 U30209 ( .A1(n27857), .A2(
        j202_soc_core_intc_core_00_rg_eimk[2]), .B1(n27758), .Y(n24982) );
  sky130_fd_sc_hd__o21ai_1 U30210 ( .A1(n24983), .A2(n27760), .B1(n24982), .Y(
        n24984) );
  sky130_fd_sc_hd__a21oi_1 U30211 ( .A1(n27860), .A2(
        j202_soc_core_intc_core_00_rg_ipr[98]), .B1(n24984), .Y(n24991) );
  sky130_fd_sc_hd__a22oi_1 U30212 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[2]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[2]), .Y(n24986) );
  sky130_fd_sc_hd__a22oi_1 U30213 ( .A1(n27852), .A2(
        j202_soc_core_intc_core_00_rg_ipr[66]), .B1(n27856), .B2(
        j202_soc_core_intc_core_00_rg_itgt[80]), .Y(n24985) );
  sky130_fd_sc_hd__o211ai_1 U30214 ( .A1(n24987), .A2(n27676), .B1(n24986), 
        .C1(n24985), .Y(n24988) );
  sky130_fd_sc_hd__a21oi_1 U30215 ( .A1(n27869), .A2(
        j202_soc_core_intc_core_00_rg_itgt[72]), .B1(n24988), .Y(n24990) );
  sky130_fd_sc_hd__a22oi_1 U30216 ( .A1(n27862), .A2(
        j202_soc_core_intc_core_00_rg_ipr[34]), .B1(n27861), .B2(
        j202_soc_core_intc_core_00_rg_itgt[88]), .Y(n24989) );
  sky130_fd_sc_hd__nand3_1 U30217 ( .A(n24991), .B(n24990), .C(n24989), .Y(
        j202_soc_core_ahb2apb_01_N130) );
  sky130_fd_sc_hd__nor2_1 U30218 ( .A(n26211), .B(n24992), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N360) );
  sky130_fd_sc_hd__nor2_1 U30219 ( .A(n26211), .B(n24993), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N359) );
  sky130_fd_sc_hd__nor2_1 U30220 ( .A(n26039), .B(n26007), .Y(n28221) );
  sky130_fd_sc_hd__nor2_1 U30221 ( .A(n28158), .B(n28126), .Y(n28129) );
  sky130_fd_sc_hd__a21oi_1 U30222 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[1]), .A2(n25026), .B1(n28129), 
        .Y(n24994) );
  sky130_fd_sc_hd__nor2_1 U30223 ( .A(n28590), .B(n24994), .Y(
        j202_soc_core_wbqspiflash_00_N739) );
  sky130_fd_sc_hd__a211o_1 U30224 ( .A1(n28221), .A2(n26116), .B1(n28590), 
        .C1(n24995), .X(j202_soc_core_wbqspiflash_00_N738) );
  sky130_fd_sc_hd__nand2_1 U30225 ( .A(n24996), .B(n29594), .Y(
        j202_soc_core_wbqspiflash_00_N743) );
  sky130_fd_sc_hd__nand2_1 U30227 ( .A(n26516), .B(n26329), .Y(n25194) );
  sky130_fd_sc_hd__o22ai_1 U30228 ( .A1(n24998), .A2(n26070), .B1(n25714), 
        .B2(n27349), .Y(n24999) );
  sky130_fd_sc_hd__a21oi_1 U30229 ( .A1(n26516), .A2(n25000), .B1(n24999), .Y(
        n25001) );
  sky130_fd_sc_hd__o21ai_1 U30230 ( .A1(n25194), .A2(n25002), .B1(n25001), .Y(
        j202_soc_core_j22_cpu_rf_N3379) );
  sky130_fd_sc_hd__and3_1 U30231 ( .A(n26155), .B(
        j202_soc_core_qspi_wb_addr[2]), .C(n26032), .X(n28078) );
  sky130_fd_sc_hd__nand2_1 U30232 ( .A(n28228), .B(n25916), .Y(n28086) );
  sky130_fd_sc_hd__nand2_1 U30233 ( .A(n25003), .B(n28237), .Y(n26018) );
  sky130_fd_sc_hd__o21ai_1 U30234 ( .A1(n28086), .A2(n26018), .B1(n28187), .Y(
        n25005) );
  sky130_fd_sc_hd__nand2_1 U30235 ( .A(n25004), .B(n26188), .Y(n28250) );
  sky130_fd_sc_hd__nand2_1 U30236 ( .A(n26035), .B(n25954), .Y(n28097) );
  sky130_fd_sc_hd__nand2b_1 U30237 ( .A_N(n28097), .B(n28058), .Y(n28083) );
  sky130_fd_sc_hd__a211oi_1 U30239 ( .A1(n28078), .A2(
        j202_soc_core_qspi_wb_addr[3]), .B1(n25005), .C1(n28238), .Y(n28265)
         );
  sky130_fd_sc_hd__nand2_1 U30240 ( .A(n26009), .B(n26255), .Y(n25900) );
  sky130_fd_sc_hd__nor2_1 U30241 ( .A(j202_soc_core_wbqspiflash_00_spif_cmd), 
        .B(j202_soc_core_wbqspiflash_00_spif_ctrl), .Y(n28207) );
  sky130_fd_sc_hd__nand2_1 U30242 ( .A(n28089), .B(n26171), .Y(n26014) );
  sky130_fd_sc_hd__a21o_1 U30243 ( .A1(n28103), .A2(n28207), .B1(n28215), .X(
        n28258) );
  sky130_fd_sc_hd__nand2_1 U30244 ( .A(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled), .B(n28258), .Y(n28075) );
  sky130_fd_sc_hd__nand2_1 U30245 ( .A(n25884), .B(n28075), .Y(n28085) );
  sky130_fd_sc_hd__a31oi_1 U30246 ( .A1(n28090), .A2(n28089), .A3(
        j202_soc_core_qspi_wb_addr[23]), .B1(n28085), .Y(n25008) );
  sky130_fd_sc_hd__nand3_1 U30247 ( .A(n28080), .B(n28079), .C(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]), .Y(n25007) );
  sky130_fd_sc_hd__nand2_1 U30248 ( .A(n26119), .B(n28079), .Y(n28108) );
  sky130_fd_sc_hd__nand2_1 U30249 ( .A(n28259), .B(
        j202_soc_core_wbqspiflash_00_spif_data[31]), .Y(n25006) );
  sky130_fd_sc_hd__nand4_1 U30250 ( .A(n28265), .B(n25008), .C(n25007), .D(
        n25006), .Y(n10506) );
  sky130_fd_sc_hd__nand2_1 U30251 ( .A(n28737), .B(n26198), .Y(n28748) );
  sky130_fd_sc_hd__nand4_1 U30252 ( .A(n28748), .B(n25010), .C(n25009), .D(
        n28747), .Y(j202_soc_core_wbqspiflash_00_lldriver_N312) );
  sky130_fd_sc_hd__a211oi_1 U30254 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[7]), .A2(n28064), .B1(
        n28058), .C1(n25014), .Y(n25013) );
  sky130_fd_sc_hd__nor2_1 U30255 ( .A(n28063), .B(n25013), .Y(
        j202_soc_core_wbqspiflash_00_N621) );
  sky130_fd_sc_hd__xnor2_1 U30256 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[8]), .B(n25014), .Y(n25015)
         );
  sky130_fd_sc_hd__a21oi_1 U30257 ( .A1(n25015), .A2(
        j202_soc_core_wbqspiflash_00_state[0]), .B1(n28063), .Y(
        j202_soc_core_wbqspiflash_00_N622) );
  sky130_fd_sc_hd__a21oi_1 U30258 ( .A1(n25016), .A2(
        j202_soc_core_wbqspiflash_00_reset_counter[9]), .B1(n28058), .Y(n25017) );
  sky130_fd_sc_hd__a21oi_1 U30259 ( .A1(n25017), .A2(n26183), .B1(n28063), .Y(
        j202_soc_core_wbqspiflash_00_N623) );
  sky130_fd_sc_hd__nor2_1 U30260 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[0]), .B(n28751), .Y(
        j202_soc_core_wbqspiflash_00_N614) );
  sky130_fd_sc_hd__xnor2_1 U30261 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[2]), .B(n28749), .Y(n25018)
         );
  sky130_fd_sc_hd__a21oi_1 U30262 ( .A1(n25018), .A2(
        j202_soc_core_wbqspiflash_00_state[0]), .B1(n28063), .Y(
        j202_soc_core_wbqspiflash_00_N616) );
  sky130_fd_sc_hd__nand2_1 U30263 ( .A(n25019), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[3]), .Y(n25021) );
  sky130_fd_sc_hd__a21oi_1 U30264 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[2]), .A2(
        j202_soc_core_wbqspiflash_00_reset_counter[3]), .B1(n28058), .Y(n25020) );
  sky130_fd_sc_hd__a31oi_1 U30265 ( .A1(n25021), .A2(n25020), .A3(n28056), 
        .B1(n28063), .Y(j202_soc_core_wbqspiflash_00_N617) );
  sky130_fd_sc_hd__nor2_1 U30266 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[8]), .B(n25022), .Y(n28094)
         );
  sky130_fd_sc_hd__nand2_1 U30267 ( .A(n28094), .B(n25023), .Y(
        j202_soc_core_wbqspiflash_00_N85) );
  sky130_fd_sc_hd__nor2_1 U30269 ( .A(n28163), .B(n27874), .Y(
        j202_soc_core_wbqspiflash_00_N669) );
  sky130_fd_sc_hd__nor2_1 U30270 ( .A(n25057), .B(n26349), .Y(n25040) );
  sky130_fd_sc_hd__nand2_1 U30271 ( .A(n25057), .B(n26325), .Y(n26671) );
  sky130_fd_sc_hd__nand2_1 U30272 ( .A(n27383), .B(n26722), .Y(n26672) );
  sky130_fd_sc_hd__nand3_1 U30273 ( .A(n26671), .B(n26326), .C(n26672), .Y(
        n25028) );
  sky130_fd_sc_hd__o21ai_1 U30274 ( .A1(n18916), .A2(n25030), .B1(n25029), .Y(
        n25039) );
  sky130_fd_sc_hd__o22ai_1 U30275 ( .A1(n25821), .A2(n26419), .B1(n26426), 
        .B2(n26418), .Y(n25038) );
  sky130_fd_sc_hd__o22ai_1 U30276 ( .A1(n25229), .A2(n26416), .B1(n25788), 
        .B2(n26427), .Y(n25031) );
  sky130_fd_sc_hd__a21oi_1 U30277 ( .A1(n26338), .A2(n27435), .B1(n25031), .Y(
        n25036) );
  sky130_fd_sc_hd__o22a_1 U30278 ( .A1(n27383), .A2(n26423), .B1(n26432), .B2(
        n26672), .X(n25032) );
  sky130_fd_sc_hd__o21ai_0 U30279 ( .A1(n26336), .A2(n26424), .B1(n25032), .Y(
        n25033) );
  sky130_fd_sc_hd__a21oi_1 U30280 ( .A1(n26341), .A2(n26718), .B1(n25033), .Y(
        n25035) );
  sky130_fd_sc_hd__nand2_1 U30281 ( .A(n26342), .B(n25061), .Y(n25034) );
  sky130_fd_sc_hd__nand4_1 U30282 ( .A(n25036), .B(n25035), .C(n26344), .D(
        n25034), .Y(n25037) );
  sky130_fd_sc_hd__or4_1 U30283 ( .A(n25040), .B(n25039), .C(n25038), .D(
        n25037), .X(n25041) );
  sky130_fd_sc_hd__a21oi_1 U30284 ( .A1(n25042), .A2(n26409), .B1(n25041), .Y(
        n25044) );
  sky130_fd_sc_hd__nor2_1 U30286 ( .A(n26946), .B(n12160), .Y(
        j202_soc_core_j22_cpu_rf_N2653) );
  sky130_fd_sc_hd__mux2i_1 U30287 ( .A0(n12160), .A1(n27276), .S(n27460), .Y(
        j202_soc_core_j22_cpu_rf_N3281) );
  sky130_fd_sc_hd__o22ai_1 U30288 ( .A1(n27276), .A2(n26378), .B1(n26449), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N3244) );
  sky130_fd_sc_hd__o22ai_1 U30289 ( .A1(n27276), .A2(n26899), .B1(n26898), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N3321) );
  sky130_fd_sc_hd__o22ai_1 U30290 ( .A1(n27276), .A2(n11141), .B1(n27124), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N2689) );
  sky130_fd_sc_hd__o22ai_1 U30291 ( .A1(n27276), .A2(n27466), .B1(n27465), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N2763) );
  sky130_fd_sc_hd__o22ai_1 U30292 ( .A1(n27276), .A2(n27209), .B1(n23039), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N2726) );
  sky130_fd_sc_hd__o22ai_1 U30293 ( .A1(n27276), .A2(n27213), .B1(n27212), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N2800) );
  sky130_fd_sc_hd__o22ai_1 U30294 ( .A1(n27276), .A2(n27215), .B1(n27214), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N2911) );
  sky130_fd_sc_hd__o22ai_1 U30295 ( .A1(n27276), .A2(n27223), .B1(n27222), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N3022) );
  sky130_fd_sc_hd__o22ai_1 U30296 ( .A1(n27276), .A2(n27226), .B1(n23079), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N3133) );
  sky130_fd_sc_hd__o22ai_1 U30297 ( .A1(n27276), .A2(n27219), .B1(n27218), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N2985) );
  sky130_fd_sc_hd__o22ai_1 U30298 ( .A1(n27276), .A2(n27228), .B1(n27227), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N3170) );
  sky130_fd_sc_hd__o22ai_1 U30299 ( .A1(n27276), .A2(n27333), .B1(n23178), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N3059) );
  sky130_fd_sc_hd__o22ai_1 U30300 ( .A1(n27276), .A2(n27221), .B1(n27220), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N2874) );
  sky130_fd_sc_hd__o22ai_1 U30301 ( .A1(n27276), .A2(n27211), .B1(n27210), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N3207) );
  sky130_fd_sc_hd__o22ai_1 U30302 ( .A1(n27276), .A2(n27217), .B1(n27216), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N2837) );
  sky130_fd_sc_hd__o22ai_1 U30303 ( .A1(n27276), .A2(n27225), .B1(n27224), 
        .B2(n12160), .Y(j202_soc_core_j22_cpu_rf_N2948) );
  sky130_fd_sc_hd__mux2i_1 U30304 ( .A0(n27276), .A1(n26325), .S(n27006), .Y(
        j202_soc_core_j22_cpu_ml_N313) );
  sky130_fd_sc_hd__a21oi_1 U30305 ( .A1(n25344), .A2(n12708), .B1(n26976), .Y(
        n25052) );
  sky130_fd_sc_hd__nand3_1 U30306 ( .A(n12356), .B(n25049), .C(n26872), .Y(
        n25051) );
  sky130_fd_sc_hd__a22oi_1 U30307 ( .A1(n25053), .A2(n26948), .B1(n12645), 
        .B2(n24650), .Y(n25054) );
  sky130_fd_sc_hd__o22ai_1 U30309 ( .A1(n27380), .A2(n26431), .B1(n25057), 
        .B2(n26412), .Y(n25068) );
  sky130_fd_sc_hd__xor2_1 U30310 ( .A(n26718), .B(n27380), .X(n26623) );
  sky130_fd_sc_hd__o22ai_1 U30311 ( .A1(n26571), .A2(n26416), .B1(n26415), 
        .B2(n26623), .Y(n25059) );
  sky130_fd_sc_hd__o22ai_1 U30312 ( .A1(n26701), .A2(n26419), .B1(n26705), 
        .B2(n26418), .Y(n25058) );
  sky130_fd_sc_hd__nor2_1 U30313 ( .A(n25059), .B(n25058), .Y(n25066) );
  sky130_fd_sc_hd__o21a_1 U30314 ( .A1(n26432), .A2(n27380), .B1(n26422), .X(
        n25060) );
  sky130_fd_sc_hd__o22ai_1 U30315 ( .A1(n26423), .A2(n25061), .B1(n26563), 
        .B2(n25060), .Y(n25062) );
  sky130_fd_sc_hd__a21oi_1 U30316 ( .A1(n25063), .A2(n25130), .B1(n25062), .Y(
        n25065) );
  sky130_fd_sc_hd__o22a_1 U30317 ( .A1(n26706), .A2(n26427), .B1(n26325), .B2(
        n26425), .X(n25064) );
  sky130_fd_sc_hd__nand4_1 U30318 ( .A(n25066), .B(n25065), .C(n25064), .D(
        n26411), .Y(n25067) );
  sky130_fd_sc_hd__nor2_1 U30319 ( .A(n25068), .B(n25067), .Y(n25072) );
  sky130_fd_sc_hd__nand2_1 U30320 ( .A(n26563), .B(n26443), .Y(n25069) );
  sky130_fd_sc_hd__nand2_1 U30321 ( .A(n25070), .B(n26409), .Y(n25071) );
  sky130_fd_sc_hd__buf_4 U30322 ( .A(n12363), .X(n25115) );
  sky130_fd_sc_hd__nor2_1 U30323 ( .A(n26946), .B(n25223), .Y(
        j202_soc_core_j22_cpu_rf_N2671) );
  sky130_fd_sc_hd__nand2_1 U30324 ( .A(n12740), .B(n27460), .Y(n25076) );
  sky130_fd_sc_hd__o22ai_1 U30326 ( .A1(n26378), .A2(n11102), .B1(n26449), 
        .B2(n25223), .Y(j202_soc_core_j22_cpu_rf_N3262) );
  sky130_fd_sc_hd__o22ai_1 U30327 ( .A1(n26899), .A2(n11102), .B1(n26898), 
        .B2(n25115), .Y(j202_soc_core_j22_cpu_rf_N3338) );
  sky130_fd_sc_hd__o22ai_1 U30328 ( .A1(n11141), .A2(n11102), .B1(n27124), 
        .B2(n25223), .Y(j202_soc_core_j22_cpu_rf_N2707) );
  sky130_fd_sc_hd__o21ai_1 U30329 ( .A1(n26951), .A2(n25223), .B1(n25078), .Y(
        j202_soc_core_j22_cpu_rf_N3374) );
  sky130_fd_sc_hd__nand2_1 U30330 ( .A(n12740), .B(n27339), .Y(n25080) );
  sky130_fd_sc_hd__o211ai_1 U30331 ( .A1(n26563), .A2(n25215), .B1(n25080), 
        .C1(n27346), .Y(j202_soc_core_j22_cpu_ml_N330) );
  sky130_fd_sc_hd__nand3_1 U30332 ( .A(n25083), .B(n25082), .C(n25081), .Y(
        n25084) );
  sky130_fd_sc_hd__a22oi_1 U30333 ( .A1(n27187), .A2(n25085), .B1(n27273), 
        .B2(n25084), .Y(n25086) );
  sky130_fd_sc_hd__nand2_1 U30334 ( .A(n27189), .B(n25086), .Y(
        j202_soc_core_j22_cpu_ml_machj[26]) );
  sky130_fd_sc_hd__o22ai_1 U30335 ( .A1(n25097), .A2(n27021), .B1(n25087), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U30336 ( .A1(n25097), .A2(n25534), .B1(n25088), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U30337 ( .A1(n25097), .A2(n27990), .B1(n25089), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U30338 ( .A1(n25097), .A2(n28535), .B1(n25090), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U30339 ( .A1(n25097), .A2(n28547), .B1(n25091), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U30340 ( .A1(n25097), .A2(n28538), .B1(n25099), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U30341 ( .A1(n25097), .A2(n28541), .B1(n25092), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U30342 ( .A1(n28544), .A2(n25097), .B1(n25093), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__nand3_1 U30343 ( .A(n25095), .B(j202_soc_core_pwrite[1]), 
        .C(n28884), .Y(n28594) );
  sky130_fd_sc_hd__nor2_1 U30344 ( .A(j202_soc_core_intc_core_00_bs_addr[7]), 
        .B(n28594), .Y(n25351) );
  sky130_fd_sc_hd__nor2_1 U30345 ( .A(n28590), .B(n25351), .Y(n25350) );
  sky130_fd_sc_hd__o22ai_1 U30346 ( .A1(n25097), .A2(n27194), .B1(n25096), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__a21oi_1 U30347 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[26]), .B1(n27758), .Y(n25098) );
  sky130_fd_sc_hd__o21ai_1 U30348 ( .A1(n25099), .A2(n27097), .B1(n25098), .Y(
        n25100) );
  sky130_fd_sc_hd__a21oi_1 U30349 ( .A1(j202_soc_core_intc_core_00_rg_ipr[58]), 
        .A2(n27862), .B1(n25100), .Y(n25105) );
  sky130_fd_sc_hd__a22o_1 U30350 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[26]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[90]), .X(n25101) );
  sky130_fd_sc_hd__a21oi_1 U30351 ( .A1(n27850), .A2(
        j202_soc_core_intc_core_00_rg_itgt[70]), .B1(n25101), .Y(n25104) );
  sky130_fd_sc_hd__a22oi_1 U30352 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[94]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[122]), .Y(n25103) );
  sky130_fd_sc_hd__nand2_1 U30353 ( .A(n27869), .B(
        j202_soc_core_intc_core_00_rg_itgt[78]), .Y(n25102) );
  sky130_fd_sc_hd__nand4_1 U30354 ( .A(n25105), .B(n25104), .C(n25103), .D(
        n25102), .Y(j202_soc_core_ahb2apb_01_N154) );
  sky130_fd_sc_hd__nand2_1 U30355 ( .A(n25107), .B(n25106), .Y(n25110) );
  sky130_fd_sc_hd__nand3_1 U30356 ( .A(n25111), .B(n25110), .C(n25109), .Y(
        j202_soc_core_ahb2aqu_00_N164) );
  sky130_fd_sc_hd__nand2_1 U30357 ( .A(n25112), .B(j202_soc_core_aquc_SEL__3_), 
        .Y(n27108) );
  sky130_fd_sc_hd__nand2_1 U30358 ( .A(n27108), .B(j202_soc_core_uart_div0[2]), 
        .Y(n25113) );
  sky130_fd_sc_hd__o22ai_1 U30360 ( .A1(n27333), .A2(n11102), .B1(n23178), 
        .B2(n25115), .Y(j202_soc_core_j22_cpu_rf_N3077) );
  sky130_fd_sc_hd__o22ai_1 U30361 ( .A1(n27466), .A2(n11102), .B1(n27465), 
        .B2(n25115), .Y(j202_soc_core_j22_cpu_rf_N2781) );
  sky130_fd_sc_hd__o22ai_1 U30362 ( .A1(n27209), .A2(n11102), .B1(n23039), 
        .B2(n25115), .Y(j202_soc_core_j22_cpu_rf_N2744) );
  sky130_fd_sc_hd__o22ai_1 U30363 ( .A1(n27221), .A2(n11102), .B1(n27220), 
        .B2(n25115), .Y(j202_soc_core_j22_cpu_rf_N2892) );
  sky130_fd_sc_hd__o22ai_1 U30364 ( .A1(n27211), .A2(n11102), .B1(n27210), 
        .B2(n25223), .Y(j202_soc_core_j22_cpu_rf_N3225) );
  sky130_fd_sc_hd__o22ai_1 U30365 ( .A1(n27213), .A2(n11102), .B1(n27212), 
        .B2(n25115), .Y(j202_soc_core_j22_cpu_rf_N2818) );
  sky130_fd_sc_hd__o22ai_1 U30366 ( .A1(n27215), .A2(n11102), .B1(n27214), 
        .B2(n25223), .Y(j202_soc_core_j22_cpu_rf_N2929) );
  sky130_fd_sc_hd__o22ai_1 U30367 ( .A1(n27223), .A2(n11661), .B1(n27222), 
        .B2(n25223), .Y(j202_soc_core_j22_cpu_rf_N3040) );
  sky130_fd_sc_hd__o22ai_1 U30368 ( .A1(n27217), .A2(n11102), .B1(n27216), 
        .B2(n25115), .Y(j202_soc_core_j22_cpu_rf_N2855) );
  sky130_fd_sc_hd__o22ai_1 U30369 ( .A1(n27225), .A2(n11102), .B1(n27224), 
        .B2(n25223), .Y(j202_soc_core_j22_cpu_rf_N2966) );
  sky130_fd_sc_hd__o22ai_1 U30370 ( .A1(n27226), .A2(n11102), .B1(n23079), 
        .B2(n25223), .Y(j202_soc_core_j22_cpu_rf_N3151) );
  sky130_fd_sc_hd__o22ai_1 U30371 ( .A1(n27219), .A2(n11102), .B1(n27218), 
        .B2(n25115), .Y(j202_soc_core_j22_cpu_rf_N3003) );
  sky130_fd_sc_hd__o22ai_1 U30372 ( .A1(n27228), .A2(n11102), .B1(n27227), 
        .B2(n25223), .Y(j202_soc_core_j22_cpu_rf_N3188) );
  sky130_fd_sc_hd__o21a_1 U30373 ( .A1(n26352), .A2(n25137), .B1(n26351), .X(
        n25120) );
  sky130_fd_sc_hd__nand2_1 U30374 ( .A(n25137), .B(n26323), .Y(n25119) );
  sky130_fd_sc_hd__o22a_1 U30375 ( .A1(n27386), .A2(n26431), .B1(n25121), .B2(
        n26412), .X(n25134) );
  sky130_fd_sc_hd__o22ai_1 U30376 ( .A1(n26701), .A2(n26427), .B1(n25788), 
        .B2(n26425), .Y(n25127) );
  sky130_fd_sc_hd__nand2_1 U30377 ( .A(n25122), .B(n25137), .Y(n26611) );
  sky130_fd_sc_hd__nand2_1 U30378 ( .A(n27386), .B(n26706), .Y(n26612) );
  sky130_fd_sc_hd__nand3_1 U30379 ( .A(n26612), .B(n26326), .C(n26611), .Y(
        n25123) );
  sky130_fd_sc_hd__o211ai_1 U30380 ( .A1(n26432), .A2(n26611), .B1(n25124), 
        .C1(n25123), .Y(n25125) );
  sky130_fd_sc_hd__o21bai_1 U30381 ( .A1(n26704), .A2(n26419), .B1_N(n25125), 
        .Y(n25126) );
  sky130_fd_sc_hd__nor2_1 U30382 ( .A(n25127), .B(n25126), .Y(n25133) );
  sky130_fd_sc_hd__o22ai_1 U30383 ( .A1(n25128), .A2(n26416), .B1(n26563), 
        .B2(n26424), .Y(n25129) );
  sky130_fd_sc_hd__a21oi_1 U30384 ( .A1(n25131), .A2(n25130), .B1(n25129), .Y(
        n25132) );
  sky130_fd_sc_hd__nand4_1 U30385 ( .A(n25134), .B(n25133), .C(n25132), .D(
        n26411), .Y(n25135) );
  sky130_fd_sc_hd__a21oi_1 U30386 ( .A1(n25136), .A2(n26409), .B1(n25135), .Y(
        n25139) );
  sky130_fd_sc_hd__nand2_1 U30387 ( .A(n12385), .B(n27192), .Y(n25141) );
  sky130_fd_sc_hd__o21ai_1 U30388 ( .A1(n27192), .A2(n25157), .B1(n25141), .Y(
        j202_soc_core_j22_cpu_rf_N3300) );
  sky130_fd_sc_hd__nand3_1 U30389 ( .A(n25144), .B(n25143), .C(n25142), .Y(
        n25145) );
  sky130_fd_sc_hd__a22oi_1 U30390 ( .A1(n27187), .A2(n22685), .B1(n27273), 
        .B2(n25145), .Y(n25146) );
  sky130_fd_sc_hd__nand2_1 U30391 ( .A(n27189), .B(n25146), .Y(
        j202_soc_core_j22_cpu_ml_machj[27]) );
  sky130_fd_sc_hd__a21oi_1 U30392 ( .A1(n25875), .A2(n25148), .B1(n26976), .Y(
        n25149) );
  sky130_fd_sc_hd__o21ai_1 U30393 ( .A1(n25150), .A2(n12917), .B1(n25149), .Y(
        j202_soc_core_j22_cpu_ml_maclj[27]) );
  sky130_fd_sc_hd__o22ai_1 U30394 ( .A1(n25151), .A2(n26070), .B1(n25714), 
        .B2(n25157), .Y(n25154) );
  sky130_fd_sc_hd__nor2_1 U30395 ( .A(n26951), .B(n25152), .Y(n25153) );
  sky130_fd_sc_hd__nor2_1 U30396 ( .A(n25154), .B(n25153), .Y(n25155) );
  sky130_fd_sc_hd__o21ai_1 U30397 ( .A1(n26951), .A2(n12488), .B1(n25155), .Y(
        j202_soc_core_j22_cpu_rf_N3375) );
  sky130_fd_sc_hd__xnor2_1 U30398 ( .A(n26061), .B(n26064), .Y(n25185) );
  sky130_fd_sc_hd__nand2b_1 U30399 ( .A_N(n26323), .B(n25159), .Y(n26405) );
  sky130_fd_sc_hd__o21ai_1 U30400 ( .A1(n26406), .A2(n26061), .B1(n26405), .Y(
        n25160) );
  sky130_fd_sc_hd__nand2_1 U30401 ( .A(n25160), .B(n26407), .Y(n25180) );
  sky130_fd_sc_hd__nand2_1 U30402 ( .A(n26077), .B(n26859), .Y(n25162) );
  sky130_fd_sc_hd__nand2_1 U30403 ( .A(n25165), .B(n26704), .Y(n26647) );
  sky130_fd_sc_hd__nand2_1 U30404 ( .A(n27399), .B(n26061), .Y(n26646) );
  sky130_fd_sc_hd__nand3_1 U30405 ( .A(n26647), .B(n26326), .C(n26646), .Y(
        n25161) );
  sky130_fd_sc_hd__o211ai_1 U30406 ( .A1(n26567), .A2(n26416), .B1(n25162), 
        .C1(n25161), .Y(n25164) );
  sky130_fd_sc_hd__o22ai_1 U30407 ( .A1(n26706), .A2(n26418), .B1(n26570), 
        .B2(n26419), .Y(n25163) );
  sky130_fd_sc_hd__nor2_1 U30408 ( .A(n25164), .B(n25163), .Y(n25174) );
  sky130_fd_sc_hd__o22a_1 U30409 ( .A1(n25165), .A2(n26431), .B1(n26790), .B2(
        n26412), .X(n25173) );
  sky130_fd_sc_hd__o22ai_1 U30410 ( .A1(n18916), .A2(n25166), .B1(n26423), 
        .B2(n27399), .Y(n25167) );
  sky130_fd_sc_hd__a21oi_1 U30411 ( .A1(n26085), .A2(n26061), .B1(n25167), .Y(
        n25168) );
  sky130_fd_sc_hd__o21ai_0 U30412 ( .A1(n26432), .A2(n26646), .B1(n25168), .Y(
        n25171) );
  sky130_fd_sc_hd__nor2_1 U30413 ( .A(n26701), .B(n26424), .Y(n25170) );
  sky130_fd_sc_hd__o22ai_1 U30414 ( .A1(n26703), .A2(n26427), .B1(n25798), 
        .B2(n26425), .Y(n25169) );
  sky130_fd_sc_hd__nor3_1 U30415 ( .A(n25171), .B(n25170), .C(n25169), .Y(
        n25172) );
  sky130_fd_sc_hd__nand4_1 U30416 ( .A(n25174), .B(n25173), .C(n26411), .D(
        n25172), .Y(n25175) );
  sky130_fd_sc_hd__a21oi_1 U30417 ( .A1(n25176), .A2(n26409), .B1(n25175), .Y(
        n25177) );
  sky130_fd_sc_hd__a21oi_1 U30419 ( .A1(n26064), .A2(n25180), .B1(n25179), .Y(
        n25184) );
  sky130_fd_sc_hd__nand2b_1 U30420 ( .A_N(n25182), .B(n25181), .Y(n25183) );
  sky130_fd_sc_hd__o211ai_1 U30421 ( .A1(n26352), .A2(n25185), .B1(n25184), 
        .C1(n25183), .Y(n26073) );
  sky130_fd_sc_hd__buf_6 U30422 ( .A(n25186), .X(n26066) );
  sky130_fd_sc_hd__o22ai_1 U30423 ( .A1(n27333), .A2(n27401), .B1(n23178), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N3074) );
  sky130_fd_sc_hd__o22ai_1 U30424 ( .A1(n27213), .A2(n27401), .B1(n27212), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N2815) );
  sky130_fd_sc_hd__o22ai_1 U30425 ( .A1(n27225), .A2(n27401), .B1(n27224), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N2963) );
  sky130_fd_sc_hd__o22ai_1 U30426 ( .A1(n26378), .A2(n27401), .B1(n26449), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N3259) );
  sky130_fd_sc_hd__o22ai_1 U30427 ( .A1(n11141), .A2(n27401), .B1(n27124), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N2704) );
  sky130_fd_sc_hd__o22ai_1 U30428 ( .A1(n27226), .A2(n27401), .B1(n23079), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N3148) );
  sky130_fd_sc_hd__o22ai_1 U30429 ( .A1(n27219), .A2(n27401), .B1(n27218), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N3000) );
  sky130_fd_sc_hd__nor2_1 U30430 ( .A(n26946), .B(n26066), .Y(
        j202_soc_core_j22_cpu_rf_N2667) );
  sky130_fd_sc_hd__o22ai_1 U30431 ( .A1(n27466), .A2(n27401), .B1(n27465), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N2778) );
  sky130_fd_sc_hd__o22ai_1 U30432 ( .A1(n27209), .A2(n27401), .B1(n23039), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N2741) );
  sky130_fd_sc_hd__o22ai_1 U30433 ( .A1(n27221), .A2(n27401), .B1(n27220), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N2889) );
  sky130_fd_sc_hd__o22ai_1 U30434 ( .A1(n27211), .A2(n27401), .B1(n27210), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N3222) );
  sky130_fd_sc_hd__o22ai_1 U30435 ( .A1(n27215), .A2(n27401), .B1(n27214), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N2926) );
  sky130_fd_sc_hd__o22ai_1 U30436 ( .A1(n27223), .A2(n27401), .B1(n27222), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N3037) );
  sky130_fd_sc_hd__o22ai_1 U30437 ( .A1(n27217), .A2(n27401), .B1(n27216), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N2852) );
  sky130_fd_sc_hd__o22ai_1 U30438 ( .A1(n27228), .A2(n27401), .B1(n27227), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N3185) );
  sky130_fd_sc_hd__nand2_1 U30439 ( .A(n25116), .B(n27460), .Y(n25187) );
  sky130_fd_sc_hd__o21ai_1 U30440 ( .A1(n27460), .A2(n25222), .B1(n25187), .Y(
        j202_soc_core_j22_cpu_rf_N3298) );
  sky130_fd_sc_hd__nor2_1 U30441 ( .A(n26946), .B(n25222), .Y(
        j202_soc_core_j22_cpu_rf_N2670) );
  sky130_fd_sc_hd__a21oi_1 U30442 ( .A1(n25191), .A2(n26516), .B1(n25190), .Y(
        n25192) );
  sky130_fd_sc_hd__o21ai_1 U30443 ( .A1(n25194), .A2(n25193), .B1(n25192), .Y(
        j202_soc_core_j22_cpu_rf_N3373) );
  sky130_fd_sc_hd__o22ai_1 U30444 ( .A1(n25203), .A2(n27021), .B1(n25195), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U30445 ( .A1(n25203), .A2(n25534), .B1(n25196), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U30446 ( .A1(n25203), .A2(n27990), .B1(n25197), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U30447 ( .A1(n25203), .A2(n28535), .B1(n25198), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U30448 ( .A1(n25203), .A2(n28547), .B1(n25199), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U30449 ( .A1(n25203), .A2(n28538), .B1(n25205), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U30450 ( .A1(n25203), .A2(n28541), .B1(n25200), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U30451 ( .A1(n28544), .A2(n25203), .B1(n25201), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U30452 ( .A1(n25203), .A2(n27194), .B1(n25202), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__a21oi_1 U30453 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[25]), .B1(n27758), .Y(n25204) );
  sky130_fd_sc_hd__a21oi_1 U30455 ( .A1(j202_soc_core_intc_core_00_rg_ipr[57]), 
        .A2(n27862), .B1(n25206), .Y(n25211) );
  sky130_fd_sc_hd__a22o_1 U30456 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[25]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[89]), .X(n25207) );
  sky130_fd_sc_hd__a21oi_1 U30457 ( .A1(n27850), .A2(
        j202_soc_core_intc_core_00_rg_itgt[38]), .B1(n25207), .Y(n25210) );
  sky130_fd_sc_hd__a22oi_1 U30458 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[62]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[121]), .Y(n25209) );
  sky130_fd_sc_hd__nand2_1 U30459 ( .A(n27869), .B(
        j202_soc_core_intc_core_00_rg_itgt[46]), .Y(n25208) );
  sky130_fd_sc_hd__nand4_1 U30460 ( .A(n25211), .B(n25210), .C(n25209), .D(
        n25208), .Y(j202_soc_core_ahb2apb_01_N153) );
  sky130_fd_sc_hd__nand2_1 U30461 ( .A(n27108), .B(j202_soc_core_uart_div0[1]), 
        .Y(n25212) );
  sky130_fd_sc_hd__o21ai_1 U30462 ( .A1(n25213), .A2(n27108), .B1(n25212), .Y(
        n135) );
  sky130_fd_sc_hd__nand2_1 U30463 ( .A(n25116), .B(n27339), .Y(n25214) );
  sky130_fd_sc_hd__o211ai_1 U30464 ( .A1(n26706), .A2(n25215), .B1(n25214), 
        .C1(n27346), .Y(j202_soc_core_j22_cpu_ml_N329) );
  sky130_fd_sc_hd__o211ai_1 U30465 ( .A1(n25219), .A2(n25218), .B1(n25217), 
        .C1(n25216), .Y(n25220) );
  sky130_fd_sc_hd__a22oi_1 U30466 ( .A1(n27187), .A2(n18656), .B1(n27273), 
        .B2(n25220), .Y(n25221) );
  sky130_fd_sc_hd__nand2_1 U30467 ( .A(n27189), .B(n25221), .Y(
        j202_soc_core_j22_cpu_ml_machj[25]) );
  sky130_fd_sc_hd__o22ai_1 U30468 ( .A1(n27575), .A2(n11102), .B1(n27574), 
        .B2(n25115), .Y(j202_soc_core_j22_cpu_rf_N3114) );
  sky130_fd_sc_hd__nand3_1 U30469 ( .A(n25226), .B(n25225), .C(n25224), .Y(
        n25228) );
  sky130_fd_sc_hd__nor2_1 U30470 ( .A(n25228), .B(n25227), .Y(n29323) );
  sky130_fd_sc_hd__mux2i_1 U30471 ( .A0(n12451), .A1(n25229), .S(n27006), .Y(
        j202_soc_core_j22_cpu_ml_N305) );
  sky130_fd_sc_hd__a21oi_1 U30472 ( .A1(n25233), .A2(n26802), .B1(n25232), .Y(
        n25234) );
  sky130_fd_sc_hd__buf_4 U30473 ( .A(n25234), .X(n26858) );
  sky130_fd_sc_hd__nor2_1 U30474 ( .A(n26946), .B(n26858), .Y(
        j202_soc_core_j22_cpu_rf_N2644) );
  sky130_fd_sc_hd__o22ai_1 U30475 ( .A1(n12451), .A2(n26378), .B1(n26449), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N3235) );
  sky130_fd_sc_hd__o22ai_1 U30476 ( .A1(n25237), .A2(n26892), .B1(n26891), 
        .B2(n25236), .Y(n25238) );
  sky130_fd_sc_hd__a21oi_1 U30477 ( .A1(n25244), .A2(n26895), .B1(n25238), .Y(
        n25239) );
  sky130_fd_sc_hd__nand2_1 U30478 ( .A(n25240), .B(n25239), .Y(
        j202_soc_core_j22_cpu_rf_N300) );
  sky130_fd_sc_hd__o22ai_1 U30479 ( .A1(n12451), .A2(n26899), .B1(n26898), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N3311) );
  sky130_fd_sc_hd__o22ai_1 U30480 ( .A1(n12451), .A2(n27575), .B1(n27574), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N3087) );
  sky130_fd_sc_hd__o22ai_1 U30481 ( .A1(n12451), .A2(n27333), .B1(n23178), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N3050) );
  sky130_fd_sc_hd__o22ai_1 U30482 ( .A1(n12451), .A2(n27219), .B1(n27218), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N2976) );
  sky130_fd_sc_hd__o22ai_1 U30483 ( .A1(n12451), .A2(n27217), .B1(n27216), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N2828) );
  sky130_fd_sc_hd__o22ai_1 U30484 ( .A1(n12451), .A2(n27228), .B1(n27227), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N3161) );
  sky130_fd_sc_hd__o22ai_1 U30485 ( .A1(n12451), .A2(n27225), .B1(n27224), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N2939) );
  sky130_fd_sc_hd__o22ai_1 U30486 ( .A1(n12451), .A2(n27466), .B1(n27465), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N2754) );
  sky130_fd_sc_hd__o22ai_1 U30487 ( .A1(n12451), .A2(n27215), .B1(n27214), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N2902) );
  sky130_fd_sc_hd__o22ai_1 U30488 ( .A1(n12451), .A2(n27223), .B1(n27222), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N3013) );
  sky130_fd_sc_hd__o22ai_1 U30489 ( .A1(n12451), .A2(n27211), .B1(n27210), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N3198) );
  sky130_fd_sc_hd__o22ai_1 U30490 ( .A1(n12451), .A2(n27221), .B1(n27220), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N2865) );
  sky130_fd_sc_hd__o22ai_1 U30491 ( .A1(n12451), .A2(n27226), .B1(n23079), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N3124) );
  sky130_fd_sc_hd__o22ai_1 U30492 ( .A1(n12451), .A2(n27213), .B1(n27212), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N2791) );
  sky130_fd_sc_hd__o22ai_1 U30493 ( .A1(n12451), .A2(n27209), .B1(n23039), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N2717) );
  sky130_fd_sc_hd__o22ai_1 U30494 ( .A1(n12451), .A2(n11141), .B1(n27124), 
        .B2(n26858), .Y(j202_soc_core_j22_cpu_rf_N2680) );
  sky130_fd_sc_hd__nor2_1 U30495 ( .A(n26951), .B(n25241), .Y(n25242) );
  sky130_fd_sc_hd__nand2_1 U30496 ( .A(n25243), .B(n25242), .Y(n25246) );
  sky130_fd_sc_hd__nand2_1 U30497 ( .A(n25246), .B(n25245), .Y(
        j202_soc_core_j22_cpu_rf_N3347) );
  sky130_fd_sc_hd__nand4_1 U30498 ( .A(n25250), .B(n25251), .C(n25249), .D(
        n25248), .Y(n25252) );
  sky130_fd_sc_hd__nand2_1 U30499 ( .A(n27273), .B(n25252), .Y(n25253) );
  sky130_fd_sc_hd__nand2_1 U30500 ( .A(n27189), .B(n25253), .Y(
        j202_soc_core_j22_cpu_ml_machj[18]) );
  sky130_fd_sc_hd__nand2_1 U30501 ( .A(n27593), .B(j202_soc_core_uart_div1[2]), 
        .Y(n25255) );
  sky130_fd_sc_hd__o21ai_1 U30502 ( .A1(n25256), .A2(n27593), .B1(n25255), .Y(
        n108) );
  sky130_fd_sc_hd__nor2_1 U30503 ( .A(n28590), .B(n28180), .Y(
        j202_soc_core_wbqspiflash_00_N715) );
  sky130_fd_sc_hd__o21ai_1 U30504 ( .A1(n27040), .A2(n27039), .B1(n26130), .Y(
        n27718) );
  sky130_fd_sc_hd__a22o_1 U30505 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[18]), .A2(n27719), .B1(n27718), 
        .B2(j202_soc_core_wbqspiflash_00_erased_sector[4]), .X(
        j202_soc_core_wbqspiflash_00_N685) );
  sky130_fd_sc_hd__nand2_1 U30506 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[18]), .Y(n25257) );
  sky130_fd_sc_hd__o21ai_1 U30507 ( .A1(n25258), .A2(n27983), .B1(n25257), .Y(
        n65) );
  sky130_fd_sc_hd__nand2_1 U30508 ( .A(n25259), .B(n27460), .Y(n25260) );
  sky130_fd_sc_hd__o22ai_1 U30510 ( .A1(n27333), .A2(n27434), .B1(n23178), 
        .B2(n12433), .Y(j202_soc_core_j22_cpu_rf_N3068) );
  sky130_fd_sc_hd__a22oi_1 U30511 ( .A1(n26948), .A2(n25261), .B1(n11764), 
        .B2(n24650), .Y(n25263) );
  sky130_fd_sc_hd__nand2_1 U30512 ( .A(n27048), .B(n26067), .Y(n25262) );
  sky130_fd_sc_hd__o211ai_1 U30513 ( .A1(n12124), .A2(n26951), .B1(n25263), 
        .C1(n25262), .Y(j202_soc_core_j22_cpu_rf_N3363) );
  sky130_fd_sc_hd__mux2i_1 U30514 ( .A0(n25276), .A1(n26567), .S(n27006), .Y(
        j202_soc_core_j22_cpu_ml_N318) );
  sky130_fd_sc_hd__o21ai_1 U30515 ( .A1(n25824), .A2(n25264), .B1(n25822), .Y(
        n25265) );
  sky130_fd_sc_hd__a31oi_1 U30516 ( .A1(n26871), .A2(n26872), .A3(n12357), 
        .B1(n25265), .Y(n25267) );
  sky130_fd_sc_hd__nand2_1 U30517 ( .A(n25267), .B(n25266), .Y(
        j202_soc_core_j22_cpu_ml_maclj[15]) );
  sky130_fd_sc_hd__o21ai_1 U30518 ( .A1(n25270), .A2(n25829), .B1(n27189), .Y(
        j202_soc_core_j22_cpu_ml_machj[15]) );
  sky130_fd_sc_hd__nand2_1 U30519 ( .A(n26948), .B(n25268), .Y(n25275) );
  sky130_fd_sc_hd__nand2_1 U30520 ( .A(n11131), .B(n29535), .Y(n25272) );
  sky130_fd_sc_hd__nand2_1 U30521 ( .A(n25270), .B(n12422), .Y(n25271) );
  sky130_fd_sc_hd__o211ai_1 U30522 ( .A1(n25273), .A2(n25272), .B1(n26516), 
        .C1(n25271), .Y(n25274) );
  sky130_fd_sc_hd__o211ai_1 U30523 ( .A1(n25714), .A2(n25276), .B1(n25275), 
        .C1(n25274), .Y(j202_soc_core_j22_cpu_rf_N3361) );
  sky130_fd_sc_hd__o22ai_1 U30524 ( .A1(n28607), .A2(n25534), .B1(n25277), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U30525 ( .A1(n28596), .A2(n25534), .B1(n25278), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U30526 ( .A1(n28614), .A2(n27194), .B1(n25283), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__nor3_1 U30527 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]), .B(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[3]), .C(n25495), .Y(n25747) );
  sky130_fd_sc_hd__nand3b_1 U30528 ( .A_N(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[4]), .B(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[6]), .C(j202_soc_core_intc_core_00_cp_intack_all_0_), .Y(n25352) );
  sky130_fd_sc_hd__nor2_1 U30529 ( .A(n28512), .B(n25352), .Y(n27196) );
  sky130_fd_sc_hd__a21oi_1 U30530 ( .A1(n25747), .A2(n27196), .B1(
        j202_soc_core_intc_core_00_rg_irqc[3]), .Y(n25281) );
  sky130_fd_sc_hd__nor2_1 U30531 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[3]), 
        .B(n25279), .Y(n25280) );
  sky130_fd_sc_hd__a31oi_1 U30532 ( .A1(n25281), .A2(
        j202_soc_core_intc_core_00_in_intreq[3]), .A3(n29594), .B1(n25280), 
        .Y(n25282) );
  sky130_fd_sc_hd__nor2_1 U30533 ( .A(n25283), .B(n25282), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N6) );
  sky130_fd_sc_hd__nor2_1 U30534 ( .A(n28590), .B(
        j202_soc_core_qspi_wb_wdat[12]), .Y(n28355) );
  sky130_fd_sc_hd__o22ai_1 U30535 ( .A1(n27154), .A2(n25284), .B1(n28355), 
        .B2(n27152), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__nand2_1 U30536 ( .A(n27459), .B(n26383), .Y(n25285) );
  sky130_fd_sc_hd__o21ai_0 U30537 ( .A1(n27461), .A2(n26899), .B1(n25285), .Y(
        j202_soc_core_j22_cpu_rf_N3324) );
  sky130_fd_sc_hd__mux2i_1 U30538 ( .A0(n27461), .A1(n26708), .S(n27006), .Y(
        j202_soc_core_j22_cpu_ml_N316) );
  sky130_fd_sc_hd__o21ai_0 U30539 ( .A1(n25824), .A2(n17585), .B1(n25822), .Y(
        n25286) );
  sky130_fd_sc_hd__nand3_1 U30540 ( .A(n25875), .B(n26978), .C(n26872), .Y(
        n25287) );
  sky130_fd_sc_hd__nand2_1 U30541 ( .A(n25288), .B(n25287), .Y(
        j202_soc_core_j22_cpu_ml_maclj[13]) );
  sky130_fd_sc_hd__nor2_1 U30542 ( .A(n25290), .B(n25289), .Y(n25295) );
  sky130_fd_sc_hd__o21ai_0 U30543 ( .A1(n25295), .A2(n27274), .B1(n27273), .Y(
        j202_soc_core_j22_cpu_ml_machj[13]) );
  sky130_fd_sc_hd__a22oi_1 U30544 ( .A1(n25291), .A2(n26948), .B1(n11611), 
        .B2(n24650), .Y(n25292) );
  sky130_fd_sc_hd__o21ai_1 U30545 ( .A1(n25335), .A2(n25295), .B1(n25294), .Y(
        j202_soc_core_j22_cpu_rf_N3359) );
  sky130_fd_sc_hd__o22ai_1 U30546 ( .A1(n28598), .A2(n25534), .B1(n25296), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__a21oi_1 U30547 ( .A1(n27361), .A2(n25415), .B1(n26085), .Y(
        n25297) );
  sky130_fd_sc_hd__nand2_1 U30548 ( .A(n25298), .B(n25297), .Y(n25299) );
  sky130_fd_sc_hd__nand2_1 U30549 ( .A(n25299), .B(n26725), .Y(n25322) );
  sky130_fd_sc_hd__o22ai_1 U30550 ( .A1(n26581), .A2(n26418), .B1(n26426), 
        .B2(n26419), .Y(n25306) );
  sky130_fd_sc_hd__nor2_1 U30551 ( .A(n26564), .B(n26349), .Y(n25305) );
  sky130_fd_sc_hd__xnor2_1 U30552 ( .A(n27361), .B(n26725), .Y(n26670) );
  sky130_fd_sc_hd__o21ai_0 U30554 ( .A1(n26670), .A2(n26415), .B1(n25303), .Y(
        n25304) );
  sky130_fd_sc_hd__nor3_1 U30555 ( .A(n25306), .B(n25305), .C(n25304), .Y(
        n25314) );
  sky130_fd_sc_hd__o22ai_1 U30556 ( .A1(n11145), .A2(n26416), .B1(n26567), 
        .B2(n26424), .Y(n25307) );
  sky130_fd_sc_hd__a21oi_1 U30557 ( .A1(n26341), .A2(n26716), .B1(n25307), .Y(
        n25313) );
  sky130_fd_sc_hd__a22oi_1 U30558 ( .A1(n25308), .A2(n26564), .B1(n26077), 
        .B2(n26508), .Y(n25310) );
  sky130_fd_sc_hd__nand2_1 U30559 ( .A(n26338), .B(n27409), .Y(n25309) );
  sky130_fd_sc_hd__o211ai_1 U30560 ( .A1(n26708), .A2(n26427), .B1(n25310), 
        .C1(n25309), .Y(n25311) );
  sky130_fd_sc_hd__a21oi_1 U30561 ( .A1(n26342), .A2(n27357), .B1(n25311), .Y(
        n25312) );
  sky130_fd_sc_hd__nand4_1 U30562 ( .A(n25314), .B(n25313), .C(n25312), .D(
        n26344), .Y(n25315) );
  sky130_fd_sc_hd__a21oi_1 U30563 ( .A1(n25316), .A2(n26409), .B1(n25315), .Y(
        n25317) );
  sky130_fd_sc_hd__o21a_1 U30564 ( .A1(n18916), .A2(n25318), .B1(n25317), .X(
        n25321) );
  sky130_fd_sc_hd__nand2_1 U30566 ( .A(n27360), .B(n25319), .Y(n25320) );
  sky130_fd_sc_hd__and3_1 U30567 ( .A(n25325), .B(n25324), .C(n25323), .X(
        n25334) );
  sky130_fd_sc_hd__o22ai_1 U30568 ( .A1(n27575), .A2(n27125), .B1(n27574), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N3101) );
  sky130_fd_sc_hd__o22ai_1 U30569 ( .A1(n27333), .A2(n27125), .B1(n23178), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N3064) );
  sky130_fd_sc_hd__o22ai_1 U30570 ( .A1(n27219), .A2(n27125), .B1(n27218), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N2990) );
  sky130_fd_sc_hd__o22ai_1 U30571 ( .A1(n27217), .A2(n27125), .B1(n27216), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N2842) );
  sky130_fd_sc_hd__o22ai_1 U30572 ( .A1(n27228), .A2(n27125), .B1(n27227), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N3175) );
  sky130_fd_sc_hd__o22ai_1 U30573 ( .A1(n27225), .A2(n27125), .B1(n27224), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N2953) );
  sky130_fd_sc_hd__o22ai_1 U30574 ( .A1(n27466), .A2(n27125), .B1(n27465), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N2768) );
  sky130_fd_sc_hd__o22ai_1 U30575 ( .A1(n27215), .A2(n27125), .B1(n27214), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N2916) );
  sky130_fd_sc_hd__o22ai_1 U30576 ( .A1(n27223), .A2(n27125), .B1(n27222), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N3027) );
  sky130_fd_sc_hd__o22ai_1 U30577 ( .A1(n27211), .A2(n27125), .B1(n27210), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N3212) );
  sky130_fd_sc_hd__o22ai_1 U30578 ( .A1(n27221), .A2(n27125), .B1(n27220), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N2879) );
  sky130_fd_sc_hd__o22ai_1 U30579 ( .A1(n27226), .A2(n27125), .B1(n23079), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N3138) );
  sky130_fd_sc_hd__o22ai_1 U30580 ( .A1(n27213), .A2(n27125), .B1(n27212), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N2805) );
  sky130_fd_sc_hd__o22ai_1 U30581 ( .A1(n26378), .A2(n27125), .B1(n26449), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N3249) );
  sky130_fd_sc_hd__o22ai_1 U30582 ( .A1(n27209), .A2(n27125), .B1(n23039), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N2731) );
  sky130_fd_sc_hd__nor2_1 U30583 ( .A(n26946), .B(n27127), .Y(
        j202_soc_core_j22_cpu_rf_N2657) );
  sky130_fd_sc_hd__o22ai_1 U30584 ( .A1(n27125), .A2(n26899), .B1(n26898), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N3325) );
  sky130_fd_sc_hd__nand2_1 U30585 ( .A(n27360), .B(n27343), .Y(n25327) );
  sky130_fd_sc_hd__o21ai_0 U30586 ( .A1(n26565), .A2(n27343), .B1(n25327), .Y(
        j202_soc_core_j22_cpu_ml_N317) );
  sky130_fd_sc_hd__a21oi_1 U30587 ( .A1(j202_soc_core_j22_cpu_ml_bufa[14]), 
        .A2(n27187), .B1(n25829), .Y(n25328) );
  sky130_fd_sc_hd__o21ai_1 U30588 ( .A1(n27274), .A2(n25334), .B1(n25328), .Y(
        j202_soc_core_j22_cpu_ml_machj[14]) );
  sky130_fd_sc_hd__o22ai_1 U30589 ( .A1(n26070), .A2(n25330), .B1(n25714), 
        .B2(n27125), .Y(n25331) );
  sky130_fd_sc_hd__a21oi_1 U30590 ( .A1(n26516), .A2(n25332), .B1(n25331), .Y(
        n25333) );
  sky130_fd_sc_hd__o21ai_1 U30591 ( .A1(n25335), .A2(n25334), .B1(n25333), .Y(
        j202_soc_core_j22_cpu_rf_N3360) );
  sky130_fd_sc_hd__mux2i_1 U30592 ( .A0(n26556), .A1(n11145), .S(n27006), .Y(
        j202_soc_core_j22_cpu_ml_N309) );
  sky130_fd_sc_hd__nor2_1 U30593 ( .A(n26946), .B(n13320), .Y(
        j202_soc_core_j22_cpu_rf_N2648) );
  sky130_fd_sc_hd__mux2i_1 U30594 ( .A0(n13320), .A1(n26556), .S(n27460), .Y(
        j202_soc_core_j22_cpu_rf_N3276) );
  sky130_fd_sc_hd__nand2_1 U30595 ( .A(n25811), .B(n29075), .Y(n25340) );
  sky130_fd_sc_hd__nand2_1 U30596 ( .A(n25341), .B(n25340), .Y(n25342) );
  sky130_fd_sc_hd__a21oi_1 U30597 ( .A1(n27882), .A2(n12617), .B1(n25342), .Y(
        n25343) );
  sky130_fd_sc_hd__o21ai_1 U30598 ( .A1(n25343), .A2(n27928), .B1(n27300), .Y(
        n10497) );
  sky130_fd_sc_hd__o22ai_1 U30599 ( .A1(n26556), .A2(n26899), .B1(n26898), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N3316) );
  sky130_fd_sc_hd__a21oi_1 U30600 ( .A1(n25344), .A2(
        j202_soc_core_j22_cpu_ml_bufa[6]), .B1(n26976), .Y(n25348) );
  sky130_fd_sc_hd__nand3_1 U30601 ( .A(n12916), .B(
        j202_soc_core_j22_cpu_ml_macl[6]), .C(n25826), .Y(n25347) );
  sky130_fd_sc_hd__nand3_1 U30602 ( .A(n12357), .B(n25345), .C(n26872), .Y(
        n25346) );
  sky130_fd_sc_hd__nand3_1 U30603 ( .A(n25348), .B(n25347), .C(n25346), .Y(
        j202_soc_core_j22_cpu_ml_maclj[6]) );
  sky130_fd_sc_hd__o22ai_1 U30604 ( .A1(n28609), .A2(n25534), .B1(n25349), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o22a_1 U30605 ( .A1(j202_soc_core_intc_core_00_rg_ie[0]), 
        .A2(n25351), .B1(n29086), .B2(n25350), .X(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__nor2_1 U30606 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[1]), .B(n25352), .Y(n25746) );
  sky130_fd_sc_hd__nor3_1 U30607 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .B(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]), .C(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[3]), .Y(n27195) );
  sky130_fd_sc_hd__a21oi_1 U30608 ( .A1(n25746), .A2(n27195), .B1(
        j202_soc_core_intc_core_00_rg_irqc[0]), .Y(n25355) );
  sky130_fd_sc_hd__nor2_1 U30609 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[0]), 
        .B(n25353), .Y(n25354) );
  sky130_fd_sc_hd__a31oi_1 U30610 ( .A1(n25355), .A2(
        j202_soc_core_intc_core_00_in_intreq[0]), .A3(n29594), .B1(n25354), 
        .Y(n25356) );
  sky130_fd_sc_hd__nor2_1 U30611 ( .A(n25357), .B(n25356), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N3) );
  sky130_fd_sc_hd__nor2_1 U30612 ( .A(n28590), .B(
        j202_soc_core_qspi_wb_wdat[0]), .Y(n27755) );
  sky130_fd_sc_hd__o22ai_1 U30613 ( .A1(n27154), .A2(n27761), .B1(n27755), 
        .B2(n27152), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U30614 ( .A1(n28603), .A2(n25534), .B1(n27677), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U30615 ( .A1(n28608), .A2(n25534), .B1(n25358), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U30616 ( .A1(n28599), .A2(n25534), .B1(n25359), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U30617 ( .A1(n26494), .A2(n25534), .B1(n26499), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U30618 ( .A1(n28605), .A2(n25534), .B1(n25360), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U30619 ( .A1(n28612), .A2(n27194), .B1(n25365), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__nor3_1 U30620 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[3]), .B(n28514), .C(n25495), .Y(n25439) );
  sky130_fd_sc_hd__a21oi_1 U30621 ( .A1(n25439), .A2(n25746), .B1(
        j202_soc_core_intc_core_00_rg_irqc[5]), .Y(n25363) );
  sky130_fd_sc_hd__nor2_1 U30622 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[5]), 
        .B(n25361), .Y(n25362) );
  sky130_fd_sc_hd__a31oi_1 U30623 ( .A1(n25363), .A2(
        j202_soc_core_intc_core_00_in_intreq[5]), .A3(n29594), .B1(n25362), 
        .Y(n25364) );
  sky130_fd_sc_hd__nor2_1 U30624 ( .A(n25365), .B(n25364), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N8) );
  sky130_fd_sc_hd__nor2_1 U30625 ( .A(n28590), .B(
        j202_soc_core_qspi_wb_wdat[20]), .Y(n28412) );
  sky130_fd_sc_hd__o22ai_1 U30626 ( .A1(n27154), .A2(n25366), .B1(n28412), 
        .B2(n27152), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U30627 ( .A1(n28613), .A2(n27194), .B1(n25371), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__nor3_1 U30628 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .B(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[3]), .C(n28514), .Y(n26479) );
  sky130_fd_sc_hd__a21oi_1 U30629 ( .A1(n26479), .A2(n25746), .B1(
        j202_soc_core_intc_core_00_rg_irqc[4]), .Y(n25369) );
  sky130_fd_sc_hd__nor2_1 U30630 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[4]), 
        .B(n25367), .Y(n25368) );
  sky130_fd_sc_hd__a31oi_1 U30631 ( .A1(n25369), .A2(
        j202_soc_core_intc_core_00_in_intreq[4]), .A3(n29594), .B1(n25368), 
        .Y(n25370) );
  sky130_fd_sc_hd__nor2_1 U30632 ( .A(n25371), .B(n25370), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N7) );
  sky130_fd_sc_hd__nor2_1 U30633 ( .A(n28590), .B(
        j202_soc_core_qspi_wb_wdat[16]), .Y(n28384) );
  sky130_fd_sc_hd__o22ai_1 U30634 ( .A1(n27154), .A2(n25372), .B1(n28384), 
        .B2(n27152), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__nand2_1 U30635 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[21]), .Y(n25373) );
  sky130_fd_sc_hd__o21ai_1 U30636 ( .A1(n25374), .A2(n27983), .B1(n25373), .Y(
        n67) );
  sky130_fd_sc_hd__o22ai_1 U30637 ( .A1(n25427), .A2(n27021), .B1(n25375), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30638 ( .A1(n25427), .A2(n27990), .B1(n25376), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30639 ( .A1(n25427), .A2(n28535), .B1(n25377), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30640 ( .A1(n25427), .A2(n28547), .B1(n25378), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30641 ( .A1(n25427), .A2(n28538), .B1(n25383), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30642 ( .A1(n25427), .A2(n28541), .B1(n25379), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30643 ( .A1(n28544), .A2(n25427), .B1(n25380), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30644 ( .A1(n25427), .A2(n27194), .B1(n25381), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__a21oi_1 U30645 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[21]), .B1(n27758), .Y(n25382) );
  sky130_fd_sc_hd__o21ai_1 U30646 ( .A1(n25383), .A2(n27097), .B1(n25382), .Y(
        n25384) );
  sky130_fd_sc_hd__a21oi_1 U30647 ( .A1(j202_soc_core_intc_core_00_rg_ipr[53]), 
        .A2(n27862), .B1(n25384), .Y(n25389) );
  sky130_fd_sc_hd__a22o_1 U30648 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[21]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[85]), .X(n25385) );
  sky130_fd_sc_hd__a21oi_1 U30649 ( .A1(n27850), .A2(
        j202_soc_core_intc_core_00_rg_itgt[37]), .B1(n25385), .Y(n25388) );
  sky130_fd_sc_hd__a22oi_1 U30650 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[61]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[117]), .Y(n25387) );
  sky130_fd_sc_hd__nand2_1 U30651 ( .A(n27869), .B(
        j202_soc_core_intc_core_00_rg_itgt[45]), .Y(n25386) );
  sky130_fd_sc_hd__nand4_1 U30652 ( .A(n25389), .B(n25388), .C(n25387), .D(
        n25386), .Y(j202_soc_core_ahb2apb_01_N149) );
  sky130_fd_sc_hd__nand2_1 U30653 ( .A(n27593), .B(j202_soc_core_uart_div1[5]), 
        .Y(n25390) );
  sky130_fd_sc_hd__o21ai_1 U30654 ( .A1(n25391), .A2(n27593), .B1(n25390), .Y(
        n110) );
  sky130_fd_sc_hd__nor2_1 U30655 ( .A(n28590), .B(n25392), .Y(
        j202_soc_core_wbqspiflash_00_N718) );
  sky130_fd_sc_hd__a22o_1 U30656 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[21]), .A2(n27719), .B1(n27718), 
        .B2(j202_soc_core_wbqspiflash_00_erased_sector[7]), .X(
        j202_soc_core_wbqspiflash_00_N688) );
  sky130_fd_sc_hd__nand2_1 U30657 ( .A(n12212), .B(n25396), .Y(n25400) );
  sky130_fd_sc_hd__a31oi_1 U30658 ( .A1(n25398), .A2(n11713), .A3(n25397), 
        .B1(n18916), .Y(n25399) );
  sky130_fd_sc_hd__nand2_1 U30659 ( .A(n25400), .B(n25399), .Y(n25422) );
  sky130_fd_sc_hd__a21oi_1 U30660 ( .A1(n27183), .A2(n26323), .B1(n26406), .Y(
        n25414) );
  sky130_fd_sc_hd__nand2_1 U30661 ( .A(n26077), .B(n26971), .Y(n25402) );
  sky130_fd_sc_hd__xor2_1 U30662 ( .A(n27183), .B(n27412), .X(n26644) );
  sky130_fd_sc_hd__nand2_1 U30663 ( .A(n26644), .B(n26326), .Y(n25401) );
  sky130_fd_sc_hd__o211ai_1 U30664 ( .A1(n27412), .A2(n26423), .B1(n25402), 
        .C1(n25401), .Y(n25405) );
  sky130_fd_sc_hd__o22ai_1 U30665 ( .A1(n26704), .A2(n26418), .B1(n25403), 
        .B2(n26419), .Y(n25404) );
  sky130_fd_sc_hd__nor2_1 U30666 ( .A(n25405), .B(n25404), .Y(n25410) );
  sky130_fd_sc_hd__o22a_1 U30667 ( .A1(n26569), .A2(n26431), .B1(n26893), .B2(
        n26412), .X(n25409) );
  sky130_fd_sc_hd__o22ai_1 U30668 ( .A1(n26417), .A2(n26427), .B1(n26703), 
        .B2(n26424), .Y(n25407) );
  sky130_fd_sc_hd__o22ai_1 U30669 ( .A1(n26708), .A2(n26416), .B1(n26577), 
        .B2(n26425), .Y(n25406) );
  sky130_fd_sc_hd__nor2_1 U30670 ( .A(n25407), .B(n25406), .Y(n25408) );
  sky130_fd_sc_hd__nand4_1 U30671 ( .A(n25410), .B(n25409), .C(n25408), .D(
        n26411), .Y(n25411) );
  sky130_fd_sc_hd__a21oi_1 U30672 ( .A1(n25412), .A2(n26409), .B1(n25411), .Y(
        n25413) );
  sky130_fd_sc_hd__o21a_1 U30673 ( .A1(n25414), .A2(n27414), .B1(n25413), .X(
        n25421) );
  sky130_fd_sc_hd__a21oi_1 U30675 ( .A1(n27412), .A2(n25415), .B1(n26085), .Y(
        n25416) );
  sky130_fd_sc_hd__a2bb2oi_1 U30676 ( .B1(n27182), .B2(n25419), .A1_N(n26570), 
        .A2_N(n25418), .Y(n25420) );
  sky130_fd_sc_hd__nand3_2 U30677 ( .A(n25421), .B(n25422), .C(n25420), .Y(
        n27190) );
  sky130_fd_sc_hd__inv_4 U30678 ( .A(n27190), .Y(n25426) );
  sky130_fd_sc_hd__o22ai_1 U30679 ( .A1(n26378), .A2(n27414), .B1(n26449), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N3257) );
  sky130_fd_sc_hd__o22ai_1 U30680 ( .A1(n27414), .A2(n26899), .B1(n26898), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N3333) );
  sky130_fd_sc_hd__nand2_1 U30681 ( .A(n27190), .B(n26516), .Y(n25425) );
  sky130_fd_sc_hd__a22oi_1 U30682 ( .A1(n25423), .A2(n26948), .B1(n29549), 
        .B2(n24650), .Y(n25424) );
  sky130_fd_sc_hd__nand2_1 U30683 ( .A(n25425), .B(n25424), .Y(
        j202_soc_core_j22_cpu_rf_N3368) );
  sky130_fd_sc_hd__o22ai_1 U30684 ( .A1(n11141), .A2(n27414), .B1(n27124), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N2702) );
  sky130_fd_sc_hd__o22ai_1 U30685 ( .A1(n27575), .A2(n27414), .B1(n27574), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N3109) );
  sky130_fd_sc_hd__o22ai_1 U30686 ( .A1(n27333), .A2(n27414), .B1(n23178), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N3072) );
  sky130_fd_sc_hd__o22ai_1 U30687 ( .A1(n27219), .A2(n27414), .B1(n27218), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N2998) );
  sky130_fd_sc_hd__o22ai_1 U30688 ( .A1(n27217), .A2(n27414), .B1(n27216), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N2850) );
  sky130_fd_sc_hd__o22ai_1 U30689 ( .A1(n27228), .A2(n27414), .B1(n27227), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N3183) );
  sky130_fd_sc_hd__o22ai_1 U30690 ( .A1(n27225), .A2(n27414), .B1(n27224), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N2961) );
  sky130_fd_sc_hd__o22ai_1 U30691 ( .A1(n27466), .A2(n27414), .B1(n27465), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N2776) );
  sky130_fd_sc_hd__o22ai_1 U30692 ( .A1(n27215), .A2(n27414), .B1(n27214), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N2924) );
  sky130_fd_sc_hd__o22ai_1 U30693 ( .A1(n27223), .A2(n27414), .B1(n27222), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N3035) );
  sky130_fd_sc_hd__o22ai_1 U30694 ( .A1(n27211), .A2(n27414), .B1(n27210), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N3220) );
  sky130_fd_sc_hd__o22ai_1 U30695 ( .A1(n27221), .A2(n27414), .B1(n27220), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N2887) );
  sky130_fd_sc_hd__o22ai_1 U30696 ( .A1(n27226), .A2(n27414), .B1(n23079), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N3146) );
  sky130_fd_sc_hd__o22ai_1 U30697 ( .A1(n27213), .A2(n27414), .B1(n27212), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N2813) );
  sky130_fd_sc_hd__o22ai_1 U30698 ( .A1(n27209), .A2(n27414), .B1(n23039), 
        .B2(n25426), .Y(j202_soc_core_j22_cpu_rf_N2739) );
  sky130_fd_sc_hd__o22ai_1 U30699 ( .A1(n25427), .A2(n25534), .B1(n19623), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U30700 ( .A1(n28602), .A2(n25534), .B1(n25428), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U30701 ( .A1(n28606), .A2(n25534), .B1(n25429), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U30702 ( .A1(n28604), .A2(n25534), .B1(n25430), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U30703 ( .A1(n28600), .A2(n25534), .B1(n25431), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U30704 ( .A1(n27028), .A2(n25534), .B1(n25432), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U30705 ( .A1(n27575), .A2(n27359), .B1(n27574), 
        .B2(n26523), .Y(j202_soc_core_j22_cpu_rf_N3119) );
  sky130_fd_sc_hd__o22ai_1 U30706 ( .A1(n27219), .A2(n27359), .B1(n27218), 
        .B2(n26523), .Y(j202_soc_core_j22_cpu_rf_N3008) );
  sky130_fd_sc_hd__o22ai_1 U30707 ( .A1(n27217), .A2(n27359), .B1(n27216), 
        .B2(n26523), .Y(j202_soc_core_j22_cpu_rf_N2860) );
  sky130_fd_sc_hd__o22ai_1 U30708 ( .A1(n27228), .A2(n27359), .B1(n27227), 
        .B2(n26523), .Y(j202_soc_core_j22_cpu_rf_N3193) );
  sky130_fd_sc_hd__o22ai_1 U30709 ( .A1(n27225), .A2(n27359), .B1(n27224), 
        .B2(n26523), .Y(j202_soc_core_j22_cpu_rf_N2971) );
  sky130_fd_sc_hd__o22ai_1 U30710 ( .A1(n27466), .A2(n27359), .B1(n27465), 
        .B2(n26523), .Y(j202_soc_core_j22_cpu_rf_N2786) );
  sky130_fd_sc_hd__o22ai_1 U30711 ( .A1(n27215), .A2(n27359), .B1(n27214), 
        .B2(n26523), .Y(j202_soc_core_j22_cpu_rf_N2934) );
  sky130_fd_sc_hd__o22ai_1 U30712 ( .A1(n27223), .A2(n27359), .B1(n27222), 
        .B2(n26523), .Y(j202_soc_core_j22_cpu_rf_N3045) );
  sky130_fd_sc_hd__o22ai_1 U30713 ( .A1(n27211), .A2(n27359), .B1(n27210), 
        .B2(n26523), .Y(j202_soc_core_j22_cpu_rf_N3230) );
  sky130_fd_sc_hd__o22ai_1 U30714 ( .A1(n27221), .A2(n27359), .B1(n27220), 
        .B2(n26523), .Y(j202_soc_core_j22_cpu_rf_N2897) );
  sky130_fd_sc_hd__o22ai_1 U30715 ( .A1(n27213), .A2(n27359), .B1(n27212), 
        .B2(n26523), .Y(j202_soc_core_j22_cpu_rf_N2823) );
  sky130_fd_sc_hd__o22ai_1 U30716 ( .A1(n27095), .A2(n25534), .B1(n27101), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U30717 ( .A1(n28611), .A2(n27194), .B1(n25437), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__a21oi_1 U30718 ( .A1(n26479), .A2(n27196), .B1(
        j202_soc_core_intc_core_00_rg_irqc[6]), .Y(n25435) );
  sky130_fd_sc_hd__nor2_1 U30719 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[6]), 
        .B(n25433), .Y(n25434) );
  sky130_fd_sc_hd__a31oi_1 U30720 ( .A1(n25435), .A2(
        j202_soc_core_intc_core_00_in_intreq[6]), .A3(n29594), .B1(n25434), 
        .Y(n25436) );
  sky130_fd_sc_hd__nor2_1 U30721 ( .A(n25437), .B(n25436), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N9) );
  sky130_fd_sc_hd__nor2_1 U30722 ( .A(n28590), .B(
        j202_soc_core_qspi_wb_wdat[24]), .Y(n28447) );
  sky130_fd_sc_hd__o22ai_1 U30723 ( .A1(n27154), .A2(n25438), .B1(n28447), 
        .B2(n27152), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U30724 ( .A1(n28610), .A2(n27194), .B1(n25444), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__a21oi_1 U30725 ( .A1(n25439), .A2(n27196), .B1(
        j202_soc_core_intc_core_00_rg_irqc[7]), .Y(n25442) );
  sky130_fd_sc_hd__nor2_1 U30726 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[7]), 
        .B(n25440), .Y(n25441) );
  sky130_fd_sc_hd__a31oi_1 U30727 ( .A1(n25442), .A2(
        j202_soc_core_intc_core_00_in_intreq[7]), .A3(n29594), .B1(n25441), 
        .Y(n25443) );
  sky130_fd_sc_hd__nor2_1 U30728 ( .A(n25444), .B(n25443), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N10) );
  sky130_fd_sc_hd__nor2_1 U30729 ( .A(n28590), .B(
        j202_soc_core_qspi_wb_wdat[28]), .Y(n28477) );
  sky130_fd_sc_hd__o22ai_1 U30730 ( .A1(n27154), .A2(n25445), .B1(n28477), 
        .B2(n27152), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U30731 ( .A1(n26959), .A2(n25534), .B1(n25446), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U30732 ( .A1(n27081), .A2(n25534), .B1(n25447), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U30733 ( .A1(n25649), .A2(n25534), .B1(n25448), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U30734 ( .A1(n28609), .A2(n27021), .B1(n25449), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o22ai_1 U30735 ( .A1(n28597), .A2(n27021), .B1(n25450), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U30736 ( .A1(n28609), .A2(n27194), .B1(n25455), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__nand2_1 U30737 ( .A(n25451), .B(n29594), .Y(n28518) );
  sky130_fd_sc_hd__o22ai_1 U30738 ( .A1(n28518), .A2(n25495), .B1(n25452), 
        .B2(n28515), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N3) );
  sky130_fd_sc_hd__nor2_1 U30739 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]), .B(n28517), .Y(n25466) );
  sky130_fd_sc_hd__nand2_1 U30740 ( .A(n25495), .B(n25466), .Y(n25475) );
  sky130_fd_sc_hd__nor3_1 U30741 ( .A(j202_soc_core_intc_core_00_rg_irqc[10]), 
        .B(n28590), .C(n25453), .Y(n25454) );
  sky130_fd_sc_hd__o21ai_1 U30742 ( .A1(n25475), .A2(n27013), .B1(n25454), .Y(
        n25457) );
  sky130_fd_sc_hd__nand2b_1 U30743 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[10]), 
        .B(n29043), .Y(n25456) );
  sky130_fd_sc_hd__a21oi_1 U30744 ( .A1(n25457), .A2(n25456), .B1(n25455), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N13) );
  sky130_fd_sc_hd__nor2_1 U30745 ( .A(n28590), .B(
        j202_soc_core_qspi_wb_wdat[8]), .Y(n28326) );
  sky130_fd_sc_hd__o22ai_1 U30746 ( .A1(n27010), .A2(n25458), .B1(n28326), 
        .B2(n27008), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U30747 ( .A1(n27021), .A2(n28599), .B1(n25459), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U30748 ( .A1(n28598), .A2(n27021), .B1(n25460), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U30749 ( .A1(n27021), .A2(n28608), .B1(n25461), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U30750 ( .A1(n28607), .A2(n27021), .B1(n25462), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U30751 ( .A1(n28596), .A2(n27021), .B1(n25463), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U30752 ( .A1(n28611), .A2(n27021), .B1(n25464), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U30753 ( .A1(n27010), .A2(n25465), .B1(n28300), 
        .B2(n27008), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U30754 ( .A1(n28601), .A2(n27194), .B1(n25469), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__nand2_1 U30755 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .B(n25466), .Y(n27014) );
  sky130_fd_sc_hd__nor3_1 U30756 ( .A(j202_soc_core_intc_core_00_rg_irqc[9]), 
        .B(n28590), .C(n25467), .Y(n25468) );
  sky130_fd_sc_hd__nand2b_1 U30758 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[9]), 
        .B(n29044), .Y(n25470) );
  sky130_fd_sc_hd__a21oi_1 U30759 ( .A1(n25471), .A2(n25470), .B1(n25469), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N12) );
  sky130_fd_sc_hd__o22ai_1 U30760 ( .A1(n27010), .A2(n25472), .B1(n27755), 
        .B2(n27008), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U30761 ( .A1(n28599), .A2(n27194), .B1(n25476), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__nor3_1 U30762 ( .A(j202_soc_core_intc_core_00_rg_irqc[8]), 
        .B(n28590), .C(n25473), .Y(n25474) );
  sky130_fd_sc_hd__nand2b_1 U30764 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[8]), 
        .B(n29045), .Y(n25477) );
  sky130_fd_sc_hd__a21oi_1 U30765 ( .A1(n25478), .A2(n25477), .B1(n25476), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N11) );
  sky130_fd_sc_hd__o22ai_1 U30766 ( .A1(n28612), .A2(n27021), .B1(n25479), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U30767 ( .A1(n28603), .A2(n27021), .B1(n25480), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22a_1 U30768 ( .A1(j202_soc_core_intc_core_00_rg_ipr[32]), 
        .A2(n25482), .B1(n29086), .B2(n25481), .X(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U30769 ( .A1(n27021), .A2(n28613), .B1(n25483), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U30770 ( .A1(n28614), .A2(n27021), .B1(n25484), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U30771 ( .A1(n28610), .A2(n27021), .B1(n25485), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U30772 ( .A1(n27095), .A2(n27021), .B1(n25486), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U30773 ( .A1(n28607), .A2(n27194), .B1(n25489), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__nor2_1 U30774 ( .A(n28514), .B(n28517), .Y(n25494) );
  sky130_fd_sc_hd__nand2_1 U30775 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .B(n25494), .Y(n25515) );
  sky130_fd_sc_hd__nor3_1 U30776 ( .A(j202_soc_core_intc_core_00_rg_irqc[15]), 
        .B(n28590), .C(n25487), .Y(n25488) );
  sky130_fd_sc_hd__nand2b_1 U30778 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[15]), 
        .B(n29046), .Y(n25490) );
  sky130_fd_sc_hd__a21oi_1 U30779 ( .A1(n25491), .A2(n25490), .B1(n25489), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N18) );
  sky130_fd_sc_hd__o22ai_1 U30780 ( .A1(n27010), .A2(n25492), .B1(n28477), 
        .B2(n27008), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U30781 ( .A1(n27010), .A2(n25493), .B1(n28447), 
        .B2(n27008), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U30782 ( .A1(n28597), .A2(n27194), .B1(n25498), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__nand2_1 U30783 ( .A(n25495), .B(n25494), .Y(n25506) );
  sky130_fd_sc_hd__nor3_1 U30784 ( .A(j202_soc_core_intc_core_00_rg_irqc[14]), 
        .B(n28590), .C(n25496), .Y(n25497) );
  sky130_fd_sc_hd__nand2b_1 U30786 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[14]), 
        .B(n29047), .Y(n25499) );
  sky130_fd_sc_hd__a21oi_1 U30787 ( .A1(n25500), .A2(n25499), .B1(n25498), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N17) );
  sky130_fd_sc_hd__o22ai_1 U30788 ( .A1(n27081), .A2(n27021), .B1(n25501), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U30789 ( .A1(n28605), .A2(n27021), .B1(n25502), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U30790 ( .A1(n26494), .A2(n27021), .B1(n25503), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U30791 ( .A1(n28608), .A2(n27194), .B1(n25507), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__nor3_1 U30792 ( .A(j202_soc_core_intc_core_00_rg_irqc[12]), 
        .B(n28590), .C(n25504), .Y(n25505) );
  sky130_fd_sc_hd__nand2b_1 U30794 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[12]), 
        .B(n29048), .Y(n25508) );
  sky130_fd_sc_hd__a21oi_1 U30795 ( .A1(n25509), .A2(n25508), .B1(n25507), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N15) );
  sky130_fd_sc_hd__o22ai_1 U30796 ( .A1(n27010), .A2(n25510), .B1(n28384), 
        .B2(n27008), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U30797 ( .A1(n27010), .A2(n25511), .B1(n28412), 
        .B2(n27008), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U30798 ( .A1(n28598), .A2(n27194), .B1(n25516), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__nor3_1 U30799 ( .A(j202_soc_core_intc_core_00_rg_irqc[13]), 
        .B(n28590), .C(n25512), .Y(n25513) );
  sky130_fd_sc_hd__nand2b_1 U30801 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[13]), 
        .B(n29049), .Y(n25517) );
  sky130_fd_sc_hd__a21oi_1 U30802 ( .A1(n25518), .A2(n25517), .B1(n25516), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N16) );
  sky130_fd_sc_hd__o22ai_1 U30803 ( .A1(n27021), .A2(n28606), .B1(n25519), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U30804 ( .A1(n27021), .A2(n28604), .B1(n25520), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U30805 ( .A1(n28611), .A2(n27990), .B1(n25521), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U30806 ( .A1(n28605), .A2(n27990), .B1(n25522), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U30807 ( .A1(n25524), .A2(n26904), .B1(n25523), 
        .B2(n26902), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N5) );
  sky130_fd_sc_hd__nand2_1 U30808 ( .A(n26814), .B(n28510), .Y(
        j202_soc_core_j22_cpu_rf_N3391) );
  sky130_fd_sc_hd__a22oi_1 U30809 ( .A1(n25529), .A2(n26948), .B1(n12493), 
        .B2(n24650), .Y(n25525) );
  sky130_fd_sc_hd__o21ai_1 U30810 ( .A1(n26951), .A2(n13320), .B1(n25525), .Y(
        j202_soc_core_j22_cpu_rf_N3351) );
  sky130_fd_sc_hd__o22ai_1 U30811 ( .A1(n26556), .A2(n27575), .B1(n27574), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N3091) );
  sky130_fd_sc_hd__o22ai_1 U30812 ( .A1(n26556), .A2(n27219), .B1(n27218), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N2980) );
  sky130_fd_sc_hd__o22ai_1 U30813 ( .A1(n26556), .A2(n27217), .B1(n27216), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N2832) );
  sky130_fd_sc_hd__o22ai_1 U30814 ( .A1(n26556), .A2(n27466), .B1(n27465), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N2758) );
  sky130_fd_sc_hd__o22ai_1 U30815 ( .A1(n26556), .A2(n27223), .B1(n27222), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N3017) );
  sky130_fd_sc_hd__o22ai_1 U30816 ( .A1(n26556), .A2(n27221), .B1(n27220), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N2869) );
  sky130_fd_sc_hd__o22ai_1 U30817 ( .A1(n26556), .A2(n27213), .B1(n27212), 
        .B2(n13320), .Y(j202_soc_core_j22_cpu_rf_N2795) );
  sky130_fd_sc_hd__nand2_1 U30818 ( .A(n12493), .B(n11157), .Y(n25531) );
  sky130_fd_sc_hd__o22ai_1 U30819 ( .A1(n11977), .A2(n26892), .B1(n26891), 
        .B2(n25527), .Y(n25528) );
  sky130_fd_sc_hd__a21oi_1 U30820 ( .A1(n25529), .A2(n26895), .B1(n25528), .Y(
        n25530) );
  sky130_fd_sc_hd__nand2_1 U30821 ( .A(n25531), .B(n25530), .Y(
        j202_soc_core_j22_cpu_rf_N304) );
  sky130_fd_sc_hd__o22ai_1 U30822 ( .A1(n28597), .A2(n25534), .B1(n25533), 
        .B2(n25532), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U30823 ( .A1(n28610), .A2(n27990), .B1(n27313), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U30824 ( .A1(n28596), .A2(n27990), .B1(n25535), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U30825 ( .A1(n28600), .A2(n27990), .B1(n25536), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U30826 ( .A1(n25538), .A2(n26904), .B1(n25537), 
        .B2(n26902), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N6) );
  sky130_fd_sc_hd__nand2_1 U30827 ( .A(n25756), .B(n26329), .Y(n25546) );
  sky130_fd_sc_hd__nand2_1 U30828 ( .A(n12455), .B(n26908), .Y(n25541) );
  sky130_fd_sc_hd__a21oi_1 U30829 ( .A1(j202_soc_core_intr_level__3_), .A2(
        n26907), .B1(n26906), .Y(n25540) );
  sky130_fd_sc_hd__nand2_1 U30830 ( .A(n25541), .B(n25540), .Y(n25542) );
  sky130_fd_sc_hd__a21oi_1 U30831 ( .A1(n24737), .A2(n25756), .B1(n25542), .Y(
        n25544) );
  sky130_fd_sc_hd__o21ai_1 U30832 ( .A1(n25546), .A2(n25545), .B1(n25544), .Y(
        j202_soc_core_j22_cpu_rf_N3392) );
  sky130_fd_sc_hd__nand2_1 U30833 ( .A(n26739), .B(n26755), .Y(n25554) );
  sky130_fd_sc_hd__a21oi_1 U30834 ( .A1(n26805), .A2(n25554), .B1(n14849), .Y(
        n25553) );
  sky130_fd_sc_hd__nor2_1 U30835 ( .A(n26727), .B(n25554), .Y(n26742) );
  sky130_fd_sc_hd__nand3_1 U30836 ( .A(n26812), .B(n26742), .C(n27347), .Y(
        n25552) );
  sky130_fd_sc_hd__nand2_1 U30837 ( .A(n25547), .B(n25557), .Y(n25550) );
  sky130_fd_sc_hd__nand3_1 U30838 ( .A(n26812), .B(n26801), .C(n25554), .Y(
        n25548) );
  sky130_fd_sc_hd__a21oi_1 U30839 ( .A1(n25557), .A2(n29535), .B1(n25548), .Y(
        n25549) );
  sky130_fd_sc_hd__nand2_1 U30840 ( .A(n25550), .B(n25549), .Y(n25551) );
  sky130_fd_sc_hd__o211ai_1 U30841 ( .A1(n25640), .A2(n25553), .B1(n25552), 
        .C1(n25551), .Y(j202_soc_core_j22_cpu_rf_N2640) );
  sky130_fd_sc_hd__a22oi_1 U30843 ( .A1(n26948), .A2(n25555), .B1(n12389), 
        .B2(n24650), .Y(n25556) );
  sky130_fd_sc_hd__a21oi_1 U30845 ( .A1(n27471), .A2(n25562), .B1(n25561), .Y(
        n25566) );
  sky130_fd_sc_hd__and3_1 U30846 ( .A(n25563), .B(
        j202_soc_core_cmt_core_00_cnt0[2]), .C(n25567), .X(n25564) );
  sky130_fd_sc_hd__a21oi_1 U30847 ( .A1(n27482), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[3]), .B1(n25564), .Y(n25565) );
  sky130_fd_sc_hd__o21ai_1 U30848 ( .A1(n25567), .A2(n25566), .B1(n25565), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[3]) );
  sky130_fd_sc_hd__nand2_1 U30849 ( .A(j202_soc_core_cmt_core_00_cnt0[2]), .B(
        j202_soc_core_cmt_core_00_cnt0[3]), .Y(n25569) );
  sky130_fd_sc_hd__nor2_1 U30850 ( .A(n25569), .B(n25568), .Y(n25570) );
  sky130_fd_sc_hd__a21oi_1 U30851 ( .A1(n26281), .A2(n25570), .B1(
        j202_soc_core_cmt_core_00_cnt0[4]), .Y(n25571) );
  sky130_fd_sc_hd__nand2_1 U30852 ( .A(n25570), .B(
        j202_soc_core_cmt_core_00_cnt0[4]), .Y(n25573) );
  sky130_fd_sc_hd__o22ai_1 U30854 ( .A1(n27473), .A2(n26986), .B1(n25571), 
        .B2(n26916), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[4])
         );
  sky130_fd_sc_hd__nand2_1 U30855 ( .A(j202_soc_core_cmt_core_00_cnt0[5]), .B(
        j202_soc_core_cmt_core_00_cnt0[6]), .Y(n25577) );
  sky130_fd_sc_hd__nor2_1 U30856 ( .A(n25577), .B(n25573), .Y(n25582) );
  sky130_fd_sc_hd__a21oi_1 U30857 ( .A1(n27471), .A2(n25572), .B1(n28619), .Y(
        n25578) );
  sky130_fd_sc_hd__nand2_1 U30858 ( .A(n26281), .B(n25574), .Y(n26919) );
  sky130_fd_sc_hd__a21oi_1 U30859 ( .A1(n25575), .A2(
        j202_soc_core_cmt_core_00_cnt0[5]), .B1(
        j202_soc_core_cmt_core_00_cnt0[6]), .Y(n25576) );
  sky130_fd_sc_hd__o22ai_1 U30860 ( .A1(n27473), .A2(n27527), .B1(n25578), 
        .B2(n25576), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[6])
         );
  sky130_fd_sc_hd__nor2_1 U30861 ( .A(n25577), .B(n26919), .Y(n25584) );
  sky130_fd_sc_hd__a22oi_1 U30862 ( .A1(n27482), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[7]), .B1(n25579), .B2(
        j202_soc_core_cmt_core_00_cnt0[7]), .Y(n25580) );
  sky130_fd_sc_hd__nand2_1 U30864 ( .A(j202_soc_core_cmt_core_00_cnt0[7]), .B(
        j202_soc_core_cmt_core_00_cnt0[8]), .Y(n25590) );
  sky130_fd_sc_hd__nand2_1 U30865 ( .A(n25582), .B(n25581), .Y(n26277) );
  sky130_fd_sc_hd__a21oi_1 U30867 ( .A1(n25584), .A2(
        j202_soc_core_cmt_core_00_cnt0[7]), .B1(
        j202_soc_core_cmt_core_00_cnt0[8]), .Y(n25585) );
  sky130_fd_sc_hd__o22ai_1 U30868 ( .A1(n27473), .A2(n27145), .B1(n25586), 
        .B2(n25585), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[8])
         );
  sky130_fd_sc_hd__a22oi_1 U30869 ( .A1(n27482), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[9]), .B1(n25587), .B2(
        j202_soc_core_cmt_core_00_cnt0[9]), .Y(n25588) );
  sky130_fd_sc_hd__o31ai_1 U30870 ( .A1(j202_soc_core_cmt_core_00_cnt0[9]), 
        .A2(n25590), .A3(n25589), .B1(n25588), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[9]) );
  sky130_fd_sc_hd__nand2_1 U30871 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[9]), .Y(n25591) );
  sky130_fd_sc_hd__o21ai_1 U30872 ( .A1(n25619), .A2(n27827), .B1(n25591), .Y(
        n28) );
  sky130_fd_sc_hd__nand3_1 U30873 ( .A(j202_soc_core_cmt_core_00_cnt1[0]), .B(
        j202_soc_core_cmt_core_00_cnt1[2]), .C(
        j202_soc_core_cmt_core_00_cnt1[1]), .Y(n25593) );
  sky130_fd_sc_hd__nor2_1 U30874 ( .A(n25592), .B(n25593), .Y(n25597) );
  sky130_fd_sc_hd__o21ai_1 U30875 ( .A1(n26301), .A2(n25597), .B1(n26300), .Y(
        n25596) );
  sky130_fd_sc_hd__a22o_1 U30877 ( .A1(n27498), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[3]), .B1(n25596), .B2(n25594), 
        .X(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[3]) );
  sky130_fd_sc_hd__nand2_1 U30878 ( .A(n25597), .B(n27489), .Y(n25598) );
  sky130_fd_sc_hd__o22ai_1 U30879 ( .A1(n27491), .A2(n26986), .B1(
        j202_soc_core_cmt_core_00_cnt1[4]), .B2(n25598), .Y(n25595) );
  sky130_fd_sc_hd__a21o_1 U30880 ( .A1(n25596), .A2(
        j202_soc_core_cmt_core_00_cnt1[4]), .B1(n25595), .X(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[4]) );
  sky130_fd_sc_hd__nand3_1 U30881 ( .A(n25597), .B(
        j202_soc_core_cmt_core_00_cnt1[4]), .C(
        j202_soc_core_cmt_core_00_cnt1[5]), .Y(n25606) );
  sky130_fd_sc_hd__a21oi_1 U30882 ( .A1(n25606), .A2(n27489), .B1(n28622), .Y(
        n25604) );
  sky130_fd_sc_hd__nor2_1 U30883 ( .A(n25599), .B(n25598), .Y(n25605) );
  sky130_fd_sc_hd__nor2_1 U30884 ( .A(j202_soc_core_cmt_core_00_cnt1[5]), .B(
        n25605), .Y(n25600) );
  sky130_fd_sc_hd__o22ai_1 U30885 ( .A1(n27491), .A2(n26924), .B1(n25604), 
        .B2(n25600), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[5])
         );
  sky130_fd_sc_hd__nor2_1 U30886 ( .A(n27527), .B(n27491), .Y(n25601) );
  sky130_fd_sc_hd__a31oi_1 U30887 ( .A1(n25605), .A2(
        j202_soc_core_cmt_core_00_cnt1[5]), .A3(n25603), .B1(n25601), .Y(
        n25602) );
  sky130_fd_sc_hd__a31oi_1 U30889 ( .A1(n25605), .A2(
        j202_soc_core_cmt_core_00_cnt1[6]), .A3(
        j202_soc_core_cmt_core_00_cnt1[5]), .B1(
        j202_soc_core_cmt_core_00_cnt1[7]), .Y(n25608) );
  sky130_fd_sc_hd__nand2_1 U30890 ( .A(j202_soc_core_cmt_core_00_cnt1[6]), .B(
        j202_soc_core_cmt_core_00_cnt1[7]), .Y(n25607) );
  sky130_fd_sc_hd__nor2_1 U30891 ( .A(n25607), .B(n25606), .Y(n25614) );
  sky130_fd_sc_hd__a21oi_1 U30892 ( .A1(n25609), .A2(n27489), .B1(n28622), .Y(
        n25612) );
  sky130_fd_sc_hd__o22ai_1 U30893 ( .A1(n27326), .A2(n27491), .B1(n25608), 
        .B2(n25612), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[7])
         );
  sky130_fd_sc_hd__nor3_1 U30894 ( .A(j202_soc_core_cmt_core_00_cnt1[8]), .B(
        n26301), .C(n25609), .Y(n25610) );
  sky130_fd_sc_hd__a21oi_1 U30895 ( .A1(n27498), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[8]), .B1(n25610), .Y(n25611) );
  sky130_fd_sc_hd__o21ai_1 U30896 ( .A1(n25613), .A2(n25612), .B1(n25611), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[8]) );
  sky130_fd_sc_hd__nand3_1 U30897 ( .A(n25614), .B(
        j202_soc_core_cmt_core_00_cnt1[8]), .C(
        j202_soc_core_cmt_core_00_cnt1[9]), .Y(n26298) );
  sky130_fd_sc_hd__nand2_1 U30899 ( .A(n26293), .B(
        j202_soc_core_cmt_core_00_cnt1[9]), .Y(n25617) );
  sky130_fd_sc_hd__nand2_1 U30900 ( .A(n27498), .B(
        j202_soc_core_cmt_core_00_wdata_cnt0[9]), .Y(n25616) );
  sky130_fd_sc_hd__nand4_1 U30901 ( .A(n26298), .B(n25614), .C(n27489), .D(
        j202_soc_core_cmt_core_00_cnt1[8]), .Y(n25615) );
  sky130_fd_sc_hd__nand3_1 U30902 ( .A(n25617), .B(n25616), .C(n25615), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[9]) );
  sky130_fd_sc_hd__nand2_1 U30903 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[9]), .Y(n25618) );
  sky130_fd_sc_hd__o21ai_1 U30904 ( .A1(n25619), .A2(n27833), .B1(n25618), .Y(
        n29) );
  sky130_fd_sc_hd__a22oi_1 U30905 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[9]), .B1(n27837), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[9]), .Y(
        n25622) );
  sky130_fd_sc_hd__nand2_1 U30906 ( .A(n27840), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[9]), .Y(
        n25621) );
  sky130_fd_sc_hd__nand2_1 U30907 ( .A(n27835), .B(
        j202_soc_core_cmt_core_00_const1[9]), .Y(n25620) );
  sky130_fd_sc_hd__nand3_1 U30908 ( .A(n25622), .B(n25621), .C(n25620), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[9]) );
  sky130_fd_sc_hd__nand2_1 U30909 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[9]), .Y(n25623) );
  sky130_fd_sc_hd__o21ai_1 U30910 ( .A1(n25624), .A2(n27983), .B1(n25623), .Y(
        n30) );
  sky130_fd_sc_hd__o22ai_1 U30911 ( .A1(n28601), .A2(n27990), .B1(n25625), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U30912 ( .A1(n28601), .A2(n28535), .B1(n25626), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U30913 ( .A1(n28601), .A2(n28547), .B1(n25627), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U30914 ( .A1(n28601), .A2(n28538), .B1(n25628), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U30915 ( .A1(n28601), .A2(n28541), .B1(n25629), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U30916 ( .A1(n28544), .A2(n28601), .B1(n25630), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__a22oi_1 U30917 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[9]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[73]), .Y(n25632) );
  sky130_fd_sc_hd__a22oi_1 U30918 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[9]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[9]), .Y(n25631) );
  sky130_fd_sc_hd__nand3_1 U30919 ( .A(n25632), .B(n25631), .C(n27865), .Y(
        n25633) );
  sky130_fd_sc_hd__a21oi_1 U30920 ( .A1(n27869), .A2(
        j202_soc_core_intc_core_00_rg_itgt[42]), .B1(n25633), .Y(n25637) );
  sky130_fd_sc_hd__a22oi_1 U30921 ( .A1(n27856), .A2(
        j202_soc_core_intc_core_00_rg_itgt[50]), .B1(n27850), .B2(
        j202_soc_core_intc_core_00_rg_itgt[34]), .Y(n25636) );
  sky130_fd_sc_hd__a22oi_1 U30922 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[58]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[105]), .Y(n25635) );
  sky130_fd_sc_hd__nand2_1 U30923 ( .A(n27862), .B(
        j202_soc_core_intc_core_00_rg_ipr[41]), .Y(n25634) );
  sky130_fd_sc_hd__nand4_1 U30924 ( .A(n25637), .B(n25636), .C(n25635), .D(
        n25634), .Y(j202_soc_core_ahb2apb_01_N137) );
  sky130_fd_sc_hd__nand2_1 U30925 ( .A(n12389), .B(n27343), .Y(n25638) );
  sky130_fd_sc_hd__o21ai_0 U30926 ( .A1(n25788), .A2(n27343), .B1(n25638), .Y(
        j202_soc_core_j22_cpu_ml_N312) );
  sky130_fd_sc_hd__o22ai_1 U30927 ( .A1(n27333), .A2(n25640), .B1(n23178), 
        .B2(n25639), .Y(j202_soc_core_j22_cpu_rf_N3058) );
  sky130_fd_sc_hd__a21oi_1 U30928 ( .A1(n25815), .A2(n25811), .B1(n11078), .Y(
        n25641) );
  sky130_fd_sc_hd__nand2_1 U30929 ( .A(n27522), .B(n25641), .Y(n10494) );
  sky130_fd_sc_hd__o22ai_1 U30931 ( .A1(n27333), .A2(n27464), .B1(n23178), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N3060) );
  sky130_fd_sc_hd__o22ai_1 U30932 ( .A1(n27219), .A2(n27464), .B1(n27218), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N2986) );
  sky130_fd_sc_hd__o22ai_1 U30933 ( .A1(n27217), .A2(n27464), .B1(n27216), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N2838) );
  sky130_fd_sc_hd__o22ai_1 U30934 ( .A1(n27228), .A2(n27464), .B1(n27227), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N3171) );
  sky130_fd_sc_hd__o22ai_1 U30935 ( .A1(n27225), .A2(n27464), .B1(n27224), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N2949) );
  sky130_fd_sc_hd__o22ai_1 U30936 ( .A1(n27215), .A2(n27464), .B1(n27214), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N2912) );
  sky130_fd_sc_hd__o22ai_1 U30937 ( .A1(n27223), .A2(n27464), .B1(n27222), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N3023) );
  sky130_fd_sc_hd__o22ai_1 U30938 ( .A1(n27211), .A2(n27464), .B1(n27210), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N3208) );
  sky130_fd_sc_hd__o22ai_1 U30939 ( .A1(n27221), .A2(n27464), .B1(n27220), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N2875) );
  sky130_fd_sc_hd__o22ai_1 U30940 ( .A1(n27226), .A2(n27464), .B1(n23079), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N3134) );
  sky130_fd_sc_hd__o22ai_1 U30941 ( .A1(n27213), .A2(n27464), .B1(n27212), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N2801) );
  sky130_fd_sc_hd__o22ai_1 U30942 ( .A1(n27209), .A2(n27464), .B1(n23039), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N2727) );
  sky130_fd_sc_hd__o22ai_1 U30943 ( .A1(n25649), .A2(n27021), .B1(n25642), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U30944 ( .A1(n25649), .A2(n27990), .B1(n25643), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U30945 ( .A1(n25649), .A2(n28535), .B1(n25644), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U30946 ( .A1(n25649), .A2(n28547), .B1(n25645), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U30947 ( .A1(n25649), .A2(n28538), .B1(n25651), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U30948 ( .A1(n25649), .A2(n28541), .B1(n25646), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U30949 ( .A1(n28544), .A2(n25649), .B1(n25647), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U30950 ( .A1(n25649), .A2(n27194), .B1(n25648), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__a21oi_1 U30951 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[27]), .B1(n27758), .Y(n25650) );
  sky130_fd_sc_hd__o21ai_1 U30952 ( .A1(n25651), .A2(n27097), .B1(n25650), .Y(
        n25652) );
  sky130_fd_sc_hd__a21oi_1 U30953 ( .A1(j202_soc_core_intc_core_00_rg_ipr[59]), 
        .A2(n27862), .B1(n25652), .Y(n25657) );
  sky130_fd_sc_hd__a22o_1 U30954 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[27]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[91]), .X(n25653) );
  sky130_fd_sc_hd__a21oi_1 U30955 ( .A1(n27850), .A2(
        j202_soc_core_intc_core_00_rg_itgt[102]), .B1(n25653), .Y(n25656) );
  sky130_fd_sc_hd__a22oi_1 U30956 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[126]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[123]), .Y(n25655) );
  sky130_fd_sc_hd__nand2_1 U30957 ( .A(n27869), .B(
        j202_soc_core_intc_core_00_rg_itgt[110]), .Y(n25654) );
  sky130_fd_sc_hd__nand4_1 U30958 ( .A(n25657), .B(n25656), .C(n25655), .D(
        n25654), .Y(j202_soc_core_ahb2apb_01_N155) );
  sky130_fd_sc_hd__nand2_1 U30959 ( .A(n27108), .B(j202_soc_core_uart_div0[3]), 
        .Y(n25658) );
  sky130_fd_sc_hd__o21ai_1 U30960 ( .A1(n25659), .A2(n27108), .B1(n25658), .Y(
        n41) );
  sky130_fd_sc_hd__a22o_1 U30961 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[27]), .A2(n27719), .B1(n27718), 
        .B2(j202_soc_core_wbqspiflash_00_quad_mode_enabled), .X(
        j202_soc_core_wbqspiflash_00_N694) );
  sky130_fd_sc_hd__nand2_1 U30962 ( .A(n11770), .B(n27460), .Y(n25660) );
  sky130_fd_sc_hd__inv_1 U30964 ( .A(n25662), .Y(n25666) );
  sky130_fd_sc_hd__nand4_1 U30965 ( .A(n25665), .B(n25666), .C(n25664), .D(
        n25663), .Y(n25668) );
  sky130_fd_sc_hd__a21oi_1 U30966 ( .A1(n25666), .A2(n29535), .B1(n26951), .Y(
        n25667) );
  sky130_fd_sc_hd__nand2_1 U30967 ( .A(n25668), .B(n25667), .Y(n25671) );
  sky130_fd_sc_hd__a22oi_1 U30968 ( .A1(n25669), .A2(n26948), .B1(n11770), 
        .B2(n24650), .Y(n25670) );
  sky130_fd_sc_hd__nand2_1 U30969 ( .A(n25671), .B(n25670), .Y(
        j202_soc_core_j22_cpu_rf_N3366) );
  sky130_fd_sc_hd__o22ai_1 U30970 ( .A1(n28600), .A2(n27021), .B1(n25672), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U30971 ( .A1(n28600), .A2(n28535), .B1(n25673), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U30972 ( .A1(n28600), .A2(n28538), .B1(n25674), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U30973 ( .A1(n28600), .A2(n28541), .B1(n25675), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U30974 ( .A1(n28600), .A2(n27194), .B1(n25689), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__nand3_1 U30975 ( .A(n25677), .B(n27604), .C(n25676), .Y(
        n25678) );
  sky130_fd_sc_hd__mux2_2 U30976 ( .A0(j202_soc_core_bldc_core_00_wdata[0]), 
        .A1(j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_), .S(
        n25678), .X(n45) );
  sky130_fd_sc_hd__nor2_1 U30977 ( .A(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_0_), .B(n29050), .Y(n25679) );
  sky130_fd_sc_hd__a211oi_1 U30978 ( .A1(n29050), .A2(n27741), .B1(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_wen), .C1(
        n25679), .Y(n44) );
  sky130_fd_sc_hd__nor2_1 U30979 ( .A(
        j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_2), .B(n25680), 
        .Y(n25681) );
  sky130_fd_sc_hd__a22oi_1 U30980 ( .A1(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_0_), .A2(n25682), .B1(n25681), .B2(
        j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1), .Y(n25683)
         );
  sky130_fd_sc_hd__o21ai_1 U30981 ( .A1(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_0_), .A2(
        n25684), .B1(n25683), .Y(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_nxt_latch_status_0_) );
  sky130_fd_sc_hd__nor2_1 U30982 ( .A(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_wen), .B(
        n25684), .Y(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_nxt_bldc_int) );
  sky130_fd_sc_hd__nand3_1 U30983 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[4]), .B(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[6]), .C(j202_soc_core_intc_core_00_cp_intack_all_0_), .Y(n25724) );
  sky130_fd_sc_hd__nor2_1 U30984 ( .A(n28512), .B(n25724), .Y(n26817) );
  sky130_fd_sc_hd__a21oi_1 U30985 ( .A1(n25747), .A2(n26817), .B1(
        j202_soc_core_intc_core_00_rg_irqc[19]), .Y(n25687) );
  sky130_fd_sc_hd__nor2_1 U30986 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[19]), 
        .B(n25685), .Y(n25686) );
  sky130_fd_sc_hd__a31oi_1 U30987 ( .A1(n25687), .A2(
        j202_soc_core_intc_core_00_in_intreq[19]), .A3(n29594), .B1(n25686), 
        .Y(n25688) );
  sky130_fd_sc_hd__nor2_1 U30988 ( .A(n25689), .B(n25688), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N22) );
  sky130_fd_sc_hd__a22oi_1 U30989 ( .A1(n27869), .A2(
        j202_soc_core_intc_core_00_rg_itgt[108]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[19]), .Y(n25691) );
  sky130_fd_sc_hd__a222oi_1 U30990 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[19]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[83]), .C1(n27861), .C2(
        j202_soc_core_intc_core_00_rg_itgt[124]), .Y(n25690) );
  sky130_fd_sc_hd__nand2_1 U30991 ( .A(n25691), .B(n25690), .Y(n25697) );
  sky130_fd_sc_hd__a21oi_1 U30993 ( .A1(n27850), .A2(
        j202_soc_core_intc_core_00_rg_itgt[100]), .B1(n25693), .Y(n25696) );
  sky130_fd_sc_hd__a22oi_1 U30994 ( .A1(n27862), .A2(
        j202_soc_core_intc_core_00_rg_ipr[51]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[115]), .Y(n25695) );
  sky130_fd_sc_hd__nand2_1 U30995 ( .A(n27856), .B(
        j202_soc_core_intc_core_00_rg_itgt[116]), .Y(n25694) );
  sky130_fd_sc_hd__nand4b_1 U30996 ( .A_N(n25697), .B(n25696), .C(n25695), .D(
        n25694), .Y(j202_soc_core_ahb2apb_01_N147) );
  sky130_fd_sc_hd__nand2_1 U30997 ( .A(n27593), .B(j202_soc_core_uart_div1[3]), 
        .Y(n25698) );
  sky130_fd_sc_hd__nor2_1 U30999 ( .A(n28590), .B(n28188), .Y(
        j202_soc_core_wbqspiflash_00_N716) );
  sky130_fd_sc_hd__a22o_1 U31000 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[19]), .A2(n27719), .B1(n27718), 
        .B2(j202_soc_core_wbqspiflash_00_erased_sector[5]), .X(
        j202_soc_core_wbqspiflash_00_N686) );
  sky130_fd_sc_hd__nand2_1 U31001 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[19]), .Y(n25700) );
  sky130_fd_sc_hd__o21ai_1 U31002 ( .A1(n25701), .A2(n27983), .B1(n25700), .Y(
        n27) );
  sky130_fd_sc_hd__a22oi_1 U31003 ( .A1(n27184), .A2(n26719), .B1(n11770), 
        .B2(n27339), .Y(n25702) );
  sky130_fd_sc_hd__nand2_1 U31004 ( .A(n27346), .B(n25702), .Y(
        j202_soc_core_j22_cpu_ml_N322) );
  sky130_fd_sc_hd__a22oi_1 U31005 ( .A1(n27187), .A2(n22951), .B1(n27273), 
        .B2(n25703), .Y(n25704) );
  sky130_fd_sc_hd__nand2_1 U31006 ( .A(n27189), .B(n25704), .Y(
        j202_soc_core_j22_cpu_ml_machj[19]) );
  sky130_fd_sc_hd__nand2_1 U31007 ( .A(n25705), .B(n27192), .Y(n25706) );
  sky130_fd_sc_hd__o21ai_0 U31008 ( .A1(n27192), .A2(n11103), .B1(n25706), .Y(
        j202_soc_core_j22_cpu_rf_N3289) );
  sky130_fd_sc_hd__o22ai_1 U31009 ( .A1(n26899), .A2(n11103), .B1(n26898), 
        .B2(n25707), .Y(j202_soc_core_j22_cpu_rf_N3328) );
  sky130_fd_sc_hd__nand4_1 U31010 ( .A(n25711), .B(n25710), .C(n25709), .D(
        n25708), .Y(n25713) );
  sky130_fd_sc_hd__a21oi_1 U31011 ( .A1(n25711), .A2(n29535), .B1(n26951), .Y(
        n25712) );
  sky130_fd_sc_hd__nand2_1 U31012 ( .A(n25713), .B(n25712), .Y(n25717) );
  sky130_fd_sc_hd__a2bb2oi_1 U31013 ( .B1(n26948), .B2(n25715), .A1_N(n25714), 
        .A2_N(n11103), .Y(n25716) );
  sky130_fd_sc_hd__nand2_1 U31014 ( .A(n25717), .B(n25716), .Y(
        j202_soc_core_j22_cpu_rf_N3364) );
  sky130_fd_sc_hd__o22ai_1 U31015 ( .A1(n28602), .A2(n27021), .B1(n25718), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U31016 ( .A1(n28602), .A2(n27990), .B1(n25719), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U31017 ( .A1(n28602), .A2(n28547), .B1(n25720), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U31018 ( .A1(n28602), .A2(n28538), .B1(n25721), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U31019 ( .A1(n28602), .A2(n28541), .B1(n25722), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U31020 ( .A1(n28602), .A2(n27194), .B1(n25729), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__nand2_1 U31021 ( .A(n27831), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[6]), .Y(n25723) );
  sky130_fd_sc_hd__o21ai_1 U31022 ( .A1(n27527), .A2(n27831), .B1(n25723), .Y(
        n103) );
  sky130_fd_sc_hd__nand3_1 U31023 ( .A(j202_soc_core_cmt_core_00_cmf1), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[6]), .C(n29593), .Y(
        n25725) );
  sky130_fd_sc_hd__nor2_1 U31024 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[1]), .B(n25724), .Y(n26480) );
  sky130_fd_sc_hd__a21oi_1 U31025 ( .A1(n26480), .A2(n25747), .B1(
        j202_soc_core_intc_core_00_rg_irqc[17]), .Y(n25727) );
  sky130_fd_sc_hd__nor2_1 U31026 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[17]), 
        .B(n25725), .Y(n25726) );
  sky130_fd_sc_hd__a31oi_1 U31027 ( .A1(n25727), .A2(
        j202_soc_core_intc_core_00_in_intreq[17]), .A3(n29594), .B1(n25726), 
        .Y(n25728) );
  sky130_fd_sc_hd__nor2_1 U31028 ( .A(n25729), .B(n25728), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N20) );
  sky130_fd_sc_hd__o22ai_1 U31029 ( .A1(n28544), .A2(n28602), .B1(n25730), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__a22oi_1 U31030 ( .A1(n27860), .A2(
        j202_soc_core_intc_core_00_rg_ipr[113]), .B1(n27869), .B2(
        j202_soc_core_intc_core_00_rg_itgt[44]), .Y(n25738) );
  sky130_fd_sc_hd__a22oi_1 U31031 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[17]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[81]), .Y(n25737) );
  sky130_fd_sc_hd__nand2_1 U31032 ( .A(n27862), .B(
        j202_soc_core_intc_core_00_rg_ipr[49]), .Y(n25736) );
  sky130_fd_sc_hd__nand2_1 U31033 ( .A(n27856), .B(
        j202_soc_core_intc_core_00_rg_itgt[52]), .Y(n25733) );
  sky130_fd_sc_hd__a22oi_1 U31034 ( .A1(n27850), .A2(
        j202_soc_core_intc_core_00_rg_itgt[36]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[17]), .Y(n25732) );
  sky130_fd_sc_hd__nand2_1 U31035 ( .A(n27864), .B(
        j202_soc_core_intc_core_00_in_intreq[17]), .Y(n25731) );
  sky130_fd_sc_hd__nand4_1 U31036 ( .A(n25733), .B(n25732), .C(n27865), .D(
        n25731), .Y(n25734) );
  sky130_fd_sc_hd__a21oi_1 U31037 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[60]), .B1(n25734), .Y(n25735) );
  sky130_fd_sc_hd__nand4_1 U31038 ( .A(n25738), .B(n25737), .C(n25736), .D(
        n25735), .Y(j202_soc_core_ahb2apb_01_N145) );
  sky130_fd_sc_hd__nand2_1 U31039 ( .A(n27593), .B(j202_soc_core_uart_div1[1]), 
        .Y(n25739) );
  sky130_fd_sc_hd__nor2_1 U31041 ( .A(n28590), .B(n25740), .Y(
        j202_soc_core_wbqspiflash_00_N714) );
  sky130_fd_sc_hd__a22o_1 U31042 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[17]), .A2(n27719), .B1(n27718), 
        .B2(j202_soc_core_wbqspiflash_00_erased_sector[3]), .X(
        j202_soc_core_wbqspiflash_00_N684) );
  sky130_fd_sc_hd__nand2_1 U31043 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[17]), .Y(n25741) );
  sky130_fd_sc_hd__mux2i_1 U31045 ( .A0(n27335), .A1(n25743), .S(n27006), .Y(
        j202_soc_core_j22_cpu_ml_N304) );
  sky130_fd_sc_hd__o21ai_1 U31046 ( .A1(n25745), .A2(n27274), .B1(n27273), .Y(
        j202_soc_core_j22_cpu_ml_machj[1]) );
  sky130_fd_sc_hd__o22ai_1 U31047 ( .A1(n28603), .A2(n27194), .B1(n25752), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__a21oi_1 U31048 ( .A1(n25747), .A2(n25746), .B1(
        j202_soc_core_intc_core_00_rg_irqc[1]), .Y(n25750) );
  sky130_fd_sc_hd__nor2_1 U31049 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[1]), 
        .B(n25748), .Y(n25749) );
  sky130_fd_sc_hd__a31oi_1 U31050 ( .A1(n25750), .A2(
        j202_soc_core_intc_core_00_in_intreq[1]), .A3(n29594), .B1(n25749), 
        .Y(n25751) );
  sky130_fd_sc_hd__nor2_1 U31051 ( .A(n25752), .B(n25751), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N4) );
  sky130_fd_sc_hd__inv_1 U31052 ( .A(n25753), .Y(n25755) );
  sky130_fd_sc_hd__o22ai_1 U31053 ( .A1(n25755), .A2(n26904), .B1(n25754), 
        .B2(n26902), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N3) );
  sky130_fd_sc_hd__a21oi_1 U31054 ( .A1(j202_soc_core_intr_level__0_), .A2(
        n26907), .B1(n26906), .Y(n25758) );
  sky130_fd_sc_hd__nand2_1 U31055 ( .A(n11704), .B(n26908), .Y(n25757) );
  sky130_fd_sc_hd__o211ai_1 U31056 ( .A1(n26911), .A2(n27208), .B1(n25758), 
        .C1(n25757), .Y(j202_soc_core_j22_cpu_rf_N3386) );
  sky130_fd_sc_hd__a22oi_1 U31057 ( .A1(n25759), .A2(n26948), .B1(n11704), 
        .B2(n24650), .Y(n25760) );
  sky130_fd_sc_hd__o21ai_0 U31058 ( .A1(n26951), .A2(n27208), .B1(n25760), .Y(
        j202_soc_core_j22_cpu_rf_N3349) );
  sky130_fd_sc_hd__o22ai_1 U31059 ( .A1(n27583), .A2(n25761), .B1(n28300), 
        .B2(n27581), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U31060 ( .A1(n28606), .A2(n27194), .B1(n25767), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__nand2_1 U31061 ( .A(n27829), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[6]), .Y(n25762) );
  sky130_fd_sc_hd__nand3_1 U31063 ( .A(j202_soc_core_cmt_core_00_cmf0), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[6]), .C(n29593), .Y(
        n25763) );
  sky130_fd_sc_hd__a21oi_1 U31064 ( .A1(n26480), .A2(n27195), .B1(
        j202_soc_core_intc_core_00_rg_irqc[16]), .Y(n25765) );
  sky130_fd_sc_hd__nor2_1 U31065 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[16]), 
        .B(n25763), .Y(n25764) );
  sky130_fd_sc_hd__a31oi_1 U31066 ( .A1(n25765), .A2(
        j202_soc_core_intc_core_00_in_intreq[16]), .A3(n29594), .B1(n25764), 
        .Y(n25766) );
  sky130_fd_sc_hd__nor2_1 U31067 ( .A(n25767), .B(n25766), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N19) );
  sky130_fd_sc_hd__o22ai_1 U31068 ( .A1(n27583), .A2(n25768), .B1(n27755), 
        .B2(n27581), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__mux2i_1 U31069 ( .A0(n25770), .A1(n26836), .S(n11700), .Y(
        n25774) );
  sky130_fd_sc_hd__o22ai_1 U31070 ( .A1(n25772), .A2(n26824), .B1(n26827), 
        .B2(n27207), .Y(n25773) );
  sky130_fd_sc_hd__mux2i_1 U31071 ( .A0(n25774), .A1(n25773), .S(n12125), .Y(
        n25777) );
  sky130_fd_sc_hd__nand3_1 U31072 ( .A(n29069), .B(n25775), .C(n26847), .Y(
        n25776) );
  sky130_fd_sc_hd__o211ai_1 U31073 ( .A1(n25777), .A2(n26904), .B1(n27018), 
        .C1(n25776), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N4) );
  sky130_fd_sc_hd__or3_1 U31074 ( .A(j202_soc_core_intr_vec__0_), .B(
        j202_soc_core_intr_vec__4_), .C(j202_soc_core_intr_vec__3_), .X(n25778) );
  sky130_fd_sc_hd__nor3_1 U31075 ( .A(j202_soc_core_intr_vec__2_), .B(
        j202_soc_core_intr_vec__6_), .C(n25778), .Y(n27918) );
  sky130_fd_sc_hd__nand2_1 U31076 ( .A(n27932), .B(n25780), .Y(n27944) );
  sky130_fd_sc_hd__a31oi_1 U31077 ( .A1(j202_soc_core_j22_cpu_opst[1]), .A2(
        n27918), .A3(n28511), .B1(n27944), .Y(
        j202_soc_core_j22_cpu_id_idec_N822) );
  sky130_fd_sc_hd__a211oi_1 U31078 ( .A1(n25783), .A2(n25782), .B1(
        j202_soc_core_intc_core_00_cp_intack_all_0_), .C1(n28518), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_req_N3) );
  sky130_fd_sc_hd__a31oi_1 U31079 ( .A1(n25785), .A2(n26318), .A3(n25784), 
        .B1(n29535), .Y(n25786) );
  sky130_fd_sc_hd__o22ai_1 U31080 ( .A1(n25789), .A2(n26416), .B1(n25788), 
        .B2(n26424), .Y(n25790) );
  sky130_fd_sc_hd__a21oi_1 U31081 ( .A1(n26341), .A2(n25871), .B1(n25790), .Y(
        n25797) );
  sky130_fd_sc_hd__nand2_1 U31082 ( .A(n25792), .B(n25791), .Y(n25794) );
  sky130_fd_sc_hd__nand2_1 U31083 ( .A(n27396), .B(n26710), .Y(n26588) );
  sky130_fd_sc_hd__o2bb2ai_1 U31084 ( .B1(n26432), .B2(n26588), .A1_N(n27045), 
        .A2_N(n26077), .Y(n25793) );
  sky130_fd_sc_hd__a21oi_1 U31085 ( .A1(n25794), .A2(n26329), .B1(n25793), .Y(
        n25796) );
  sky130_fd_sc_hd__o22a_1 U31086 ( .A1(n26325), .A2(n26418), .B1(n11145), .B2(
        n26419), .X(n25795) );
  sky130_fd_sc_hd__nand4_1 U31087 ( .A(n25797), .B(n25796), .C(n25795), .D(
        n26344), .Y(n25804) );
  sky130_fd_sc_hd__nor2_1 U31088 ( .A(n26710), .B(n27396), .Y(n26668) );
  sky130_fd_sc_hd__nor3_1 U31089 ( .A(n26415), .B(n26668), .C(n26667), .Y(
        n25800) );
  sky130_fd_sc_hd__nor2_1 U31090 ( .A(n25798), .B(n26427), .Y(n25799) );
  sky130_fd_sc_hd__a211o_1 U31091 ( .A1(n26338), .A2(n27455), .B1(n25800), 
        .C1(n25799), .X(n25801) );
  sky130_fd_sc_hd__a21oi_1 U31092 ( .A1(n26342), .A2(n27392), .B1(n25801), .Y(
        n25803) );
  sky130_fd_sc_hd__mux2_2 U31093 ( .A0(n26423), .A1(n26349), .S(n27396), .X(
        n25802) );
  sky130_fd_sc_hd__nand3b_1 U31094 ( .A_N(n25804), .B(n25803), .C(n25802), .Y(
        n25805) );
  sky130_fd_sc_hd__a21oi_1 U31095 ( .A1(n25806), .A2(n26409), .B1(n25805), .Y(
        n25808) );
  sky130_fd_sc_hd__o21ai_0 U31096 ( .A1(n26352), .A2(n26710), .B1(n26351), .Y(
        n25807) );
  sky130_fd_sc_hd__nand3_1 U31097 ( .A(n25811), .B(n27980), .C(n12617), .Y(
        n25812) );
  sky130_fd_sc_hd__nand2_1 U31098 ( .A(n25813), .B(n25812), .Y(n25814) );
  sky130_fd_sc_hd__nand3_1 U31099 ( .A(n13186), .B(n25817), .C(n25816), .Y(
        n10495) );
  sky130_fd_sc_hd__nand2_1 U31100 ( .A(n27395), .B(n27343), .Y(n25820) );
  sky130_fd_sc_hd__o21ai_0 U31101 ( .A1(n25821), .A2(n27343), .B1(n25820), .Y(
        j202_soc_core_j22_cpu_ml_N311) );
  sky130_fd_sc_hd__o21ai_1 U31102 ( .A1(n25824), .A2(n25823), .B1(n25822), .Y(
        n25825) );
  sky130_fd_sc_hd__a31oi_1 U31103 ( .A1(n25873), .A2(n26872), .A3(n12356), 
        .B1(n25825), .Y(n25828) );
  sky130_fd_sc_hd__nand2_1 U31104 ( .A(n25828), .B(n25827), .Y(
        j202_soc_core_j22_cpu_ml_maclj[8]) );
  sky130_fd_sc_hd__a21oi_1 U31105 ( .A1(n25830), .A2(n27187), .B1(n25829), .Y(
        n25831) );
  sky130_fd_sc_hd__o21ai_1 U31106 ( .A1(n27274), .A2(n25832), .B1(n25831), .Y(
        j202_soc_core_j22_cpu_ml_machj[8]) );
  sky130_fd_sc_hd__nand2_1 U31107 ( .A(n25810), .B(n27192), .Y(n25833) );
  sky130_fd_sc_hd__nand3_1 U31108 ( .A(n25834), .B(n26755), .C(n26782), .Y(
        n26777) );
  sky130_fd_sc_hd__nand2b_1 U31109 ( .A_N(n27334), .B(n26777), .Y(n25846) );
  sky130_fd_sc_hd__nor2_1 U31110 ( .A(n26777), .B(n14849), .Y(n25840) );
  sky130_fd_sc_hd__nor2_1 U31111 ( .A(n25840), .B(n26803), .Y(n25842) );
  sky130_fd_sc_hd__xnor2_1 U31112 ( .A(j202_soc_core_j22_cpu_rfuo_sr__q_), .B(
        n26859), .Y(n25839) );
  sky130_fd_sc_hd__xor2_1 U31113 ( .A(n25839), .B(n26745), .X(n26686) );
  sky130_fd_sc_hd__a22oi_1 U31114 ( .A1(n26742), .A2(n26859), .B1(n26686), 
        .B2(n16492), .Y(n25841) );
  sky130_fd_sc_hd__a2bb2oi_1 U31115 ( .B1(n25842), .B2(n27395), .A1_N(n25841), 
        .A2_N(n25847), .Y(n25843) );
  sky130_fd_sc_hd__o21a_1 U31116 ( .A1(n11559), .A2(n25846), .B1(n25843), .X(
        n25844) );
  sky130_fd_sc_hd__o21ai_1 U31117 ( .A1(n25846), .A2(n25845), .B1(n25844), .Y(
        j202_soc_core_j22_cpu_rf_N2638) );
  sky130_fd_sc_hd__nand2_1 U31118 ( .A(n26814), .B(n25847), .Y(
        j202_soc_core_j22_cpu_rf_N2637) );
  sky130_fd_sc_hd__nand2_1 U31119 ( .A(n25810), .B(n26516), .Y(n25850) );
  sky130_fd_sc_hd__a22oi_1 U31120 ( .A1(n26948), .A2(n25848), .B1(n27395), 
        .B2(n24650), .Y(n25849) );
  sky130_fd_sc_hd__nand2_1 U31121 ( .A(n25850), .B(n25849), .Y(
        j202_soc_core_j22_cpu_rf_N3354) );
  sky130_fd_sc_hd__a22oi_1 U31122 ( .A1(n25851), .A2(n26948), .B1(n12647), 
        .B2(n24650), .Y(n25852) );
  sky130_fd_sc_hd__o22ai_1 U31124 ( .A1(n27021), .A2(n25858), .B1(n25854), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U31125 ( .A1(n25858), .A2(n27990), .B1(n25862), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U31126 ( .A1(n27757), .A2(n25855), .B1(n28447), 
        .B2(n27754), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U31127 ( .A1(n27583), .A2(n25860), .B1(n28447), 
        .B2(n27581), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U31128 ( .A1(n28541), .A2(n25858), .B1(n25856), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U31129 ( .A1(n25858), .A2(n27194), .B1(n25857), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__a21oi_1 U31130 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[24]), .B1(n27758), .Y(n25859) );
  sky130_fd_sc_hd__a21oi_1 U31132 ( .A1(j202_soc_core_intc_core_00_rg_ipr[56]), 
        .A2(n27862), .B1(n25861), .Y(n25868) );
  sky130_fd_sc_hd__o22ai_1 U31133 ( .A1(n25863), .A2(n27676), .B1(n27312), 
        .B2(n25862), .Y(n25864) );
  sky130_fd_sc_hd__a21oi_1 U31134 ( .A1(j202_soc_core_intc_core_00_rg_itgt[6]), 
        .A2(n27850), .B1(n25864), .Y(n25867) );
  sky130_fd_sc_hd__a22oi_1 U31135 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[30]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[120]), .Y(n25866) );
  sky130_fd_sc_hd__nand2_1 U31136 ( .A(n27869), .B(
        j202_soc_core_intc_core_00_rg_itgt[14]), .Y(n25865) );
  sky130_fd_sc_hd__nand4_1 U31137 ( .A(n25868), .B(n25867), .C(n25866), .D(
        n25865), .Y(j202_soc_core_ahb2apb_01_N152) );
  sky130_fd_sc_hd__nand2_1 U31138 ( .A(n27108), .B(j202_soc_core_uart_div0[0]), 
        .Y(n25869) );
  sky130_fd_sc_hd__a22oi_1 U31140 ( .A1(n27184), .A2(n25871), .B1(n12647), 
        .B2(n27339), .Y(n25872) );
  sky130_fd_sc_hd__nand2_1 U31141 ( .A(n27346), .B(n25872), .Y(
        j202_soc_core_j22_cpu_ml_N328) );
  sky130_fd_sc_hd__a21oi_1 U31142 ( .A1(n25875), .A2(n25874), .B1(n26976), .Y(
        n25876) );
  sky130_fd_sc_hd__o21ai_1 U31143 ( .A1(n25877), .A2(n12917), .B1(n25876), .Y(
        j202_soc_core_j22_cpu_ml_maclj[24]) );
  sky130_fd_sc_hd__nand2_1 U31144 ( .A(n25878), .B(n27192), .Y(n25879) );
  sky130_fd_sc_hd__o21ai_0 U31145 ( .A1(n27192), .A2(n27394), .B1(n25879), .Y(
        j202_soc_core_j22_cpu_rf_N3297) );
  sky130_fd_sc_hd__nand4_1 U31146 ( .A(n29055), .B(n26147), .C(n26171), .D(
        n28116), .Y(n25896) );
  sky130_fd_sc_hd__nand3_1 U31147 ( .A(n25882), .B(n25881), .C(n25880), .Y(
        n25883) );
  sky130_fd_sc_hd__nand2_1 U31148 ( .A(n25883), .B(j202_soc_core_qspi_wb_cyc), 
        .Y(n26250) );
  sky130_fd_sc_hd__o21ai_1 U31149 ( .A1(j202_soc_core_wbqspiflash_00_state[4]), 
        .A2(n25961), .B1(n25884), .Y(n25889) );
  sky130_fd_sc_hd__a21oi_1 U31150 ( .A1(n25890), .A2(n26141), .B1(n28250), .Y(
        n25888) );
  sky130_fd_sc_hd__nor2_1 U31151 ( .A(n25993), .B(n26012), .Y(n25905) );
  sky130_fd_sc_hd__nor4_1 U31153 ( .A(n25889), .B(n25888), .C(n25905), .D(
        n25887), .Y(n25893) );
  sky130_fd_sc_hd__nand2_1 U31154 ( .A(n25958), .B(n25891), .Y(n25986) );
  sky130_fd_sc_hd__nand2_1 U31156 ( .A(n25893), .B(n25892), .Y(n25894) );
  sky130_fd_sc_hd__a31oi_1 U31157 ( .A1(n26250), .A2(n26009), .A3(
        j202_soc_core_wbqspiflash_00_state[2]), .B1(n25894), .Y(n25895) );
  sky130_fd_sc_hd__o22ai_1 U31158 ( .A1(n25896), .A2(n25993), .B1(n28590), 
        .B2(n25895), .Y(j202_soc_core_wbqspiflash_00_N727) );
  sky130_fd_sc_hd__nand3_1 U31159 ( .A(n25898), .B(n28207), .C(n25973), .Y(
        n25899) );
  sky130_fd_sc_hd__and4_1 U31160 ( .A(n25901), .B(n26050), .C(n25900), .D(
        n25899), .X(n25903) );
  sky130_fd_sc_hd__nor2_1 U31161 ( .A(n26014), .B(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled), .Y(n26034) );
  sky130_fd_sc_hd__a21oi_1 U31162 ( .A1(n28230), .A2(n26034), .B1(n26185), .Y(
        n25902) );
  sky130_fd_sc_hd__a31oi_1 U31163 ( .A1(n25903), .A2(n25902), .A3(n28083), 
        .B1(n28590), .Y(j202_soc_core_wbqspiflash_00_N737) );
  sky130_fd_sc_hd__nand2_1 U31164 ( .A(n26191), .B(n26255), .Y(n28098) );
  sky130_fd_sc_hd__nand3_1 U31165 ( .A(n28098), .B(n28187), .C(n28217), .Y(
        n26123) );
  sky130_fd_sc_hd__nand3_1 U31166 ( .A(n26042), .B(n28058), .C(
        j202_soc_core_wbqspiflash_00_state[4]), .Y(n28208) );
  sky130_fd_sc_hd__nand2_1 U31167 ( .A(n25996), .B(
        j202_soc_core_wbqspiflash_00_state[2]), .Y(n26173) );
  sky130_fd_sc_hd__nand2_1 U31168 ( .A(n28100), .B(n28067), .Y(n25904) );
  sky130_fd_sc_hd__nand2_1 U31169 ( .A(n26173), .B(n25904), .Y(n26027) );
  sky130_fd_sc_hd__nor2_1 U31170 ( .A(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled), .B(n28115), .Y(n25912) );
  sky130_fd_sc_hd__nor2_1 U31171 ( .A(n28222), .B(n25988), .Y(n26011) );
  sky130_fd_sc_hd__nand2_1 U31172 ( .A(n26188), .B(n26189), .Y(n28212) );
  sky130_fd_sc_hd__o21ai_1 U31173 ( .A1(n28089), .A2(n25924), .B1(n28212), .Y(
        n25909) );
  sky130_fd_sc_hd__nand2_1 U31174 ( .A(n28237), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .Y(n28252) );
  sky130_fd_sc_hd__nor2_1 U31175 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .B(n28252), .Y(n25969)
         );
  sky130_fd_sc_hd__a21oi_1 U31176 ( .A1(n28207), .A2(n25973), .B1(n25969), .Y(
        n25960) );
  sky130_fd_sc_hd__nand2_1 U31177 ( .A(io_out[8]), .B(n25944), .Y(n26140) );
  sky130_fd_sc_hd__nor3_1 U31178 ( .A(n25960), .B(n28208), .C(n26140), .Y(
        n25908) );
  sky130_fd_sc_hd__nand2_1 U31179 ( .A(n25955), .B(n26042), .Y(n25985) );
  sky130_fd_sc_hd__nand3_1 U31180 ( .A(n25906), .B(n26165), .C(n28236), .Y(
        n26020) );
  sky130_fd_sc_hd__nor2_1 U31181 ( .A(j202_soc_core_wbqspiflash_00_state[1]), 
        .B(n26020), .Y(n25907) );
  sky130_fd_sc_hd__nor4_1 U31182 ( .A(n28099), .B(n25909), .C(n25908), .D(
        n25907), .Y(n25910) );
  sky130_fd_sc_hd__o21ai_1 U31183 ( .A1(n26011), .A2(n28213), .B1(n25910), .Y(
        n25911) );
  sky130_fd_sc_hd__nor4_1 U31184 ( .A(n26123), .B(n26027), .C(n25912), .D(
        n25911), .Y(n25913) );
  sky130_fd_sc_hd__nor2_1 U31185 ( .A(n28590), .B(n25913), .Y(
        j202_soc_core_wbqspiflash_00_N736) );
  sky130_fd_sc_hd__nor2_1 U31186 ( .A(n26000), .B(n26250), .Y(n25947) );
  sky130_fd_sc_hd__nand2_1 U31187 ( .A(n28080), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n25914) );
  sky130_fd_sc_hd__o22ai_1 U31188 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), 
        .A2(j202_soc_core_wbqspiflash_00_state[2]), .B1(io_out[8]), .B2(n25914), .Y(n25915) );
  sky130_fd_sc_hd__a22oi_1 U31189 ( .A1(n25916), .A2(n25915), .B1(
        j202_soc_core_wbqspiflash_00_spi_spd), .B2(n28260), .Y(n25919) );
  sky130_fd_sc_hd__nor3_1 U31190 ( .A(j202_soc_core_wbqspiflash_00_spi_in[28]), 
        .B(j202_soc_core_wbqspiflash_00_spi_in[30]), .C(n28268), .Y(n25917) );
  sky130_fd_sc_hd__nand4_1 U31191 ( .A(n28080), .B(n26009), .C(
        j202_soc_core_wbqspiflash_00_spi_in[29]), .D(n25917), .Y(n25918) );
  sky130_fd_sc_hd__nand3_1 U31192 ( .A(n25919), .B(n28108), .C(n25918), .Y(
        n25945) );
  sky130_fd_sc_hd__nor2_1 U31193 ( .A(n25921), .B(n26115), .Y(n26137) );
  sky130_fd_sc_hd__nor2_1 U31195 ( .A(n25982), .B(n26122), .Y(n25922) );
  sky130_fd_sc_hd__nor2_1 U31196 ( .A(n25922), .B(n25921), .Y(n25923) );
  sky130_fd_sc_hd__nor3_1 U31197 ( .A(n28590), .B(n26137), .C(n25923), .Y(
        n25925) );
  sky130_fd_sc_hd__o211ai_1 U31198 ( .A1(n25944), .A2(n28232), .B1(n25925), 
        .C1(n25924), .Y(n25934) );
  sky130_fd_sc_hd__nand2_1 U31199 ( .A(n26244), .B(j202_soc_core_qspi_wb_cyc), 
        .Y(n26243) );
  sky130_fd_sc_hd__o22ai_1 U31200 ( .A1(n28063), .A2(n26183), .B1(n26128), 
        .B2(n26242), .Y(n25933) );
  sky130_fd_sc_hd__nand2_1 U31201 ( .A(n26189), .B(n26255), .Y(n25927) );
  sky130_fd_sc_hd__nand2_1 U31202 ( .A(n25926), .B(n25980), .Y(n25957) );
  sky130_fd_sc_hd__nand3_1 U31203 ( .A(n28229), .B(
        j202_soc_core_wbqspiflash_00_state[1]), .C(
        j202_soc_core_wbqspiflash_00_state[4]), .Y(n25999) );
  sky130_fd_sc_hd__a31oi_1 U31204 ( .A1(n25927), .A2(n25957), .A3(n25999), 
        .B1(n26167), .Y(n25932) );
  sky130_fd_sc_hd__nor2_1 U31205 ( .A(n25928), .B(n26007), .Y(n28066) );
  sky130_fd_sc_hd__nor2_1 U31206 ( .A(j202_soc_core_wbqspiflash_00_spi_len[0]), 
        .B(j202_soc_core_wbqspiflash_00_spi_len[1]), .Y(n26217) );
  sky130_fd_sc_hd__a21oi_1 U31207 ( .A1(n26217), .A2(
        j202_soc_core_wbqspiflash_00_spi_valid), .B1(n25929), .Y(n26120) );
  sky130_fd_sc_hd__nor2_1 U31208 ( .A(n26120), .B(n28103), .Y(n25930) );
  sky130_fd_sc_hd__o22ai_1 U31209 ( .A1(n26198), .A2(n26114), .B1(n25930), 
        .B2(n26140), .Y(n25931) );
  sky130_fd_sc_hd__nor4_1 U31210 ( .A(n25934), .B(n25933), .C(n25932), .D(
        n25931), .Y(n25942) );
  sky130_fd_sc_hd__nor2_1 U31211 ( .A(n26476), .B(n28083), .Y(n25936) );
  sky130_fd_sc_hd__nor3_1 U31212 ( .A(j202_soc_core_wbqspiflash_00_spi_busy), 
        .B(io_out[8]), .C(n28098), .Y(n25935) );
  sky130_fd_sc_hd__nand2_1 U31213 ( .A(j202_soc_core_wbqspiflash_00_spi_len[1]), .B(j202_soc_core_wbqspiflash_00_spi_len[0]), .Y(n26232) );
  sky130_fd_sc_hd__o21ai_1 U31214 ( .A1(n25936), .A2(n25935), .B1(n26227), .Y(
        n25940) );
  sky130_fd_sc_hd__nor3_1 U31215 ( .A(j202_soc_core_qspi_wb_addr[2]), .B(
        n26171), .C(n26029), .Y(n25937) );
  sky130_fd_sc_hd__nand4_1 U31217 ( .A(n25942), .B(n25941), .C(n25940), .D(
        n25939), .Y(n25943) );
  sky130_fd_sc_hd__a21oi_1 U31218 ( .A1(n25945), .A2(n25944), .B1(n25943), .Y(
        n25946) );
  sky130_fd_sc_hd__o21ai_1 U31219 ( .A1(n26251), .A2(n25947), .B1(n25946), .Y(
        j202_soc_core_wbqspiflash_00_N723) );
  sky130_fd_sc_hd__nor2_1 U31220 ( .A(n28590), .B(n26155), .Y(n26477) );
  sky130_fd_sc_hd__o22ai_1 U31221 ( .A1(
        j202_soc_core_wbqspiflash_00_spif_data[28]), .A2(n28086), .B1(n29054), 
        .B2(n26477), .Y(j202_soc_core_wbqspiflash_00_N722) );
  sky130_fd_sc_hd__nand2_1 U31222 ( .A(n28249), .B(n25948), .Y(n26144) );
  sky130_fd_sc_hd__a31oi_1 U31223 ( .A1(n26155), .A2(n26147), .A3(n25949), 
        .B1(n28590), .Y(n25950) );
  sky130_fd_sc_hd__o31ai_1 U31224 ( .A1(n27040), .A2(n25951), .A3(n26144), 
        .B1(n25950), .Y(j202_soc_core_wbqspiflash_00_N721) );
  sky130_fd_sc_hd__nor2_1 U31225 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[5]), .B(
        j202_soc_core_wbqspiflash_00_spif_data[6]), .Y(n25952) );
  sky130_fd_sc_hd__o21ai_1 U31226 ( .A1(
        j202_soc_core_wbqspiflash_00_last_status[5]), .A2(
        j202_soc_core_wbqspiflash_00_last_status[6]), .B1(n25952), .Y(n25994)
         );
  sky130_fd_sc_hd__o211ai_1 U31227 ( .A1(n25955), .A2(n25994), .B1(n25954), 
        .C1(n25953), .Y(n25956) );
  sky130_fd_sc_hd__nand4_1 U31228 ( .A(n26050), .B(n26251), .C(n25957), .D(
        n25956), .Y(n25979) );
  sky130_fd_sc_hd__a31oi_1 U31229 ( .A1(
        j202_soc_core_wbqspiflash_00_write_in_progress), .A2(n26017), .A3(
        n26467), .B1(n25985), .Y(n25959) );
  sky130_fd_sc_hd__nand2_1 U31230 ( .A(n25959), .B(n25958), .Y(n25968) );
  sky130_fd_sc_hd__nor2_1 U31231 ( .A(n26255), .B(n28243), .Y(n26048) );
  sky130_fd_sc_hd__nand3_1 U31232 ( .A(n25960), .B(n26048), .C(n28058), .Y(
        n25967) );
  sky130_fd_sc_hd__nor2_1 U31234 ( .A(n26127), .B(n26128), .Y(n26021) );
  sky130_fd_sc_hd__clkinv_1 U31235 ( .A(n26021), .Y(n25962) );
  sky130_fd_sc_hd__a21oi_1 U31236 ( .A1(n26035), .A2(n25962), .B1(n26007), .Y(
        n25964) );
  sky130_fd_sc_hd__nor2_1 U31237 ( .A(j202_soc_core_wbqspiflash_00_state[4]), 
        .B(j202_soc_core_wbqspiflash_00_state[3]), .Y(n25963) );
  sky130_fd_sc_hd__nand3b_1 U31238 ( .A_N(n28231), .B(n28229), .C(n25963), .Y(
        n28211) );
  sky130_fd_sc_hd__nor2_1 U31239 ( .A(n25984), .B(n28211), .Y(n28261) );
  sky130_fd_sc_hd__nor3_1 U31240 ( .A(n25965), .B(n25964), .C(n28261), .Y(
        n25966) );
  sky130_fd_sc_hd__o211ai_1 U31241 ( .A1(n25969), .A2(n25968), .B1(n25967), 
        .C1(n25966), .Y(n25978) );
  sky130_fd_sc_hd__nor2_1 U31242 ( .A(
        j202_soc_core_wbqspiflash_00_write_protect), .B(n10959), .Y(n25970) );
  sky130_fd_sc_hd__and3_1 U31243 ( .A(n26149), .B(n25970), .C(n26171), .X(
        n26033) );
  sky130_fd_sc_hd__a21oi_1 U31244 ( .A1(n28116), .A2(n25971), .B1(n26012), .Y(
        n25975) );
  sky130_fd_sc_hd__o22ai_1 U31245 ( .A1(n26029), .A2(n26154), .B1(n25973), 
        .B2(n26014), .Y(n25974) );
  sky130_fd_sc_hd__nor3_1 U31246 ( .A(n26033), .B(n25975), .C(n25974), .Y(
        n25976) );
  sky130_fd_sc_hd__nor2_1 U31247 ( .A(n25976), .B(n26013), .Y(n25977) );
  sky130_fd_sc_hd__o31a_1 U31248 ( .A1(n25979), .A2(n25978), .A3(n25977), .B1(
        n29593), .X(j202_soc_core_wbqspiflash_00_N725) );
  sky130_fd_sc_hd__nor2_1 U31249 ( .A(n25980), .B(n26174), .Y(n25981) );
  sky130_fd_sc_hd__nor2_1 U31250 ( .A(n25982), .B(n25981), .Y(n28551) );
  sky130_fd_sc_hd__nand2_1 U31251 ( .A(n28199), .B(
        j202_soc_core_wbqspiflash_00_spif_data[6]), .Y(n28196) );
  sky130_fd_sc_hd__o21ai_1 U31252 ( .A1(n27549), .A2(n28551), .B1(n28196), .Y(
        j202_soc_core_wbqspiflash_00_N612) );
  sky130_fd_sc_hd__o21ai_1 U31253 ( .A1(n28590), .A2(n26114), .B1(n25983), .Y(
        j202_soc_core_wbqspiflash_00_N750) );
  sky130_fd_sc_hd__nand2_1 U31254 ( .A(n28199), .B(
        j202_soc_core_wbqspiflash_00_spif_data[5]), .Y(n28190) );
  sky130_fd_sc_hd__o21ai_1 U31255 ( .A1(n26945), .A2(n28551), .B1(n28190), .Y(
        j202_soc_core_wbqspiflash_00_N611) );
  sky130_fd_sc_hd__nand2b_1 U31256 ( .A_N(n25985), .B(n25984), .Y(n28235) );
  sky130_fd_sc_hd__a21oi_1 U31257 ( .A1(n26017), .A2(n26467), .B1(n25986), .Y(
        n25987) );
  sky130_fd_sc_hd__nor2_1 U31258 ( .A(n28235), .B(n25987), .Y(n26005) );
  sky130_fd_sc_hd__a21oi_1 U31259 ( .A1(n26149), .A2(
        j202_soc_core_wbqspiflash_00_write_in_progress), .B1(n25988), .Y(
        n25990) );
  sky130_fd_sc_hd__nand2_1 U31260 ( .A(n26173), .B(n26174), .Y(n26247) );
  sky130_fd_sc_hd__nand2b_1 U31262 ( .A_N(n25993), .B(n25992), .Y(n28245) );
  sky130_fd_sc_hd__nand2_1 U31263 ( .A(n28199), .B(n25995), .Y(n25998) );
  sky130_fd_sc_hd__nand2_1 U31264 ( .A(n25996), .B(n26017), .Y(n25997) );
  sky130_fd_sc_hd__nand4_1 U31265 ( .A(n28245), .B(n25999), .C(n25998), .D(
        n25997), .Y(n26003) );
  sky130_fd_sc_hd__nand4_1 U31266 ( .A(n26042), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .C(j202_soc_core_qspi_wb_cyc), 
        .D(j202_soc_core_wbqspiflash_00_state[4]), .Y(n26001) );
  sky130_fd_sc_hd__nor2_1 U31267 ( .A(n26001), .B(n26124), .Y(n26002) );
  sky130_fd_sc_hd__nor4_1 U31268 ( .A(n26005), .B(n26004), .C(n26003), .D(
        n26002), .Y(n26006) );
  sky130_fd_sc_hd__nor2_1 U31269 ( .A(n28590), .B(n26006), .Y(
        j202_soc_core_wbqspiflash_00_N728) );
  sky130_fd_sc_hd__nor2_1 U31270 ( .A(n26255), .B(n26007), .Y(n26051) );
  sky130_fd_sc_hd__o31ai_1 U31272 ( .A1(n26012), .A2(n26011), .A3(n26013), 
        .B1(n26010), .Y(n26026) );
  sky130_fd_sc_hd__nand2_1 U31273 ( .A(n26016), .B(n26015), .Y(n28123) );
  sky130_fd_sc_hd__nand3_1 U31274 ( .A(n26018), .B(n28251), .C(n26048), .Y(
        n26019) );
  sky130_fd_sc_hd__nand3_1 U31275 ( .A(n28123), .B(n26020), .C(n26019), .Y(
        n26025) );
  sky130_fd_sc_hd__a31oi_1 U31276 ( .A1(n26053), .A2(n26021), .A3(n28110), 
        .B1(n26191), .Y(n26023) );
  sky130_fd_sc_hd__nand3_1 U31277 ( .A(n26023), .B(n26050), .C(n26022), .Y(
        n26024) );
  sky130_fd_sc_hd__nor4_1 U31278 ( .A(n26027), .B(n26026), .C(n26025), .D(
        n26024), .Y(n26028) );
  sky130_fd_sc_hd__nor2_1 U31279 ( .A(n28590), .B(n26028), .Y(
        j202_soc_core_wbqspiflash_00_N726) );
  sky130_fd_sc_hd__nand3_1 U31280 ( .A(n26030), .B(n28106), .C(n26171), .Y(
        n26038) );
  sky130_fd_sc_hd__nand2_1 U31281 ( .A(n28106), .B(
        j202_soc_core_qspi_wb_addr[2]), .Y(n26031) );
  sky130_fd_sc_hd__mux2i_1 U31282 ( .A0(n26147), .A1(n26032), .S(n26031), .Y(
        n26037) );
  sky130_fd_sc_hd__nor2_1 U31283 ( .A(n26034), .B(n26033), .Y(n26036) );
  sky130_fd_sc_hd__nand2_1 U31284 ( .A(n26035), .B(n28058), .Y(n28224) );
  sky130_fd_sc_hd__a31oi_1 U31285 ( .A1(n26038), .A2(n26037), .A3(n26036), 
        .B1(n28224), .Y(n26045) );
  sky130_fd_sc_hd__a211oi_1 U31286 ( .A1(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled), .A2(n28207), .B1(
        j202_soc_core_wbqspiflash_00_state[0]), .C1(n26039), .Y(n26044) );
  sky130_fd_sc_hd__a21oi_1 U31287 ( .A1(n26041), .A2(n28252), .B1(n26040), .Y(
        n26043) );
  sky130_fd_sc_hd__o31ai_1 U31288 ( .A1(n26045), .A2(n26044), .A3(n26043), 
        .B1(n26042), .Y(n26058) );
  sky130_fd_sc_hd__nor2_1 U31289 ( .A(n26046), .B(n28224), .Y(n26047) );
  sky130_fd_sc_hd__a31oi_1 U31290 ( .A1(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled), .A2(n28229), .A3(
        n26048), .B1(n26047), .Y(n26057) );
  sky130_fd_sc_hd__nor4_1 U31291 ( .A(n26052), .B(n28119), .C(n26051), .D(
        n28261), .Y(n26056) );
  sky130_fd_sc_hd__nor2_1 U31292 ( .A(n26128), .B(
        j202_soc_core_wbqspiflash_00_spi_spd), .Y(n26054) );
  sky130_fd_sc_hd__nand4_1 U31294 ( .A(n26058), .B(n26057), .C(n26056), .D(
        n26055), .Y(n26059) );
  sky130_fd_sc_hd__a31oi_1 U31295 ( .A1(n26250), .A2(n28079), .A3(n26161), 
        .B1(n26059), .Y(n26060) );
  sky130_fd_sc_hd__nor2_1 U31296 ( .A(n28590), .B(n26060), .Y(
        j202_soc_core_wbqspiflash_00_N724) );
  sky130_fd_sc_hd__a22oi_1 U31297 ( .A1(n27184), .A2(n26061), .B1(n11589), 
        .B2(n27339), .Y(n26062) );
  sky130_fd_sc_hd__nand2_1 U31298 ( .A(n27346), .B(n26062), .Y(
        j202_soc_core_j22_cpu_ml_N327) );
  sky130_fd_sc_hd__a22oi_1 U31299 ( .A1(n27187), .A2(n22029), .B1(n27273), 
        .B2(n26068), .Y(n26063) );
  sky130_fd_sc_hd__nand2_1 U31300 ( .A(n27189), .B(n26063), .Y(
        j202_soc_core_j22_cpu_ml_machj[23]) );
  sky130_fd_sc_hd__o22ai_1 U31301 ( .A1(n27575), .A2(n27401), .B1(n27574), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N3111) );
  sky130_fd_sc_hd__nand2_1 U31302 ( .A(n11589), .B(n27460), .Y(n26065) );
  sky130_fd_sc_hd__o22ai_1 U31304 ( .A1(n27401), .A2(n26899), .B1(n26898), 
        .B2(n26066), .Y(j202_soc_core_j22_cpu_rf_N3335) );
  sky130_fd_sc_hd__nand2_1 U31305 ( .A(n26068), .B(n26067), .Y(n26075) );
  sky130_fd_sc_hd__o22ai_1 U31306 ( .A1(n26071), .A2(n26070), .B1(n25714), 
        .B2(n27401), .Y(n26072) );
  sky130_fd_sc_hd__a21oi_1 U31307 ( .A1(n26073), .A2(n26516), .B1(n26072), .Y(
        n26074) );
  sky130_fd_sc_hd__nand2_1 U31308 ( .A(n26075), .B(n26074), .Y(
        j202_soc_core_j22_cpu_rf_N3370) );
  sky130_fd_sc_hd__nand2_1 U31309 ( .A(n26510), .B(n26802), .Y(n26103) );
  sky130_fd_sc_hd__o21ai_1 U31310 ( .A1(n26406), .A2(n26508), .B1(n26405), .Y(
        n26076) );
  sky130_fd_sc_hd__nand2_1 U31311 ( .A(n26076), .B(n26407), .Y(n26098) );
  sky130_fd_sc_hd__nand2_1 U31312 ( .A(n26082), .B(n26703), .Y(n26655) );
  sky130_fd_sc_hd__nand2_1 U31313 ( .A(n27405), .B(n26508), .Y(n26656) );
  sky130_fd_sc_hd__nand3_1 U31314 ( .A(n26655), .B(n26326), .C(n26656), .Y(
        n26079) );
  sky130_fd_sc_hd__nand2_1 U31315 ( .A(n26077), .B(n26716), .Y(n26078) );
  sky130_fd_sc_hd__o211ai_1 U31316 ( .A1(n11145), .A2(n26425), .B1(n26079), 
        .C1(n26078), .Y(n26081) );
  sky130_fd_sc_hd__o22ai_1 U31317 ( .A1(n26417), .A2(n26419), .B1(n26701), 
        .B2(n26418), .Y(n26080) );
  sky130_fd_sc_hd__nor2_1 U31318 ( .A(n26081), .B(n26080), .Y(n26092) );
  sky130_fd_sc_hd__o22a_1 U31319 ( .A1(n26082), .A2(n26431), .B1(n11977), .B2(
        n26412), .X(n26091) );
  sky130_fd_sc_hd__o22ai_1 U31320 ( .A1(n18916), .A2(n26083), .B1(n26423), 
        .B2(n27405), .Y(n26084) );
  sky130_fd_sc_hd__a21oi_1 U31321 ( .A1(n26085), .A2(n26508), .B1(n26084), .Y(
        n26086) );
  sky130_fd_sc_hd__o21ai_0 U31322 ( .A1(n26432), .A2(n26656), .B1(n26086), .Y(
        n26089) );
  sky130_fd_sc_hd__nor2_1 U31323 ( .A(n26704), .B(n26424), .Y(n26088) );
  sky130_fd_sc_hd__o22ai_1 U31324 ( .A1(n26565), .A2(n26416), .B1(n26570), 
        .B2(n26427), .Y(n26087) );
  sky130_fd_sc_hd__nor3_1 U31325 ( .A(n26089), .B(n26088), .C(n26087), .Y(
        n26090) );
  sky130_fd_sc_hd__nand4_1 U31326 ( .A(n26092), .B(n26091), .C(n26411), .D(
        n26090), .Y(n26095) );
  sky130_fd_sc_hd__nor2_1 U31327 ( .A(n18916), .B(n26093), .Y(n26094) );
  sky130_fd_sc_hd__a211oi_1 U31328 ( .A1(n26096), .A2(n26409), .B1(n26095), 
        .C1(n26094), .Y(n26097) );
  sky130_fd_sc_hd__a21boi_1 U31329 ( .A1(n26507), .A2(n26098), .B1_N(n26097), 
        .Y(n26099) );
  sky130_fd_sc_hd__nand2_1 U31330 ( .A(n26105), .B(n27192), .Y(n26104) );
  sky130_fd_sc_hd__o22ai_1 U31332 ( .A1(n27407), .A2(n26899), .B1(n26898), 
        .B2(n12391), .Y(j202_soc_core_j22_cpu_rf_N3334) );
  sky130_fd_sc_hd__o22ai_1 U31333 ( .A1(n26378), .A2(n27407), .B1(n26449), 
        .B2(n12391), .Y(j202_soc_core_j22_cpu_rf_N3258) );
  sky130_fd_sc_hd__o22ai_1 U31334 ( .A1(n11141), .A2(n27407), .B1(n27124), 
        .B2(n12391), .Y(j202_soc_core_j22_cpu_rf_N2703) );
  sky130_fd_sc_hd__nand4_1 U31335 ( .A(n26108), .B(n11464), .C(n26107), .D(
        n26106), .Y(n26110) );
  sky130_fd_sc_hd__a21oi_1 U31336 ( .A1(n11464), .A2(n29535), .B1(n26951), .Y(
        n26109) );
  sky130_fd_sc_hd__nand2_1 U31337 ( .A(n26110), .B(n26109), .Y(n26113) );
  sky130_fd_sc_hd__a22oi_1 U31338 ( .A1(n26111), .A2(n26948), .B1(n26507), 
        .B2(n24650), .Y(n26112) );
  sky130_fd_sc_hd__nand2_1 U31339 ( .A(n26113), .B(n26112), .Y(
        j202_soc_core_j22_cpu_rf_N3369) );
  sky130_fd_sc_hd__o22ai_1 U31340 ( .A1(n27575), .A2(n27407), .B1(n27574), 
        .B2(n12391), .Y(j202_soc_core_j22_cpu_rf_N3110) );
  sky130_fd_sc_hd__o22ai_1 U31341 ( .A1(n27333), .A2(n27407), .B1(n23178), 
        .B2(n12392), .Y(j202_soc_core_j22_cpu_rf_N3073) );
  sky130_fd_sc_hd__o22ai_1 U31342 ( .A1(n27219), .A2(n27407), .B1(n27218), 
        .B2(n12392), .Y(j202_soc_core_j22_cpu_rf_N2999) );
  sky130_fd_sc_hd__o22ai_1 U31343 ( .A1(n27217), .A2(n27407), .B1(n27216), 
        .B2(n12391), .Y(j202_soc_core_j22_cpu_rf_N2851) );
  sky130_fd_sc_hd__o22ai_1 U31344 ( .A1(n27228), .A2(n27407), .B1(n27227), 
        .B2(n12392), .Y(j202_soc_core_j22_cpu_rf_N3184) );
  sky130_fd_sc_hd__o22ai_1 U31345 ( .A1(n27225), .A2(n27407), .B1(n27224), 
        .B2(n12392), .Y(j202_soc_core_j22_cpu_rf_N2962) );
  sky130_fd_sc_hd__o22ai_1 U31346 ( .A1(n27215), .A2(n27407), .B1(n27214), 
        .B2(n12391), .Y(j202_soc_core_j22_cpu_rf_N2925) );
  sky130_fd_sc_hd__o22ai_1 U31347 ( .A1(n27223), .A2(n27407), .B1(n27222), 
        .B2(n12392), .Y(j202_soc_core_j22_cpu_rf_N3036) );
  sky130_fd_sc_hd__o22ai_1 U31348 ( .A1(n27211), .A2(n27407), .B1(n27210), 
        .B2(n12392), .Y(j202_soc_core_j22_cpu_rf_N3221) );
  sky130_fd_sc_hd__o22ai_1 U31349 ( .A1(n27221), .A2(n27407), .B1(n27220), 
        .B2(n12392), .Y(j202_soc_core_j22_cpu_rf_N2888) );
  sky130_fd_sc_hd__o22ai_1 U31350 ( .A1(n27226), .A2(n27407), .B1(n23079), 
        .B2(n12391), .Y(j202_soc_core_j22_cpu_rf_N3147) );
  sky130_fd_sc_hd__o22ai_1 U31351 ( .A1(n27213), .A2(n27407), .B1(n27212), 
        .B2(n12392), .Y(j202_soc_core_j22_cpu_rf_N2814) );
  sky130_fd_sc_hd__o22ai_1 U31352 ( .A1(n27209), .A2(n27407), .B1(n23039), 
        .B2(n12392), .Y(j202_soc_core_j22_cpu_rf_N2740) );
  sky130_fd_sc_hd__nand2_1 U31353 ( .A(n26114), .B(n28232), .Y(n26163) );
  sky130_fd_sc_hd__o22ai_1 U31355 ( .A1(j202_soc_core_wbqspiflash_00_spi_valid), .A2(n27039), .B1(n26116), .B2(n26115), .Y(n26117) );
  sky130_fd_sc_hd__or4_1 U31356 ( .A(n26120), .B(n26119), .C(n26118), .D(
        n26117), .X(n26121) );
  sky130_fd_sc_hd__nor4_1 U31357 ( .A(n26123), .B(n26163), .C(n26122), .D(
        n26121), .Y(n26126) );
  sky130_fd_sc_hd__o22ai_1 U31358 ( .A1(n26126), .A2(n26125), .B1(n26251), 
        .B2(n26124), .Y(n26133) );
  sky130_fd_sc_hd__a21oi_1 U31359 ( .A1(n26128), .A2(
        j202_soc_core_wbqspiflash_00_spif_req), .B1(n26127), .Y(n26129) );
  sky130_fd_sc_hd__o22ai_1 U31360 ( .A1(n26131), .A2(n26130), .B1(n26242), 
        .B2(n26129), .Y(n26132) );
  sky130_fd_sc_hd__a21o_1 U31361 ( .A1(n26133), .A2(j202_soc_core_qspi_wb_cyc), 
        .B1(n26132), .X(n10505) );
  sky130_fd_sc_hd__a21oi_1 U31362 ( .A1(n27040), .A2(n26135), .B1(n26134), .Y(
        n26136) );
  sky130_fd_sc_hd__a21oi_1 U31363 ( .A1(j202_soc_core_wbqspiflash_00_spif_cmd), 
        .A2(j202_soc_core_wbqspiflash_00_write_protect), .B1(n26136), .Y(
        n26145) );
  sky130_fd_sc_hd__a21oi_1 U31364 ( .A1(n26138), .A2(n28119), .B1(n26137), .Y(
        n26139) );
  sky130_fd_sc_hd__o31a_1 U31365 ( .A1(n26141), .A2(n26140), .A3(n28250), .B1(
        n26139), .X(n26143) );
  sky130_fd_sc_hd__o211ai_1 U31366 ( .A1(n26145), .A2(n26144), .B1(n26143), 
        .C1(n26142), .Y(n26146) );
  sky130_fd_sc_hd__nand3_1 U31367 ( .A(n26146), .B(
        j202_soc_core_wbqspiflash_00_spif_req), .C(n29593), .Y(n26160) );
  sky130_fd_sc_hd__a21oi_1 U31368 ( .A1(n29593), .A2(n26148), .B1(n29055), .Y(
        n26151) );
  sky130_fd_sc_hd__nand4_1 U31369 ( .A(n26149), .B(n10958), .C(
        j202_soc_core_wbqspiflash_00_write_protect), .D(n12142), .Y(n26150) );
  sky130_fd_sc_hd__a211oi_1 U31371 ( .A1(n26154), .A2(n10959), .B1(n10539), 
        .C1(n26153), .Y(n26156) );
  sky130_fd_sc_hd__o21ai_1 U31372 ( .A1(n26157), .A2(n26156), .B1(n26155), .Y(
        n26158) );
  sky130_fd_sc_hd__nand3_1 U31373 ( .A(n26160), .B(n26159), .C(n26158), .Y(
        j202_soc_core_wbqspiflash_00_N730) );
  sky130_fd_sc_hd__nand2_1 U31374 ( .A(n26161), .B(n29594), .Y(n26475) );
  sky130_fd_sc_hd__nand2_1 U31375 ( .A(n26163), .B(n26162), .Y(
        j202_soc_core_wbqspiflash_00_N729) );
  sky130_fd_sc_hd__a21oi_1 U31376 ( .A1(n26165), .A2(n26164), .B1(n26191), .Y(
        n26166) );
  sky130_fd_sc_hd__nor2_1 U31377 ( .A(n26167), .B(n26166), .Y(n26168) );
  sky130_fd_sc_hd__nor3_1 U31378 ( .A(n26170), .B(n26169), .C(n26168), .Y(
        n26179) );
  sky130_fd_sc_hd__a211oi_1 U31379 ( .A1(j202_soc_core_ahb2wbqspi_00_stb_o), 
        .A2(j202_soc_core_qspi_wb_cyc), .B1(n26171), .C1(n28096), .Y(n26172)
         );
  sky130_fd_sc_hd__a211oi_1 U31380 ( .A1(n28100), .A2(n26248), .B1(n28066), 
        .C1(n26172), .Y(n26178) );
  sky130_fd_sc_hd__nor3_1 U31381 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(j202_soc_core_wbqspiflash_00_spi_busy), .C(n26174), .Y(n26176) );
  sky130_fd_sc_hd__nor4_1 U31382 ( .A(n28234), .B(n26176), .C(n26175), .D(
        n28248), .Y(n26177) );
  sky130_fd_sc_hd__nand4_1 U31383 ( .A(n26179), .B(n26178), .C(n26177), .D(
        n28098), .Y(n26180) );
  sky130_fd_sc_hd__a31oi_1 U31384 ( .A1(n26181), .A2(n28099), .A3(n28089), 
        .B1(n26180), .Y(n26182) );
  sky130_fd_sc_hd__nor2_1 U31385 ( .A(n28590), .B(n26182), .Y(
        j202_soc_core_wbqspiflash_00_N734) );
  sky130_fd_sc_hd__nand3_1 U31386 ( .A(n26184), .B(n29593), .C(n26183), .Y(
        j202_soc_core_wbqspiflash_00_N733) );
  sky130_fd_sc_hd__nand3_1 U31387 ( .A(n26185), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .C(
        j202_soc_core_wbqspiflash_00_spi_busy), .Y(n26186) );
  sky130_fd_sc_hd__nand2_1 U31389 ( .A(n26188), .B(
        j202_soc_core_wbqspiflash_00_spi_busy), .Y(n26257) );
  sky130_fd_sc_hd__a21oi_1 U31390 ( .A1(n26189), .A2(n26257), .B1(n28066), .Y(
        n26190) );
  sky130_fd_sc_hd__nand3_1 U31391 ( .A(n28250), .B(n26190), .C(n26252), .Y(
        n26193) );
  sky130_fd_sc_hd__nor3_1 U31392 ( .A(n26193), .B(n26192), .C(n26191), .Y(
        n28102) );
  sky130_fd_sc_hd__a21oi_1 U31393 ( .A1(n28102), .A2(n26195), .B1(n28590), .Y(
        j202_soc_core_wbqspiflash_00_N746) );
  sky130_fd_sc_hd__nand2_1 U31394 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B(n28649), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N423) );
  sky130_fd_sc_hd__nand2_1 U31395 ( .A(n26214), .B(n28110), .Y(n26207) );
  sky130_fd_sc_hd__o211ai_1 U31396 ( .A1(n26197), .A2(n26196), .B1(n26207), 
        .C1(n26205), .Y(j202_soc_core_wbqspiflash_00_lldriver_N425) );
  sky130_fd_sc_hd__nor2_1 U31397 ( .A(n26198), .B(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .Y(n28641) );
  sky130_fd_sc_hd__nor2_1 U31398 ( .A(n26199), .B(n28641), .Y(n26241) );
  sky130_fd_sc_hd__nand2_1 U31399 ( .A(n26241), .B(n26201), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N424) );
  sky130_fd_sc_hd__nor2_1 U31400 ( .A(n28109), .B(n26202), .Y(n28636) );
  sky130_fd_sc_hd__nor2_1 U31401 ( .A(n28109), .B(n26260), .Y(n26234) );
  sky130_fd_sc_hd__nor3_1 U31402 ( .A(n28636), .B(n26203), .C(n26234), .Y(
        DP_OP_1508J1_126_2326_n6) );
  sky130_fd_sc_hd__nand2_1 U31403 ( .A(n26207), .B(n13300), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N426) );
  sky130_fd_sc_hd__nand2_1 U31404 ( .A(U7_RSOP_1495_C3_DATA3_2), .B(n28743), 
        .Y(n26208) );
  sky130_fd_sc_hd__nand3_1 U31405 ( .A(n26208), .B(n26211), .C(n26225), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N427) );
  sky130_fd_sc_hd__nor2_1 U31406 ( .A(n29056), .B(n28743), .Y(n26231) );
  sky130_fd_sc_hd__o22ai_1 U31407 ( .A1(n26211), .A2(
        j202_soc_core_wbqspiflash_00_spi_len[0]), .B1(n26210), .B2(n26209), 
        .Y(n26212) );
  sky130_fd_sc_hd__nor2_1 U31408 ( .A(n26212), .B(DP_OP_1508J1_126_2326_n3), 
        .Y(n26219) );
  sky130_fd_sc_hd__a21oi_1 U31409 ( .A1(DP_OP_1508J1_126_2326_n3), .A2(n26212), 
        .B1(n26219), .Y(n26216) );
  sky130_fd_sc_hd__nor2_1 U31410 ( .A(j202_soc_core_wbqspiflash_00_spi_len[0]), 
        .B(j202_soc_core_wbqspiflash_00_lldriver_N311), .Y(n26213) );
  sky130_fd_sc_hd__a21oi_1 U31411 ( .A1(n26214), .A2(
        j202_soc_core_wbqspiflash_00_spi_len[0]), .B1(n26213), .Y(n26215) );
  sky130_fd_sc_hd__nor2_1 U31413 ( .A(n26217), .B(n26227), .Y(n26218) );
  sky130_fd_sc_hd__nand2_1 U31414 ( .A(n28727), .B(n26218), .Y(n26224) );
  sky130_fd_sc_hd__a22oi_1 U31415 ( .A1(n26218), .A2(n29056), .B1(n28743), 
        .B2(j202_soc_core_wbqspiflash_00_lldriver_spi_len[4]), .Y(n26220) );
  sky130_fd_sc_hd__nand2_1 U31416 ( .A(n26219), .B(n26220), .Y(n26229) );
  sky130_fd_sc_hd__a21oi_1 U31417 ( .A1(n26229), .A2(n26219), .B1(n26231), .Y(
        n26222) );
  sky130_fd_sc_hd__nand2_1 U31418 ( .A(n26229), .B(n26220), .Y(n26221) );
  sky130_fd_sc_hd__nand2_1 U31419 ( .A(n26222), .B(n26221), .Y(n26223) );
  sky130_fd_sc_hd__o211ai_1 U31420 ( .A1(n26226), .A2(n26225), .B1(n26224), 
        .C1(n26223), .Y(j202_soc_core_wbqspiflash_00_lldriver_N429) );
  sky130_fd_sc_hd__a22oi_1 U31421 ( .A1(n26227), .A2(n29056), .B1(n28743), 
        .B2(j202_soc_core_wbqspiflash_00_lldriver_spi_len[5]), .Y(n26228) );
  sky130_fd_sc_hd__xnor2_1 U31422 ( .A(n26229), .B(n26228), .Y(n26230) );
  sky130_fd_sc_hd__o22ai_1 U31423 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .A2(n26232), .B1(n26231), 
        .B2(n26230), .Y(j202_soc_core_wbqspiflash_00_lldriver_N430) );
  sky130_fd_sc_hd__nor4_1 U31424 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[3]), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[4]), .C(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[5]), .D(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[1]), .Y(n26238) );
  sky130_fd_sc_hd__nand2_1 U31425 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[0]), .B(n26233), .Y(
        n26236) );
  sky130_fd_sc_hd__nand2_1 U31426 ( .A(n26234), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[2]), .Y(n26235) );
  sky130_fd_sc_hd__o22ai_1 U31427 ( .A1(n26236), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[2]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[0]), .B2(n26235), .Y(
        n26237) );
  sky130_fd_sc_hd__a21oi_1 U31428 ( .A1(n26238), .A2(n26237), .B1(n28642), .Y(
        n26239) );
  sky130_fd_sc_hd__nand3_1 U31429 ( .A(n26241), .B(n26240), .C(n26239), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N307) );
  sky130_fd_sc_hd__a22oi_1 U31431 ( .A1(n26248), .A2(n26247), .B1(n26246), 
        .B2(n26245), .Y(n26249) );
  sky130_fd_sc_hd__o21ai_1 U31432 ( .A1(n26251), .A2(n26250), .B1(n26249), .Y(
        j202_soc_core_wbqspiflash_00_N590) );
  sky130_fd_sc_hd__a21oi_1 U31434 ( .A1(j202_soc_core_wbqspiflash_00_state[3]), 
        .A2(n26254), .B1(n26253), .Y(n26259) );
  sky130_fd_sc_hd__a21oi_1 U31435 ( .A1(n28229), .A2(n26255), .B1(
        j202_soc_core_wbqspiflash_00_state[1]), .Y(n26256) );
  sky130_fd_sc_hd__a21oi_1 U31437 ( .A1(n26259), .A2(n26258), .B1(n28590), .Y(
        j202_soc_core_wbqspiflash_00_N745) );
  sky130_fd_sc_hd__nor2_1 U31438 ( .A(n26261), .B(n28747), .Y(n28589) );
  sky130_fd_sc_hd__nor2_1 U31439 ( .A(j202_soc_core_wbqspiflash_00_spi_hold), 
        .B(n28748), .Y(n28645) );
  sky130_fd_sc_hd__or4_1 U31440 ( .A(n26262), .B(n28589), .C(n28727), .D(
        n28645), .X(j202_soc_core_wbqspiflash_00_lldriver_N308) );
  sky130_fd_sc_hd__o22ai_1 U31441 ( .A1(n28608), .A2(n27990), .B1(n26263), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U31442 ( .A1(n27757), .A2(n26264), .B1(n28355), 
        .B2(n27754), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U31443 ( .A1(n27583), .A2(n26265), .B1(n28355), 
        .B2(n27581), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U31444 ( .A1(n28541), .A2(n28608), .B1(n26266), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__a22oi_1 U31445 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[12]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[76]), .Y(n26268) );
  sky130_fd_sc_hd__a22oi_1 U31446 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[12]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[12]), .Y(n26267) );
  sky130_fd_sc_hd__nand3_1 U31447 ( .A(n26268), .B(n26267), .C(n27865), .Y(
        n26269) );
  sky130_fd_sc_hd__a21oi_1 U31448 ( .A1(j202_soc_core_intc_core_00_rg_itgt[11]), .A2(n27869), .B1(n26269), .Y(n26273) );
  sky130_fd_sc_hd__a22oi_1 U31449 ( .A1(n27856), .A2(
        j202_soc_core_intc_core_00_rg_itgt[19]), .B1(n27850), .B2(
        j202_soc_core_intc_core_00_rg_itgt[3]), .Y(n26272) );
  sky130_fd_sc_hd__a22oi_1 U31450 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[27]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[108]), .Y(n26271) );
  sky130_fd_sc_hd__nand2_1 U31451 ( .A(n27862), .B(
        j202_soc_core_intc_core_00_rg_ipr[44]), .Y(n26270) );
  sky130_fd_sc_hd__nand4_1 U31452 ( .A(n26273), .B(n26272), .C(n26271), .D(
        n26270), .Y(j202_soc_core_ahb2apb_01_N140) );
  sky130_fd_sc_hd__nand2_1 U31453 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[12]), .Y(n26274) );
  sky130_fd_sc_hd__o21ai_1 U31454 ( .A1(n26275), .A2(n27983), .B1(n26274), .Y(
        n60) );
  sky130_fd_sc_hd__nand2_1 U31455 ( .A(j202_soc_core_cmt_core_00_cnt0[10]), 
        .B(j202_soc_core_cmt_core_00_cnt0[9]), .Y(n26276) );
  sky130_fd_sc_hd__nor2_1 U31456 ( .A(n26276), .B(n26277), .Y(n26282) );
  sky130_fd_sc_hd__a21oi_1 U31457 ( .A1(n26278), .A2(
        j202_soc_core_cmt_core_00_cnt0[9]), .B1(
        j202_soc_core_cmt_core_00_cnt0[10]), .Y(n26280) );
  sky130_fd_sc_hd__a22oi_1 U31458 ( .A1(n27482), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[10]), .B1(n28619), .B2(
        j202_soc_core_cmt_core_00_cnt0[10]), .Y(n26279) );
  sky130_fd_sc_hd__o31ai_1 U31459 ( .A1(n26282), .A2(n26288), .A3(n26280), 
        .B1(n26279), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[10])
         );
  sky130_fd_sc_hd__a21oi_1 U31460 ( .A1(n26281), .A2(n26282), .B1(
        j202_soc_core_cmt_core_00_cnt0[11]), .Y(n26286) );
  sky130_fd_sc_hd__nand2_1 U31461 ( .A(n26282), .B(
        j202_soc_core_cmt_core_00_cnt0[11]), .Y(n26287) );
  sky130_fd_sc_hd__a21oi_1 U31462 ( .A1(n26285), .A2(n26284), .B1(n26283), .Y(
        n27469) );
  sky130_fd_sc_hd__o22ai_1 U31463 ( .A1(n27473), .A2(n27237), .B1(n26286), 
        .B2(n26290), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[11])
         );
  sky130_fd_sc_hd__nor2_1 U31464 ( .A(n26288), .B(n26287), .Y(n27468) );
  sky130_fd_sc_hd__a22oi_1 U31465 ( .A1(n27482), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[12]), .B1(n27468), .B2(n26291), 
        .Y(n26289) );
  sky130_fd_sc_hd__o21ai_1 U31466 ( .A1(n26291), .A2(n26290), .B1(n26289), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[12]) );
  sky130_fd_sc_hd__nand2_1 U31467 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[12]), .Y(n26292) );
  sky130_fd_sc_hd__o21ai_1 U31468 ( .A1(n26307), .A2(n27827), .B1(n26292), .Y(
        n127) );
  sky130_fd_sc_hd__nand2_1 U31469 ( .A(n26293), .B(
        j202_soc_core_cmt_core_00_cnt1[10]), .Y(n26296) );
  sky130_fd_sc_hd__nor3_1 U31470 ( .A(j202_soc_core_cmt_core_00_cnt1[10]), .B(
        n26301), .C(n26298), .Y(n26294) );
  sky130_fd_sc_hd__a21oi_1 U31471 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[10]), .A2(n27498), .B1(n26294), 
        .Y(n26295) );
  sky130_fd_sc_hd__nand2_1 U31472 ( .A(n26296), .B(n26295), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[10]) );
  sky130_fd_sc_hd__a31oi_1 U31473 ( .A1(n26297), .A2(n27489), .A3(
        j202_soc_core_cmt_core_00_cnt1[10]), .B1(
        j202_soc_core_cmt_core_00_cnt1[11]), .Y(n26302) );
  sky130_fd_sc_hd__nand2_1 U31474 ( .A(j202_soc_core_cmt_core_00_cnt1[10]), 
        .B(j202_soc_core_cmt_core_00_cnt1[11]), .Y(n26299) );
  sky130_fd_sc_hd__nor2_1 U31475 ( .A(n26299), .B(n26298), .Y(n27487) );
  sky130_fd_sc_hd__o21ai_1 U31476 ( .A1(n26301), .A2(n27487), .B1(n26300), .Y(
        n27488) );
  sky130_fd_sc_hd__o22ai_1 U31477 ( .A1(n27491), .A2(n27237), .B1(n26302), 
        .B2(n26304), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[11])
         );
  sky130_fd_sc_hd__nand2_1 U31478 ( .A(n27487), .B(n27489), .Y(n27492) );
  sky130_fd_sc_hd__a2bb2oi_1 U31479 ( .B1(n27498), .B2(
        j202_soc_core_cmt_core_00_wdata_cnt0[12]), .A1_N(
        j202_soc_core_cmt_core_00_cnt1[12]), .A2_N(n27492), .Y(n26303) );
  sky130_fd_sc_hd__o21ai_1 U31480 ( .A1(n26305), .A2(n26304), .B1(n26303), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[12]) );
  sky130_fd_sc_hd__nand2_1 U31481 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[12]), .Y(n26306) );
  sky130_fd_sc_hd__o21ai_1 U31482 ( .A1(n26307), .A2(n27833), .B1(n26306), .Y(
        n121) );
  sky130_fd_sc_hd__a22oi_1 U31483 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[12]), .B1(n27837), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[12]), 
        .Y(n26310) );
  sky130_fd_sc_hd__nand2_1 U31484 ( .A(n27840), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[12]), 
        .Y(n26309) );
  sky130_fd_sc_hd__nand2_1 U31485 ( .A(n27835), .B(
        j202_soc_core_cmt_core_00_const1[12]), .Y(n26308) );
  sky130_fd_sc_hd__nand3_1 U31486 ( .A(n26310), .B(n26309), .C(n26308), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[12]) );
  sky130_fd_sc_hd__a31oi_1 U31487 ( .A1(n26319), .A2(n26318), .A3(n26317), 
        .B1(n29535), .Y(n26320) );
  sky130_fd_sc_hd__nand2_1 U31488 ( .A(n26324), .B(n26422), .Y(n26358) );
  sky130_fd_sc_hd__o22ai_1 U31489 ( .A1(n26325), .A2(n26419), .B1(n26565), 
        .B2(n26418), .Y(n26335) );
  sky130_fd_sc_hd__nand2_1 U31490 ( .A(n26413), .B(n26426), .Y(n26664) );
  sky130_fd_sc_hd__nand2_1 U31491 ( .A(n27372), .B(n26709), .Y(n26663) );
  sky130_fd_sc_hd__nand3_1 U31492 ( .A(n26664), .B(n26326), .C(n26663), .Y(
        n26332) );
  sky130_fd_sc_hd__nand2_1 U31493 ( .A(n26328), .B(n26327), .Y(n26330) );
  sky130_fd_sc_hd__nand2_1 U31494 ( .A(n26330), .B(n26329), .Y(n26331) );
  sky130_fd_sc_hd__o211ai_1 U31495 ( .A1(n26417), .A2(n26333), .B1(n26332), 
        .C1(n26331), .Y(n26334) );
  sky130_fd_sc_hd__nor2_1 U31496 ( .A(n26335), .B(n26334), .Y(n26348) );
  sky130_fd_sc_hd__o22ai_1 U31497 ( .A1(n27007), .A2(n26416), .B1(n26336), 
        .B2(n26427), .Y(n26337) );
  sky130_fd_sc_hd__a21oi_1 U31498 ( .A1(n26338), .A2(n27422), .B1(n26337), .Y(
        n26346) );
  sky130_fd_sc_hd__o22a_1 U31499 ( .A1(n26423), .A2(n27372), .B1(n26432), .B2(
        n26663), .X(n26339) );
  sky130_fd_sc_hd__o21ai_0 U31500 ( .A1(n26708), .A2(n26424), .B1(n26339), .Y(
        n26340) );
  sky130_fd_sc_hd__a21oi_1 U31501 ( .A1(n26341), .A2(n26414), .B1(n26340), .Y(
        n26345) );
  sky130_fd_sc_hd__nand2_1 U31502 ( .A(n26342), .B(n27368), .Y(n26343) );
  sky130_fd_sc_hd__and4_1 U31503 ( .A(n26346), .B(n26345), .C(n26344), .D(
        n26343), .X(n26347) );
  sky130_fd_sc_hd__o211ai_1 U31504 ( .A1(n26413), .A2(n26349), .B1(n26348), 
        .C1(n26347), .Y(n26350) );
  sky130_fd_sc_hd__a21oi_1 U31505 ( .A1(n26387), .A2(n26409), .B1(n26350), .Y(
        n26355) );
  sky130_fd_sc_hd__o21ai_1 U31506 ( .A1(n26352), .A2(n26709), .B1(n26351), .Y(
        n26353) );
  sky130_fd_sc_hd__nand2_1 U31507 ( .A(n27371), .B(n26353), .Y(n26354) );
  sky130_fd_sc_hd__nand2_1 U31508 ( .A(n26393), .B(n26360), .Y(n26361) );
  sky130_fd_sc_hd__o21ai_1 U31509 ( .A1(n27209), .A2(n26395), .B1(n26361), .Y(
        j202_soc_core_j22_cpu_rf_N2728) );
  sky130_fd_sc_hd__nand2_1 U31510 ( .A(n26393), .B(n26362), .Y(n26363) );
  sky130_fd_sc_hd__o21ai_1 U31511 ( .A1(n27213), .A2(n26395), .B1(n26363), .Y(
        j202_soc_core_j22_cpu_rf_N2802) );
  sky130_fd_sc_hd__nand2_1 U31512 ( .A(n26393), .B(n27215), .Y(n26364) );
  sky130_fd_sc_hd__o21ai_1 U31513 ( .A1(n27215), .A2(n26395), .B1(n26364), .Y(
        j202_soc_core_j22_cpu_rf_N2913) );
  sky130_fd_sc_hd__nand2_1 U31514 ( .A(n26393), .B(n27223), .Y(n26365) );
  sky130_fd_sc_hd__o21ai_1 U31515 ( .A1(n27223), .A2(n26395), .B1(n26365), .Y(
        j202_soc_core_j22_cpu_rf_N3024) );
  sky130_fd_sc_hd__nand2_1 U31516 ( .A(n26393), .B(n25819), .Y(n26366) );
  sky130_fd_sc_hd__nand2_1 U31518 ( .A(n26393), .B(n27225), .Y(n26367) );
  sky130_fd_sc_hd__o21ai_1 U31519 ( .A1(n27225), .A2(n26395), .B1(n26367), .Y(
        j202_soc_core_j22_cpu_rf_N2950) );
  sky130_fd_sc_hd__nand2_1 U31520 ( .A(n26393), .B(n11141), .Y(n26368) );
  sky130_fd_sc_hd__o21ai_1 U31521 ( .A1(n11141), .A2(n26395), .B1(n26368), .Y(
        j202_soc_core_j22_cpu_rf_N2691) );
  sky130_fd_sc_hd__nand2_1 U31522 ( .A(n26393), .B(n26369), .Y(n26370) );
  sky130_fd_sc_hd__o21ai_1 U31523 ( .A1(n27219), .A2(n26395), .B1(n26370), .Y(
        j202_soc_core_j22_cpu_rf_N2987) );
  sky130_fd_sc_hd__nand2_1 U31524 ( .A(n26393), .B(n26371), .Y(n26372) );
  sky130_fd_sc_hd__nand2_1 U31525 ( .A(n26393), .B(n25818), .Y(n26373) );
  sky130_fd_sc_hd__o21ai_1 U31526 ( .A1(n27466), .A2(n26395), .B1(n26373), .Y(
        j202_soc_core_j22_cpu_rf_N2765) );
  sky130_fd_sc_hd__nand2_1 U31527 ( .A(n26393), .B(n26374), .Y(n26375) );
  sky130_fd_sc_hd__nand2_1 U31528 ( .A(n26393), .B(n27211), .Y(n26376) );
  sky130_fd_sc_hd__o21ai_1 U31529 ( .A1(n27211), .A2(n26395), .B1(n26376), .Y(
        j202_soc_core_j22_cpu_rf_N3209) );
  sky130_fd_sc_hd__nand2_1 U31530 ( .A(n26393), .B(n26378), .Y(n26377) );
  sky130_fd_sc_hd__o21ai_1 U31531 ( .A1(n26378), .A2(n26395), .B1(n26377), .Y(
        j202_soc_core_j22_cpu_rf_N3246) );
  sky130_fd_sc_hd__nand2_1 U31532 ( .A(n26393), .B(n26379), .Y(n26380) );
  sky130_fd_sc_hd__o21ai_1 U31533 ( .A1(n27226), .A2(n26395), .B1(n26380), .Y(
        j202_soc_core_j22_cpu_rf_N3135) );
  sky130_fd_sc_hd__nand2_1 U31534 ( .A(n26393), .B(n27228), .Y(n26381) );
  sky130_fd_sc_hd__o21ai_1 U31535 ( .A1(n27228), .A2(n26395), .B1(n26381), .Y(
        j202_soc_core_j22_cpu_rf_N3172) );
  sky130_fd_sc_hd__mux2i_1 U31536 ( .A0(n26395), .A1(n26426), .S(n27006), .Y(
        j202_soc_core_j22_cpu_ml_N315) );
  sky130_fd_sc_hd__mux2i_1 U31537 ( .A0(n26382), .A1(n26395), .S(n27460), .Y(
        j202_soc_core_j22_cpu_rf_N3283) );
  sky130_fd_sc_hd__nand2_1 U31538 ( .A(n26393), .B(n26383), .Y(n26384) );
  sky130_fd_sc_hd__o21ai_0 U31539 ( .A1(n26395), .A2(n26899), .B1(n26384), .Y(
        j202_soc_core_j22_cpu_rf_N3323) );
  sky130_fd_sc_hd__nand2_1 U31540 ( .A(n26393), .B(n26516), .Y(n26386) );
  sky130_fd_sc_hd__a22oi_1 U31541 ( .A1(n26390), .A2(n26948), .B1(n27371), 
        .B2(n24650), .Y(n26385) );
  sky130_fd_sc_hd__nand2_1 U31542 ( .A(n26386), .B(n26385), .Y(
        j202_soc_core_j22_cpu_rf_N3358) );
  sky130_fd_sc_hd__nand2_1 U31543 ( .A(n27371), .B(n11157), .Y(n26392) );
  sky130_fd_sc_hd__o22ai_1 U31544 ( .A1(n26413), .A2(n26892), .B1(n26891), 
        .B2(n26388), .Y(n26389) );
  sky130_fd_sc_hd__a21oi_1 U31545 ( .A1(n26390), .A2(n26895), .B1(n26389), .Y(
        n26391) );
  sky130_fd_sc_hd__nand2_1 U31546 ( .A(n26392), .B(n26391), .Y(
        j202_soc_core_j22_cpu_rf_N310) );
  sky130_fd_sc_hd__nand2_1 U31547 ( .A(n26393), .B(n11109), .Y(n26394) );
  sky130_fd_sc_hd__o21ai_1 U31548 ( .A1(n27575), .A2(n26395), .B1(n26394), .Y(
        j202_soc_core_j22_cpu_rf_N3098) );
  sky130_fd_sc_hd__a31oi_1 U31549 ( .A1(n26402), .A2(n11713), .A3(n26401), 
        .B1(n18916), .Y(n26403) );
  sky130_fd_sc_hd__o21ai_1 U31550 ( .A1(n26406), .A2(n26414), .B1(n26405), .Y(
        n26408) );
  sky130_fd_sc_hd__nand2_1 U31551 ( .A(n26408), .B(n26407), .Y(n26442) );
  sky130_fd_sc_hd__nand2_1 U31552 ( .A(n26410), .B(n26409), .Y(n26440) );
  sky130_fd_sc_hd__xnor2_1 U31554 ( .A(n26414), .B(n27368), .Y(n26622) );
  sky130_fd_sc_hd__o22ai_1 U31555 ( .A1(n26417), .A2(n26416), .B1(n26415), 
        .B2(n26622), .Y(n26421) );
  sky130_fd_sc_hd__o22ai_1 U31556 ( .A1(n26563), .A2(n26419), .B1(n26578), 
        .B2(n26418), .Y(n26420) );
  sky130_fd_sc_hd__nor2_1 U31557 ( .A(n26421), .B(n26420), .Y(n26436) );
  sky130_fd_sc_hd__o22ai_1 U31558 ( .A1(n26423), .A2(n27368), .B1(n26422), 
        .B2(n26705), .Y(n26430) );
  sky130_fd_sc_hd__nor2_1 U31559 ( .A(n26702), .B(n26424), .Y(n26429) );
  sky130_fd_sc_hd__o22ai_1 U31560 ( .A1(n26707), .A2(n26427), .B1(n26426), 
        .B2(n26425), .Y(n26428) );
  sky130_fd_sc_hd__nor3_1 U31561 ( .A(n26430), .B(n26429), .C(n26428), .Y(
        n26435) );
  sky130_fd_sc_hd__nand2_1 U31563 ( .A(n26433), .B(n27368), .Y(n26434) );
  sky130_fd_sc_hd__nand3_1 U31564 ( .A(n26436), .B(n26435), .C(n26434), .Y(
        n26437) );
  sky130_fd_sc_hd__nor2_1 U31565 ( .A(n26438), .B(n26437), .Y(n26439) );
  sky130_fd_sc_hd__nand2_1 U31566 ( .A(n26440), .B(n26439), .Y(n26441) );
  sky130_fd_sc_hd__a21oi_1 U31567 ( .A1(n26557), .A2(n26442), .B1(n26441), .Y(
        n26445) );
  sky130_fd_sc_hd__a22oi_1 U31568 ( .A1(n26446), .A2(n26948), .B1(n26557), 
        .B2(n24650), .Y(n26447) );
  sky130_fd_sc_hd__nand2_1 U31569 ( .A(n26448), .B(n26447), .Y(
        j202_soc_core_j22_cpu_rf_N3376) );
  sky130_fd_sc_hd__o22ai_1 U31571 ( .A1(n27219), .A2(n27370), .B1(n27218), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N3006) );
  sky130_fd_sc_hd__o22ai_1 U31572 ( .A1(n27217), .A2(n27370), .B1(n27216), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N2858) );
  sky130_fd_sc_hd__o22ai_1 U31573 ( .A1(n27228), .A2(n27370), .B1(n27227), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N3191) );
  sky130_fd_sc_hd__o22ai_1 U31574 ( .A1(n27225), .A2(n27370), .B1(n27224), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N2969) );
  sky130_fd_sc_hd__o22ai_1 U31575 ( .A1(n27466), .A2(n27370), .B1(n27465), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N2784) );
  sky130_fd_sc_hd__o22ai_1 U31576 ( .A1(n27215), .A2(n27370), .B1(n27214), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N2932) );
  sky130_fd_sc_hd__o22ai_1 U31577 ( .A1(n27223), .A2(n27370), .B1(n27222), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N3043) );
  sky130_fd_sc_hd__o22ai_1 U31578 ( .A1(n27211), .A2(n27370), .B1(n27210), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N3228) );
  sky130_fd_sc_hd__o22ai_1 U31579 ( .A1(n27221), .A2(n27370), .B1(n27220), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N2895) );
  sky130_fd_sc_hd__o22ai_1 U31580 ( .A1(n27226), .A2(n27370), .B1(n23079), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N3154) );
  sky130_fd_sc_hd__o22ai_1 U31581 ( .A1(n27213), .A2(n27370), .B1(n27212), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N2821) );
  sky130_fd_sc_hd__o22ai_1 U31582 ( .A1(n26378), .A2(n27370), .B1(n26449), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N3265) );
  sky130_fd_sc_hd__o22ai_1 U31583 ( .A1(n27209), .A2(n27370), .B1(n23039), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N2747) );
  sky130_fd_sc_hd__o22ai_1 U31584 ( .A1(n11141), .A2(n27370), .B1(n27124), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N2710) );
  sky130_fd_sc_hd__o22ai_1 U31585 ( .A1(n27370), .A2(n26899), .B1(n26898), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N3340) );
  sky130_fd_sc_hd__o22ai_1 U31586 ( .A1(n27021), .A2(n26456), .B1(n26451), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U31587 ( .A1(n26456), .A2(n27990), .B1(n26452), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U31588 ( .A1(n27757), .A2(n26453), .B1(n28477), 
        .B2(n27754), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U31589 ( .A1(n27583), .A2(n26458), .B1(n28477), 
        .B2(n27581), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U31590 ( .A1(n28541), .A2(n26456), .B1(n26454), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U31591 ( .A1(n26456), .A2(n27194), .B1(n26455), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__a21oi_1 U31592 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[28]), .B1(n27758), .Y(n26457) );
  sky130_fd_sc_hd__o21ai_1 U31593 ( .A1(n26458), .A2(n27097), .B1(n26457), .Y(
        n26459) );
  sky130_fd_sc_hd__a21oi_1 U31594 ( .A1(n27862), .A2(
        j202_soc_core_intc_core_00_rg_ipr[60]), .B1(n26459), .Y(n26464) );
  sky130_fd_sc_hd__a22o_1 U31595 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[28]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[92]), .X(n26460) );
  sky130_fd_sc_hd__a21oi_1 U31596 ( .A1(j202_soc_core_intc_core_00_rg_itgt[7]), 
        .A2(n27850), .B1(n26460), .Y(n26463) );
  sky130_fd_sc_hd__a22oi_1 U31597 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[31]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[124]), .Y(n26462) );
  sky130_fd_sc_hd__nand2_1 U31598 ( .A(n27869), .B(
        j202_soc_core_intc_core_00_rg_itgt[15]), .Y(n26461) );
  sky130_fd_sc_hd__nand4_1 U31599 ( .A(n26464), .B(n26463), .C(n26462), .D(
        n26461), .Y(j202_soc_core_ahb2apb_01_N156) );
  sky130_fd_sc_hd__nand2_1 U31600 ( .A(n27108), .B(j202_soc_core_uart_div0[4]), 
        .Y(n26465) );
  sky130_fd_sc_hd__o21ai_1 U31601 ( .A1(n26466), .A2(n27108), .B1(n26465), .Y(
        n42) );
  sky130_fd_sc_hd__a22o_1 U31602 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[28]), .A2(n27719), .B1(n27718), 
        .B2(n26467), .X(j202_soc_core_wbqspiflash_00_N695) );
  sky130_fd_sc_hd__o21ai_0 U31603 ( .A1(n27192), .A2(n27370), .B1(n26468), .Y(
        j202_soc_core_j22_cpu_rf_N3302) );
  sky130_fd_sc_hd__o22ai_1 U31604 ( .A1(n27333), .A2(n27370), .B1(n23178), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N3080) );
  sky130_fd_sc_hd__o22ai_1 U31605 ( .A1(n27466), .A2(n24546), .B1(n27465), 
        .B2(n26470), .Y(j202_soc_core_j22_cpu_rf_N2774) );
  sky130_fd_sc_hd__nand2_1 U31606 ( .A(n26717), .B(n27184), .Y(n26471) );
  sky130_fd_sc_hd__o211ai_1 U31607 ( .A1(n24546), .A2(n26861), .B1(n26471), 
        .C1(n27346), .Y(j202_soc_core_j22_cpu_ml_N324) );
  sky130_fd_sc_hd__a22oi_1 U31608 ( .A1(n27187), .A2(
        j202_soc_core_j22_cpu_ml_bufa[20]), .B1(n27273), .B2(n26472), .Y(
        n26473) );
  sky130_fd_sc_hd__nand2_1 U31609 ( .A(n27189), .B(n26473), .Y(
        j202_soc_core_j22_cpu_ml_machj[20]) );
  sky130_fd_sc_hd__o22ai_1 U31610 ( .A1(n28604), .A2(n27194), .B1(n26485), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__nor2_1 U31611 ( .A(n26475), .B(n26474), .Y(
        j202_soc_core_wbqspiflash_00_N741) );
  sky130_fd_sc_hd__a21oi_1 U31612 ( .A1(n28148), .A2(
        j202_soc_core_wbqspiflash_00_write_in_progress), .B1(n26476), .Y(
        n26478) );
  sky130_fd_sc_hd__a21oi_1 U31614 ( .A1(n26480), .A2(n26479), .B1(
        j202_soc_core_intc_core_00_rg_irqc[20]), .Y(n26483) );
  sky130_fd_sc_hd__nor2_1 U31615 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[20]), 
        .B(n26481), .Y(n26482) );
  sky130_fd_sc_hd__a31oi_1 U31616 ( .A1(n26483), .A2(
        j202_soc_core_intc_core_00_in_intreq[20]), .A3(n29594), .B1(n26482), 
        .Y(n26484) );
  sky130_fd_sc_hd__nor2_1 U31617 ( .A(n26485), .B(n26484), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N23) );
  sky130_fd_sc_hd__o22ai_1 U31618 ( .A1(n27583), .A2(n26486), .B1(n28384), 
        .B2(n27581), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__nand2_1 U31619 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[22]), .Y(n26487) );
  sky130_fd_sc_hd__o21ai_1 U31620 ( .A1(n26488), .A2(n27983), .B1(n26487), .Y(
        n68) );
  sky130_fd_sc_hd__o22ai_1 U31621 ( .A1(n26494), .A2(n27990), .B1(n26498), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U31622 ( .A1(n26494), .A2(n28535), .B1(n26489), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U31623 ( .A1(n26494), .A2(n28547), .B1(n26490), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U31624 ( .A1(n26494), .A2(n28538), .B1(n26496), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U31625 ( .A1(n26494), .A2(n28541), .B1(n26491), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U31626 ( .A1(n28544), .A2(n26494), .B1(n26492), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U31627 ( .A1(n26494), .A2(n27194), .B1(n26493), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__a21oi_1 U31628 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[22]), .B1(n27758), .Y(n26495) );
  sky130_fd_sc_hd__o21ai_1 U31629 ( .A1(n26496), .A2(n27097), .B1(n26495), .Y(
        n26497) );
  sky130_fd_sc_hd__a21oi_1 U31630 ( .A1(j202_soc_core_intc_core_00_rg_ipr[54]), 
        .A2(n27862), .B1(n26497), .Y(n26504) );
  sky130_fd_sc_hd__o22ai_1 U31631 ( .A1(n26499), .A2(n27676), .B1(n27312), 
        .B2(n26498), .Y(n26500) );
  sky130_fd_sc_hd__a21oi_1 U31632 ( .A1(n27850), .A2(
        j202_soc_core_intc_core_00_rg_itgt[69]), .B1(n26500), .Y(n26503) );
  sky130_fd_sc_hd__a22oi_1 U31633 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[93]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[118]), .Y(n26502) );
  sky130_fd_sc_hd__nand2_1 U31634 ( .A(n27869), .B(
        j202_soc_core_intc_core_00_rg_itgt[77]), .Y(n26501) );
  sky130_fd_sc_hd__nand4_1 U31635 ( .A(n26504), .B(n26503), .C(n26502), .D(
        n26501), .Y(j202_soc_core_ahb2apb_01_N150) );
  sky130_fd_sc_hd__nand2_1 U31636 ( .A(n27593), .B(j202_soc_core_uart_div1[6]), 
        .Y(n26505) );
  sky130_fd_sc_hd__o21ai_1 U31637 ( .A1(n26506), .A2(n27593), .B1(n26505), .Y(
        n74) );
  sky130_fd_sc_hd__a22oi_1 U31638 ( .A1(n27184), .A2(n26508), .B1(n26507), 
        .B2(n27339), .Y(n26509) );
  sky130_fd_sc_hd__nand2_1 U31639 ( .A(n27346), .B(n26509), .Y(
        j202_soc_core_j22_cpu_ml_N326) );
  sky130_fd_sc_hd__a22oi_1 U31640 ( .A1(n27187), .A2(n12725), .B1(n27273), 
        .B2(n26510), .Y(n26511) );
  sky130_fd_sc_hd__nand2_1 U31641 ( .A(n27189), .B(n26511), .Y(
        j202_soc_core_j22_cpu_ml_machj[22]) );
  sky130_fd_sc_hd__o22ai_1 U31642 ( .A1(n27466), .A2(n27407), .B1(n27465), 
        .B2(n12391), .Y(j202_soc_core_j22_cpu_rf_N2777) );
  sky130_fd_sc_hd__o21ai_0 U31644 ( .A1(n18916), .A2(n26515), .B1(n26514), .Y(
        n26517) );
  sky130_fd_sc_hd__a22oi_1 U31646 ( .A1(n26520), .A2(n26948), .B1(n11771), 
        .B2(n24650), .Y(n26521) );
  sky130_fd_sc_hd__nand2_1 U31647 ( .A(n26522), .B(n26521), .Y(
        j202_soc_core_j22_cpu_rf_N3378) );
  sky130_fd_sc_hd__nand4b_1 U31648 ( .A_N(n11669), .B(n12399), .C(n29513), .D(
        n26524), .Y(n26527) );
  sky130_fd_sc_hd__nor3_1 U31649 ( .A(n12616), .B(n29517), .C(n26527), .Y(
        n26547) );
  sky130_fd_sc_hd__nor2_1 U31650 ( .A(n26529), .B(n26528), .Y(n26534) );
  sky130_fd_sc_hd__nand2_1 U31651 ( .A(n26532), .B(n26539), .Y(n26533) );
  sky130_fd_sc_hd__o211a_2 U31652 ( .A1(n26548), .A2(n26534), .B1(n26783), 
        .C1(n26533), .X(n26546) );
  sky130_fd_sc_hd__nand4_1 U31653 ( .A(n26538), .B(n12359), .C(n26536), .D(
        n26535), .Y(n26540) );
  sky130_fd_sc_hd__nand2_1 U31654 ( .A(n26540), .B(n26539), .Y(n26541) );
  sky130_fd_sc_hd__nand3_1 U31655 ( .A(n26543), .B(n26542), .C(n26541), .Y(
        n26544) );
  sky130_fd_sc_hd__nor2_1 U31656 ( .A(n12120), .B(n26544), .Y(n26545) );
  sky130_fd_sc_hd__o211ai_1 U31657 ( .A1(n26548), .A2(n26547), .B1(n26546), 
        .C1(n26545), .Y(n26549) );
  sky130_fd_sc_hd__nor2_1 U31658 ( .A(n12647), .B(n26549), .Y(n26562) );
  sky130_fd_sc_hd__nor2_1 U31659 ( .A(n11704), .B(n12645), .Y(n26561) );
  sky130_fd_sc_hd__nor3_1 U31660 ( .A(n27442), .B(n12417), .C(n26554), .Y(
        n26560) );
  sky130_fd_sc_hd__nand4_1 U31661 ( .A(n26556), .B(n12451), .C(n27417), .D(
        n26555), .Y(n26558) );
  sky130_fd_sc_hd__nor2_1 U31662 ( .A(n26558), .B(n26557), .Y(n26559) );
  sky130_fd_sc_hd__nand4_1 U31663 ( .A(n26562), .B(n26561), .C(n26560), .D(
        n26559), .Y(n26599) );
  sky130_fd_sc_hd__o22ai_1 U31664 ( .A1(n27380), .A2(n26563), .B1(n27375), 
        .B2(n26707), .Y(n26576) );
  sky130_fd_sc_hd__o22ai_1 U31665 ( .A1(n26567), .A2(n26566), .B1(n26565), 
        .B2(n26564), .Y(n26575) );
  sky130_fd_sc_hd__o22ai_1 U31666 ( .A1(n26570), .A2(n26569), .B1(n26568), 
        .B2(n26705), .Y(n26574) );
  sky130_fd_sc_hd__o22ai_1 U31667 ( .A1(n27341), .A2(n26885), .B1(n26572), 
        .B2(n26571), .Y(n26573) );
  sky130_fd_sc_hd__nor4_1 U31668 ( .A(n26576), .B(n26575), .C(n26574), .D(
        n26573), .Y(n26597) );
  sky130_fd_sc_hd__nand2_1 U31669 ( .A(n26672), .B(n26746), .Y(n26587) );
  sky130_fd_sc_hd__o22ai_1 U31670 ( .A1(n26791), .A2(n27007), .B1(n26893), 
        .B2(n26577), .Y(n26586) );
  sky130_fd_sc_hd__o22ai_1 U31671 ( .A1(n26581), .A2(n26580), .B1(n26579), 
        .B2(n26578), .Y(n26585) );
  sky130_fd_sc_hd__o22ai_1 U31672 ( .A1(n11145), .A2(n11977), .B1(n26708), 
        .B2(n26582), .Y(n26584) );
  sky130_fd_sc_hd__nor4_1 U31673 ( .A(n26587), .B(n26586), .C(n26585), .D(
        n26584), .Y(n26596) );
  sky130_fd_sc_hd__nand4_1 U31674 ( .A(n26634), .B(n26632), .C(n26673), .D(
        n26650), .Y(n26594) );
  sky130_fd_sc_hd__nand4_1 U31675 ( .A(n26611), .B(n26663), .C(n26615), .D(
        n26613), .Y(n26593) );
  sky130_fd_sc_hd__nand4_1 U31676 ( .A(n26656), .B(n26657), .C(n26648), .D(
        n26646), .Y(n26592) );
  sky130_fd_sc_hd__a21oi_1 U31677 ( .A1(n27377), .A2(n26720), .B1(n26605), .Y(
        n26590) );
  sky130_fd_sc_hd__nand4_1 U31678 ( .A(n26590), .B(n26589), .C(n26627), .D(
        n26588), .Y(n26591) );
  sky130_fd_sc_hd__nor4_1 U31679 ( .A(n26594), .B(n26593), .C(n26592), .D(
        n26591), .Y(n26595) );
  sky130_fd_sc_hd__nand3_1 U31680 ( .A(n26597), .B(n26596), .C(n26595), .Y(
        n26598) );
  sky130_fd_sc_hd__mux2i_1 U31681 ( .A0(n26599), .A1(n26598), .S(
        j202_soc_core_j22_cpu_exuop_EXU_[0]), .Y(n26800) );
  sky130_fd_sc_hd__a22oi_1 U31682 ( .A1(n26912), .A2(n26711), .B1(n12493), 
        .B2(n26600), .Y(n26602) );
  sky130_fd_sc_hd__nand2_1 U31683 ( .A(n26602), .B(n26601), .Y(n26685) );
  sky130_fd_sc_hd__a22oi_1 U31684 ( .A1(n12417), .A2(n26723), .B1(n26603), 
        .B2(n27442), .Y(n26609) );
  sky130_fd_sc_hd__nor2_1 U31685 ( .A(n26605), .B(n26604), .Y(n26608) );
  sky130_fd_sc_hd__nand2_1 U31686 ( .A(n11704), .B(n26712), .Y(n26607) );
  sky130_fd_sc_hd__nand4_1 U31687 ( .A(n26609), .B(n26608), .C(n26607), .D(
        n26606), .Y(n26684) );
  sky130_fd_sc_hd__xor2_1 U31688 ( .A(n26610), .B(n26745), .X(n26689) );
  sky130_fd_sc_hd__xor2_1 U31689 ( .A(n26883), .B(n26689), .X(n26699) );
  sky130_fd_sc_hd__nand2_1 U31690 ( .A(n26612), .B(n26611), .Y(n26619) );
  sky130_fd_sc_hd__nand2_1 U31691 ( .A(n26614), .B(n26613), .Y(n26618) );
  sky130_fd_sc_hd__nand2_1 U31692 ( .A(n26616), .B(n26615), .Y(n26617) );
  sky130_fd_sc_hd__nand4_1 U31693 ( .A(n26700), .B(n26619), .C(n26618), .D(
        n26617), .Y(n26625) );
  sky130_fd_sc_hd__nor2_1 U31694 ( .A(n26621), .B(n26620), .Y(n26624) );
  sky130_fd_sc_hd__nand4b_1 U31695 ( .A_N(n26625), .B(n26624), .C(n26623), .D(
        n26622), .Y(n26764) );
  sky130_fd_sc_hd__nand2_1 U31696 ( .A(n26626), .B(n26746), .Y(n26630) );
  sky130_fd_sc_hd__nand2_1 U31697 ( .A(n26628), .B(n26627), .Y(n26629) );
  sky130_fd_sc_hd__nand3_1 U31698 ( .A(n26631), .B(n26630), .C(n26629), .Y(
        n26643) );
  sky130_fd_sc_hd__nand2_1 U31699 ( .A(n26633), .B(n26632), .Y(n26637) );
  sky130_fd_sc_hd__nand2_1 U31700 ( .A(n26635), .B(n26634), .Y(n26636) );
  sky130_fd_sc_hd__nand2_1 U31701 ( .A(n26637), .B(n26636), .Y(n26639) );
  sky130_fd_sc_hd__nor2_1 U31702 ( .A(n26639), .B(n26638), .Y(n26641) );
  sky130_fd_sc_hd__nor2_1 U31703 ( .A(n26645), .B(n26644), .Y(n26662) );
  sky130_fd_sc_hd__nand2_1 U31704 ( .A(n26647), .B(n26646), .Y(n26654) );
  sky130_fd_sc_hd__nand2_1 U31705 ( .A(n26649), .B(n26648), .Y(n26653) );
  sky130_fd_sc_hd__nand2_1 U31706 ( .A(n26651), .B(n26650), .Y(n26652) );
  sky130_fd_sc_hd__and3_1 U31707 ( .A(n26654), .B(n26653), .C(n26652), .X(
        n26661) );
  sky130_fd_sc_hd__a22oi_1 U31708 ( .A1(n26658), .A2(n26657), .B1(n26656), 
        .B2(n26655), .Y(n26660) );
  sky130_fd_sc_hd__nand4_1 U31709 ( .A(n26662), .B(n26661), .C(n26660), .D(
        n26659), .Y(n26763) );
  sky130_fd_sc_hd__nand2_1 U31710 ( .A(n26664), .B(n26663), .Y(n26666) );
  sky130_fd_sc_hd__o211ai_1 U31711 ( .A1(n26668), .A2(n26667), .B1(n26666), 
        .C1(n26665), .Y(n26678) );
  sky130_fd_sc_hd__nand2_1 U31712 ( .A(n26670), .B(n26669), .Y(n26677) );
  sky130_fd_sc_hd__a22oi_1 U31713 ( .A1(n26674), .A2(n26673), .B1(n26672), 
        .B2(n26671), .Y(n26676) );
  sky130_fd_sc_hd__and4_1 U31714 ( .A(n26764), .B(n26753), .C(n26763), .D(
        n26754), .X(n26680) );
  sky130_fd_sc_hd__nand2_1 U31715 ( .A(n26738), .B(n26682), .Y(n26756) );
  sky130_fd_sc_hd__nand2_1 U31716 ( .A(n26682), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n26774) );
  sky130_fd_sc_hd__nand2b_1 U31717 ( .A_N(n26774), .B(n26679), .Y(n26697) );
  sky130_fd_sc_hd__o22ai_1 U31718 ( .A1(n26680), .A2(n26756), .B1(n26697), 
        .B2(n26745), .Y(n26681) );
  sky130_fd_sc_hd__a31oi_1 U31719 ( .A1(n26699), .A2(n26682), .A3(n26755), 
        .B1(n26681), .Y(n26683) );
  sky130_fd_sc_hd__xnor2_1 U31720 ( .A(j202_soc_core_j22_cpu_rfuo_sr__m_), .B(
        n26686), .Y(n26688) );
  sky130_fd_sc_hd__nand2_1 U31721 ( .A(n26775), .B(n26755), .Y(n26779) );
  sky130_fd_sc_hd__clkinv_1 U31722 ( .A(n26779), .Y(n26687) );
  sky130_fd_sc_hd__nand2_1 U31723 ( .A(n26688), .B(n26687), .Y(n26696) );
  sky130_fd_sc_hd__nand3_1 U31724 ( .A(n26692), .B(n26691), .C(n26690), .Y(
        n26695) );
  sky130_fd_sc_hd__nand3_1 U31725 ( .A(n26745), .B(n26693), .C(n26727), .Y(
        n26694) );
  sky130_fd_sc_hd__a31oi_1 U31726 ( .A1(n26696), .A2(n26695), .A3(n26694), 
        .B1(n26781), .Y(n26773) );
  sky130_fd_sc_hd__clkinv_1 U31727 ( .A(n26697), .Y(n26698) );
  sky130_fd_sc_hd__nand3_1 U31728 ( .A(n26699), .B(n26776), .C(n26698), .Y(
        n26771) );
  sky130_fd_sc_hd__nand4_1 U31729 ( .A(n26704), .B(n26703), .C(n26702), .D(
        n26701), .Y(n26737) );
  sky130_fd_sc_hd__nand4_1 U31730 ( .A(n26708), .B(n26707), .C(n26706), .D(
        n26705), .Y(n26736) );
  sky130_fd_sc_hd__nor4_1 U31731 ( .A(n26712), .B(n26711), .C(n26710), .D(
        n26709), .Y(n26715) );
  sky130_fd_sc_hd__nand4_1 U31732 ( .A(n26715), .B(n26714), .C(n26713), .D(
        n11145), .Y(n26735) );
  sky130_fd_sc_hd__nor4_1 U31733 ( .A(n26719), .B(n26718), .C(n26717), .D(
        n26716), .Y(n26733) );
  sky130_fd_sc_hd__nor4_1 U31734 ( .A(n26723), .B(n26722), .C(n26721), .D(
        n26720), .Y(n26732) );
  sky130_fd_sc_hd__nor4_1 U31735 ( .A(n26727), .B(n26726), .C(n26725), .D(
        n26724), .Y(n26731) );
  sky130_fd_sc_hd__nor4_1 U31736 ( .A(n26729), .B(n26728), .C(n27045), .D(
        n27183), .Y(n26730) );
  sky130_fd_sc_hd__nand4_1 U31737 ( .A(n26733), .B(n26732), .C(n26731), .D(
        n26730), .Y(n26734) );
  sky130_fd_sc_hd__or4_1 U31738 ( .A(n26737), .B(n26736), .C(n26735), .D(
        n26734), .X(n26741) );
  sky130_fd_sc_hd__nand2_1 U31739 ( .A(n26739), .B(n26738), .Y(n26785) );
  sky130_fd_sc_hd__nor2_1 U31740 ( .A(n26785), .B(n26859), .Y(n26740) );
  sky130_fd_sc_hd__a22oi_1 U31741 ( .A1(n26743), .A2(n26742), .B1(n26741), 
        .B2(n26740), .Y(n26770) );
  sky130_fd_sc_hd__o21ai_0 U31743 ( .A1(n27455), .A2(n27341), .B1(n26746), .Y(
        n26748) );
  sky130_fd_sc_hd__nand2_1 U31744 ( .A(n26748), .B(n26747), .Y(n26751) );
  sky130_fd_sc_hd__nand2_1 U31745 ( .A(n26750), .B(n26749), .Y(n26794) );
  sky130_fd_sc_hd__a21o_1 U31746 ( .A1(n26752), .A2(n26751), .B1(n26794), .X(
        n26769) );
  sky130_fd_sc_hd__o21ai_1 U31747 ( .A1(n26758), .A2(n26757), .B1(n26756), .Y(
        n26759) );
  sky130_fd_sc_hd__nand2_1 U31748 ( .A(n26759), .B(n26776), .Y(n26786) );
  sky130_fd_sc_hd__clkinv_1 U31749 ( .A(n26786), .Y(n26760) );
  sky130_fd_sc_hd__and3_1 U31750 ( .A(n26762), .B(n26761), .C(n26760), .X(
        n26767) );
  sky130_fd_sc_hd__nand3_1 U31751 ( .A(n26767), .B(n26766), .C(n26765), .Y(
        n26768) );
  sky130_fd_sc_hd__nand4_1 U31752 ( .A(n26771), .B(n26770), .C(n26769), .D(
        n26768), .Y(n26772) );
  sky130_fd_sc_hd__o21bai_1 U31753 ( .A1(n26776), .A2(n26775), .B1_N(n26774), 
        .Y(n26778) );
  sky130_fd_sc_hd__nand2_1 U31754 ( .A(n26778), .B(n26777), .Y(n26789) );
  sky130_fd_sc_hd__o22ai_1 U31755 ( .A1(n26781), .A2(n26780), .B1(
        j202_soc_core_j22_cpu_exuop_EXU_[3]), .B2(n26779), .Y(n26788) );
  sky130_fd_sc_hd__nand2_1 U31756 ( .A(n26783), .B(n26782), .Y(n26784) );
  sky130_fd_sc_hd__nand3_1 U31757 ( .A(n26786), .B(n26785), .C(n26784), .Y(
        n26787) );
  sky130_fd_sc_hd__nor3_1 U31758 ( .A(n26789), .B(n26788), .C(n26787), .Y(
        n26797) );
  sky130_fd_sc_hd__nor2_1 U31759 ( .A(n27443), .B(n27409), .Y(n26793) );
  sky130_fd_sc_hd__nand4_1 U31760 ( .A(n26793), .B(n26792), .C(n26791), .D(
        n26790), .Y(n26795) );
  sky130_fd_sc_hd__a21o_1 U31761 ( .A1(n26795), .A2(
        j202_soc_core_j22_cpu_exuop_EXU_[3]), .B1(n26794), .X(n26796) );
  sky130_fd_sc_hd__a21o_1 U31762 ( .A1(n26797), .A2(n26796), .B1(n14849), .X(
        n26813) );
  sky130_fd_sc_hd__nand3_1 U31764 ( .A(n26812), .B(n26802), .C(n26801), .Y(
        n26808) );
  sky130_fd_sc_hd__a22oi_1 U31765 ( .A1(n26805), .A2(n12417), .B1(n26804), 
        .B2(n26803), .Y(n26806) );
  sky130_fd_sc_hd__nand2_1 U31767 ( .A(n26809), .B(n26813), .Y(n26810) );
  sky130_fd_sc_hd__o211ai_1 U31768 ( .A1(n26812), .A2(n27064), .B1(n26811), 
        .C1(n26810), .Y(j202_soc_core_j22_cpu_rf_N2626) );
  sky130_fd_sc_hd__nand2_1 U31769 ( .A(n26814), .B(n26813), .Y(
        j202_soc_core_j22_cpu_rf_N2625) );
  sky130_fd_sc_hd__a22oi_1 U31770 ( .A1(j202_soc_core_j22_cpu_pc[0]), .A2(
        n26948), .B1(n12417), .B2(n24650), .Y(n26815) );
  sky130_fd_sc_hd__o21ai_1 U31771 ( .A1(n26951), .A2(n27063), .B1(n26815), .Y(
        j202_soc_core_j22_cpu_rf_N3345) );
  sky130_fd_sc_hd__o22ai_1 U31772 ( .A1(n27064), .A2(n27575), .B1(n27574), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N3085) );
  sky130_fd_sc_hd__o22ai_1 U31773 ( .A1(n27064), .A2(n27219), .B1(n27218), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N2974) );
  sky130_fd_sc_hd__o22ai_1 U31774 ( .A1(n27064), .A2(n27217), .B1(n27216), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N2826) );
  sky130_fd_sc_hd__o22ai_1 U31775 ( .A1(n27064), .A2(n27228), .B1(n27227), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N3159) );
  sky130_fd_sc_hd__o22ai_1 U31776 ( .A1(n27064), .A2(n27225), .B1(n27224), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N2937) );
  sky130_fd_sc_hd__o22ai_1 U31777 ( .A1(n27064), .A2(n27466), .B1(n27465), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N2752) );
  sky130_fd_sc_hd__o22ai_1 U31778 ( .A1(n27064), .A2(n27215), .B1(n27214), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N2900) );
  sky130_fd_sc_hd__o22ai_1 U31779 ( .A1(n27064), .A2(n27223), .B1(n27222), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N3011) );
  sky130_fd_sc_hd__o22ai_1 U31780 ( .A1(n27064), .A2(n27211), .B1(n27210), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N3196) );
  sky130_fd_sc_hd__o22ai_1 U31781 ( .A1(n27064), .A2(n27221), .B1(n27220), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N2863) );
  sky130_fd_sc_hd__o22ai_1 U31782 ( .A1(n27064), .A2(n27226), .B1(n23079), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N3122) );
  sky130_fd_sc_hd__o22ai_1 U31783 ( .A1(n27064), .A2(n27213), .B1(n27212), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N2789) );
  sky130_fd_sc_hd__o22ai_1 U31784 ( .A1(n27064), .A2(n27209), .B1(n23039), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N2715) );
  sky130_fd_sc_hd__o22ai_1 U31785 ( .A1(n27583), .A2(n26816), .B1(n28326), 
        .B2(n27581), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U31786 ( .A1(n28605), .A2(n27194), .B1(n26822), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__a21oi_1 U31787 ( .A1(n27195), .A2(n26817), .B1(
        j202_soc_core_intc_core_00_rg_irqc[18]), .Y(n26820) );
  sky130_fd_sc_hd__nor2_1 U31788 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[18]), 
        .B(n26818), .Y(n26819) );
  sky130_fd_sc_hd__a31oi_1 U31789 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[18]), .A2(n26820), .A3(n29594), 
        .B1(n26819), .Y(n26821) );
  sky130_fd_sc_hd__nor2_1 U31790 ( .A(n26822), .B(n26821), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N21) );
  sky130_fd_sc_hd__a22oi_1 U31791 ( .A1(n26826), .A2(n26825), .B1(n26824), 
        .B2(n26823), .Y(n26833) );
  sky130_fd_sc_hd__mux2i_1 U31792 ( .A0(n26830), .A1(n26829), .S(n26828), .Y(
        n26832) );
  sky130_fd_sc_hd__mux2i_1 U31793 ( .A0(n26833), .A1(n26832), .S(n26831), .Y(
        n26857) );
  sky130_fd_sc_hd__nand2_1 U31794 ( .A(n26834), .B(n12125), .Y(n27206) );
  sky130_fd_sc_hd__mux2i_1 U31795 ( .A0(n26838), .A1(n26837), .S(n26836), .Y(
        n26845) );
  sky130_fd_sc_hd__mux2i_1 U31796 ( .A0(n26842), .A1(n26841), .S(n26840), .Y(
        n26844) );
  sky130_fd_sc_hd__mux2i_1 U31797 ( .A0(n26845), .A1(n26844), .S(n26843), .Y(
        n26855) );
  sky130_fd_sc_hd__nor2_1 U31798 ( .A(n26848), .B(n26847), .Y(n26853) );
  sky130_fd_sc_hd__o21ai_1 U31799 ( .A1(n26850), .A2(n26849), .B1(n12142), .Y(
        n26852) );
  sky130_fd_sc_hd__nor4_1 U31800 ( .A(n26853), .B(n27204), .C(n26852), .D(
        n26851), .Y(n26854) );
  sky130_fd_sc_hd__o21ai_1 U31801 ( .A1(n26857), .A2(n27206), .B1(n26856), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N3) );
  sky130_fd_sc_hd__mux2i_1 U31802 ( .A0(n26858), .A1(n12451), .S(n27460), .Y(
        j202_soc_core_j22_cpu_rf_N3272) );
  sky130_fd_sc_hd__nand2_1 U31803 ( .A(n26859), .B(n27184), .Y(n26860) );
  sky130_fd_sc_hd__o211ai_1 U31804 ( .A1(n27349), .A2(n26861), .B1(n26860), 
        .C1(n27346), .Y(j202_soc_core_j22_cpu_ml_N335) );
  sky130_fd_sc_hd__nand2_1 U31805 ( .A(n12706), .B(n26862), .Y(n26868) );
  sky130_fd_sc_hd__nand2_1 U31806 ( .A(n26864), .B(n26863), .Y(n26866) );
  sky130_fd_sc_hd__a31oi_1 U31807 ( .A1(n26868), .A2(n26867), .A3(n26866), 
        .B1(n26865), .Y(n26869) );
  sky130_fd_sc_hd__a21oi_1 U31808 ( .A1(n22487), .A2(n27187), .B1(n26869), .Y(
        n26870) );
  sky130_fd_sc_hd__nand2_1 U31809 ( .A(n27189), .B(n26870), .Y(
        j202_soc_core_j22_cpu_ml_machj[31]) );
  sky130_fd_sc_hd__nand2_1 U31810 ( .A(n26873), .B(n26872), .Y(n26876) );
  sky130_fd_sc_hd__a31oi_1 U31811 ( .A1(n26876), .A2(n26875), .A3(n26874), 
        .B1(n26878), .Y(n26877) );
  sky130_fd_sc_hd__a21oi_1 U31812 ( .A1(n23247), .A2(n26878), .B1(n26877), .Y(
        n26879) );
  sky130_fd_sc_hd__nand3_1 U31813 ( .A(n26880), .B(n26879), .C(n27273), .Y(
        j202_soc_core_j22_cpu_ml_maclj[31]) );
  sky130_fd_sc_hd__nand2_1 U31814 ( .A(n26881), .B(n27192), .Y(n26882) );
  sky130_fd_sc_hd__o21ai_0 U31815 ( .A1(n27192), .A2(n27349), .B1(n26882), .Y(
        j202_soc_core_j22_cpu_rf_N3305) );
  sky130_fd_sc_hd__o22ai_1 U31816 ( .A1(n26885), .A2(n26892), .B1(n26891), 
        .B2(n26884), .Y(n26886) );
  sky130_fd_sc_hd__a21oi_1 U31817 ( .A1(n26887), .A2(n26895), .B1(n26886), .Y(
        n26888) );
  sky130_fd_sc_hd__o21ai_0 U31818 ( .A1(n26897), .A2(n27349), .B1(n26888), .Y(
        j202_soc_core_j22_cpu_rf_N329) );
  sky130_fd_sc_hd__o22ai_1 U31819 ( .A1(n26893), .A2(n26892), .B1(n26891), 
        .B2(n26890), .Y(n26894) );
  sky130_fd_sc_hd__a21oi_1 U31820 ( .A1(n26913), .A2(n26895), .B1(n26894), .Y(
        n26896) );
  sky130_fd_sc_hd__o21ai_0 U31821 ( .A1(n26897), .A2(n27417), .B1(n26896), .Y(
        j202_soc_core_j22_cpu_rf_N303) );
  sky130_fd_sc_hd__o22ai_1 U31822 ( .A1(n27417), .A2(n26899), .B1(n26898), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N3315) );
  sky130_fd_sc_hd__o22ai_1 U31823 ( .A1(n27417), .A2(n11141), .B1(n27124), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N2683) );
  sky130_fd_sc_hd__o22ai_1 U31824 ( .A1(n28612), .A2(n27990), .B1(n26900), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U31825 ( .A1(n26905), .A2(n26904), .B1(n26903), 
        .B2(n26902), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N4) );
  sky130_fd_sc_hd__a21oi_1 U31826 ( .A1(j202_soc_core_intr_level__1_), .A2(
        n26907), .B1(n26906), .Y(n26910) );
  sky130_fd_sc_hd__nand2_1 U31827 ( .A(n12504), .B(n26908), .Y(n26909) );
  sky130_fd_sc_hd__o211ai_1 U31828 ( .A1(n26911), .A2(n26915), .B1(n26910), 
        .C1(n26909), .Y(j202_soc_core_j22_cpu_rf_N3388) );
  sky130_fd_sc_hd__a22oi_1 U31829 ( .A1(n26913), .A2(n26948), .B1(n12504), 
        .B2(n24650), .Y(n26914) );
  sky130_fd_sc_hd__o21ai_1 U31830 ( .A1(n26951), .A2(n26915), .B1(n26914), .Y(
        j202_soc_core_j22_cpu_rf_N3350) );
  sky130_fd_sc_hd__o22ai_1 U31831 ( .A1(n27417), .A2(n27575), .B1(n27574), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N3090) );
  sky130_fd_sc_hd__o22ai_1 U31832 ( .A1(n27417), .A2(n27333), .B1(n23178), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N3053) );
  sky130_fd_sc_hd__o22ai_1 U31833 ( .A1(n27417), .A2(n27219), .B1(n27218), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N2979) );
  sky130_fd_sc_hd__o22ai_1 U31834 ( .A1(n27417), .A2(n27217), .B1(n27216), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N2831) );
  sky130_fd_sc_hd__o22ai_1 U31835 ( .A1(n27417), .A2(n27228), .B1(n27227), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N3164) );
  sky130_fd_sc_hd__o22ai_1 U31836 ( .A1(n27417), .A2(n27466), .B1(n27465), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N2757) );
  sky130_fd_sc_hd__o22ai_1 U31837 ( .A1(n27417), .A2(n27215), .B1(n27214), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N2905) );
  sky130_fd_sc_hd__o22ai_1 U31838 ( .A1(n27417), .A2(n27223), .B1(n27222), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N3016) );
  sky130_fd_sc_hd__o22ai_1 U31839 ( .A1(n27417), .A2(n27221), .B1(n27220), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N2868) );
  sky130_fd_sc_hd__o22ai_1 U31840 ( .A1(n27417), .A2(n27226), .B1(n23079), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N3127) );
  sky130_fd_sc_hd__o22ai_1 U31841 ( .A1(n27417), .A2(n27213), .B1(n27212), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N2794) );
  sky130_fd_sc_hd__o22ai_1 U31842 ( .A1(n27417), .A2(n27209), .B1(n23039), 
        .B2(n26915), .Y(j202_soc_core_j22_cpu_rf_N2720) );
  sky130_fd_sc_hd__a22oi_1 U31843 ( .A1(n27482), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[5]), .B1(n26917), .B2(
        j202_soc_core_cmt_core_00_cnt0[5]), .Y(n26918) );
  sky130_fd_sc_hd__o21ai_1 U31844 ( .A1(j202_soc_core_cmt_core_00_cnt0[5]), 
        .A2(n26919), .B1(n26918), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[5]) );
  sky130_fd_sc_hd__nand2_1 U31845 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[5]), .Y(n26920) );
  sky130_fd_sc_hd__o21ai_1 U31846 ( .A1(n26924), .A2(n27827), .B1(n26920), .Y(
        n101) );
  sky130_fd_sc_hd__nand2_1 U31847 ( .A(n27829), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[5]), .Y(n26921) );
  sky130_fd_sc_hd__o21ai_1 U31848 ( .A1(n26924), .A2(n27829), .B1(n26921), .Y(
        n99) );
  sky130_fd_sc_hd__nand2_1 U31849 ( .A(n27831), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[5]), .Y(n26922) );
  sky130_fd_sc_hd__o21ai_1 U31850 ( .A1(n26924), .A2(n27831), .B1(n26922), .Y(
        n100) );
  sky130_fd_sc_hd__nand2_1 U31851 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[5]), .Y(n26923) );
  sky130_fd_sc_hd__o21ai_1 U31852 ( .A1(n26924), .A2(n27833), .B1(n26923), .Y(
        n102) );
  sky130_fd_sc_hd__a22oi_1 U31853 ( .A1(n27836), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[5]), .B1(n27835), .B2(
        j202_soc_core_cmt_core_00_const1[5]), .Y(n26928) );
  sky130_fd_sc_hd__a22oi_1 U31854 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[5]), .B1(n27837), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[5]), .Y(
        n26927) );
  sky130_fd_sc_hd__nand2_1 U31855 ( .A(n27839), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[5]), .Y(n26926) );
  sky130_fd_sc_hd__nand2_1 U31856 ( .A(n27840), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[5]), .Y(
        n26925) );
  sky130_fd_sc_hd__nand4_1 U31857 ( .A(n26928), .B(n26927), .C(n26926), .D(
        n26925), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[5]) );
  sky130_fd_sc_hd__nand2_1 U31858 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[5]), .Y(n26929) );
  sky130_fd_sc_hd__o21ai_1 U31859 ( .A1(n26930), .A2(n27983), .B1(n26929), .Y(
        n54) );
  sky130_fd_sc_hd__o22ai_1 U31860 ( .A1(n28612), .A2(n28535), .B1(n26937), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U31861 ( .A1(n28612), .A2(n28526), .B1(n26931), 
        .B2(n28524), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U31862 ( .A1(n28612), .A2(n28547), .B1(n26932), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U31863 ( .A1(n28612), .A2(n28538), .B1(n26933), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U31864 ( .A1(n28612), .A2(n28541), .B1(n26934), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U31865 ( .A1(n28544), .A2(n28612), .B1(n26935), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__a21oi_1 U31866 ( .A1(n27857), .A2(
        j202_soc_core_intc_core_00_rg_eimk[5]), .B1(n27758), .Y(n26936) );
  sky130_fd_sc_hd__o21ai_1 U31867 ( .A1(n26937), .A2(n27760), .B1(n26936), .Y(
        n26938) );
  sky130_fd_sc_hd__a21oi_1 U31868 ( .A1(n27860), .A2(
        j202_soc_core_intc_core_00_rg_ipr[101]), .B1(n26938), .Y(n26944) );
  sky130_fd_sc_hd__a22oi_1 U31869 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[5]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[5]), .Y(n26940) );
  sky130_fd_sc_hd__a22oi_1 U31870 ( .A1(n27852), .A2(
        j202_soc_core_intc_core_00_rg_ipr[69]), .B1(n27856), .B2(
        j202_soc_core_intc_core_00_rg_itgt[49]), .Y(n26939) );
  sky130_fd_sc_hd__o211ai_1 U31871 ( .A1(n24056), .A2(n27676), .B1(n26940), 
        .C1(n26939), .Y(n26941) );
  sky130_fd_sc_hd__a21oi_1 U31872 ( .A1(n27869), .A2(
        j202_soc_core_intc_core_00_rg_itgt[41]), .B1(n26941), .Y(n26943) );
  sky130_fd_sc_hd__a22oi_1 U31873 ( .A1(n27862), .A2(
        j202_soc_core_intc_core_00_rg_ipr[37]), .B1(n27861), .B2(
        j202_soc_core_intc_core_00_rg_itgt[57]), .Y(n26942) );
  sky130_fd_sc_hd__nand3_1 U31874 ( .A(n26944), .B(n26943), .C(n26942), .Y(
        j202_soc_core_ahb2apb_01_N133) );
  sky130_fd_sc_hd__nor2_1 U31875 ( .A(n26945), .B(n27874), .Y(
        j202_soc_core_wbqspiflash_00_N672) );
  sky130_fd_sc_hd__nor2_1 U31876 ( .A(n26946), .B(n11047), .Y(
        j202_soc_core_j22_cpu_rf_N2674) );
  sky130_fd_sc_hd__nand2_1 U31877 ( .A(n11612), .B(n27460), .Y(n26947) );
  sky130_fd_sc_hd__o21ai_1 U31878 ( .A1(n27460), .A2(n11047), .B1(n26947), .Y(
        j202_soc_core_j22_cpu_rf_N3303) );
  sky130_fd_sc_hd__a22oi_1 U31879 ( .A1(n26949), .A2(n26948), .B1(n11612), 
        .B2(n24650), .Y(n26950) );
  sky130_fd_sc_hd__o21ai_1 U31880 ( .A1(n26951), .A2(n11047), .B1(n26950), .Y(
        j202_soc_core_j22_cpu_rf_N3377) );
  sky130_fd_sc_hd__o22ai_1 U31881 ( .A1(n26959), .A2(n27021), .B1(n26952), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U31882 ( .A1(n26959), .A2(n27990), .B1(n26953), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U31883 ( .A1(n26959), .A2(n28535), .B1(n26954), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U31884 ( .A1(n26959), .A2(n28547), .B1(n26955), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U31885 ( .A1(n26959), .A2(n28538), .B1(n26961), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U31886 ( .A1(n26959), .A2(n28541), .B1(n26956), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U31887 ( .A1(n28544), .A2(n26959), .B1(n26957), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U31888 ( .A1(n26959), .A2(n27194), .B1(n26958), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__a21oi_1 U31889 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[29]), .B1(n27758), .Y(n26960) );
  sky130_fd_sc_hd__o21ai_1 U31890 ( .A1(n26961), .A2(n27097), .B1(n26960), .Y(
        n26962) );
  sky130_fd_sc_hd__a21oi_1 U31891 ( .A1(j202_soc_core_intc_core_00_rg_ipr[61]), 
        .A2(n27862), .B1(n26962), .Y(n26967) );
  sky130_fd_sc_hd__a22o_1 U31892 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[29]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[93]), .X(n26963) );
  sky130_fd_sc_hd__a21oi_1 U31893 ( .A1(n27850), .A2(
        j202_soc_core_intc_core_00_rg_itgt[39]), .B1(n26963), .Y(n26966) );
  sky130_fd_sc_hd__a22oi_1 U31894 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[63]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[125]), .Y(n26965) );
  sky130_fd_sc_hd__nand2_1 U31895 ( .A(n27869), .B(
        j202_soc_core_intc_core_00_rg_itgt[47]), .Y(n26964) );
  sky130_fd_sc_hd__nand4_1 U31896 ( .A(n26967), .B(n26966), .C(n26965), .D(
        n26964), .Y(j202_soc_core_ahb2apb_01_N157) );
  sky130_fd_sc_hd__nand2_1 U31897 ( .A(n27108), .B(j202_soc_core_uart_div0[5]), 
        .Y(n26968) );
  sky130_fd_sc_hd__o21ai_1 U31898 ( .A1(n26969), .A2(n27108), .B1(n26968), .Y(
        n72) );
  sky130_fd_sc_hd__a22o_1 U31899 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[29]), .A2(n27719), .B1(n27718), 
        .B2(j202_soc_core_wbqspiflash_00_spi_busy), .X(
        j202_soc_core_wbqspiflash_00_N696) );
  sky130_fd_sc_hd__a22oi_1 U31900 ( .A1(n27184), .A2(n26971), .B1(n11612), 
        .B2(n27339), .Y(n26972) );
  sky130_fd_sc_hd__nand2_1 U31901 ( .A(n27346), .B(n26972), .Y(
        j202_soc_core_j22_cpu_ml_N333) );
  sky130_fd_sc_hd__and3_1 U31902 ( .A(n26975), .B(n26974), .C(n26973), .X(
        n26980) );
  sky130_fd_sc_hd__o21ai_1 U31903 ( .A1(n26981), .A2(n26980), .B1(n26979), .Y(
        j202_soc_core_j22_cpu_ml_maclj[29]) );
  sky130_fd_sc_hd__nand2_1 U31904 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[4]), .Y(n26982) );
  sky130_fd_sc_hd__nand2_1 U31906 ( .A(n27829), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[4]), .Y(n26983) );
  sky130_fd_sc_hd__o21ai_1 U31907 ( .A1(n26986), .A2(n27829), .B1(n26983), .Y(
        n95) );
  sky130_fd_sc_hd__nand2_1 U31908 ( .A(n27831), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[4]), .Y(n26984) );
  sky130_fd_sc_hd__o21ai_1 U31909 ( .A1(n26986), .A2(n27831), .B1(n26984), .Y(
        n96) );
  sky130_fd_sc_hd__nand2_1 U31910 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[4]), .Y(n26985) );
  sky130_fd_sc_hd__o21ai_1 U31911 ( .A1(n26986), .A2(n27833), .B1(n26985), .Y(
        n98) );
  sky130_fd_sc_hd__a22oi_1 U31912 ( .A1(n27836), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[4]), .B1(n27835), .B2(
        j202_soc_core_cmt_core_00_const1[4]), .Y(n26990) );
  sky130_fd_sc_hd__a22oi_1 U31913 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[4]), .B1(n27837), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[4]), .Y(
        n26989) );
  sky130_fd_sc_hd__nand2_1 U31914 ( .A(n27839), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[4]), .Y(n26988) );
  sky130_fd_sc_hd__nand2_1 U31915 ( .A(n27840), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[4]), .Y(
        n26987) );
  sky130_fd_sc_hd__nand4_1 U31916 ( .A(n26990), .B(n26989), .C(n26988), .D(
        n26987), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[4]) );
  sky130_fd_sc_hd__nand2_1 U31917 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[4]), .Y(n26991) );
  sky130_fd_sc_hd__o21ai_1 U31918 ( .A1(n26992), .A2(n27983), .B1(n26991), .Y(
        n53) );
  sky130_fd_sc_hd__o22ai_1 U31919 ( .A1(n28613), .A2(n28526), .B1(n26993), 
        .B2(n28524), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U31920 ( .A1(n27757), .A2(n26994), .B1(n28300), 
        .B2(n27754), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U31921 ( .A1(n28541), .A2(n28613), .B1(n26995), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__a21oi_1 U31922 ( .A1(n27857), .A2(
        j202_soc_core_intc_core_00_rg_eimk[4]), .B1(n27758), .Y(n26996) );
  sky130_fd_sc_hd__o21ai_1 U31923 ( .A1(n26997), .A2(n27760), .B1(n26996), .Y(
        n26998) );
  sky130_fd_sc_hd__a21oi_1 U31924 ( .A1(n27860), .A2(
        j202_soc_core_intc_core_00_rg_ipr[100]), .B1(n26998), .Y(n27005) );
  sky130_fd_sc_hd__a22oi_1 U31925 ( .A1(n27852), .A2(
        j202_soc_core_intc_core_00_rg_ipr[68]), .B1(n27856), .B2(
        j202_soc_core_intc_core_00_rg_itgt[17]), .Y(n27001) );
  sky130_fd_sc_hd__a22oi_1 U31926 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[4]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[4]), .Y(n27000) );
  sky130_fd_sc_hd__nand2_1 U31927 ( .A(n27851), .B(
        j202_soc_core_intc_core_00_rg_ipr[4]), .Y(n26999) );
  sky130_fd_sc_hd__nand3_1 U31928 ( .A(n27001), .B(n27000), .C(n26999), .Y(
        n27002) );
  sky130_fd_sc_hd__a21oi_1 U31929 ( .A1(j202_soc_core_intc_core_00_rg_itgt[9]), 
        .A2(n27869), .B1(n27002), .Y(n27004) );
  sky130_fd_sc_hd__a22oi_1 U31930 ( .A1(n27862), .A2(
        j202_soc_core_intc_core_00_rg_ipr[36]), .B1(n27861), .B2(
        j202_soc_core_intc_core_00_rg_itgt[25]), .Y(n27003) );
  sky130_fd_sc_hd__nand3_1 U31931 ( .A(n27005), .B(n27004), .C(n27003), .Y(
        j202_soc_core_ahb2apb_01_N132) );
  sky130_fd_sc_hd__nor2_1 U31932 ( .A(n28178), .B(n27874), .Y(
        j202_soc_core_wbqspiflash_00_N671) );
  sky130_fd_sc_hd__mux2i_1 U31933 ( .A0(n27234), .A1(n27007), .S(n27006), .Y(
        j202_soc_core_j22_cpu_ml_N307) );
  sky130_fd_sc_hd__o22ai_1 U31934 ( .A1(n27010), .A2(n27009), .B1(n28355), 
        .B2(n27008), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U31935 ( .A1(n28596), .A2(n27194), .B1(n27015), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__nor3_1 U31936 ( .A(j202_soc_core_intc_core_00_rg_irqc[11]), 
        .B(n28590), .C(n27011), .Y(n27012) );
  sky130_fd_sc_hd__nand2b_1 U31938 ( .A_N(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[11]), 
        .B(n29060), .Y(n27016) );
  sky130_fd_sc_hd__a21oi_1 U31939 ( .A1(n27017), .A2(n27016), .B1(n27015), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N14) );
  sky130_fd_sc_hd__nand2_1 U31940 ( .A(n27206), .B(n27018), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N6) );
  sky130_fd_sc_hd__o22ai_1 U31941 ( .A1(n27028), .A2(n27021), .B1(n27020), 
        .B2(n27019), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U31942 ( .A1(n27028), .A2(n27990), .B1(n27022), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U31943 ( .A1(n27028), .A2(n28535), .B1(n27023), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U31944 ( .A1(n27028), .A2(n28547), .B1(n27024), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U31945 ( .A1(n27028), .A2(n28538), .B1(n27030), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U31946 ( .A1(n27028), .A2(n28541), .B1(n27025), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U31947 ( .A1(n28544), .A2(n27028), .B1(n27026), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U31948 ( .A1(n27028), .A2(n27194), .B1(n27027), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__a21oi_1 U31949 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[23]), .B1(n27758), .Y(n27029) );
  sky130_fd_sc_hd__o21ai_1 U31950 ( .A1(n27030), .A2(n27097), .B1(n27029), .Y(
        n27031) );
  sky130_fd_sc_hd__a21oi_1 U31951 ( .A1(j202_soc_core_intc_core_00_rg_ipr[55]), 
        .A2(n27862), .B1(n27031), .Y(n27036) );
  sky130_fd_sc_hd__a22o_1 U31952 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[23]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[87]), .X(n27032) );
  sky130_fd_sc_hd__a21oi_1 U31953 ( .A1(n27850), .A2(
        j202_soc_core_intc_core_00_rg_itgt[101]), .B1(n27032), .Y(n27035) );
  sky130_fd_sc_hd__a22oi_1 U31954 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[125]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[119]), .Y(n27034) );
  sky130_fd_sc_hd__nand2_1 U31955 ( .A(n27869), .B(
        j202_soc_core_intc_core_00_rg_itgt[109]), .Y(n27033) );
  sky130_fd_sc_hd__nand4_1 U31956 ( .A(n27036), .B(n27035), .C(n27034), .D(
        n27033), .Y(j202_soc_core_ahb2apb_01_N151) );
  sky130_fd_sc_hd__a22oi_1 U31957 ( .A1(
        j202_soc_core_wbqspiflash_00_write_in_progress), .A2(n27037), .B1(
        j202_soc_core_wbqspiflash_00_spi_out[31]), .B2(n27719), .Y(n27038) );
  sky130_fd_sc_hd__o31ai_1 U31958 ( .A1(n27040), .A2(n27039), .A3(n28148), 
        .B1(n27038), .Y(j202_soc_core_wbqspiflash_00_N698) );
  sky130_fd_sc_hd__nand2_1 U31959 ( .A(n27042), .B(
        j202_soc_core_qspi_wb_wdat[31]), .Y(n27041) );
  sky130_fd_sc_hd__a22oi_1 U31961 ( .A1(n27184), .A2(n27045), .B1(n11764), 
        .B2(n27339), .Y(n27046) );
  sky130_fd_sc_hd__nand2_1 U31962 ( .A(n27346), .B(n27046), .Y(
        j202_soc_core_j22_cpu_ml_N319) );
  sky130_fd_sc_hd__a22oi_1 U31963 ( .A1(n27187), .A2(n12577), .B1(n27048), 
        .B2(n27047), .Y(n27049) );
  sky130_fd_sc_hd__nand2_1 U31964 ( .A(n27189), .B(n27049), .Y(
        j202_soc_core_j22_cpu_ml_machj[16]) );
  sky130_fd_sc_hd__nand2_1 U31965 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[16]), .Y(n27050) );
  sky130_fd_sc_hd__o21ai_1 U31966 ( .A1(n27051), .A2(n27983), .B1(n27050), .Y(
        n64) );
  sky130_fd_sc_hd__o22ai_1 U31967 ( .A1(n27757), .A2(n27052), .B1(n28384), 
        .B2(n27754), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U31968 ( .A1(n28541), .A2(n28606), .B1(n27053), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__a22oi_1 U31969 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[16]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[80]), .Y(n27055) );
  sky130_fd_sc_hd__a22oi_1 U31970 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[16]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[16]), .Y(n27054) );
  sky130_fd_sc_hd__nand3_1 U31971 ( .A(n27055), .B(n27054), .C(n27865), .Y(
        n27056) );
  sky130_fd_sc_hd__a21oi_1 U31972 ( .A1(j202_soc_core_intc_core_00_rg_itgt[12]), .A2(n27869), .B1(n27056), .Y(n27060) );
  sky130_fd_sc_hd__a22oi_1 U31973 ( .A1(n27856), .A2(
        j202_soc_core_intc_core_00_rg_itgt[20]), .B1(n27850), .B2(
        j202_soc_core_intc_core_00_rg_itgt[4]), .Y(n27059) );
  sky130_fd_sc_hd__a22oi_1 U31974 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[28]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[112]), .Y(n27058) );
  sky130_fd_sc_hd__nand2_1 U31975 ( .A(n27862), .B(
        j202_soc_core_intc_core_00_rg_ipr[48]), .Y(n27057) );
  sky130_fd_sc_hd__nand4_1 U31976 ( .A(n27060), .B(n27059), .C(n27058), .D(
        n27057), .Y(j202_soc_core_ahb2apb_01_N144) );
  sky130_fd_sc_hd__nand2_1 U31977 ( .A(n27593), .B(j202_soc_core_uart_div1[0]), 
        .Y(n27061) );
  sky130_fd_sc_hd__o21ai_1 U31978 ( .A1(n27062), .A2(n27593), .B1(n27061), .Y(
        n70) );
  sky130_fd_sc_hd__nor2_1 U31979 ( .A(n28590), .B(n28165), .Y(
        j202_soc_core_wbqspiflash_00_N713) );
  sky130_fd_sc_hd__a22o_1 U31980 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[16]), .A2(n27719), .B1(n27718), 
        .B2(j202_soc_core_wbqspiflash_00_erased_sector[2]), .X(
        j202_soc_core_wbqspiflash_00_N683) );
  sky130_fd_sc_hd__o22ai_1 U31981 ( .A1(n27064), .A2(n27333), .B1(n23178), 
        .B2(n27063), .Y(j202_soc_core_j22_cpu_rf_N3048) );
  sky130_fd_sc_hd__mux2i_1 U31982 ( .A0(n27063), .A1(n27064), .S(n27460), .Y(
        j202_soc_core_j22_cpu_rf_N3270) );
  sky130_fd_sc_hd__clkinv_1 U31983 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[0]), 
        .Y(n27068) );
  sky130_fd_sc_hd__nor2_1 U31984 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[1]), 
        .B(n27068), .Y(n27071) );
  sky130_fd_sc_hd__clkinv_1 U31985 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[1]), 
        .Y(n27065) );
  sky130_fd_sc_hd__nor2_1 U31986 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[0]), 
        .B(n27065), .Y(n27069) );
  sky130_fd_sc_hd__a21oi_1 U31987 ( .A1(j202_soc_core_intc_core_00_bs_addr[1]), 
        .A2(n27071), .B1(n27069), .Y(n27067) );
  sky130_fd_sc_hd__o31ai_1 U31988 ( .A1(j202_soc_core_intc_core_00_bs_addr[1]), 
        .A2(j202_soc_core_ahb2apb_01_hsize_buf[0]), .A3(n27074), .B1(n27067), 
        .Y(n10747) );
  sky130_fd_sc_hd__o21ai_0 U31989 ( .A1(j202_soc_core_ahb2apb_01_hsize_buf[0]), 
        .A2(n28880), .B1(n27067), .Y(n10748) );
  sky130_fd_sc_hd__nand2_1 U31990 ( .A(j202_soc_core_intc_core_00_bs_addr[1]), 
        .B(n27068), .Y(n27073) );
  sky130_fd_sc_hd__a21oi_1 U31991 ( .A1(n27071), .A2(n27070), .B1(n27069), .Y(
        n27072) );
  sky130_fd_sc_hd__o21ai_0 U31992 ( .A1(j202_soc_core_intc_core_00_bs_addr[0]), 
        .A2(n27073), .B1(n27072), .Y(n10746) );
  sky130_fd_sc_hd__o21ai_0 U31993 ( .A1(n27074), .A2(n27073), .B1(n27072), .Y(
        n10745) );
  sky130_fd_sc_hd__o22ai_1 U31994 ( .A1(n27081), .A2(n27990), .B1(n27075), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U31995 ( .A1(n27081), .A2(n28535), .B1(n27076), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U31996 ( .A1(n27081), .A2(n28547), .B1(n27077), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U31997 ( .A1(n27081), .A2(n28538), .B1(n27083), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U31998 ( .A1(n27081), .A2(n28541), .B1(n27078), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U31999 ( .A1(n27081), .A2(n28544), .B1(n27079), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o22ai_1 U32000 ( .A1(n27081), .A2(n27194), .B1(n27080), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__a21oi_1 U32001 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[31]), .B1(n27758), .Y(n27082) );
  sky130_fd_sc_hd__o21ai_1 U32002 ( .A1(n27083), .A2(n27097), .B1(n27082), .Y(
        n27084) );
  sky130_fd_sc_hd__a21oi_1 U32003 ( .A1(j202_soc_core_intc_core_00_rg_ipr[63]), 
        .A2(n27862), .B1(n27084), .Y(n27089) );
  sky130_fd_sc_hd__a22o_1 U32004 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[31]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[95]), .X(n27085) );
  sky130_fd_sc_hd__a21oi_1 U32005 ( .A1(n27850), .A2(
        j202_soc_core_intc_core_00_rg_itgt[103]), .B1(n27085), .Y(n27088) );
  sky130_fd_sc_hd__a22oi_1 U32006 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[127]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[127]), .Y(n27087) );
  sky130_fd_sc_hd__nand2_1 U32007 ( .A(n27869), .B(
        j202_soc_core_intc_core_00_rg_itgt[111]), .Y(n27086) );
  sky130_fd_sc_hd__nand4_1 U32008 ( .A(n27089), .B(n27088), .C(n27087), .D(
        n27086), .Y(j202_soc_core_ahb2apb_01_N159) );
  sky130_fd_sc_hd__o22ai_1 U32009 ( .A1(n27095), .A2(n27990), .B1(n27100), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U32010 ( .A1(n27095), .A2(n28535), .B1(n27090), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U32011 ( .A1(n27095), .A2(n28547), .B1(n27091), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U32012 ( .A1(n27095), .A2(n28538), .B1(n27098), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U32013 ( .A1(n27095), .A2(n28541), .B1(n27092), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U32014 ( .A1(n28544), .A2(n27095), .B1(n27093), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U32015 ( .A1(n27095), .A2(n27194), .B1(n27094), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__a21oi_1 U32016 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[30]), .B1(n27758), .Y(n27096) );
  sky130_fd_sc_hd__o21ai_1 U32017 ( .A1(n27098), .A2(n27097), .B1(n27096), .Y(
        n27099) );
  sky130_fd_sc_hd__a21oi_1 U32018 ( .A1(j202_soc_core_intc_core_00_rg_ipr[62]), 
        .A2(n27862), .B1(n27099), .Y(n27106) );
  sky130_fd_sc_hd__o22ai_1 U32019 ( .A1(n27101), .A2(n27676), .B1(n27312), 
        .B2(n27100), .Y(n27102) );
  sky130_fd_sc_hd__a21oi_1 U32020 ( .A1(n27850), .A2(
        j202_soc_core_intc_core_00_rg_itgt[71]), .B1(n27102), .Y(n27105) );
  sky130_fd_sc_hd__a22oi_1 U32021 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[95]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[126]), .Y(n27104) );
  sky130_fd_sc_hd__nand2_1 U32022 ( .A(n27869), .B(
        j202_soc_core_intc_core_00_rg_itgt[79]), .Y(n27103) );
  sky130_fd_sc_hd__nand4_1 U32023 ( .A(n27106), .B(n27105), .C(n27104), .D(
        n27103), .Y(j202_soc_core_ahb2apb_01_N158) );
  sky130_fd_sc_hd__nand2_1 U32024 ( .A(n27108), .B(j202_soc_core_uart_div0[6]), 
        .Y(n27107) );
  sky130_fd_sc_hd__nor2_1 U32026 ( .A(n28590), .B(n27110), .Y(
        j202_soc_core_wbqspiflash_00_N717) );
  sky130_fd_sc_hd__nor2_1 U32027 ( .A(n28590), .B(n28150), .Y(
        j202_soc_core_wbqspiflash_00_N711) );
  sky130_fd_sc_hd__nor2_1 U32028 ( .A(n28590), .B(n27111), .Y(
        j202_soc_core_wbqspiflash_00_N712) );
  sky130_fd_sc_hd__xor2_1 U32029 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[1]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]), .X(n27115) );
  sky130_fd_sc_hd__xor2_1 U32030 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[2]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .X(n27114) );
  sky130_fd_sc_hd__xor2_1 U32031 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[7]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]), .X(n27113) );
  sky130_fd_sc_hd__xor2_1 U32032 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[0]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]), .X(n27112) );
  sky130_fd_sc_hd__nor4_1 U32033 ( .A(n27115), .B(n27114), .C(n27113), .D(
        n27112), .Y(n27121) );
  sky130_fd_sc_hd__xor2_1 U32034 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[4]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]), .X(n27117) );
  sky130_fd_sc_hd__xor2_1 U32035 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[3]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .X(n27116) );
  sky130_fd_sc_hd__nor3_1 U32036 ( .A(n27117), .B(n27116), .C(n28232), .Y(
        n27120) );
  sky130_fd_sc_hd__xnor2_1 U32037 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[5]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]), .Y(n27119) );
  sky130_fd_sc_hd__xnor2_1 U32038 ( .A(
        j202_soc_core_wbqspiflash_00_erased_sector[6]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .Y(n27118) );
  sky130_fd_sc_hd__nand4_1 U32039 ( .A(n27121), .B(n27120), .C(n27119), .D(
        n27118), .Y(n27122) );
  sky130_fd_sc_hd__nand2_1 U32040 ( .A(n27123), .B(n27122), .Y(
        j202_soc_core_wbqspiflash_00_N719) );
  sky130_fd_sc_hd__a22o_1 U32041 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[30]), .A2(n27719), .B1(n27718), 
        .B2(j202_soc_core_wbqspiflash_00_dirty_sector), .X(
        j202_soc_core_wbqspiflash_00_N697) );
  sky130_fd_sc_hd__o22ai_1 U32042 ( .A1(n11141), .A2(n27125), .B1(n27124), 
        .B2(n27127), .Y(j202_soc_core_j22_cpu_rf_N2694) );
  sky130_fd_sc_hd__nand2_1 U32043 ( .A(n27360), .B(n27460), .Y(n27126) );
  sky130_fd_sc_hd__nand3_1 U32045 ( .A(n29065), .B(n27129), .C(n29064), .Y(
        n27130) );
  sky130_fd_sc_hd__inv_1 U32046 ( .A(n27130), .Y(j202_soc_core_ahb2aqu_00_N98)
         );
  sky130_fd_sc_hd__a21oi_1 U32047 ( .A1(n27137), .A2(n27141), .B1(n27131), .Y(
        n94) );
  sky130_fd_sc_hd__a21oi_1 U32049 ( .A1(n27134), .A2(n27133), .B1(n29355), .Y(
        n130) );
  sky130_fd_sc_hd__nor2_1 U32050 ( .A(n27137), .B(n27135), .Y(n27136) );
  sky130_fd_sc_hd__a21oi_1 U32051 ( .A1(n27140), .A2(n27137), .B1(n27136), .Y(
        n27139) );
  sky130_fd_sc_hd__o211ai_1 U32052 ( .A1(j202_soc_core_uart_TOP_rx_fifo_wp[0]), 
        .A2(n27140), .B1(n27139), .C1(n27138), .Y(n27142) );
  sky130_fd_sc_hd__nor2_1 U32053 ( .A(n28590), .B(n27142), .Y(
        j202_soc_core_uart_TOP_rx_fifo_N42) );
  sky130_fd_sc_hd__nand3_1 U32054 ( .A(n27142), .B(n29593), .C(n27141), .Y(
        j202_soc_core_uart_TOP_rx_fifo_N41) );
  sky130_fd_sc_hd__nand2_1 U32055 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[8]), .Y(n27143) );
  sky130_fd_sc_hd__o21ai_1 U32056 ( .A1(n27145), .A2(n27827), .B1(n27143), .Y(
        n116) );
  sky130_fd_sc_hd__nand2_1 U32057 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[8]), .Y(n27144) );
  sky130_fd_sc_hd__o21ai_1 U32058 ( .A1(n27145), .A2(n27833), .B1(n27144), .Y(
        n117) );
  sky130_fd_sc_hd__a22oi_1 U32059 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[8]), .B1(n27837), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[8]), .Y(
        n27148) );
  sky130_fd_sc_hd__nand2_1 U32060 ( .A(n27840), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[8]), .Y(
        n27147) );
  sky130_fd_sc_hd__nand2_1 U32061 ( .A(n27835), .B(
        j202_soc_core_cmt_core_00_const1[8]), .Y(n27146) );
  sky130_fd_sc_hd__nand3_1 U32062 ( .A(n27148), .B(n27147), .C(n27146), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[8]) );
  sky130_fd_sc_hd__nand2_1 U32063 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[8]), .Y(n27149) );
  sky130_fd_sc_hd__o21ai_1 U32064 ( .A1(n27150), .A2(n27983), .B1(n27149), .Y(
        n57) );
  sky130_fd_sc_hd__o22ai_1 U32065 ( .A1(n28599), .A2(n27990), .B1(n27151), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U32066 ( .A1(n27154), .A2(n27153), .B1(n28326), 
        .B2(n27152), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U32067 ( .A1(n27757), .A2(n27155), .B1(n28326), 
        .B2(n27754), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U32068 ( .A1(n28541), .A2(n28599), .B1(n27156), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__a22oi_1 U32069 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[8]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[72]), .Y(n27158) );
  sky130_fd_sc_hd__a22oi_1 U32070 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[8]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[8]), .Y(n27157) );
  sky130_fd_sc_hd__nand3_1 U32071 ( .A(n27158), .B(n27157), .C(n27865), .Y(
        n27159) );
  sky130_fd_sc_hd__a21oi_1 U32072 ( .A1(j202_soc_core_intc_core_00_rg_itgt[10]), .A2(n27869), .B1(n27159), .Y(n27163) );
  sky130_fd_sc_hd__a22oi_1 U32073 ( .A1(n27856), .A2(
        j202_soc_core_intc_core_00_rg_itgt[18]), .B1(n27850), .B2(
        j202_soc_core_intc_core_00_rg_itgt[2]), .Y(n27162) );
  sky130_fd_sc_hd__a22oi_1 U32074 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[26]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[104]), .Y(n27161) );
  sky130_fd_sc_hd__nand2_1 U32075 ( .A(n27862), .B(
        j202_soc_core_intc_core_00_rg_ipr[40]), .Y(n27160) );
  sky130_fd_sc_hd__nand4_1 U32076 ( .A(n27163), .B(n27162), .C(n27161), .D(
        n27160), .Y(j202_soc_core_ahb2apb_01_N136) );
  sky130_fd_sc_hd__nand4_1 U32077 ( .A(n27167), .B(n27166), .C(n27165), .D(
        n27164), .Y(n10536) );
  sky130_fd_sc_hd__nand3_1 U32078 ( .A(n27171), .B(n27686), .C(n27170), .Y(
        n27172) );
  sky130_fd_sc_hd__nand2_1 U32079 ( .A(n27174), .B(n27173), .Y(n27179) );
  sky130_fd_sc_hd__nand4_1 U32080 ( .A(n27177), .B(n27176), .C(n27175), .D(
        n27942), .Y(n27178) );
  sky130_fd_sc_hd__a21oi_1 U32081 ( .A1(n27179), .A2(n27980), .B1(n27178), .Y(
        n27180) );
  sky130_fd_sc_hd__nand2_1 U32082 ( .A(n27181), .B(n27180), .Y(n10583) );
  sky130_fd_sc_hd__a22oi_1 U32083 ( .A1(n27184), .A2(n27183), .B1(n29549), 
        .B2(n27339), .Y(n27185) );
  sky130_fd_sc_hd__nand2_1 U32084 ( .A(n27346), .B(n27185), .Y(
        j202_soc_core_j22_cpu_ml_N325) );
  sky130_fd_sc_hd__a22oi_1 U32085 ( .A1(n27187), .A2(n22112), .B1(n27273), 
        .B2(n27186), .Y(n27188) );
  sky130_fd_sc_hd__nand2_1 U32086 ( .A(n27189), .B(n27188), .Y(
        j202_soc_core_j22_cpu_ml_machj[21]) );
  sky130_fd_sc_hd__nand2_1 U32087 ( .A(n27190), .B(n27192), .Y(n27191) );
  sky130_fd_sc_hd__o22ai_1 U32089 ( .A1(n28615), .A2(n27194), .B1(n27201), 
        .B2(n27193), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__a21oi_1 U32090 ( .A1(n27196), .A2(n27195), .B1(
        j202_soc_core_intc_core_00_rg_irqc[2]), .Y(n27199) );
  sky130_fd_sc_hd__nor2_1 U32091 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[2]), 
        .B(n27197), .Y(n27198) );
  sky130_fd_sc_hd__a31oi_1 U32092 ( .A1(n27199), .A2(
        j202_soc_core_intc_core_00_in_intreq[2]), .A3(n29594), .B1(n27198), 
        .Y(n27200) );
  sky130_fd_sc_hd__nor2_1 U32093 ( .A(n27201), .B(n27200), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N5) );
  sky130_fd_sc_hd__a22oi_1 U32094 ( .A1(n29069), .A2(n27204), .B1(n27203), 
        .B2(n11700), .Y(n27205) );
  sky130_fd_sc_hd__o21ai_1 U32095 ( .A1(n27207), .A2(n27206), .B1(n27205), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N5) );
  sky130_fd_sc_hd__o22ai_1 U32096 ( .A1(n27234), .A2(n27333), .B1(n23178), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N3052) );
  sky130_fd_sc_hd__o22ai_1 U32097 ( .A1(n27234), .A2(n27466), .B1(n27465), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N2756) );
  sky130_fd_sc_hd__o22ai_1 U32098 ( .A1(n27234), .A2(n27209), .B1(n23039), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N2719) );
  sky130_fd_sc_hd__o22ai_1 U32099 ( .A1(n27234), .A2(n27211), .B1(n27210), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N3200) );
  sky130_fd_sc_hd__o22ai_1 U32100 ( .A1(n27234), .A2(n27213), .B1(n27212), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N2793) );
  sky130_fd_sc_hd__o22ai_1 U32101 ( .A1(n27234), .A2(n27215), .B1(n27214), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N2904) );
  sky130_fd_sc_hd__o22ai_1 U32102 ( .A1(n27234), .A2(n27217), .B1(n27216), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N2830) );
  sky130_fd_sc_hd__o22ai_1 U32103 ( .A1(n27234), .A2(n27219), .B1(n27218), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N2978) );
  sky130_fd_sc_hd__o22ai_1 U32104 ( .A1(n27234), .A2(n27221), .B1(n27220), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N2867) );
  sky130_fd_sc_hd__o22ai_1 U32105 ( .A1(n27234), .A2(n27223), .B1(n27222), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N3015) );
  sky130_fd_sc_hd__o22ai_1 U32106 ( .A1(n27234), .A2(n27225), .B1(n27224), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N2941) );
  sky130_fd_sc_hd__o22ai_1 U32107 ( .A1(n27234), .A2(n27226), .B1(n23079), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N3126) );
  sky130_fd_sc_hd__o22ai_1 U32108 ( .A1(n27234), .A2(n27228), .B1(n27227), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N3163) );
  sky130_fd_sc_hd__o22ai_1 U32109 ( .A1(n13271), .A2(n27297), .B1(n27230), 
        .B2(n27229), .Y(n27231) );
  sky130_fd_sc_hd__o21ai_1 U32110 ( .A1(n27928), .A2(n27233), .B1(n27300), .Y(
        n10499) );
  sky130_fd_sc_hd__o22ai_1 U32111 ( .A1(n27234), .A2(n27575), .B1(n27574), 
        .B2(n27208), .Y(j202_soc_core_j22_cpu_rf_N3089) );
  sky130_fd_sc_hd__nand2_1 U32112 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[11]), .Y(n27235) );
  sky130_fd_sc_hd__o21ai_1 U32113 ( .A1(n27237), .A2(n27827), .B1(n27235), .Y(
        n126) );
  sky130_fd_sc_hd__nand2_1 U32114 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[11]), .Y(n27236) );
  sky130_fd_sc_hd__a22oi_1 U32116 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[11]), .B1(n27837), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[11]), 
        .Y(n27240) );
  sky130_fd_sc_hd__nand2_1 U32117 ( .A(n27840), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[11]), 
        .Y(n27239) );
  sky130_fd_sc_hd__nand2_1 U32118 ( .A(n27835), .B(
        j202_soc_core_cmt_core_00_const1[11]), .Y(n27238) );
  sky130_fd_sc_hd__nand3_1 U32119 ( .A(n27240), .B(n27239), .C(n27238), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[11]) );
  sky130_fd_sc_hd__nand2_1 U32120 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[11]), .Y(n27241) );
  sky130_fd_sc_hd__o21ai_1 U32121 ( .A1(n27242), .A2(n27983), .B1(n27241), .Y(
        n59) );
  sky130_fd_sc_hd__o22ai_1 U32122 ( .A1(n28596), .A2(n28535), .B1(n27243), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U32123 ( .A1(n28596), .A2(n28547), .B1(n27244), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__clkinv_1 U32124 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[114]), .Y(n27245) );
  sky130_fd_sc_hd__o22ai_1 U32125 ( .A1(n28596), .A2(n28538), .B1(n27245), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U32126 ( .A1(n28544), .A2(n28596), .B1(n27246), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__a22oi_1 U32127 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[11]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[107]), .Y(n27248) );
  sky130_fd_sc_hd__nand2_1 U32128 ( .A(n27864), .B(
        j202_soc_core_intc_core_00_in_intreq[11]), .Y(n27247) );
  sky130_fd_sc_hd__nand3_1 U32129 ( .A(n27865), .B(n27248), .C(n27247), .Y(
        n27253) );
  sky130_fd_sc_hd__a22o_1 U32130 ( .A1(n27856), .A2(
        j202_soc_core_intc_core_00_rg_itgt[114]), .B1(n27850), .B2(
        j202_soc_core_intc_core_00_rg_itgt[98]), .X(n27249) );
  sky130_fd_sc_hd__a21oi_1 U32131 ( .A1(j202_soc_core_intc_core_00_rg_ipr[43]), 
        .A2(n27862), .B1(n27249), .Y(n27252) );
  sky130_fd_sc_hd__a22oi_1 U32132 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[122]), .B1(n27869), .B2(
        j202_soc_core_intc_core_00_rg_itgt[106]), .Y(n27251) );
  sky130_fd_sc_hd__a22oi_1 U32133 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[11]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[75]), .Y(n27250) );
  sky130_fd_sc_hd__nand4b_1 U32134 ( .A_N(n27253), .B(n27252), .C(n27251), .D(
        n27250), .Y(j202_soc_core_ahb2apb_01_N139) );
  sky130_fd_sc_hd__nand3b_1 U32135 ( .A_N(n27880), .B(n11642), .C(n12437), .Y(
        n27254) );
  sky130_fd_sc_hd__a21oi_1 U32136 ( .A1(n27255), .A2(n29071), .B1(n27254), .Y(
        n27262) );
  sky130_fd_sc_hd__nor2_1 U32138 ( .A(n27257), .B(n12712), .Y(n27793) );
  sky130_fd_sc_hd__nand3_1 U32139 ( .A(n27262), .B(n27793), .C(n12117), .Y(
        n27263) );
  sky130_fd_sc_hd__nand2_1 U32140 ( .A(n27263), .B(n27980), .Y(n27266) );
  sky130_fd_sc_hd__nand4_1 U32141 ( .A(n27266), .B(n27572), .C(n27265), .D(
        n27947), .Y(n10591) );
  sky130_fd_sc_hd__nor2_1 U32142 ( .A(n27268), .B(n27267), .Y(
        j202_soc_core_j22_cpu_ma_N54) );
  sky130_fd_sc_hd__nand2_1 U32143 ( .A(n27269), .B(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[2]), .Y(n27270) );
  sky130_fd_sc_hd__o211ai_1 U32144 ( .A1(n27338), .A2(n27272), .B1(n27271), 
        .C1(n27270), .Y(j202_soc_core_j22_cpu_ml_N154) );
  sky130_fd_sc_hd__nand2_1 U32146 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[10]), .Y(n27277) );
  sky130_fd_sc_hd__o21ai_1 U32147 ( .A1(n27279), .A2(n27827), .B1(n27277), .Y(
        n125) );
  sky130_fd_sc_hd__nand2_1 U32148 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[10]), .Y(n27278) );
  sky130_fd_sc_hd__o21ai_1 U32149 ( .A1(n27279), .A2(n27833), .B1(n27278), .Y(
        n119) );
  sky130_fd_sc_hd__a22oi_1 U32150 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[10]), .B1(n27837), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[10]), 
        .Y(n27282) );
  sky130_fd_sc_hd__nand2_1 U32151 ( .A(n27840), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[10]), 
        .Y(n27281) );
  sky130_fd_sc_hd__nand2_1 U32152 ( .A(n27835), .B(
        j202_soc_core_cmt_core_00_const1[10]), .Y(n27280) );
  sky130_fd_sc_hd__nand3_1 U32153 ( .A(n27282), .B(n27281), .C(n27280), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[10]) );
  sky130_fd_sc_hd__o22ai_1 U32154 ( .A1(n28609), .A2(n27990), .B1(n27283), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o22ai_1 U32155 ( .A1(n28609), .A2(n28535), .B1(n27284), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o22ai_1 U32156 ( .A1(n28609), .A2(n28547), .B1(n27285), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o22ai_1 U32157 ( .A1(n28609), .A2(n28538), .B1(n27286), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o22ai_1 U32158 ( .A1(n28609), .A2(n28541), .B1(n27287), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o22ai_1 U32159 ( .A1(n28544), .A2(n28609), .B1(n27288), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__a22oi_1 U32160 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[10]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[74]), .Y(n27290) );
  sky130_fd_sc_hd__a22oi_1 U32161 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[10]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[10]), .Y(n27289) );
  sky130_fd_sc_hd__nand3_1 U32162 ( .A(n27290), .B(n27289), .C(n27865), .Y(
        n27291) );
  sky130_fd_sc_hd__a21oi_1 U32163 ( .A1(n27869), .A2(
        j202_soc_core_intc_core_00_rg_itgt[74]), .B1(n27291), .Y(n27295) );
  sky130_fd_sc_hd__a22oi_1 U32164 ( .A1(n27856), .A2(
        j202_soc_core_intc_core_00_rg_itgt[82]), .B1(n27850), .B2(
        j202_soc_core_intc_core_00_rg_itgt[66]), .Y(n27294) );
  sky130_fd_sc_hd__a22oi_1 U32165 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[90]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[106]), .Y(n27293) );
  sky130_fd_sc_hd__nand2_1 U32166 ( .A(n27862), .B(
        j202_soc_core_intc_core_00_rg_ipr[42]), .Y(n27292) );
  sky130_fd_sc_hd__nand4_1 U32167 ( .A(n27295), .B(n27294), .C(n27293), .D(
        n27292), .Y(j202_soc_core_ahb2apb_01_N138) );
  sky130_fd_sc_hd__o21ai_1 U32168 ( .A1(n27298), .A2(n27297), .B1(n27296), .Y(
        n27299) );
  sky130_fd_sc_hd__a21oi_1 U32169 ( .A1(n29072), .A2(n27882), .B1(n27299), .Y(
        n27301) );
  sky130_fd_sc_hd__o21ai_1 U32170 ( .A1(n27301), .A2(n27928), .B1(n27300), .Y(
        n10498) );
  sky130_fd_sc_hd__o22ai_1 U32171 ( .A1(n28610), .A2(n28535), .B1(n27302), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U32172 ( .A1(n28610), .A2(n28547), .B1(n27303), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U32173 ( .A1(n28610), .A2(n28538), .B1(n27304), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U32174 ( .A1(n28610), .A2(n28541), .B1(n27305), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__a22oi_1 U32175 ( .A1(n27308), .A2(
        j202_soc_core_intc_core_00_rg_eimk[7]), .B1(n27307), .B2(
        j202_soc_core_intc_core_00_rg_itgt[105]), .Y(n27310) );
  sky130_fd_sc_hd__o22ai_1 U32176 ( .A1(n27310), .A2(n28590), .B1(n27309), 
        .B2(n27764), .Y(n27315) );
  sky130_fd_sc_hd__a21oi_1 U32177 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[7]), .B1(n27758), .Y(n27311) );
  sky130_fd_sc_hd__o21ai_1 U32178 ( .A1(n27313), .A2(n27312), .B1(n27311), .Y(
        n27314) );
  sky130_fd_sc_hd__a211oi_1 U32179 ( .A1(j202_soc_core_intc_core_00_rg_ipr[7]), 
        .A2(n27851), .B1(n27315), .C1(n27314), .Y(n27319) );
  sky130_fd_sc_hd__a22oi_1 U32180 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[121]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[103]), .Y(n27318) );
  sky130_fd_sc_hd__a22oi_1 U32181 ( .A1(n27856), .A2(
        j202_soc_core_intc_core_00_rg_itgt[113]), .B1(n27850), .B2(
        j202_soc_core_intc_core_00_rg_itgt[97]), .Y(n27317) );
  sky130_fd_sc_hd__nand2_1 U32182 ( .A(n27862), .B(
        j202_soc_core_intc_core_00_rg_ipr[39]), .Y(n27316) );
  sky130_fd_sc_hd__nand4_1 U32183 ( .A(n27319), .B(n27318), .C(n27317), .D(
        n27316), .Y(j202_soc_core_ahb2apb_01_N135) );
  sky130_fd_sc_hd__nand2_1 U32184 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[7]), .Y(n27320) );
  sky130_fd_sc_hd__o21ai_1 U32185 ( .A1(n27326), .A2(n27827), .B1(n27320), .Y(
        n106) );
  sky130_fd_sc_hd__nand2_1 U32187 ( .A(n27322), .B(n27321), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_nxt_latch_status_0_) );
  sky130_fd_sc_hd__nand2_1 U32189 ( .A(n27324), .B(n27323), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_nxt_latch_status_0_) );
  sky130_fd_sc_hd__nand2_1 U32190 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[7]), .Y(n27325) );
  sky130_fd_sc_hd__a22oi_1 U32192 ( .A1(n27836), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_0_), .B1(
        n27835), .B2(j202_soc_core_cmt_core_00_const1[7]), .Y(n27330) );
  sky130_fd_sc_hd__a22oi_1 U32193 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[7]), .B1(n27837), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[7]), .Y(
        n27329) );
  sky130_fd_sc_hd__nand2_1 U32194 ( .A(n27839), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_0_), .Y(
        n27328) );
  sky130_fd_sc_hd__nand2_1 U32195 ( .A(n27840), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[7]), .Y(
        n27327) );
  sky130_fd_sc_hd__nand4_1 U32196 ( .A(n27330), .B(n27329), .C(n27328), .D(
        n27327), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[7]) );
  sky130_fd_sc_hd__nor2_1 U32197 ( .A(n28200), .B(n27874), .Y(
        j202_soc_core_wbqspiflash_00_N674) );
  sky130_fd_sc_hd__nand2_1 U32198 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[7]), .Y(n27331) );
  sky130_fd_sc_hd__o21ai_1 U32199 ( .A1(n27332), .A2(n27983), .B1(n27331), .Y(
        n56) );
  sky130_fd_sc_hd__o22ai_1 U32200 ( .A1(n27335), .A2(n27333), .B1(n23178), 
        .B2(n29565), .Y(j202_soc_core_j22_cpu_rf_N3049) );
  sky130_fd_sc_hd__mux2i_1 U32201 ( .A0(n29565), .A1(n27335), .S(n27334), .Y(
        j202_soc_core_j22_cpu_rf_N2628) );
  sky130_fd_sc_hd__o21ai_1 U32202 ( .A1(n27338), .A2(n27337), .B1(n27336), .Y(
        j202_soc_core_j22_cpu_ml_N193) );
  sky130_fd_sc_hd__nand3_1 U32203 ( .A(n27340), .B(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[3]), .C(n27339), .Y(n27345) );
  sky130_fd_sc_hd__or3_1 U32204 ( .A(n27343), .B(n27342), .C(n27341), .X(
        n27344) );
  sky130_fd_sc_hd__nand3_1 U32205 ( .A(n27346), .B(n27345), .C(n27344), .Y(
        j202_soc_core_j22_cpu_ml_N336) );
  sky130_fd_sc_hd__nand2_1 U32206 ( .A(n27347), .B(n27446), .Y(n27348) );
  sky130_fd_sc_hd__o211ai_1 U32207 ( .A1(n27349), .A2(n27450), .B1(n27348), 
        .C1(n27448), .Y(j202_soc_core_j22_cpu_ml_N370) );
  sky130_fd_sc_hd__mux2i_1 U32208 ( .A0(n27441), .A1(n27350), .S(n27456), .Y(
        n27353) );
  sky130_fd_sc_hd__nand3_1 U32209 ( .A(n27354), .B(n27351), .C(n27454), .Y(
        n27352) );
  sky130_fd_sc_hd__nand2_1 U32210 ( .A(n27353), .B(n27352), .Y(
        j202_soc_core_j22_cpu_ml_N429) );
  sky130_fd_sc_hd__nand2b_1 U32211 ( .A_N(n27456), .B(n27438), .Y(n27418) );
  sky130_fd_sc_hd__a22oi_1 U32212 ( .A1(j202_soc_core_j22_cpu_ml_bufb[31]), 
        .A2(n27456), .B1(n27354), .B2(n27454), .Y(n27355) );
  sky130_fd_sc_hd__o21ai_1 U32213 ( .A1(n27418), .A2(n27356), .B1(n27355), .Y(
        j202_soc_core_j22_cpu_ml_N427) );
  sky130_fd_sc_hd__nand2_1 U32214 ( .A(n27357), .B(n27446), .Y(n27358) );
  sky130_fd_sc_hd__o211ai_1 U32215 ( .A1(n27359), .A2(n27450), .B1(n27358), 
        .C1(n27448), .Y(j202_soc_core_j22_cpu_ml_N369) );
  sky130_fd_sc_hd__nand2_1 U32216 ( .A(n27360), .B(n27452), .Y(n27363) );
  sky130_fd_sc_hd__a22oi_1 U32217 ( .A1(j202_soc_core_j22_cpu_ml_bufb[30]), 
        .A2(n27456), .B1(n27361), .B2(n27454), .Y(n27362) );
  sky130_fd_sc_hd__nand2_1 U32218 ( .A(n27363), .B(n27362), .Y(
        j202_soc_core_j22_cpu_ml_N426) );
  sky130_fd_sc_hd__nand2_1 U32219 ( .A(n11611), .B(n27452), .Y(n27367) );
  sky130_fd_sc_hd__a22oi_1 U32220 ( .A1(j202_soc_core_j22_cpu_ml_bufb[29]), 
        .A2(n27456), .B1(n27365), .B2(n27454), .Y(n27366) );
  sky130_fd_sc_hd__nand2_1 U32221 ( .A(n27367), .B(n27366), .Y(
        j202_soc_core_j22_cpu_ml_N425) );
  sky130_fd_sc_hd__nand2_1 U32222 ( .A(n27368), .B(n27446), .Y(n27369) );
  sky130_fd_sc_hd__o211ai_1 U32223 ( .A1(n27370), .A2(n27450), .B1(n27369), 
        .C1(n27448), .Y(j202_soc_core_j22_cpu_ml_N367) );
  sky130_fd_sc_hd__nand2_1 U32224 ( .A(n27371), .B(n27452), .Y(n27374) );
  sky130_fd_sc_hd__a22oi_1 U32225 ( .A1(j202_soc_core_j22_cpu_ml_bufb[28]), 
        .A2(n27456), .B1(n27372), .B2(n27454), .Y(n27373) );
  sky130_fd_sc_hd__nand2_1 U32226 ( .A(n27374), .B(n27373), .Y(
        j202_soc_core_j22_cpu_ml_N424) );
  sky130_fd_sc_hd__o22ai_1 U32227 ( .A1(n27375), .A2(n27438), .B1(n27450), 
        .B2(n25157), .Y(n27376) );
  sky130_fd_sc_hd__nand2_1 U32228 ( .A(n11766), .B(n27452), .Y(n27379) );
  sky130_fd_sc_hd__a22oi_1 U32229 ( .A1(j202_soc_core_j22_cpu_ml_bufb[27]), 
        .A2(n27456), .B1(n27377), .B2(n27454), .Y(n27378) );
  sky130_fd_sc_hd__nand2_1 U32230 ( .A(n27379), .B(n27378), .Y(
        j202_soc_core_j22_cpu_ml_N423) );
  sky130_fd_sc_hd__o22ai_1 U32231 ( .A1(n27380), .A2(n27438), .B1(n27450), 
        .B2(n11102), .Y(n27381) );
  sky130_fd_sc_hd__nand2_1 U32232 ( .A(n12645), .B(n27452), .Y(n27385) );
  sky130_fd_sc_hd__a22oi_1 U32233 ( .A1(j202_soc_core_j22_cpu_ml_bufb[26]), 
        .A2(n27456), .B1(n27383), .B2(n27454), .Y(n27384) );
  sky130_fd_sc_hd__nand2_1 U32234 ( .A(n27385), .B(n27384), .Y(
        j202_soc_core_j22_cpu_ml_N422) );
  sky130_fd_sc_hd__nand2_1 U32235 ( .A(n12389), .B(n27452), .Y(n27391) );
  sky130_fd_sc_hd__a22oi_1 U32236 ( .A1(j202_soc_core_j22_cpu_ml_bufb[25]), 
        .A2(n27456), .B1(n27389), .B2(n27454), .Y(n27390) );
  sky130_fd_sc_hd__nand2_1 U32237 ( .A(n27391), .B(n27390), .Y(
        j202_soc_core_j22_cpu_ml_N421) );
  sky130_fd_sc_hd__nand2_1 U32238 ( .A(n27392), .B(n27446), .Y(n27393) );
  sky130_fd_sc_hd__o211ai_1 U32239 ( .A1(n27394), .A2(n27450), .B1(n27393), 
        .C1(n27448), .Y(j202_soc_core_j22_cpu_ml_N363) );
  sky130_fd_sc_hd__nand2_1 U32240 ( .A(n27395), .B(n27452), .Y(n27398) );
  sky130_fd_sc_hd__a22oi_1 U32241 ( .A1(j202_soc_core_j22_cpu_ml_bufb[24]), 
        .A2(n27456), .B1(n27396), .B2(n27454), .Y(n27397) );
  sky130_fd_sc_hd__nand2_1 U32242 ( .A(n27398), .B(n27397), .Y(
        j202_soc_core_j22_cpu_ml_N420) );
  sky130_fd_sc_hd__nand2_1 U32243 ( .A(n27399), .B(n27446), .Y(n27400) );
  sky130_fd_sc_hd__o211ai_1 U32244 ( .A1(n27401), .A2(n27450), .B1(n27400), 
        .C1(n27448), .Y(j202_soc_core_j22_cpu_ml_N362) );
  sky130_fd_sc_hd__nand2_1 U32245 ( .A(n12455), .B(n27452), .Y(n27404) );
  sky130_fd_sc_hd__a22oi_1 U32246 ( .A1(j202_soc_core_j22_cpu_ml_bufb[23]), 
        .A2(n27456), .B1(n27402), .B2(n27454), .Y(n27403) );
  sky130_fd_sc_hd__nand2_1 U32247 ( .A(n27404), .B(n27403), .Y(
        j202_soc_core_j22_cpu_ml_N419) );
  sky130_fd_sc_hd__nand2_1 U32248 ( .A(n27405), .B(n27446), .Y(n27406) );
  sky130_fd_sc_hd__o211ai_1 U32249 ( .A1(n27407), .A2(n27450), .B1(n27406), 
        .C1(n27448), .Y(j202_soc_core_j22_cpu_ml_N361) );
  sky130_fd_sc_hd__nand2_1 U32250 ( .A(n12493), .B(n27452), .Y(n27411) );
  sky130_fd_sc_hd__a22oi_1 U32251 ( .A1(j202_soc_core_j22_cpu_ml_bufb[22]), 
        .A2(n27456), .B1(n27409), .B2(n27454), .Y(n27410) );
  sky130_fd_sc_hd__nand2_1 U32252 ( .A(n27411), .B(n27410), .Y(
        j202_soc_core_j22_cpu_ml_N418) );
  sky130_fd_sc_hd__nand2_1 U32253 ( .A(n27412), .B(n27446), .Y(n27413) );
  sky130_fd_sc_hd__o211ai_1 U32254 ( .A1(n27414), .A2(n27450), .B1(n27413), 
        .C1(n27448), .Y(j202_soc_core_j22_cpu_ml_N360) );
  sky130_fd_sc_hd__a22oi_1 U32255 ( .A1(j202_soc_core_j22_cpu_ml_bufb[21]), 
        .A2(n27456), .B1(n27415), .B2(n27454), .Y(n27416) );
  sky130_fd_sc_hd__nand2_1 U32257 ( .A(n27419), .B(n27446), .Y(n27420) );
  sky130_fd_sc_hd__o211ai_1 U32258 ( .A1(n24546), .A2(n27450), .B1(n27420), 
        .C1(n27448), .Y(j202_soc_core_j22_cpu_ml_N359) );
  sky130_fd_sc_hd__nand2_1 U32259 ( .A(n11704), .B(n27452), .Y(n27424) );
  sky130_fd_sc_hd__a22oi_1 U32260 ( .A1(j202_soc_core_j22_cpu_ml_bufb[20]), 
        .A2(n27456), .B1(n27422), .B2(n27454), .Y(n27423) );
  sky130_fd_sc_hd__nand2_1 U32261 ( .A(n27424), .B(n27423), .Y(
        j202_soc_core_j22_cpu_ml_N416) );
  sky130_fd_sc_hd__nand2_1 U32262 ( .A(n27425), .B(n27446), .Y(n27426) );
  sky130_fd_sc_hd__o211ai_1 U32263 ( .A1(n27427), .A2(n27450), .B1(n27426), 
        .C1(n27448), .Y(j202_soc_core_j22_cpu_ml_N357) );
  sky130_fd_sc_hd__nand2_1 U32264 ( .A(n12120), .B(n27452), .Y(n27431) );
  sky130_fd_sc_hd__a22oi_1 U32265 ( .A1(j202_soc_core_j22_cpu_ml_bufb[19]), 
        .A2(n27456), .B1(n27429), .B2(n27454), .Y(n27430) );
  sky130_fd_sc_hd__nand2_1 U32266 ( .A(n27431), .B(n27430), .Y(
        j202_soc_core_j22_cpu_ml_N415) );
  sky130_fd_sc_hd__nand2_1 U32267 ( .A(n27432), .B(n27446), .Y(n27433) );
  sky130_fd_sc_hd__o211ai_1 U32268 ( .A1(n27434), .A2(n27450), .B1(n27433), 
        .C1(n27448), .Y(j202_soc_core_j22_cpu_ml_N356) );
  sky130_fd_sc_hd__a22oi_1 U32269 ( .A1(j202_soc_core_j22_cpu_ml_bufb[18]), 
        .A2(n27456), .B1(n27435), .B2(n27454), .Y(n27436) );
  sky130_fd_sc_hd__nand2_1 U32270 ( .A(n27437), .B(n27436), .Y(
        j202_soc_core_j22_cpu_ml_N414) );
  sky130_fd_sc_hd__o22ai_1 U32271 ( .A1(n27439), .A2(n27438), .B1(n27450), 
        .B2(n11103), .Y(n27440) );
  sky130_fd_sc_hd__nand2_1 U32272 ( .A(n27442), .B(n27452), .Y(n27445) );
  sky130_fd_sc_hd__a22oi_1 U32273 ( .A1(j202_soc_core_j22_cpu_ml_bufb[17]), 
        .A2(n27456), .B1(n27443), .B2(n27454), .Y(n27444) );
  sky130_fd_sc_hd__nand2_1 U32274 ( .A(n27445), .B(n27444), .Y(
        j202_soc_core_j22_cpu_ml_N413) );
  sky130_fd_sc_hd__nand2_1 U32275 ( .A(n27447), .B(n27446), .Y(n27449) );
  sky130_fd_sc_hd__o211ai_1 U32276 ( .A1(n27451), .A2(n27450), .B1(n27449), 
        .C1(n27448), .Y(j202_soc_core_j22_cpu_ml_N354) );
  sky130_fd_sc_hd__nand2_1 U32277 ( .A(n12417), .B(n27452), .Y(n27458) );
  sky130_fd_sc_hd__a22oi_1 U32278 ( .A1(j202_soc_core_j22_cpu_ml_bufb[16]), 
        .A2(n27456), .B1(n27455), .B2(n27454), .Y(n27457) );
  sky130_fd_sc_hd__nand2_1 U32279 ( .A(n27458), .B(n27457), .Y(
        j202_soc_core_j22_cpu_ml_N412) );
  sky130_fd_sc_hd__mux2i_1 U32280 ( .A0(n27462), .A1(n27461), .S(n27460), .Y(
        j202_soc_core_j22_cpu_rf_N3284) );
  sky130_fd_sc_hd__o22ai_1 U32281 ( .A1(n27466), .A2(n27464), .B1(n27465), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N2764) );
  sky130_fd_sc_hd__o22ai_1 U32282 ( .A1(n27467), .A2(n27466), .B1(n27465), 
        .B2(n11120), .Y(j202_soc_core_j22_cpu_rf_N2760) );
  sky130_fd_sc_hd__nand2_1 U32283 ( .A(n27468), .B(
        j202_soc_core_cmt_core_00_cnt0[12]), .Y(n27474) );
  sky130_fd_sc_hd__nand2_1 U32284 ( .A(j202_soc_core_cmt_core_00_cnt0[12]), 
        .B(j202_soc_core_cmt_core_00_cnt0[13]), .Y(n27470) );
  sky130_fd_sc_hd__a21o_1 U32285 ( .A1(n27471), .A2(n27470), .B1(n27469), .X(
        n27479) );
  sky130_fd_sc_hd__o21ai_1 U32286 ( .A1(j202_soc_core_cmt_core_00_cnt0[13]), 
        .A2(n27481), .B1(n27479), .Y(n27472) );
  sky130_fd_sc_hd__nor3_1 U32288 ( .A(j202_soc_core_cmt_core_00_cnt0[14]), .B(
        n27475), .C(n27474), .Y(n27478) );
  sky130_fd_sc_hd__a21oi_1 U32289 ( .A1(n27482), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[14]), .B1(n27478), .Y(n27477) );
  sky130_fd_sc_hd__nand2_1 U32290 ( .A(n27479), .B(
        j202_soc_core_cmt_core_00_cnt0[14]), .Y(n27476) );
  sky130_fd_sc_hd__nand2_1 U32291 ( .A(n27477), .B(n27476), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[14]) );
  sky130_fd_sc_hd__nand4_1 U32293 ( .A(n27481), .B(
        j202_soc_core_cmt_core_00_cnt0[13]), .C(
        j202_soc_core_cmt_core_00_cnt0[14]), .D(n27480), .Y(n27484) );
  sky130_fd_sc_hd__nand2_1 U32294 ( .A(n27482), .B(
        j202_soc_core_cmt_core_00_wdata_cnt0[15]), .Y(n27483) );
  sky130_fd_sc_hd__nand3_1 U32295 ( .A(n27485), .B(n27484), .C(n27483), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[15]) );
  sky130_fd_sc_hd__nand2_1 U32296 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[15]), .Y(n27486) );
  sky130_fd_sc_hd__o21ai_1 U32297 ( .A1(n27503), .A2(n27827), .B1(n27486), .Y(
        n124) );
  sky130_fd_sc_hd__a31oi_1 U32298 ( .A1(n27487), .A2(
        j202_soc_core_cmt_core_00_cnt1[12]), .A3(n27489), .B1(
        j202_soc_core_cmt_core_00_cnt1[13]), .Y(n27490) );
  sky130_fd_sc_hd__nand2_1 U32299 ( .A(j202_soc_core_cmt_core_00_cnt1[12]), 
        .B(j202_soc_core_cmt_core_00_cnt1[13]), .Y(n27493) );
  sky130_fd_sc_hd__a21oi_1 U32300 ( .A1(n27489), .A2(n27493), .B1(n27488), .Y(
        n27500) );
  sky130_fd_sc_hd__o22ai_1 U32301 ( .A1(n27799), .A2(n27491), .B1(n27490), 
        .B2(n27500), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[13])
         );
  sky130_fd_sc_hd__nor2_1 U32302 ( .A(n27493), .B(n27492), .Y(n27497) );
  sky130_fd_sc_hd__a22oi_1 U32303 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[14]), .A2(n27498), .B1(n27497), 
        .B2(n27495), .Y(n27494) );
  sky130_fd_sc_hd__o21ai_1 U32304 ( .A1(n27495), .A2(n27500), .B1(n27494), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[14]) );
  sky130_fd_sc_hd__xnor2_1 U32305 ( .A(j202_soc_core_cmt_core_00_cnt1[15]), 
        .B(n27495), .Y(n27496) );
  sky130_fd_sc_hd__a22oi_1 U32306 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[15]), .A2(n27498), .B1(n27497), 
        .B2(n27496), .Y(n27499) );
  sky130_fd_sc_hd__nand2_1 U32308 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[15]), .Y(n27502) );
  sky130_fd_sc_hd__o21ai_1 U32309 ( .A1(n27503), .A2(n27833), .B1(n27502), .Y(
        n118) );
  sky130_fd_sc_hd__a22oi_1 U32310 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[15]), .B1(n27837), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[15]), 
        .Y(n27506) );
  sky130_fd_sc_hd__nand2_1 U32311 ( .A(n27840), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[15]), 
        .Y(n27505) );
  sky130_fd_sc_hd__nand2_1 U32312 ( .A(n27835), .B(
        j202_soc_core_cmt_core_00_const1[15]), .Y(n27504) );
  sky130_fd_sc_hd__nand3_1 U32313 ( .A(n27506), .B(n27505), .C(n27504), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[15]) );
  sky130_fd_sc_hd__nand2_1 U32314 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[15]), .Y(n27507) );
  sky130_fd_sc_hd__o21ai_1 U32315 ( .A1(n27508), .A2(n27983), .B1(n27507), .Y(
        n63) );
  sky130_fd_sc_hd__o22ai_1 U32316 ( .A1(n28607), .A2(n27990), .B1(n27509), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U32317 ( .A1(n28607), .A2(n28535), .B1(n27510), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U32318 ( .A1(n28607), .A2(n28547), .B1(n27511), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U32319 ( .A1(n28607), .A2(n28538), .B1(n27512), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U32320 ( .A1(n28607), .A2(n28541), .B1(n27513), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U32321 ( .A1(n28544), .A2(n28607), .B1(n27514), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__a22oi_1 U32322 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[15]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[79]), .Y(n27516) );
  sky130_fd_sc_hd__a22oi_1 U32323 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[15]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[15]), .Y(n27515) );
  sky130_fd_sc_hd__nand3_1 U32324 ( .A(n27516), .B(n27515), .C(n27865), .Y(
        n27517) );
  sky130_fd_sc_hd__a21oi_1 U32325 ( .A1(n27869), .A2(
        j202_soc_core_intc_core_00_rg_itgt[107]), .B1(n27517), .Y(n27521) );
  sky130_fd_sc_hd__a22oi_1 U32326 ( .A1(n27856), .A2(
        j202_soc_core_intc_core_00_rg_itgt[115]), .B1(n27850), .B2(
        j202_soc_core_intc_core_00_rg_itgt[99]), .Y(n27520) );
  sky130_fd_sc_hd__a22oi_1 U32327 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[123]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[111]), .Y(n27519) );
  sky130_fd_sc_hd__nand2_1 U32328 ( .A(n27862), .B(
        j202_soc_core_intc_core_00_rg_ipr[47]), .Y(n27518) );
  sky130_fd_sc_hd__nand4_1 U32329 ( .A(n27521), .B(n27520), .C(n27519), .D(
        n27518), .Y(j202_soc_core_ahb2apb_01_N143) );
  sky130_fd_sc_hd__a22o_1 U32330 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[15]), .A2(n27719), .B1(n27718), 
        .B2(j202_soc_core_wbqspiflash_00_erased_sector[1]), .X(
        j202_soc_core_wbqspiflash_00_N682) );
  sky130_fd_sc_hd__nand2_1 U32331 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[6]), .Y(n27525) );
  sky130_fd_sc_hd__o21ai_1 U32332 ( .A1(n27527), .A2(n27827), .B1(n27525), .Y(
        n104) );
  sky130_fd_sc_hd__nand2_1 U32333 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[6]), .Y(n27526) );
  sky130_fd_sc_hd__o21ai_1 U32334 ( .A1(n27527), .A2(n27833), .B1(n27526), .Y(
        n105) );
  sky130_fd_sc_hd__a22oi_1 U32335 ( .A1(n27836), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[6]), .B1(n27835), .B2(
        j202_soc_core_cmt_core_00_const1[6]), .Y(n27531) );
  sky130_fd_sc_hd__a22oi_1 U32336 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[6]), .B1(n27837), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[6]), .Y(
        n27530) );
  sky130_fd_sc_hd__nand2_1 U32337 ( .A(n27839), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[6]), .Y(n27529) );
  sky130_fd_sc_hd__nand2_1 U32338 ( .A(n27840), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[6]), .Y(
        n27528) );
  sky130_fd_sc_hd__nand4_1 U32339 ( .A(n27531), .B(n27530), .C(n27529), .D(
        n27528), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[6]) );
  sky130_fd_sc_hd__nand2_1 U32340 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[6]), .Y(n27532) );
  sky130_fd_sc_hd__o21ai_1 U32341 ( .A1(n27533), .A2(n27983), .B1(n27532), .Y(
        n55) );
  sky130_fd_sc_hd__o22ai_1 U32342 ( .A1(n28611), .A2(n28535), .B1(n27540), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U32343 ( .A1(n28611), .A2(n28526), .B1(n27534), 
        .B2(n28524), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U32344 ( .A1(n28611), .A2(n28547), .B1(n27535), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U32345 ( .A1(n28611), .A2(n28538), .B1(n27536), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U32346 ( .A1(n28611), .A2(n28541), .B1(n27537), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U32347 ( .A1(n28544), .A2(n28611), .B1(n27538), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__a21oi_1 U32348 ( .A1(n27857), .A2(
        j202_soc_core_intc_core_00_rg_eimk[6]), .B1(n27758), .Y(n27539) );
  sky130_fd_sc_hd__a21oi_1 U32350 ( .A1(n27860), .A2(
        j202_soc_core_intc_core_00_rg_ipr[102]), .B1(n27541), .Y(n27548) );
  sky130_fd_sc_hd__a22oi_1 U32351 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[6]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[6]), .Y(n27543) );
  sky130_fd_sc_hd__a22oi_1 U32352 ( .A1(n27852), .A2(
        j202_soc_core_intc_core_00_rg_ipr[70]), .B1(n27856), .B2(
        j202_soc_core_intc_core_00_rg_itgt[81]), .Y(n27542) );
  sky130_fd_sc_hd__o211ai_1 U32353 ( .A1(n27544), .A2(n27676), .B1(n27543), 
        .C1(n27542), .Y(n27545) );
  sky130_fd_sc_hd__a21oi_1 U32354 ( .A1(n27869), .A2(
        j202_soc_core_intc_core_00_rg_itgt[73]), .B1(n27545), .Y(n27547) );
  sky130_fd_sc_hd__a22oi_1 U32355 ( .A1(n27862), .A2(
        j202_soc_core_intc_core_00_rg_ipr[38]), .B1(n27861), .B2(
        j202_soc_core_intc_core_00_rg_itgt[89]), .Y(n27546) );
  sky130_fd_sc_hd__nand3_1 U32356 ( .A(n27548), .B(n27547), .C(n27546), .Y(
        j202_soc_core_ahb2apb_01_N134) );
  sky130_fd_sc_hd__nor2_1 U32357 ( .A(n27549), .B(n27874), .Y(
        j202_soc_core_wbqspiflash_00_N673) );
  sky130_fd_sc_hd__nand2_1 U32358 ( .A(n27551), .B(n12731), .Y(n27552) );
  sky130_fd_sc_hd__a21oi_1 U32359 ( .A1(n27555), .A2(n13180), .B1(n27554), .Y(
        n27570) );
  sky130_fd_sc_hd__nand2_1 U32360 ( .A(n27556), .B(n29532), .Y(n27557) );
  sky130_fd_sc_hd__nand2_1 U32361 ( .A(n27559), .B(n27558), .Y(n27560) );
  sky130_fd_sc_hd__a21oi_1 U32362 ( .A1(n27595), .A2(n29075), .B1(n27562), .Y(
        n27569) );
  sky130_fd_sc_hd__o211ai_1 U32363 ( .A1(n12658), .A2(n27565), .B1(n27564), 
        .C1(n27563), .Y(n27567) );
  sky130_fd_sc_hd__nor2_1 U32364 ( .A(n27568), .B(n27567), .Y(n27597) );
  sky130_fd_sc_hd__nand2_1 U32365 ( .A(n27573), .B(n27572), .Y(n10594) );
  sky130_fd_sc_hd__o22ai_1 U32366 ( .A1(n27576), .A2(n27575), .B1(n27574), 
        .B2(n24644), .Y(j202_soc_core_j22_cpu_rf_N3088) );
  sky130_fd_sc_hd__nand2_1 U32367 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[20]), .Y(n27577) );
  sky130_fd_sc_hd__o21ai_1 U32368 ( .A1(n27578), .A2(n27983), .B1(n27577), .Y(
        n66) );
  sky130_fd_sc_hd__o22ai_1 U32369 ( .A1(n28604), .A2(n27990), .B1(n27579), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U32370 ( .A1(n27757), .A2(n27580), .B1(n28412), 
        .B2(n27754), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U32371 ( .A1(n27583), .A2(n27582), .B1(n28412), 
        .B2(n27581), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U32372 ( .A1(n28541), .A2(n28604), .B1(n27584), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__a22oi_1 U32373 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[20]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[84]), .Y(n27586) );
  sky130_fd_sc_hd__a22oi_1 U32374 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[20]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[20]), .Y(n27585) );
  sky130_fd_sc_hd__nand3_1 U32375 ( .A(n27586), .B(n27585), .C(n27865), .Y(
        n27587) );
  sky130_fd_sc_hd__a21oi_1 U32376 ( .A1(j202_soc_core_intc_core_00_rg_itgt[13]), .A2(n27869), .B1(n27587), .Y(n27591) );
  sky130_fd_sc_hd__a22oi_1 U32377 ( .A1(n27856), .A2(
        j202_soc_core_intc_core_00_rg_itgt[21]), .B1(n27850), .B2(
        j202_soc_core_intc_core_00_rg_itgt[5]), .Y(n27590) );
  sky130_fd_sc_hd__a22oi_1 U32378 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[29]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[116]), .Y(n27589) );
  sky130_fd_sc_hd__nand2_1 U32379 ( .A(n27862), .B(
        j202_soc_core_intc_core_00_rg_ipr[52]), .Y(n27588) );
  sky130_fd_sc_hd__nand4_1 U32380 ( .A(n27591), .B(n27590), .C(n27589), .D(
        n27588), .Y(j202_soc_core_ahb2apb_01_N148) );
  sky130_fd_sc_hd__nand2_1 U32381 ( .A(n27593), .B(j202_soc_core_uart_div1[4]), 
        .Y(n27592) );
  sky130_fd_sc_hd__o21ai_1 U32382 ( .A1(n27594), .A2(n27593), .B1(n27592), .Y(
        n109) );
  sky130_fd_sc_hd__a22o_1 U32383 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[20]), .A2(n27719), .B1(n27718), 
        .B2(j202_soc_core_wbqspiflash_00_erased_sector[6]), .X(
        j202_soc_core_wbqspiflash_00_N687) );
  sky130_fd_sc_hd__nand2_1 U32384 ( .A(n27597), .B(n27596), .Y(n27598) );
  sky130_fd_sc_hd__nand2_1 U32385 ( .A(n27598), .B(n27980), .Y(n27600) );
  sky130_fd_sc_hd__nand2_1 U32386 ( .A(n27600), .B(n27599), .Y(n10599) );
  sky130_fd_sc_hd__a31oi_1 U32387 ( .A1(n27823), .A2(n29593), .A3(n27602), 
        .B1(n27601), .Y(n10541) );
  sky130_fd_sc_hd__nand2_1 U32388 ( .A(n27604), .B(n27603), .Y(n27724) );
  sky130_fd_sc_hd__nand2_1 U32389 ( .A(n27724), .B(
        j202_soc_core_bldc_core_00_adc_en), .Y(n27605) );
  sky130_fd_sc_hd__o21ai_1 U32390 ( .A1(n27618), .A2(n27724), .B1(n27605), .Y(
        n39) );
  sky130_fd_sc_hd__nand2_1 U32391 ( .A(n29076), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[1]), .Y(n27606) );
  sky130_fd_sc_hd__nand2_1 U32393 ( .A(n27728), .B(
        j202_soc_core_bldc_core_00_comm[1]), .Y(n27608) );
  sky130_fd_sc_hd__o21ai_1 U32394 ( .A1(n27618), .A2(n27728), .B1(n27608), .Y(
        n40) );
  sky130_fd_sc_hd__nand2_1 U32395 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[1]), .Y(n27609) );
  sky130_fd_sc_hd__o21ai_1 U32396 ( .A1(n27611), .A2(n27827), .B1(n27609), .Y(
        n35) );
  sky130_fd_sc_hd__nand2_1 U32397 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[1]), .Y(n27610) );
  sky130_fd_sc_hd__o21ai_1 U32398 ( .A1(n27611), .A2(n27833), .B1(n27610), .Y(
        n36) );
  sky130_fd_sc_hd__a22oi_1 U32399 ( .A1(n27839), .A2(
        j202_soc_core_cmt_core_00_cks0[1]), .B1(n27840), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[1]), .Y(
        n27616) );
  sky130_fd_sc_hd__a22oi_1 U32400 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[1]), .B1(n27835), .B2(
        j202_soc_core_cmt_core_00_const1[1]), .Y(n27615) );
  sky130_fd_sc_hd__and3_1 U32401 ( .A(n27733), .B(
        j202_soc_core_cmt_core_00_str1), .C(n27732), .X(n27612) );
  sky130_fd_sc_hd__a21oi_1 U32402 ( .A1(n27837), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[1]), 
        .B1(n27612), .Y(n27614) );
  sky130_fd_sc_hd__nand2_1 U32403 ( .A(n27836), .B(
        j202_soc_core_cmt_core_00_cks1[1]), .Y(n27613) );
  sky130_fd_sc_hd__nand4_1 U32404 ( .A(n27616), .B(n27615), .C(n27614), .D(
        n27613), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[1]) );
  sky130_fd_sc_hd__nand2_1 U32405 ( .A(n27740), .B(
        j202_soc_core_bldc_core_00_pwm_period[1]), .Y(n27617) );
  sky130_fd_sc_hd__o21ai_1 U32406 ( .A1(n27618), .A2(n27740), .B1(n27617), .Y(
        n38) );
  sky130_fd_sc_hd__nand2_1 U32407 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[0]), 
        .B(j202_soc_core_ahb2apb_02_hsize_buf[1]), .Y(
        j202_soc_core_ahb2apb_02_N123) );
  sky130_fd_sc_hd__clkinv_1 U32408 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[0]), 
        .Y(n27627) );
  sky130_fd_sc_hd__nand2_1 U32409 ( .A(n27629), .B(n27627), .Y(n27626) );
  sky130_fd_sc_hd__nor2_1 U32410 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[1]), 
        .B(n27627), .Y(n27630) );
  sky130_fd_sc_hd__clkinv_1 U32411 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[1]), 
        .Y(n27624) );
  sky130_fd_sc_hd__nor2_1 U32412 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[0]), 
        .B(n27624), .Y(n27628) );
  sky130_fd_sc_hd__a21oi_1 U32413 ( .A1(j202_soc_core_gpio_core_00_reg_addr[1]), .A2(n27630), .B1(n27628), .Y(n27625) );
  sky130_fd_sc_hd__o21ai_0 U32414 ( .A1(j202_soc_core_gpio_core_00_reg_addr[0]), .A2(n27626), .B1(n27625), .Y(n10907) );
  sky130_fd_sc_hd__o21ai_0 U32415 ( .A1(n27626), .A2(n27633), .B1(n27625), .Y(
        n10906) );
  sky130_fd_sc_hd__nand2_1 U32416 ( .A(j202_soc_core_gpio_core_00_reg_addr[1]), 
        .B(n27627), .Y(n27632) );
  sky130_fd_sc_hd__a21oi_1 U32417 ( .A1(n27630), .A2(n27629), .B1(n27628), .Y(
        n27631) );
  sky130_fd_sc_hd__o21ai_0 U32418 ( .A1(j202_soc_core_gpio_core_00_reg_addr[0]), .A2(n27632), .B1(n27631), .Y(n10905) );
  sky130_fd_sc_hd__o21ai_0 U32419 ( .A1(n27633), .A2(n27632), .B1(n27631), .Y(
        n10904) );
  sky130_fd_sc_hd__a21oi_1 U32420 ( .A1(n12142), .A2(n28273), .B1(n28476), .Y(
        n27646) );
  sky130_fd_sc_hd__o22ai_1 U32421 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[1]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]), .B1(n27642), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[1]), .Y(n27643)
         );
  sky130_fd_sc_hd__a21oi_1 U32422 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[1]), .B1(n27643), 
        .Y(n27644) );
  sky130_fd_sc_hd__nand4_1 U32423 ( .A(n27644), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[1]), .C(n29594), .D(
        io_oeb[1]), .Y(n27645) );
  sky130_fd_sc_hd__nor3_2 U32425 ( .A(j202_soc_core_gpio_core_00_reg_addr[3]), 
        .B(n27660), .C(n27658), .Y(n28869) );
  sky130_fd_sc_hd__or3_1 U32426 ( .A(j202_soc_core_gpio_core_00_reg_addr[2]), 
        .B(n27651), .C(n27660), .X(n27653) );
  sky130_fd_sc_hd__nor3_2 U32427 ( .A(j202_soc_core_gpio_core_00_reg_addr[4]), 
        .B(j202_soc_core_gpio_core_00_reg_addr[3]), .C(n27653), .Y(n28873) );
  sky130_fd_sc_hd__a22oi_1 U32428 ( .A1(n28869), .A2(la_data_out[1]), .B1(
        n28873), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]), 
        .Y(n27664) );
  sky130_fd_sc_hd__nand2_1 U32429 ( .A(n28876), .B(gpio_en_o[1]), .Y(n27663)
         );
  sky130_fd_sc_hd__a22oi_1 U32430 ( .A1(n28875), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[1]), .B1(n28874), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[1]), .Y(n27662) );
  sky130_fd_sc_hd__nand2_1 U32431 ( .A(n13289), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[1]), .Y(n27661) );
  sky130_fd_sc_hd__nand4_1 U32432 ( .A(n27664), .B(n27663), .C(n27662), .D(
        n27661), .Y(j202_soc_core_ahb2apb_02_N129) );
  sky130_fd_sc_hd__o22ai_1 U32433 ( .A1(n28603), .A2(n27990), .B1(n27665), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U32434 ( .A1(n28603), .A2(n28535), .B1(n27672), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U32435 ( .A1(n28603), .A2(n28526), .B1(n27666), 
        .B2(n28524), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U32436 ( .A1(n28603), .A2(n28547), .B1(n27667), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U32437 ( .A1(n28603), .A2(n28538), .B1(n27668), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U32438 ( .A1(n28603), .A2(n28541), .B1(n27669), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U32439 ( .A1(n28544), .A2(n28603), .B1(n27670), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__a21oi_1 U32440 ( .A1(n27857), .A2(
        j202_soc_core_intc_core_00_rg_eimk[1]), .B1(n27758), .Y(n27671) );
  sky130_fd_sc_hd__o21ai_1 U32441 ( .A1(n27672), .A2(n27760), .B1(n27671), .Y(
        n27673) );
  sky130_fd_sc_hd__a21oi_1 U32442 ( .A1(n27860), .A2(
        j202_soc_core_intc_core_00_rg_ipr[97]), .B1(n27673), .Y(n27681) );
  sky130_fd_sc_hd__a22oi_1 U32443 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[1]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[1]), .Y(n27675) );
  sky130_fd_sc_hd__a22oi_1 U32444 ( .A1(n27852), .A2(
        j202_soc_core_intc_core_00_rg_ipr[65]), .B1(n27856), .B2(
        j202_soc_core_intc_core_00_rg_itgt[48]), .Y(n27674) );
  sky130_fd_sc_hd__o211ai_1 U32445 ( .A1(n27677), .A2(n27676), .B1(n27675), 
        .C1(n27674), .Y(n27678) );
  sky130_fd_sc_hd__a21oi_1 U32446 ( .A1(n27869), .A2(
        j202_soc_core_intc_core_00_rg_itgt[40]), .B1(n27678), .Y(n27680) );
  sky130_fd_sc_hd__a22oi_1 U32447 ( .A1(n27862), .A2(
        j202_soc_core_intc_core_00_rg_ipr[33]), .B1(n27861), .B2(
        j202_soc_core_intc_core_00_rg_itgt[56]), .Y(n27679) );
  sky130_fd_sc_hd__nand3_1 U32448 ( .A(n27681), .B(n27680), .C(n27679), .Y(
        j202_soc_core_ahb2apb_01_N129) );
  sky130_fd_sc_hd__nor2_1 U32449 ( .A(n27682), .B(n27874), .Y(
        j202_soc_core_wbqspiflash_00_N668) );
  sky130_fd_sc_hd__nor3_1 U32450 ( .A(n27689), .B(n27688), .C(n27687), .Y(
        n27693) );
  sky130_fd_sc_hd__nand2_1 U32451 ( .A(n27694), .B(n27980), .Y(n27696) );
  sky130_fd_sc_hd__nand2_1 U32452 ( .A(n27696), .B(n27695), .Y(n10597) );
  sky130_fd_sc_hd__nand2_1 U32453 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[14]), .Y(n27697) );
  sky130_fd_sc_hd__o21ai_1 U32454 ( .A1(n27699), .A2(n27827), .B1(n27697), .Y(
        n129) );
  sky130_fd_sc_hd__nand2_1 U32455 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[14]), .Y(n27698) );
  sky130_fd_sc_hd__o21ai_1 U32456 ( .A1(n27699), .A2(n27833), .B1(n27698), .Y(
        n123) );
  sky130_fd_sc_hd__a22oi_1 U32457 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[14]), .B1(n27837), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[14]), 
        .Y(n27702) );
  sky130_fd_sc_hd__nand2_1 U32458 ( .A(n27840), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[14]), 
        .Y(n27701) );
  sky130_fd_sc_hd__nand2_1 U32459 ( .A(n27835), .B(
        j202_soc_core_cmt_core_00_const1[14]), .Y(n27700) );
  sky130_fd_sc_hd__nand3_1 U32460 ( .A(n27702), .B(n27701), .C(n27700), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[14]) );
  sky130_fd_sc_hd__nand2_1 U32461 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[14]), .Y(n27703) );
  sky130_fd_sc_hd__o21ai_1 U32462 ( .A1(n27704), .A2(n27983), .B1(n27703), .Y(
        n62) );
  sky130_fd_sc_hd__o22ai_1 U32463 ( .A1(n28597), .A2(n27990), .B1(n27705), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U32464 ( .A1(n28597), .A2(n28535), .B1(n27706), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U32465 ( .A1(n28597), .A2(n28547), .B1(n27707), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U32466 ( .A1(n28597), .A2(n28538), .B1(n27708), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U32467 ( .A1(n28597), .A2(n28541), .B1(n27709), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U32468 ( .A1(n28544), .A2(n28597), .B1(n27710), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__a22oi_1 U32469 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[14]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[78]), .Y(n27712) );
  sky130_fd_sc_hd__a22oi_1 U32470 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[14]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[14]), .Y(n27711) );
  sky130_fd_sc_hd__nand3_1 U32471 ( .A(n27712), .B(n27711), .C(n27865), .Y(
        n27713) );
  sky130_fd_sc_hd__a21oi_1 U32472 ( .A1(n27869), .A2(
        j202_soc_core_intc_core_00_rg_itgt[75]), .B1(n27713), .Y(n27717) );
  sky130_fd_sc_hd__a22oi_1 U32473 ( .A1(n27856), .A2(
        j202_soc_core_intc_core_00_rg_itgt[83]), .B1(n27850), .B2(
        j202_soc_core_intc_core_00_rg_itgt[67]), .Y(n27716) );
  sky130_fd_sc_hd__a22oi_1 U32474 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[91]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[110]), .Y(n27715) );
  sky130_fd_sc_hd__nand2_1 U32475 ( .A(n27862), .B(
        j202_soc_core_intc_core_00_rg_ipr[46]), .Y(n27714) );
  sky130_fd_sc_hd__nand4_1 U32476 ( .A(n27717), .B(n27716), .C(n27715), .D(
        n27714), .Y(j202_soc_core_ahb2apb_01_N142) );
  sky130_fd_sc_hd__a22o_1 U32477 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[14]), .A2(n27719), .B1(n27718), 
        .B2(j202_soc_core_wbqspiflash_00_erased_sector[0]), .X(
        j202_soc_core_wbqspiflash_00_N681) );
  sky130_fd_sc_hd__nand2_1 U32479 ( .A(n27724), .B(
        j202_soc_core_bldc_core_00_pwm_en), .Y(n27723) );
  sky130_fd_sc_hd__o21ai_1 U32480 ( .A1(n27741), .A2(n27724), .B1(n27723), .Y(
        n48) );
  sky130_fd_sc_hd__nand2_1 U32481 ( .A(n29076), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[0]), .Y(n27725) );
  sky130_fd_sc_hd__o21ai_1 U32482 ( .A1(n29076), .A2(n27726), .B1(n27725), .Y(
        n137) );
  sky130_fd_sc_hd__nand2_1 U32483 ( .A(n27728), .B(
        j202_soc_core_bldc_core_00_comm[0]), .Y(n27727) );
  sky130_fd_sc_hd__nand2_1 U32485 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[0]), .Y(n27729) );
  sky130_fd_sc_hd__o21ai_1 U32486 ( .A1(n27731), .A2(n27827), .B1(n27729), .Y(
        n83) );
  sky130_fd_sc_hd__nand2_1 U32487 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[0]), .Y(n27730) );
  sky130_fd_sc_hd__o21ai_1 U32488 ( .A1(n27731), .A2(n27833), .B1(n27730), .Y(
        n84) );
  sky130_fd_sc_hd__a22oi_1 U32489 ( .A1(n27839), .A2(
        j202_soc_core_cmt_core_00_cks0[0]), .B1(n27840), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[0]), .Y(
        n27738) );
  sky130_fd_sc_hd__a22oi_1 U32490 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[0]), .B1(n27835), .B2(
        j202_soc_core_cmt_core_00_const1[0]), .Y(n27737) );
  sky130_fd_sc_hd__and3_1 U32491 ( .A(n27733), .B(
        j202_soc_core_cmt_core_00_str0), .C(n27732), .X(n27734) );
  sky130_fd_sc_hd__a21oi_1 U32492 ( .A1(n27837), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[0]), 
        .B1(n27734), .Y(n27736) );
  sky130_fd_sc_hd__nand2_1 U32493 ( .A(n27836), .B(
        j202_soc_core_cmt_core_00_cks1[0]), .Y(n27735) );
  sky130_fd_sc_hd__nand4_1 U32494 ( .A(n27738), .B(n27737), .C(n27736), .D(
        n27735), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[0]) );
  sky130_fd_sc_hd__nand2_1 U32495 ( .A(n27740), .B(
        j202_soc_core_bldc_core_00_pwm_period[0]), .Y(n27739) );
  sky130_fd_sc_hd__o21ai_1 U32496 ( .A1(n27741), .A2(n27740), .B1(n27739), .Y(
        n50) );
  sky130_fd_sc_hd__nor2_1 U32497 ( .A(n28590), .B(n27742), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N3) );
  sky130_fd_sc_hd__a21oi_1 U32498 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[0]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[0]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[0]), .Y(n27746) );
  sky130_fd_sc_hd__o21ai_1 U32499 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[0]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[0]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[0]), .Y(n27743) );
  sky130_fd_sc_hd__nand4_1 U32500 ( .A(n27743), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[0]), .C(io_oeb[0]), .D(
        n12142), .Y(n27745) );
  sky130_fd_sc_hd__o21ai_1 U32502 ( .A1(n27746), .A2(n27745), .B1(n27744), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N40) );
  sky130_fd_sc_hd__a22oi_1 U32503 ( .A1(n28869), .A2(la_data_out[0]), .B1(
        n28873), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[0]), 
        .Y(n27750) );
  sky130_fd_sc_hd__nand2_1 U32504 ( .A(n28876), .B(gpio_en_o[0]), .Y(n27749)
         );
  sky130_fd_sc_hd__a22oi_1 U32505 ( .A1(n28875), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[0]), .B1(n28874), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[0]), .Y(n27748) );
  sky130_fd_sc_hd__nand2_1 U32506 ( .A(n13289), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[0]), .Y(n27747) );
  sky130_fd_sc_hd__nand4_1 U32507 ( .A(n27750), .B(n27749), .C(n27748), .D(
        n27747), .Y(j202_soc_core_ahb2apb_02_N128) );
  sky130_fd_sc_hd__o22a_1 U32508 ( .A1(j202_soc_core_intc_core_00_rg_ipr[64]), 
        .A2(n27752), .B1(n29086), .B2(n27751), .X(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U32509 ( .A1(n28881), .A2(n28526), .B1(n27753), 
        .B2(n28524), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U32510 ( .A1(n27757), .A2(n27756), .B1(n27755), 
        .B2(n27754), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__a21oi_1 U32511 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[0]), .B1(n27758), .Y(n27759) );
  sky130_fd_sc_hd__o21ai_1 U32512 ( .A1(n27761), .A2(n27760), .B1(n27759), .Y(
        n27762) );
  sky130_fd_sc_hd__a21oi_1 U32513 ( .A1(j202_soc_core_intc_core_00_rg_ipr[32]), 
        .A2(n27862), .B1(n27762), .Y(n27770) );
  sky130_fd_sc_hd__a22oi_1 U32514 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[24]), .B1(n27869), .B2(
        j202_soc_core_intc_core_00_rg_itgt[8]), .Y(n27769) );
  sky130_fd_sc_hd__a22oi_1 U32515 ( .A1(j202_soc_core_intc_core_00_rg_itgt[16]), .A2(n27856), .B1(n27860), .B2(j202_soc_core_intc_core_00_rg_ipr[96]), .Y(
        n27763) );
  sky130_fd_sc_hd__o21ai_1 U32516 ( .A1(n27765), .A2(n27764), .B1(n27763), .Y(
        n27766) );
  sky130_fd_sc_hd__a21oi_1 U32517 ( .A1(n27857), .A2(
        j202_soc_core_intc_core_00_rg_eimk[0]), .B1(n27766), .Y(n27768) );
  sky130_fd_sc_hd__a22oi_1 U32518 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[0]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[64]), .Y(n27767) );
  sky130_fd_sc_hd__nand4_1 U32519 ( .A(n27770), .B(n27769), .C(n27768), .D(
        n27767), .Y(j202_soc_core_ahb2apb_01_N128) );
  sky130_fd_sc_hd__nor2_1 U32520 ( .A(n28148), .B(n27874), .Y(
        j202_soc_core_wbqspiflash_00_N667) );
  sky130_fd_sc_hd__nand2b_1 U32521 ( .A_N(n27956), .B(n27771), .Y(n27778) );
  sky130_fd_sc_hd__nand2_1 U32522 ( .A(n27773), .B(n27772), .Y(n27775) );
  sky130_fd_sc_hd__nand2_1 U32524 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[13]), .Y(n27797) );
  sky130_fd_sc_hd__o21ai_1 U32525 ( .A1(n27799), .A2(n27827), .B1(n27797), .Y(
        n128) );
  sky130_fd_sc_hd__nand2_1 U32526 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[13]), .Y(n27798) );
  sky130_fd_sc_hd__o21ai_1 U32527 ( .A1(n27799), .A2(n27833), .B1(n27798), .Y(
        n122) );
  sky130_fd_sc_hd__a22oi_1 U32528 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[13]), .B1(n27837), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[13]), 
        .Y(n27802) );
  sky130_fd_sc_hd__nand2_1 U32529 ( .A(n27840), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[13]), 
        .Y(n27801) );
  sky130_fd_sc_hd__nand2_1 U32530 ( .A(n27835), .B(
        j202_soc_core_cmt_core_00_const1[13]), .Y(n27800) );
  sky130_fd_sc_hd__nand3_1 U32531 ( .A(n27802), .B(n27801), .C(n27800), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[13]) );
  sky130_fd_sc_hd__nand2_1 U32532 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[13]), .Y(n27803) );
  sky130_fd_sc_hd__o21ai_1 U32533 ( .A1(n27804), .A2(n27983), .B1(n27803), .Y(
        n61) );
  sky130_fd_sc_hd__o22ai_1 U32534 ( .A1(n28598), .A2(n27990), .B1(n27805), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U32535 ( .A1(n28598), .A2(n28535), .B1(n27806), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U32536 ( .A1(n28598), .A2(n28547), .B1(n27807), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__clkinv_1 U32537 ( .A(j202_soc_core_intc_core_00_rg_itgt[51]), .Y(n27808) );
  sky130_fd_sc_hd__o22ai_1 U32538 ( .A1(n28598), .A2(n28538), .B1(n27808), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U32539 ( .A1(n28544), .A2(n28598), .B1(n27809), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__a22oi_1 U32540 ( .A1(n27863), .A2(
        j202_soc_core_intc_core_00_rg_ie[13]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[109]), .Y(n27811) );
  sky130_fd_sc_hd__nand2_1 U32541 ( .A(n27864), .B(
        j202_soc_core_intc_core_00_in_intreq[13]), .Y(n27810) );
  sky130_fd_sc_hd__nand3_1 U32542 ( .A(n27865), .B(n27811), .C(n27810), .Y(
        n27816) );
  sky130_fd_sc_hd__a22o_1 U32543 ( .A1(n27856), .A2(
        j202_soc_core_intc_core_00_rg_itgt[51]), .B1(n27850), .B2(
        j202_soc_core_intc_core_00_rg_itgt[35]), .X(n27812) );
  sky130_fd_sc_hd__a21oi_1 U32544 ( .A1(j202_soc_core_intc_core_00_rg_ipr[45]), 
        .A2(n27862), .B1(n27812), .Y(n27815) );
  sky130_fd_sc_hd__a22oi_1 U32545 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[59]), .B1(n27869), .B2(
        j202_soc_core_intc_core_00_rg_itgt[43]), .Y(n27814) );
  sky130_fd_sc_hd__a22oi_1 U32546 ( .A1(n27851), .A2(
        j202_soc_core_intc_core_00_rg_ipr[13]), .B1(n27852), .B2(
        j202_soc_core_intc_core_00_rg_ipr[77]), .Y(n27813) );
  sky130_fd_sc_hd__nand4b_1 U32547 ( .A_N(n27816), .B(n27815), .C(n27814), .D(
        n27813), .Y(j202_soc_core_ahb2apb_01_N141) );
  sky130_fd_sc_hd__o21ai_1 U32548 ( .A1(j202_soc_core_j22_cpu_opst[2]), .A2(
        j202_soc_core_j22_cpu_opst[4]), .B1(j202_soc_core_j22_cpu_opst[1]), 
        .Y(n27818) );
  sky130_fd_sc_hd__o21ai_1 U32549 ( .A1(j202_soc_core_j22_cpu_opst[1]), .A2(
        n27901), .B1(n27818), .Y(n27819) );
  sky130_fd_sc_hd__nor2_1 U32550 ( .A(n27819), .B(n27956), .Y(n27940) );
  sky130_fd_sc_hd__nor2_1 U32551 ( .A(n27940), .B(n27820), .Y(n27821) );
  sky130_fd_sc_hd__o211ai_1 U32552 ( .A1(n27928), .A2(n27822), .B1(n27821), 
        .C1(n13303), .Y(n10503) );
  sky130_fd_sc_hd__nand2_1 U32553 ( .A(n27823), .B(
        j202_soc_core_ahbcs_6__HREADY_), .Y(n27825) );
  sky130_fd_sc_hd__o21ai_1 U32554 ( .A1(n27825), .A2(n27824), .B1(n12142), .Y(
        n10540) );
  sky130_fd_sc_hd__nand2_1 U32555 ( .A(n27827), .B(
        j202_soc_core_cmt_core_00_const0[3]), .Y(n27826) );
  sky130_fd_sc_hd__o21ai_1 U32556 ( .A1(n27834), .A2(n27827), .B1(n27826), .Y(
        n114) );
  sky130_fd_sc_hd__nand2_1 U32557 ( .A(n27829), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[3]), .Y(n27828) );
  sky130_fd_sc_hd__o21ai_1 U32558 ( .A1(n27834), .A2(n27829), .B1(n27828), .Y(
        n112) );
  sky130_fd_sc_hd__nand2_1 U32559 ( .A(n27831), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[3]), .Y(n27830) );
  sky130_fd_sc_hd__o21ai_1 U32560 ( .A1(n27834), .A2(n27831), .B1(n27830), .Y(
        n113) );
  sky130_fd_sc_hd__nand2_1 U32561 ( .A(n27833), .B(
        j202_soc_core_cmt_core_00_const1[3]), .Y(n27832) );
  sky130_fd_sc_hd__a22oi_1 U32563 ( .A1(n27836), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[3]), .B1(n27835), .B2(
        j202_soc_core_cmt_core_00_const1[3]), .Y(n27844) );
  sky130_fd_sc_hd__a22oi_1 U32564 ( .A1(n27838), .A2(
        j202_soc_core_cmt_core_00_const0[3]), .B1(n27837), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[3]), .Y(
        n27843) );
  sky130_fd_sc_hd__nand2_1 U32565 ( .A(n27839), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[3]), .Y(n27842) );
  sky130_fd_sc_hd__nand2_1 U32566 ( .A(n27840), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[3]), .Y(
        n27841) );
  sky130_fd_sc_hd__nand4_1 U32567 ( .A(n27844), .B(n27843), .C(n27842), .D(
        n27841), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[3]) );
  sky130_fd_sc_hd__nand2_1 U32568 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[3]), .Y(n27845) );
  sky130_fd_sc_hd__o21ai_1 U32569 ( .A1(n27846), .A2(n27983), .B1(n27845), .Y(
        n52) );
  sky130_fd_sc_hd__o22ai_1 U32570 ( .A1(n28614), .A2(n28547), .B1(n27847), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U32571 ( .A1(n28614), .A2(n28541), .B1(n27848), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U32572 ( .A1(n28544), .A2(n28614), .B1(n27849), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__nand2_1 U32573 ( .A(n27850), .B(
        j202_soc_core_intc_core_00_rg_itgt[96]), .Y(n27855) );
  sky130_fd_sc_hd__nand2_1 U32574 ( .A(n27851), .B(
        j202_soc_core_intc_core_00_rg_ipr[3]), .Y(n27854) );
  sky130_fd_sc_hd__nand2_1 U32575 ( .A(n27852), .B(
        j202_soc_core_intc_core_00_rg_ipr[67]), .Y(n27853) );
  sky130_fd_sc_hd__and3_1 U32576 ( .A(n27855), .B(n27854), .C(n27853), .X(
        n27859) );
  sky130_fd_sc_hd__a22oi_1 U32577 ( .A1(n27857), .A2(
        j202_soc_core_intc_core_00_rg_eimk[3]), .B1(n27856), .B2(
        j202_soc_core_intc_core_00_rg_itgt[112]), .Y(n27858) );
  sky130_fd_sc_hd__nand2_1 U32578 ( .A(n27859), .B(n27858), .Y(n27872) );
  sky130_fd_sc_hd__a22oi_1 U32579 ( .A1(n27861), .A2(
        j202_soc_core_intc_core_00_rg_itgt[120]), .B1(n27860), .B2(
        j202_soc_core_intc_core_00_rg_ipr[99]), .Y(n27871) );
  sky130_fd_sc_hd__nand2_1 U32580 ( .A(n27862), .B(
        j202_soc_core_intc_core_00_rg_ipr[35]), .Y(n27867) );
  sky130_fd_sc_hd__a22oi_1 U32581 ( .A1(n27864), .A2(
        j202_soc_core_intc_core_00_in_intreq[3]), .B1(n27863), .B2(
        j202_soc_core_intc_core_00_rg_ie[3]), .Y(n27866) );
  sky130_fd_sc_hd__nand3_1 U32582 ( .A(n27867), .B(n27866), .C(n27865), .Y(
        n27868) );
  sky130_fd_sc_hd__a21oi_1 U32583 ( .A1(n27869), .A2(
        j202_soc_core_intc_core_00_rg_itgt[104]), .B1(n27868), .Y(n27870) );
  sky130_fd_sc_hd__nand3b_1 U32584 ( .A_N(n27872), .B(n27871), .C(n27870), .Y(
        j202_soc_core_ahb2apb_01_N131) );
  sky130_fd_sc_hd__nor2_1 U32585 ( .A(n26211), .B(n27873), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N361) );
  sky130_fd_sc_hd__nor2_1 U32586 ( .A(n28552), .B(n27874), .Y(
        j202_soc_core_wbqspiflash_00_N670) );
  sky130_fd_sc_hd__nand2_1 U32588 ( .A(n12655), .B(n27877), .Y(n27879) );
  sky130_fd_sc_hd__nor3_1 U32589 ( .A(n12511), .B(n27879), .C(n27880), .Y(
        n27885) );
  sky130_fd_sc_hd__nand2_1 U32590 ( .A(n12466), .B(n27887), .Y(n10582) );
  sky130_fd_sc_hd__nand3_1 U32591 ( .A(n27898), .B(n27980), .C(n12677), .Y(
        n27899) );
  sky130_fd_sc_hd__a21oi_1 U32592 ( .A1(n27932), .A2(n27901), .B1(n27900), .Y(
        n27902) );
  sky130_fd_sc_hd__nand2_1 U32593 ( .A(n27905), .B(n27904), .Y(n27907) );
  sky130_fd_sc_hd__nor2_1 U32594 ( .A(n27907), .B(n27906), .Y(n27927) );
  sky130_fd_sc_hd__nand4_1 U32595 ( .A(n27912), .B(n27911), .C(n27910), .D(
        n27909), .Y(n27913) );
  sky130_fd_sc_hd__nand3_1 U32596 ( .A(n26812), .B(n27917), .C(n27916), .Y(
        n27921) );
  sky130_fd_sc_hd__nand2_1 U32597 ( .A(n27950), .B(n27921), .Y(n27977) );
  sky130_fd_sc_hd__nand2_1 U32598 ( .A(n27918), .B(j202_soc_core_intr_vec__1_), 
        .Y(n27920) );
  sky130_fd_sc_hd__a21oi_1 U32599 ( .A1(n27927), .A2(n27920), .B1(n27919), .Y(
        n27975) );
  sky130_fd_sc_hd__nand2_1 U32601 ( .A(n27975), .B(n27922), .Y(n27973) );
  sky130_fd_sc_hd__nand2_1 U32602 ( .A(n27923), .B(n27973), .Y(n10567) );
  sky130_fd_sc_hd__a21oi_1 U32603 ( .A1(n27925), .A2(n11134), .B1(n27924), .Y(
        n27926) );
  sky130_fd_sc_hd__nand2_1 U32604 ( .A(n12393), .B(n27926), .Y(n27929) );
  sky130_fd_sc_hd__nor2_1 U32605 ( .A(n27928), .B(n27927), .Y(n27933) );
  sky130_fd_sc_hd__nand2_1 U32606 ( .A(n27929), .B(n27933), .Y(n27937) );
  sky130_fd_sc_hd__a21oi_1 U32607 ( .A1(n27932), .A2(n27931), .B1(n27930), .Y(
        n27936) );
  sky130_fd_sc_hd__nand2_1 U32608 ( .A(n27934), .B(n27933), .Y(n27935) );
  sky130_fd_sc_hd__nand3_1 U32609 ( .A(n27937), .B(n27936), .C(n27935), .Y(
        n10570) );
  sky130_fd_sc_hd__nand2_1 U32610 ( .A(n27940), .B(n27978), .Y(n27941) );
  sky130_fd_sc_hd__o21bai_1 U32611 ( .A1(n27958), .A2(n27957), .B1_N(n12556), 
        .Y(n27943) );
  sky130_fd_sc_hd__nand2_1 U32612 ( .A(n27943), .B(n27980), .Y(n27953) );
  sky130_fd_sc_hd__nand3_1 U32613 ( .A(n27953), .B(n27954), .C(n27944), .Y(
        n27945) );
  sky130_fd_sc_hd__nand2_1 U32614 ( .A(n27945), .B(n27970), .Y(n27946) );
  sky130_fd_sc_hd__nand2_1 U32615 ( .A(n27946), .B(n27973), .Y(n10566) );
  sky130_fd_sc_hd__nand4_1 U32616 ( .A(n27953), .B(n27952), .C(n27951), .D(
        n27950), .Y(n27962) );
  sky130_fd_sc_hd__o21a_1 U32617 ( .A1(n27956), .A2(n27955), .B1(n27954), .X(
        n27960) );
  sky130_fd_sc_hd__nand3_1 U32618 ( .A(n11105), .B(n27980), .C(n27958), .Y(
        n27959) );
  sky130_fd_sc_hd__nand3_1 U32619 ( .A(n27961), .B(n27960), .C(n27959), .Y(
        n27971) );
  sky130_fd_sc_hd__nor2_1 U32620 ( .A(n27962), .B(n27971), .Y(n27963) );
  sky130_fd_sc_hd__nand2_1 U32621 ( .A(n27976), .B(n27963), .Y(n10569) );
  sky130_fd_sc_hd__nand2_1 U32622 ( .A(n12390), .B(n11642), .Y(n27966) );
  sky130_fd_sc_hd__nand2_1 U32623 ( .A(n27966), .B(n27980), .Y(n27968) );
  sky130_fd_sc_hd__nand2_1 U32624 ( .A(n27968), .B(n27967), .Y(n10587) );
  sky130_fd_sc_hd__o21ai_1 U32625 ( .A1(n27972), .A2(n27971), .B1(n27970), .Y(
        n27974) );
  sky130_fd_sc_hd__nand2_1 U32626 ( .A(n27974), .B(n27973), .Y(
        j202_soc_core_j22_cpu_id_idec_N894) );
  sky130_fd_sc_hd__nand2_1 U32627 ( .A(n27983), .B(
        j202_soc_core_bldc_core_00_wdata[10]), .Y(n27982) );
  sky130_fd_sc_hd__nand2_1 U32629 ( .A(n28581), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[11]), .Y(n27987) );
  sky130_fd_sc_hd__nand2_1 U32630 ( .A(n27985), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .Y(n27986) );
  sky130_fd_sc_hd__xor2_1 U32631 ( .A(n27987), .B(n27986), .X(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[11]) );
  sky130_fd_sc_hd__o22ai_1 U32632 ( .A1(n28614), .A2(n27990), .B1(n27989), 
        .B2(n27988), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__nand4_1 U32633 ( .A(n27993), .B(j202_soc_core_uart_sio_ce), 
        .C(n27992), .D(n27991), .Y(n27994) );
  sky130_fd_sc_hd__nand2_1 U32634 ( .A(n27994), .B(n12142), .Y(
        j202_soc_core_uart_TOP_N16) );
  sky130_fd_sc_hd__nand2_1 U32635 ( .A(n12142), .B(n28564), .Y(n10679) );
  sky130_fd_sc_hd__nand2b_1 U32636 ( .A_N(j202_soc_core_uart_TOP_rxd_s), .B(
        j202_soc_core_uart_TOP_rxd_r), .Y(n27995) );
  sky130_fd_sc_hd__o211ai_1 U32637 ( .A1(j202_soc_core_uart_TOP_rx_go), .A2(
        n27995), .B1(n28000), .C1(n29593), .Y(j202_soc_core_uart_TOP_N85) );
  sky130_fd_sc_hd__a21oi_1 U32638 ( .A1(n28623), .A2(
        j202_soc_core_uart_TOP_rx_bit_cnt[1]), .B1(n27996), .Y(n27997) );
  sky130_fd_sc_hd__o21ai_1 U32639 ( .A1(n28000), .A2(n27997), .B1(n12142), .Y(
        j202_soc_core_uart_TOP_N87) );
  sky130_fd_sc_hd__xor2_1 U32640 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[3]), 
        .B(n27998), .X(n27999) );
  sky130_fd_sc_hd__o21ai_1 U32641 ( .A1(n28000), .A2(n27999), .B1(n12142), .Y(
        j202_soc_core_uart_TOP_N89) );
  sky130_fd_sc_hd__nand2_1 U32642 ( .A(j202_soc_core_uart_TOP_tx_bit_cnt[0]), 
        .B(j202_soc_core_uart_TOP_tx_bit_cnt[1]), .Y(n28007) );
  sky130_fd_sc_hd__nand2_1 U32644 ( .A(n29080), .B(n28001), .Y(n28005) );
  sky130_fd_sc_hd__nor2_1 U32645 ( .A(n28002), .B(n28005), .Y(
        j202_soc_core_uart_TOP_N59) );
  sky130_fd_sc_hd__nand2_1 U32646 ( .A(n28781), .B(n12142), .Y(
        j202_soc_core_uart_TOP_N57) );
  sky130_fd_sc_hd__and3_1 U32648 ( .A(j202_soc_core_uart_TOP_tx_bit_cnt[0]), 
        .B(j202_soc_core_uart_TOP_tx_bit_cnt[1]), .C(
        j202_soc_core_uart_TOP_tx_bit_cnt[2]), .X(n28006) );
  sky130_fd_sc_hd__xnor2_1 U32649 ( .A(j202_soc_core_uart_TOP_tx_bit_cnt[3]), 
        .B(n28006), .Y(n28004) );
  sky130_fd_sc_hd__o21ai_1 U32650 ( .A1(n28005), .A2(n28004), .B1(n12142), .Y(
        j202_soc_core_uart_TOP_N61) );
  sky130_fd_sc_hd__a211oi_1 U32651 ( .A1(n28007), .A2(n28625), .B1(n28006), 
        .C1(n28005), .Y(j202_soc_core_uart_TOP_N60) );
  sky130_fd_sc_hd__nand2_1 U32652 ( .A(n28008), .B(n12142), .Y(
        j202_soc_core_uart_BRG_N55) );
  sky130_fd_sc_hd__nor2_1 U32653 ( .A(j202_soc_core_uart_BRG_cnt[1]), .B(
        n28009), .Y(n28010) );
  sky130_fd_sc_hd__nor2_1 U32654 ( .A(n28010), .B(n29082), .Y(n28011) );
  sky130_fd_sc_hd__nor2_1 U32655 ( .A(n29090), .B(n28011), .Y(
        j202_soc_core_uart_BRG_N57) );
  sky130_fd_sc_hd__nand2_1 U32656 ( .A(j202_soc_core_uart_BRG_ps[1]), .B(
        j202_soc_core_uart_BRG_ps[0]), .Y(n28014) );
  sky130_fd_sc_hd__o21ai_1 U32657 ( .A1(j202_soc_core_uart_BRG_ps[1]), .A2(
        j202_soc_core_uart_BRG_ps[0]), .B1(n28014), .Y(n28013) );
  sky130_fd_sc_hd__nand2_1 U32658 ( .A(n28012), .B(n12142), .Y(n28034) );
  sky130_fd_sc_hd__nor2_1 U32659 ( .A(n28013), .B(n28034), .Y(
        j202_soc_core_uart_BRG_N13) );
  sky130_fd_sc_hd__nor2_1 U32660 ( .A(j202_soc_core_uart_BRG_ps[0]), .B(n28034), .Y(j202_soc_core_uart_BRG_N12) );
  sky130_fd_sc_hd__nor2_1 U32661 ( .A(n28015), .B(n28014), .Y(n28019) );
  sky130_fd_sc_hd__o21ai_1 U32662 ( .A1(n28017), .A2(
        j202_soc_core_uart_BRG_ps[2]), .B1(n28016), .Y(n28018) );
  sky130_fd_sc_hd__nor2_1 U32663 ( .A(n28018), .B(n28034), .Y(
        j202_soc_core_uart_BRG_N14) );
  sky130_fd_sc_hd__nand2_1 U32664 ( .A(j202_soc_core_uart_BRG_ps[3]), .B(
        n28019), .Y(n28021) );
  sky130_fd_sc_hd__nor2_1 U32666 ( .A(n28020), .B(n28034), .Y(
        j202_soc_core_uart_BRG_N15) );
  sky130_fd_sc_hd__nor2_1 U32667 ( .A(n28022), .B(n28021), .Y(n28026) );
  sky130_fd_sc_hd__o21ai_1 U32668 ( .A1(n28024), .A2(
        j202_soc_core_uart_BRG_ps[4]), .B1(n28023), .Y(n28025) );
  sky130_fd_sc_hd__nor2_1 U32669 ( .A(n28025), .B(n28034), .Y(
        j202_soc_core_uart_BRG_N16) );
  sky130_fd_sc_hd__nand2_1 U32670 ( .A(j202_soc_core_uart_BRG_ps[5]), .B(
        n28026), .Y(n28028) );
  sky130_fd_sc_hd__o21ai_1 U32671 ( .A1(j202_soc_core_uart_BRG_ps[5]), .A2(
        n28026), .B1(n28028), .Y(n28027) );
  sky130_fd_sc_hd__nor2_1 U32672 ( .A(n28027), .B(n28034), .Y(
        j202_soc_core_uart_BRG_N17) );
  sky130_fd_sc_hd__nor2_1 U32673 ( .A(n28029), .B(n28028), .Y(n28628) );
  sky130_fd_sc_hd__o21ai_1 U32674 ( .A1(n28031), .A2(
        j202_soc_core_uart_BRG_ps[6]), .B1(n28030), .Y(n28032) );
  sky130_fd_sc_hd__nor2_1 U32675 ( .A(n28032), .B(n28034), .Y(
        j202_soc_core_uart_BRG_N18) );
  sky130_fd_sc_hd__nand2_1 U32676 ( .A(j202_soc_core_uart_BRG_br_cnt[1]), .B(
        j202_soc_core_uart_BRG_br_cnt[0]), .Y(n28054) );
  sky130_fd_sc_hd__nor2_1 U32677 ( .A(n28040), .B(n28054), .Y(n28039) );
  sky130_fd_sc_hd__nand2_1 U32678 ( .A(j202_soc_core_uart_BRG_br_cnt[3]), .B(
        n28039), .Y(n28042) );
  sky130_fd_sc_hd__o21ai_1 U32679 ( .A1(j202_soc_core_uart_BRG_br_cnt[3]), 
        .A2(n28039), .B1(n28042), .Y(n28033) );
  sky130_fd_sc_hd__nand3_1 U32680 ( .A(n28035), .B(
        j202_soc_core_uart_BRG_ps_clr), .C(n29593), .Y(n28629) );
  sky130_fd_sc_hd__nor2_1 U32681 ( .A(n28033), .B(n28629), .Y(
        j202_soc_core_uart_BRG_N38) );
  sky130_fd_sc_hd__nand2_1 U32682 ( .A(n28626), .B(n28035), .Y(n10678) );
  sky130_fd_sc_hd__nor2_1 U32683 ( .A(j202_soc_core_uart_BRG_br_cnt[0]), .B(
        n28629), .Y(j202_soc_core_uart_BRG_N35) );
  sky130_fd_sc_hd__nor2_1 U32684 ( .A(n28043), .B(n28042), .Y(n28041) );
  sky130_fd_sc_hd__nand2_1 U32685 ( .A(j202_soc_core_uart_BRG_br_cnt[5]), .B(
        n28041), .Y(n28037) );
  sky130_fd_sc_hd__nor2_1 U32686 ( .A(n28036), .B(n28037), .Y(n28632) );
  sky130_fd_sc_hd__a211oi_1 U32687 ( .A1(n28036), .A2(n28037), .B1(n28632), 
        .C1(n28629), .Y(j202_soc_core_uart_BRG_N41) );
  sky130_fd_sc_hd__nor2_1 U32689 ( .A(n28038), .B(n28629), .Y(
        j202_soc_core_uart_BRG_N40) );
  sky130_fd_sc_hd__a211oi_1 U32690 ( .A1(n28040), .A2(n28054), .B1(n28039), 
        .C1(n28629), .Y(j202_soc_core_uart_BRG_N37) );
  sky130_fd_sc_hd__a211oi_1 U32691 ( .A1(n28043), .A2(n28042), .B1(n28041), 
        .C1(n28629), .Y(j202_soc_core_uart_BRG_N39) );
  sky130_fd_sc_hd__xnor2_1 U32692 ( .A(j202_soc_core_uart_div1[2]), .B(
        j202_soc_core_uart_BRG_br_cnt[2]), .Y(n28047) );
  sky130_fd_sc_hd__xnor2_1 U32693 ( .A(j202_soc_core_uart_div1[4]), .B(
        j202_soc_core_uart_BRG_br_cnt[4]), .Y(n28046) );
  sky130_fd_sc_hd__xnor2_1 U32694 ( .A(j202_soc_core_uart_div1[6]), .B(
        j202_soc_core_uart_BRG_br_cnt[6]), .Y(n28045) );
  sky130_fd_sc_hd__xnor2_1 U32695 ( .A(j202_soc_core_uart_div1[7]), .B(
        j202_soc_core_uart_BRG_br_cnt[7]), .Y(n28044) );
  sky130_fd_sc_hd__nand4_1 U32696 ( .A(n28047), .B(n28046), .C(n28045), .D(
        n28044), .Y(n28053) );
  sky130_fd_sc_hd__xnor2_1 U32697 ( .A(j202_soc_core_uart_div1[1]), .B(
        j202_soc_core_uart_BRG_br_cnt[1]), .Y(n28051) );
  sky130_fd_sc_hd__xnor2_1 U32698 ( .A(j202_soc_core_uart_div1[5]), .B(
        j202_soc_core_uart_BRG_br_cnt[5]), .Y(n28050) );
  sky130_fd_sc_hd__xnor2_1 U32699 ( .A(j202_soc_core_uart_div1[3]), .B(
        j202_soc_core_uart_BRG_br_cnt[3]), .Y(n28049) );
  sky130_fd_sc_hd__xnor2_1 U32700 ( .A(j202_soc_core_uart_div1[0]), .B(
        j202_soc_core_uart_BRG_br_cnt[0]), .Y(n28048) );
  sky130_fd_sc_hd__nand4_1 U32701 ( .A(n28051), .B(n28050), .C(n28049), .D(
        n28048), .Y(n28052) );
  sky130_fd_sc_hd__nor2_1 U32702 ( .A(n28053), .B(n28052), .Y(
        j202_soc_core_uart_BRG_N47) );
  sky130_fd_sc_hd__o21ai_1 U32703 ( .A1(j202_soc_core_uart_BRG_br_cnt[1]), 
        .A2(j202_soc_core_uart_BRG_br_cnt[0]), .B1(n28054), .Y(n28055) );
  sky130_fd_sc_hd__nor2_1 U32704 ( .A(n28055), .B(n28629), .Y(
        j202_soc_core_uart_BRG_N36) );
  sky130_fd_sc_hd__nand2_1 U32705 ( .A(n28056), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[4]), .Y(n28057) );
  sky130_fd_sc_hd__a31oi_1 U32706 ( .A1(n28057), .A2(
        j202_soc_core_wbqspiflash_00_state[0]), .A3(n28059), .B1(n28063), .Y(
        j202_soc_core_wbqspiflash_00_N618) );
  sky130_fd_sc_hd__a211oi_1 U32707 ( .A1(n28059), .A2(
        j202_soc_core_wbqspiflash_00_reset_counter[5]), .B1(n28058), .C1(
        n28061), .Y(n28060) );
  sky130_fd_sc_hd__nor2_1 U32708 ( .A(n28063), .B(n28060), .Y(
        j202_soc_core_wbqspiflash_00_N619) );
  sky130_fd_sc_hd__nand2_1 U32709 ( .A(n28062), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[6]), .Y(n28065) );
  sky130_fd_sc_hd__a31oi_1 U32710 ( .A1(n28065), .A2(
        j202_soc_core_wbqspiflash_00_state[0]), .A3(n28064), .B1(n28063), .Y(
        j202_soc_core_wbqspiflash_00_N620) );
  sky130_fd_sc_hd__a21oi_1 U32711 ( .A1(n28067), .A2(n28100), .B1(n28066), .Y(
        n28082) );
  sky130_fd_sc_hd__nand2_1 U32712 ( .A(n28237), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .Y(n28087) );
  sky130_fd_sc_hd__o22ai_1 U32713 ( .A1(n28086), .A2(n28087), .B1(n28069), 
        .B2(n28068), .Y(n28070) );
  sky130_fd_sc_hd__nor2_1 U32714 ( .A(n28078), .B(n28070), .Y(n28072) );
  sky130_fd_sc_hd__nand2_1 U32715 ( .A(n28259), .B(
        j202_soc_core_wbqspiflash_00_spif_data[28]), .Y(n28071) );
  sky130_fd_sc_hd__nand4_1 U32716 ( .A(n28073), .B(n28082), .C(n28072), .D(
        n28071), .Y(n28074) );
  sky130_fd_sc_hd__a211o_1 U32717 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]), .B1(n28172), .C1(n28074), .X(n10509) );
  sky130_fd_sc_hd__a22oi_1 U32718 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[30]), .Y(n28076) );
  sky130_fd_sc_hd__nand4_1 U32719 ( .A(n28083), .B(n28076), .C(n28187), .D(
        n28075), .Y(n28077) );
  sky130_fd_sc_hd__a21o_1 U32720 ( .A1(n28261), .A2(
        j202_soc_core_qspi_wb_addr[22]), .B1(n28077), .X(n10507) );
  sky130_fd_sc_hd__nand3_1 U32721 ( .A(n28080), .B(n28079), .C(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]), .Y(n28081) );
  sky130_fd_sc_hd__nand3_1 U32722 ( .A(n28083), .B(n28082), .C(n28081), .Y(
        n28084) );
  sky130_fd_sc_hd__a211oi_1 U32723 ( .A1(n28259), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[29]), .B1(n28085), .C1(n28084), 
        .Y(n28092) );
  sky130_fd_sc_hd__nor3_1 U32724 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .B(n28087), .C(n28086), 
        .Y(n28088) );
  sky130_fd_sc_hd__a31oi_1 U32725 ( .A1(n28090), .A2(n28089), .A3(
        j202_soc_core_qspi_wb_addr[21]), .B1(n28088), .Y(n28091) );
  sky130_fd_sc_hd__o211ai_1 U32726 ( .A1(j202_soc_core_qspi_wb_addr[3]), .A2(
        n28093), .B1(n28092), .C1(n28091), .Y(n10508) );
  sky130_fd_sc_hd__nand2_1 U32727 ( .A(n28095), .B(n28094), .Y(
        j202_soc_core_wbqspiflash_00_N86) );
  sky130_fd_sc_hd__nand3_1 U32728 ( .A(n28098), .B(n28097), .C(n28096), .Y(
        j202_soc_core_wbqspiflash_00_N594) );
  sky130_fd_sc_hd__a21oi_1 U32729 ( .A1(n28100), .A2(
        j202_soc_core_wbqspiflash_00_state[4]), .B1(n28099), .Y(n28101) );
  sky130_fd_sc_hd__a21oi_1 U32730 ( .A1(n28102), .A2(n28101), .B1(n28590), .Y(
        j202_soc_core_wbqspiflash_00_N747) );
  sky130_fd_sc_hd__nor2_1 U32731 ( .A(n28127), .B(n28108), .Y(
        j202_soc_core_wbqspiflash_00_N628) );
  sky130_fd_sc_hd__nor2_1 U32732 ( .A(n28652), .B(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N391) );
  sky130_fd_sc_hd__nand2_1 U32733 ( .A(n28207), .B(n28103), .Y(n28104) );
  sky130_fd_sc_hd__nand2_1 U32734 ( .A(n28232), .B(n28104), .Y(n28201) );
  sky130_fd_sc_hd__a22oi_1 U32735 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .A2(n28201), .B1(n28259), 
        .B2(j202_soc_core_wbqspiflash_00_spif_data[3]), .Y(n28105) );
  sky130_fd_sc_hd__o21ai_1 U32736 ( .A1(n28106), .A2(n28115), .B1(n28105), .Y(
        n10534) );
  sky130_fd_sc_hd__a222oi_1 U32737 ( .A1(n28201), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[4]), .B1(n28215), .B2(
        j202_soc_core_qspi_wb_addr[4]), .C1(n28259), .C2(
        j202_soc_core_wbqspiflash_00_spif_data[4]), .Y(n28107) );
  sky130_fd_sc_hd__nor2_1 U32738 ( .A(n28158), .B(n28108), .Y(
        j202_soc_core_wbqspiflash_00_N629) );
  sky130_fd_sc_hd__nand2_1 U32739 ( .A(n28743), .B(n28109), .Y(n28738) );
  sky130_fd_sc_hd__nand2_1 U32740 ( .A(n28737), .B(n28110), .Y(n28740) );
  sky130_fd_sc_hd__a22oi_1 U32741 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[0]), .B1(n28719), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[0]), .Y(n28111) );
  sky130_fd_sc_hd__o21ai_1 U32742 ( .A1(n28655), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B1(n28111), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N392) );
  sky130_fd_sc_hd__a22oi_1 U32743 ( .A1(n28201), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[5]), .B1(n28119), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[5]), .Y(n28112) );
  sky130_fd_sc_hd__nor2_1 U32744 ( .A(n28260), .B(n28261), .Y(n28120) );
  sky130_fd_sc_hd__o211ai_1 U32745 ( .A1(n28123), .A2(n28113), .B1(n28112), 
        .C1(n28120), .Y(n10532) );
  sky130_fd_sc_hd__a22oi_1 U32746 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .A2(n28201), .B1(n28259), 
        .B2(j202_soc_core_wbqspiflash_00_spif_data[2]), .Y(n28114) );
  sky130_fd_sc_hd__o21ai_1 U32747 ( .A1(n28116), .A2(n28115), .B1(n28114), .Y(
        n10535) );
  sky130_fd_sc_hd__a22oi_1 U32748 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[1]), .B1(n28719), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[1]), .Y(n28117) );
  sky130_fd_sc_hd__o21ai_1 U32749 ( .A1(n28658), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B1(n28117), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N393) );
  sky130_fd_sc_hd__a222oi_1 U32750 ( .A1(n28201), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[6]), .B1(n28215), .B2(
        j202_soc_core_qspi_wb_addr[6]), .C1(n28259), .C2(
        j202_soc_core_wbqspiflash_00_spif_data[6]), .Y(n28118) );
  sky130_fd_sc_hd__a22oi_1 U32751 ( .A1(n28201), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[7]), .B1(n28119), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[7]), .Y(n28121) );
  sky130_fd_sc_hd__o211ai_1 U32752 ( .A1(n28123), .A2(n28122), .B1(n28121), 
        .C1(n28120), .Y(n10530) );
  sky130_fd_sc_hd__a22oi_1 U32753 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[8]), .A2(n28201), .B1(n28259), 
        .B2(j202_soc_core_wbqspiflash_00_spif_data[8]), .Y(n28125) );
  sky130_fd_sc_hd__nand2_1 U32754 ( .A(n28215), .B(
        j202_soc_core_qspi_wb_addr[8]), .Y(n28124) );
  sky130_fd_sc_hd__o211ai_1 U32755 ( .A1(n28127), .A2(n28126), .B1(n28125), 
        .C1(n28124), .Y(n10529) );
  sky130_fd_sc_hd__a22o_1 U32756 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[9]), .A2(n28201), .B1(n28259), 
        .B2(j202_soc_core_wbqspiflash_00_spif_data[9]), .X(n28128) );
  sky130_fd_sc_hd__a211o_1 U32757 ( .A1(j202_soc_core_qspi_wb_addr[9]), .A2(
        n28215), .B1(n28129), .C1(n28128), .X(n10528) );
  sky130_fd_sc_hd__a22oi_1 U32758 ( .A1(n28261), .A2(
        j202_soc_core_qspi_wb_addr[2]), .B1(n28215), .B2(
        j202_soc_core_qspi_wb_addr[10]), .Y(n28132) );
  sky130_fd_sc_hd__a22oi_1 U32759 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[10]), .Y(n28131) );
  sky130_fd_sc_hd__a22oi_1 U32760 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[10]), .A2(n28201), .B1(n28221), .B2(j202_soc_core_wbqspiflash_00_spif_data[2]), .Y(n28130) );
  sky130_fd_sc_hd__nand3_1 U32761 ( .A(n28132), .B(n28131), .C(n28130), .Y(
        n10527) );
  sky130_fd_sc_hd__a22oi_1 U32762 ( .A1(n28261), .A2(
        j202_soc_core_qspi_wb_addr[3]), .B1(n28215), .B2(
        j202_soc_core_qspi_wb_addr[11]), .Y(n28135) );
  sky130_fd_sc_hd__a22oi_1 U32763 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[11]), .Y(n28134) );
  sky130_fd_sc_hd__a22oi_1 U32764 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[11]), .A2(n28201), .B1(n28221), .B2(j202_soc_core_wbqspiflash_00_spif_data[3]), .Y(n28133) );
  sky130_fd_sc_hd__nand3_1 U32765 ( .A(n28135), .B(n28134), .C(n28133), .Y(
        n10526) );
  sky130_fd_sc_hd__a22oi_1 U32766 ( .A1(n28261), .A2(
        j202_soc_core_qspi_wb_addr[4]), .B1(n28215), .B2(
        j202_soc_core_qspi_wb_addr[12]), .Y(n28138) );
  sky130_fd_sc_hd__a22oi_1 U32767 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[4]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[12]), .Y(n28137) );
  sky130_fd_sc_hd__a22oi_1 U32768 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[12]), .A2(n28201), .B1(n28221), .B2(j202_soc_core_wbqspiflash_00_spif_data[4]), .Y(n28136) );
  sky130_fd_sc_hd__nand3_1 U32769 ( .A(n28138), .B(n28137), .C(n28136), .Y(
        n10525) );
  sky130_fd_sc_hd__a22oi_1 U32770 ( .A1(n28261), .A2(
        j202_soc_core_qspi_wb_addr[5]), .B1(n28215), .B2(
        j202_soc_core_qspi_wb_addr[13]), .Y(n28141) );
  sky130_fd_sc_hd__a22oi_1 U32771 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[5]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[13]), .Y(n28140) );
  sky130_fd_sc_hd__a22oi_1 U32772 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[13]), .A2(n28201), .B1(n28221), .B2(j202_soc_core_wbqspiflash_00_spif_data[5]), .Y(n28139) );
  sky130_fd_sc_hd__nand3_1 U32773 ( .A(n28141), .B(n28140), .C(n28139), .Y(
        n10524) );
  sky130_fd_sc_hd__a22oi_1 U32774 ( .A1(n28261), .A2(
        j202_soc_core_qspi_wb_addr[6]), .B1(n28215), .B2(
        j202_soc_core_qspi_wb_addr[14]), .Y(n28144) );
  sky130_fd_sc_hd__a22oi_1 U32775 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[6]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[14]), .Y(n28143) );
  sky130_fd_sc_hd__a22oi_1 U32776 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]), .A2(n28201), .B1(n28221), .B2(j202_soc_core_wbqspiflash_00_spif_data[6]), .Y(n28142) );
  sky130_fd_sc_hd__nand3_1 U32777 ( .A(n28144), .B(n28143), .C(n28142), .Y(
        n10523) );
  sky130_fd_sc_hd__a22oi_1 U32778 ( .A1(n28261), .A2(
        j202_soc_core_qspi_wb_addr[7]), .B1(n28215), .B2(
        j202_soc_core_qspi_wb_addr[15]), .Y(n28147) );
  sky130_fd_sc_hd__a22oi_1 U32779 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[7]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[15]), .Y(n28146) );
  sky130_fd_sc_hd__a22oi_1 U32780 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[15]), .A2(n28201), .B1(n28221), .B2(j202_soc_core_wbqspiflash_00_spif_data[7]), .Y(n28145) );
  sky130_fd_sc_hd__nand3_1 U32781 ( .A(n28147), .B(n28146), .C(n28145), .Y(
        n10522) );
  sky130_fd_sc_hd__nand2_1 U32782 ( .A(n28199), .B(
        j202_soc_core_wbqspiflash_00_spif_data[0]), .Y(n28153) );
  sky130_fd_sc_hd__o21ai_1 U32783 ( .A1(n28148), .A2(n28551), .B1(n28153), .Y(
        j202_soc_core_wbqspiflash_00_N605) );
  sky130_fd_sc_hd__a22oi_1 U32784 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]), .A2(n28201), .B1(n28221), .B2(j202_soc_core_wbqspiflash_00_last_status[0]), .Y(n28149) );
  sky130_fd_sc_hd__o21ai_1 U32785 ( .A1(n28150), .A2(n28187), .B1(n28149), .Y(
        n28151) );
  sky130_fd_sc_hd__a21oi_1 U32786 ( .A1(n28215), .A2(
        j202_soc_core_qspi_wb_addr[16]), .B1(n28151), .Y(n28155) );
  sky130_fd_sc_hd__a22oi_1 U32787 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[8]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[16]), .Y(n28154) );
  sky130_fd_sc_hd__nand2_1 U32788 ( .A(n28261), .B(
        j202_soc_core_qspi_wb_addr[8]), .Y(n28152) );
  sky130_fd_sc_hd__nand4_1 U32789 ( .A(n28155), .B(n28154), .C(n28153), .D(
        n28152), .Y(n10521) );
  sky130_fd_sc_hd__a22o_1 U32790 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[9]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[17]), .X(n28156) );
  sky130_fd_sc_hd__a21oi_1 U32791 ( .A1(n28221), .A2(
        j202_soc_core_wbqspiflash_00_last_status[1]), .B1(n28156), .Y(n28162)
         );
  sky130_fd_sc_hd__nor2_1 U32792 ( .A(n28158), .B(n28157), .Y(n28548) );
  sky130_fd_sc_hd__a21oi_1 U32793 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]), .A2(n28201), .B1(n28548), .Y(n28161) );
  sky130_fd_sc_hd__a22oi_1 U32794 ( .A1(n28261), .A2(
        j202_soc_core_qspi_wb_addr[9]), .B1(n28215), .B2(
        j202_soc_core_qspi_wb_addr[17]), .Y(n28160) );
  sky130_fd_sc_hd__nand2_1 U32795 ( .A(n28172), .B(
        j202_soc_core_wbqspiflash_00_spif_data[15]), .Y(n28159) );
  sky130_fd_sc_hd__nand4_1 U32796 ( .A(n28162), .B(n28161), .C(n28160), .D(
        n28159), .Y(n10520) );
  sky130_fd_sc_hd__nand2_1 U32797 ( .A(n28199), .B(
        j202_soc_core_wbqspiflash_00_spif_data[2]), .Y(n28168) );
  sky130_fd_sc_hd__o21ai_1 U32798 ( .A1(n28163), .A2(n28551), .B1(n28168), .Y(
        j202_soc_core_wbqspiflash_00_N607) );
  sky130_fd_sc_hd__a22oi_1 U32799 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .A2(n28201), .B1(n28221), .B2(j202_soc_core_wbqspiflash_00_last_status[2]), .Y(n28164) );
  sky130_fd_sc_hd__o21ai_1 U32800 ( .A1(n28165), .A2(n28187), .B1(n28164), .Y(
        n28166) );
  sky130_fd_sc_hd__a21oi_1 U32801 ( .A1(n28215), .A2(
        j202_soc_core_qspi_wb_addr[18]), .B1(n28166), .Y(n28170) );
  sky130_fd_sc_hd__a22oi_1 U32802 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[10]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[18]), .Y(n28169) );
  sky130_fd_sc_hd__nand2_1 U32803 ( .A(n28261), .B(
        j202_soc_core_qspi_wb_addr[10]), .Y(n28167) );
  sky130_fd_sc_hd__nand4_1 U32804 ( .A(n28170), .B(n28169), .C(n28168), .D(
        n28167), .Y(n10519) );
  sky130_fd_sc_hd__nand2_1 U32805 ( .A(n28199), .B(
        j202_soc_core_wbqspiflash_00_spif_data[3]), .Y(n28550) );
  sky130_fd_sc_hd__a21oi_1 U32806 ( .A1(n28221), .A2(
        j202_soc_core_wbqspiflash_00_last_status[3]), .B1(n28171), .Y(n28177)
         );
  sky130_fd_sc_hd__a22oi_1 U32807 ( .A1(n28261), .A2(
        j202_soc_core_qspi_wb_addr[11]), .B1(n28172), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[17]), .Y(n28176) );
  sky130_fd_sc_hd__a22o_1 U32808 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[11]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[19]), .X(n28173) );
  sky130_fd_sc_hd__a21oi_1 U32809 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .A2(n28201), .B1(n28173), .Y(n28175) );
  sky130_fd_sc_hd__nand2_1 U32810 ( .A(n28215), .B(
        j202_soc_core_qspi_wb_addr[19]), .Y(n28174) );
  sky130_fd_sc_hd__nand4_1 U32811 ( .A(n28177), .B(n28176), .C(n28175), .D(
        n28174), .Y(n10518) );
  sky130_fd_sc_hd__nand2_1 U32812 ( .A(n28199), .B(
        j202_soc_core_wbqspiflash_00_spif_data[4]), .Y(n28182) );
  sky130_fd_sc_hd__o21ai_1 U32813 ( .A1(n28178), .A2(n28551), .B1(n28182), .Y(
        j202_soc_core_wbqspiflash_00_N609) );
  sky130_fd_sc_hd__a22oi_1 U32814 ( .A1(n28221), .A2(
        j202_soc_core_wbqspiflash_00_last_status[4]), .B1(n28201), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]), .Y(n28179) );
  sky130_fd_sc_hd__a21oi_1 U32816 ( .A1(n28215), .A2(
        j202_soc_core_qspi_wb_addr[20]), .B1(n28181), .Y(n28185) );
  sky130_fd_sc_hd__nand2_1 U32817 ( .A(n28261), .B(
        j202_soc_core_qspi_wb_addr[12]), .Y(n28184) );
  sky130_fd_sc_hd__a22oi_1 U32818 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[12]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[20]), .Y(n28183) );
  sky130_fd_sc_hd__nand4_1 U32819 ( .A(n28185), .B(n28184), .C(n28183), .D(
        n28182), .Y(n10517) );
  sky130_fd_sc_hd__a22oi_1 U32820 ( .A1(n28221), .A2(
        j202_soc_core_wbqspiflash_00_last_status[5]), .B1(n28201), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]), .Y(n28186) );
  sky130_fd_sc_hd__o21ai_1 U32821 ( .A1(n28188), .A2(n28187), .B1(n28186), .Y(
        n28189) );
  sky130_fd_sc_hd__a21oi_1 U32822 ( .A1(n28215), .A2(
        j202_soc_core_qspi_wb_addr[21]), .B1(n28189), .Y(n28193) );
  sky130_fd_sc_hd__nand2_1 U32823 ( .A(n28261), .B(
        j202_soc_core_qspi_wb_addr[13]), .Y(n28192) );
  sky130_fd_sc_hd__a22oi_1 U32824 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[13]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[21]), .Y(n28191) );
  sky130_fd_sc_hd__nand4_1 U32825 ( .A(n28193), .B(n28192), .C(n28191), .D(
        n28190), .Y(n10516) );
  sky130_fd_sc_hd__a22o_1 U32826 ( .A1(n28221), .A2(
        j202_soc_core_wbqspiflash_00_last_status[6]), .B1(n28201), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .X(n28194) );
  sky130_fd_sc_hd__a21oi_1 U32827 ( .A1(n28261), .A2(
        j202_soc_core_qspi_wb_addr[14]), .B1(n28194), .Y(n28198) );
  sky130_fd_sc_hd__a22oi_1 U32828 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[22]), .Y(n28197) );
  sky130_fd_sc_hd__nand2_1 U32829 ( .A(n28215), .B(
        j202_soc_core_qspi_wb_addr[22]), .Y(n28195) );
  sky130_fd_sc_hd__nand4_1 U32830 ( .A(n28198), .B(n28197), .C(n28196), .D(
        n28195), .Y(n10515) );
  sky130_fd_sc_hd__nand2_1 U32831 ( .A(n28199), .B(
        j202_soc_core_wbqspiflash_00_spif_data[7]), .Y(n28204) );
  sky130_fd_sc_hd__o21ai_1 U32832 ( .A1(n28200), .A2(n28551), .B1(n28204), .Y(
        j202_soc_core_wbqspiflash_00_N613) );
  sky130_fd_sc_hd__a22o_1 U32833 ( .A1(n28221), .A2(
        j202_soc_core_wbqspiflash_00_last_status[7]), .B1(n28201), .B2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]), .X(n28202) );
  sky130_fd_sc_hd__a21oi_1 U32834 ( .A1(n28261), .A2(
        j202_soc_core_qspi_wb_addr[15]), .B1(n28202), .Y(n28206) );
  sky130_fd_sc_hd__a22oi_1 U32835 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[15]), .B1(n28259), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[23]), .Y(n28205) );
  sky130_fd_sc_hd__nand2_1 U32836 ( .A(n28215), .B(
        j202_soc_core_qspi_wb_addr[23]), .Y(n28203) );
  sky130_fd_sc_hd__nand4_1 U32837 ( .A(n28206), .B(n28205), .C(n28204), .D(
        n28203), .Y(n10514) );
  sky130_fd_sc_hd__a211o_1 U32838 ( .A1(n28210), .A2(n28209), .B1(
        j202_soc_core_wbqspiflash_00_state[2]), .C1(n28208), .X(n28219) );
  sky130_fd_sc_hd__nand3_1 U32839 ( .A(n28213), .B(n28212), .C(n28751), .Y(
        n28246) );
  sky130_fd_sc_hd__a21o_1 U32840 ( .A1(n28254), .A2(
        j202_soc_core_qspi_wb_addr[16]), .B1(n28246), .X(n28214) );
  sky130_fd_sc_hd__a211oi_1 U32841 ( .A1(n28249), .A2(n28237), .B1(n28215), 
        .C1(n28214), .Y(n28218) );
  sky130_fd_sc_hd__nand2_1 U32842 ( .A(n28260), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]), .Y(n28216) );
  sky130_fd_sc_hd__nand4_1 U32843 ( .A(n28219), .B(n28218), .C(n28217), .D(
        n28216), .Y(n28220) );
  sky130_fd_sc_hd__a211o_1 U32844 ( .A1(n28259), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[24]), .B1(n28221), .C1(n28220), 
        .X(n10513) );
  sky130_fd_sc_hd__o21ai_1 U32845 ( .A1(n10958), .A2(n28223), .B1(
        j202_soc_core_ahb2wbqspi_00_stb_o), .Y(n28226) );
  sky130_fd_sc_hd__a21oi_1 U32846 ( .A1(n28226), .A2(n28225), .B1(n28224), .Y(
        n28227) );
  sky130_fd_sc_hd__a21oi_1 U32847 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]), .A2(n28228), .B1(n28227), .Y(n28244) );
  sky130_fd_sc_hd__nand4b_1 U32848 ( .A_N(n28231), .B(n28230), .C(n28229), .D(
        j202_soc_core_qspi_wb_addr[17]), .Y(n28233) );
  sky130_fd_sc_hd__nand2_1 U32849 ( .A(n28233), .B(n28232), .Y(n28241) );
  sky130_fd_sc_hd__o2bb2ai_1 U32850 ( .B1(
        j202_soc_core_wbqspiflash_00_spif_ctrl), .B2(n28250), .A1_N(n28234), 
        .A2_N(j202_soc_core_wbqspiflash_00_spif_data[25]), .Y(n28240) );
  sky130_fd_sc_hd__a21oi_1 U32851 ( .A1(n28237), .A2(n28236), .B1(n28235), .Y(
        n28239) );
  sky130_fd_sc_hd__nor4_1 U32852 ( .A(n28241), .B(n28240), .C(n28239), .D(
        n28238), .Y(n28242) );
  sky130_fd_sc_hd__o21ai_1 U32853 ( .A1(n28244), .A2(n28243), .B1(n28242), .Y(
        n10512) );
  sky130_fd_sc_hd__nor4_1 U32854 ( .A(n28249), .B(n28248), .C(n28247), .D(
        n28246), .Y(n28257) );
  sky130_fd_sc_hd__a21oi_1 U32855 ( .A1(n28252), .A2(n28251), .B1(n28250), .Y(
        n28253) );
  sky130_fd_sc_hd__a21oi_1 U32856 ( .A1(n28259), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[26]), .B1(n28253), .Y(n28256)
         );
  sky130_fd_sc_hd__a22oi_1 U32857 ( .A1(n28260), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .B1(n28254), .B2(
        j202_soc_core_qspi_wb_addr[18]), .Y(n28255) );
  sky130_fd_sc_hd__nand3_1 U32858 ( .A(n28257), .B(n28256), .C(n28255), .Y(
        n10511) );
  sky130_fd_sc_hd__a21oi_1 U32859 ( .A1(n28259), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[27]), .B1(n28258), .Y(n28264)
         );
  sky130_fd_sc_hd__nand2_1 U32860 ( .A(n28260), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .Y(n28263) );
  sky130_fd_sc_hd__nand2_1 U32861 ( .A(n28261), .B(
        j202_soc_core_qspi_wb_addr[19]), .Y(n28262) );
  sky130_fd_sc_hd__nand4_1 U32862 ( .A(n28265), .B(n28264), .C(n28263), .D(
        n28262), .Y(n10510) );
  sky130_fd_sc_hd__a22oi_1 U32863 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[30]), .B1(n28733), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[27]), .Y(n28267) );
  sky130_fd_sc_hd__a22oi_1 U32864 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[30]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[27]), .B2(n28734), .Y(n28266) );
  sky130_fd_sc_hd__o211ai_1 U32865 ( .A1(n28268), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B1(n28267), .C1(n28266), 
        .Y(j202_soc_core_wbqspiflash_00_lldriver_N422) );
  sky130_fd_sc_hd__o22ai_1 U32866 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[30]), .B1(n28901), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[27]), .Y(n28269) );
  sky130_fd_sc_hd__nor2_1 U32867 ( .A(n26211), .B(n28269), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N389) );
  sky130_fd_sc_hd__nand2_1 U32868 ( .A(n28281), .B(j202_soc_core_uart_din_i[0]), .Y(n28270) );
  sky130_fd_sc_hd__o21ai_1 U32869 ( .A1(n28271), .A2(n28281), .B1(n28270), .Y(
        n85) );
  sky130_fd_sc_hd__nand2_1 U32870 ( .A(n28281), .B(j202_soc_core_uart_din_i[1]), .Y(n28272) );
  sky130_fd_sc_hd__o21ai_1 U32871 ( .A1(n28273), .A2(n28281), .B1(n28272), .Y(
        n37) );
  sky130_fd_sc_hd__nand2_1 U32872 ( .A(n28281), .B(j202_soc_core_uart_din_i[2]), .Y(n28274) );
  sky130_fd_sc_hd__o21ai_1 U32873 ( .A1(n28283), .A2(n28281), .B1(n28274), .Y(
        n79) );
  sky130_fd_sc_hd__nand2_1 U32874 ( .A(n28281), .B(j202_soc_core_uart_din_i[3]), .Y(n28275) );
  sky130_fd_sc_hd__nand2_1 U32876 ( .A(n28281), .B(j202_soc_core_uart_din_i[4]), .Y(n28276) );
  sky130_fd_sc_hd__o21ai_1 U32877 ( .A1(n28277), .A2(n28281), .B1(n28276), .Y(
        n91) );
  sky130_fd_sc_hd__nand2_1 U32878 ( .A(n28281), .B(j202_soc_core_uart_din_i[5]), .Y(n28278) );
  sky130_fd_sc_hd__o21ai_1 U32879 ( .A1(n28304), .A2(n28281), .B1(n28278), .Y(
        n90) );
  sky130_fd_sc_hd__nand2_1 U32880 ( .A(n28281), .B(j202_soc_core_uart_din_i[6]), .Y(n28279) );
  sky130_fd_sc_hd__o21ai_1 U32881 ( .A1(n28311), .A2(n28281), .B1(n28279), .Y(
        n89) );
  sky130_fd_sc_hd__nand2_1 U32882 ( .A(n28281), .B(j202_soc_core_uart_din_i[7]), .Y(n28280) );
  sky130_fd_sc_hd__nor2_1 U32884 ( .A(n28590), .B(n28282), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N4) );
  sky130_fd_sc_hd__nand2_1 U32885 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[18]), .Y(n28399) );
  sky130_fd_sc_hd__nand2_1 U32886 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[19]), .Y(n28407) );
  sky130_fd_sc_hd__nand2_1 U32887 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[20]), .Y(n28414) );
  sky130_fd_sc_hd__nand2_1 U32888 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[21]), .Y(n28424) );
  sky130_fd_sc_hd__nand2_1 U32889 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[22]), .Y(n28432) );
  sky130_fd_sc_hd__nand2_1 U32890 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[25]), .Y(n28454) );
  sky130_fd_sc_hd__nand2_1 U32891 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[26]), .Y(n28462) );
  sky130_fd_sc_hd__nand2_1 U32892 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[27]), .Y(n28470) );
  sky130_fd_sc_hd__nand2_1 U32893 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[29]), .Y(n28488) );
  sky130_fd_sc_hd__nand2_1 U32894 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[30]), .Y(n28496) );
  sky130_fd_sc_hd__nand2_1 U32895 ( .A(n12142), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[31]), .Y(n28504) );
  sky130_fd_sc_hd__a21oi_1 U32896 ( .A1(n29593), .A2(n28283), .B1(n28476), .Y(
        n28288) );
  sky130_fd_sc_hd__o22ai_1 U32897 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[2]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[2]), .B1(n28284), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[2]), .Y(n28285)
         );
  sky130_fd_sc_hd__a21oi_1 U32898 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[2]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[2]), .B1(n28285), 
        .Y(n28286) );
  sky130_fd_sc_hd__nand4_1 U32899 ( .A(n28286), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[2]), .C(n29594), .D(
        io_oeb[2]), .Y(n28287) );
  sky130_fd_sc_hd__nor2_1 U32901 ( .A(n28590), .B(n28290), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N6) );
  sky130_fd_sc_hd__a21oi_1 U32902 ( .A1(n12142), .A2(n28291), .B1(n28476), .Y(
        n28296) );
  sky130_fd_sc_hd__a21oi_1 U32904 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[3]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[3]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]), .Y(n28292) );
  sky130_fd_sc_hd__nor2b_1 U32905 ( .B_N(n28293), .A(n28292), .Y(n28294) );
  sky130_fd_sc_hd__nand4_1 U32906 ( .A(n28294), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[3]), .C(n29594), .D(
        io_oeb[3]), .Y(n28295) );
  sky130_fd_sc_hd__o21ai_1 U32907 ( .A1(n28297), .A2(n28296), .B1(n28295), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N43) );
  sky130_fd_sc_hd__a21oi_1 U32908 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[4]), .A2(n29594), .B1(
        n29083), .Y(n28303) );
  sky130_fd_sc_hd__o2bb2ai_1 U32909 ( .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[4]), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[4]), .A1_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[4]), .A2_N(n28298), 
        .Y(n28299) );
  sky130_fd_sc_hd__nand3_1 U32910 ( .A(n28299), .B(io_oeb[4]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[4]), .Y(n28302) );
  sky130_fd_sc_hd__o21ai_1 U32912 ( .A1(n28303), .A2(n28302), .B1(n28301), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N44) );
  sky130_fd_sc_hd__a21oi_1 U32913 ( .A1(n12142), .A2(n28304), .B1(n28476), .Y(
        n28309) );
  sky130_fd_sc_hd__o22ai_1 U32914 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[5]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]), .B1(n28305), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[5]), .Y(n28306)
         );
  sky130_fd_sc_hd__a21oi_1 U32915 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[5]), .B1(n28306), 
        .Y(n28307) );
  sky130_fd_sc_hd__nand4_1 U32916 ( .A(n28307), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[5]), .C(n29594), .D(
        io_oeb[7]), .Y(n28308) );
  sky130_fd_sc_hd__o21ai_1 U32917 ( .A1(n28310), .A2(n28309), .B1(n28308), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N45) );
  sky130_fd_sc_hd__a21oi_1 U32918 ( .A1(n29593), .A2(n28311), .B1(n28476), .Y(
        n28316) );
  sky130_fd_sc_hd__o22ai_1 U32919 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[6]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]), .B1(n28312), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[6]), .Y(n28313)
         );
  sky130_fd_sc_hd__a21oi_1 U32920 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[6]), .B1(n28313), 
        .Y(n28314) );
  sky130_fd_sc_hd__nand4_1 U32921 ( .A(n28314), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[6]), .C(n29594), .D(
        io_oeb[26]), .Y(n28315) );
  sky130_fd_sc_hd__o21ai_1 U32922 ( .A1(n28317), .A2(n28316), .B1(n28315), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N46) );
  sky130_fd_sc_hd__a21oi_1 U32923 ( .A1(n29593), .A2(n28318), .B1(n28476), .Y(
        n28323) );
  sky130_fd_sc_hd__o22ai_1 U32924 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[7]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]), .B1(n28319), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[7]), .Y(n28320)
         );
  sky130_fd_sc_hd__a21oi_1 U32925 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[7]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]), .B1(n28320), 
        .Y(n28321) );
  sky130_fd_sc_hd__nand4_1 U32926 ( .A(n28321), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[7]), .C(n29594), .D(
        io_oeb[27]), .Y(n28322) );
  sky130_fd_sc_hd__o21ai_1 U32927 ( .A1(n28324), .A2(n28323), .B1(n28322), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N47) );
  sky130_fd_sc_hd__nor2_1 U32928 ( .A(n28590), .B(n28325), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N11) );
  sky130_fd_sc_hd__a21oi_1 U32931 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[8]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[8]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]), .Y(n28327) );
  sky130_fd_sc_hd__nor2b_1 U32932 ( .B_N(n28328), .A(n28327), .Y(n28329) );
  sky130_fd_sc_hd__nand4_1 U32933 ( .A(n28329), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[8]), .C(n29594), .D(
        io_oeb[28]), .Y(n28330) );
  sky130_fd_sc_hd__nand2_1 U32934 ( .A(n28331), .B(n28330), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N48) );
  sky130_fd_sc_hd__a21oi_1 U32935 ( .A1(n29593), .A2(n28332), .B1(n28476), .Y(
        n28337) );
  sky130_fd_sc_hd__clkinv_1 U32936 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[9]), .Y(n28333) );
  sky130_fd_sc_hd__o221ai_1 U32937 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[9]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[9]), .B1(n28333), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[9]), .C1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[9]), .Y(n28334) );
  sky130_fd_sc_hd__a21oi_1 U32938 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[9]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[9]), .B1(n28334), 
        .Y(n28335) );
  sky130_fd_sc_hd__nand3_1 U32939 ( .A(n28335), .B(n12142), .C(io_oeb[29]), 
        .Y(n28336) );
  sky130_fd_sc_hd__o21ai_1 U32940 ( .A1(n28338), .A2(n28337), .B1(n28336), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N49) );
  sky130_fd_sc_hd__a21oi_1 U32941 ( .A1(n29593), .A2(n28339), .B1(n28476), .Y(
        n28344) );
  sky130_fd_sc_hd__o22ai_1 U32942 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[10]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[10]), .B1(n28340), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[10]), .Y(n28341)
         );
  sky130_fd_sc_hd__a21oi_1 U32943 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[10]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[10]), .B1(n28341), 
        .Y(n28342) );
  sky130_fd_sc_hd__nand4_1 U32944 ( .A(n28342), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[10]), .C(n29594), .D(
        io_oeb[30]), .Y(n28343) );
  sky130_fd_sc_hd__o21ai_1 U32945 ( .A1(n28345), .A2(n28344), .B1(n28343), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N50) );
  sky130_fd_sc_hd__a21oi_1 U32946 ( .A1(n29593), .A2(n28346), .B1(n28476), .Y(
        n28351) );
  sky130_fd_sc_hd__o22ai_1 U32947 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[11]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[11]), .B1(n28347), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[11]), .Y(n28348)
         );
  sky130_fd_sc_hd__a21oi_1 U32948 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[11]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[11]), .B1(n28348), 
        .Y(n28349) );
  sky130_fd_sc_hd__nand4_1 U32949 ( .A(n28349), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[11]), .C(n29593), .D(
        io_oeb[31]), .Y(n28350) );
  sky130_fd_sc_hd__a21oi_1 U32951 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[12]), .A2(n29594), .B1(
        n29084), .Y(n28358) );
  sky130_fd_sc_hd__a21oi_1 U32952 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[12]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[12]), .B1(
        gpio_en_o[12]), .Y(n28353) );
  sky130_fd_sc_hd__o211ai_1 U32953 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[12]), .A2(n28354), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_ier[12]), .C1(n28353), .Y(
        n28357) );
  sky130_fd_sc_hd__o21ai_1 U32955 ( .A1(n28358), .A2(n28357), .B1(n28356), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N52) );
  sky130_fd_sc_hd__nor2_1 U32956 ( .A(n28590), .B(n28359), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N16) );
  sky130_fd_sc_hd__a21oi_1 U32957 ( .A1(n29593), .A2(n28360), .B1(n28476), .Y(
        n28365) );
  sky130_fd_sc_hd__a21oi_1 U32959 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[13]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[13]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13]), .Y(n28361) );
  sky130_fd_sc_hd__nor2b_1 U32960 ( .B_N(n28362), .A(n28361), .Y(n28363) );
  sky130_fd_sc_hd__nand4_1 U32961 ( .A(n28363), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[13]), .C(n29593), .D(
        io_oeb[33]), .Y(n28364) );
  sky130_fd_sc_hd__o21ai_1 U32962 ( .A1(n28366), .A2(n28365), .B1(n28364), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N53) );
  sky130_fd_sc_hd__a21oi_1 U32963 ( .A1(n29593), .A2(n28367), .B1(n28476), .Y(
        n28372) );
  sky130_fd_sc_hd__o22ai_1 U32964 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[14]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14]), .B1(n28368), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[14]), .Y(n28369)
         );
  sky130_fd_sc_hd__a21oi_1 U32965 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[14]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14]), .B1(n28369), 
        .Y(n28370) );
  sky130_fd_sc_hd__nand4_1 U32966 ( .A(n28370), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[14]), .C(n29594), .D(
        io_oeb[34]), .Y(n28371) );
  sky130_fd_sc_hd__o21ai_1 U32967 ( .A1(n28373), .A2(n28372), .B1(n28371), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N54) );
  sky130_fd_sc_hd__a21oi_1 U32968 ( .A1(n29593), .A2(n28374), .B1(n28476), .Y(
        n28379) );
  sky130_fd_sc_hd__o22ai_1 U32969 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[15]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15]), .B1(n28375), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[15]), .Y(n28376)
         );
  sky130_fd_sc_hd__a21oi_1 U32970 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[15]), .B1(n28376), 
        .Y(n28377) );
  sky130_fd_sc_hd__nand4_1 U32971 ( .A(n28377), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[15]), .C(n29594), .D(
        io_oeb[35]), .Y(n28378) );
  sky130_fd_sc_hd__nor2_1 U32973 ( .A(n28590), .B(n28381), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N19) );
  sky130_fd_sc_hd__a21oi_1 U32974 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[16]), .B1(n28590), 
        .Y(n28382) );
  sky130_fd_sc_hd__o21ai_1 U32975 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[16]), .B1(n28382), .Y(
        n28387) );
  sky130_fd_sc_hd__o211ai_1 U32976 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[16]), .A2(n28383), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_ier[16]), .C1(io_oeb[36]), 
        .Y(n28386) );
  sky130_fd_sc_hd__o21ai_1 U32977 ( .A1(n28384), .A2(n28476), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[16]), .Y(n28385) );
  sky130_fd_sc_hd__nor2_1 U32979 ( .A(n28590), .B(n28388), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N20) );
  sky130_fd_sc_hd__a21oi_1 U32980 ( .A1(n12142), .A2(n28389), .B1(n28476), .Y(
        n28394) );
  sky130_fd_sc_hd__a21oi_1 U32981 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[17]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[17]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[17]), .Y(n28392) );
  sky130_fd_sc_hd__nor2_1 U32982 ( .A(n28590), .B(gpio_en_o[17]), .Y(n28391)
         );
  sky130_fd_sc_hd__o21ai_1 U32983 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[17]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[17]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[17]), .Y(n28390) );
  sky130_fd_sc_hd__nand4b_1 U32984 ( .A_N(n28392), .B(n28391), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[17]), .D(n28390), .Y(
        n28393) );
  sky130_fd_sc_hd__o21ai_1 U32985 ( .A1(n28395), .A2(n28394), .B1(n28393), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N57) );
  sky130_fd_sc_hd__a21oi_1 U32986 ( .A1(n28396), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[18]), .B1(
        gpio_en_o[18]), .Y(n28397) );
  sky130_fd_sc_hd__nand2_1 U32987 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[18]), .B(n28397), .Y(
        n28398) );
  sky130_fd_sc_hd__a21oi_1 U32988 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[18]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[18]), .B1(n28398), .Y(
        n28403) );
  sky130_fd_sc_hd__o21ai_1 U32989 ( .A1(n28590), .A2(n28400), .B1(n28399), .Y(
        n28402) );
  sky130_fd_sc_hd__a22o_1 U32991 ( .A1(n28403), .A2(n28402), .B1(n28401), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[18]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N58) );
  sky130_fd_sc_hd__a21oi_1 U32992 ( .A1(n28404), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[19]), .B1(
        gpio_en_o[19]), .Y(n28405) );
  sky130_fd_sc_hd__nand2_1 U32993 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[19]), .B(n28405), .Y(
        n28406) );
  sky130_fd_sc_hd__a21oi_1 U32994 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[19]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[19]), .B1(n28406), .Y(
        n28411) );
  sky130_fd_sc_hd__o21ai_1 U32995 ( .A1(n28590), .A2(n28408), .B1(n28407), .Y(
        n28410) );
  sky130_fd_sc_hd__a22o_1 U32997 ( .A1(n28411), .A2(n28410), .B1(n28409), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[19]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N59) );
  sky130_fd_sc_hd__o21ai_1 U32998 ( .A1(n28412), .A2(n28476), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[20]), .Y(n28420) );
  sky130_fd_sc_hd__a21oi_1 U33000 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[20]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[20]), .B1(n28413), 
        .Y(n28418) );
  sky130_fd_sc_hd__nand3_1 U33002 ( .A(n28418), .B(n28417), .C(n28416), .Y(
        n28419) );
  sky130_fd_sc_hd__nand2_1 U33003 ( .A(n28420), .B(n28419), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N60) );
  sky130_fd_sc_hd__a21oi_1 U33004 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[21]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[21]), .B1(gpio_en_o[21]), 
        .Y(n28421) );
  sky130_fd_sc_hd__nand2_1 U33005 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[21]), .B(n28421), .Y(
        n28422) );
  sky130_fd_sc_hd__a21oi_1 U33006 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[21]), .A2(n28423), 
        .B1(n28422), .Y(n28428) );
  sky130_fd_sc_hd__o21ai_1 U33007 ( .A1(n28590), .A2(n28425), .B1(n28424), .Y(
        n28427) );
  sky130_fd_sc_hd__o21ai_1 U33008 ( .A1(n28590), .A2(
        j202_soc_core_qspi_wb_wdat[21]), .B1(n28506), .Y(n28426) );
  sky130_fd_sc_hd__a22o_1 U33009 ( .A1(n28428), .A2(n28427), .B1(n28426), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[21]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N61) );
  sky130_fd_sc_hd__a21oi_1 U33010 ( .A1(n28429), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[22]), .B1(
        gpio_en_o[22]), .Y(n28430) );
  sky130_fd_sc_hd__nand2_1 U33011 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[22]), .B(n28430), .Y(
        n28431) );
  sky130_fd_sc_hd__a21oi_1 U33012 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[22]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[22]), .B1(n28431), .Y(
        n28436) );
  sky130_fd_sc_hd__o21ai_1 U33013 ( .A1(n28590), .A2(n28433), .B1(n28432), .Y(
        n28435) );
  sky130_fd_sc_hd__a22o_1 U33015 ( .A1(n28436), .A2(n28435), .B1(n28434), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[22]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N62) );
  sky130_fd_sc_hd__a21oi_1 U33016 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[23]), .A2(n29594), 
        .B1(n29085), .Y(n28437) );
  sky130_fd_sc_hd__nor2_1 U33017 ( .A(gpio_en_o[23]), .B(n28437), .Y(n28442)
         );
  sky130_fd_sc_hd__a21oi_1 U33019 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[23]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[23]), .B1(n28439), 
        .Y(n28441) );
  sky130_fd_sc_hd__o21ai_1 U33020 ( .A1(n28590), .A2(
        j202_soc_core_qspi_wb_wdat[23]), .B1(n28506), .Y(n28440) );
  sky130_fd_sc_hd__a22o_1 U33021 ( .A1(n28442), .A2(n28441), .B1(n28440), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[23]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N63) );
  sky130_fd_sc_hd__nor2_1 U33022 ( .A(n28590), .B(n28443), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N27) );
  sky130_fd_sc_hd__nand2_1 U33023 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[24]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[24]), .Y(n28444) );
  sky130_fd_sc_hd__o211ai_1 U33024 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[24]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[24]), .B1(n29594), 
        .C1(n28444), .Y(n28450) );
  sky130_fd_sc_hd__clkinv_1 U33025 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[24]), .Y(n28446) );
  sky130_fd_sc_hd__o211ai_1 U33026 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[24]), .A2(n28446), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[24]), .C1(n28445), .Y(
        n28449) );
  sky130_fd_sc_hd__o21ai_1 U33027 ( .A1(n28447), .A2(n28476), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[24]), .Y(n28448) );
  sky130_fd_sc_hd__o21ai_1 U33028 ( .A1(n28450), .A2(n28449), .B1(n28448), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N64) );
  sky130_fd_sc_hd__a21oi_1 U33029 ( .A1(n28451), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[25]), .B1(
        gpio_en_o[25]), .Y(n28452) );
  sky130_fd_sc_hd__nand2_1 U33030 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[25]), .B(n28452), .Y(
        n28453) );
  sky130_fd_sc_hd__a21oi_1 U33031 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[25]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[25]), .B1(n28453), .Y(
        n28458) );
  sky130_fd_sc_hd__o21ai_1 U33032 ( .A1(n28590), .A2(n28455), .B1(n28454), .Y(
        n28457) );
  sky130_fd_sc_hd__a22o_1 U33034 ( .A1(n28458), .A2(n28457), .B1(n28456), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[25]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N65) );
  sky130_fd_sc_hd__a21oi_1 U33035 ( .A1(n28459), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[26]), .B1(
        gpio_en_o[26]), .Y(n28460) );
  sky130_fd_sc_hd__nand2_1 U33036 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[26]), .B(n28460), .Y(
        n28461) );
  sky130_fd_sc_hd__a21oi_1 U33037 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[26]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[26]), .B1(n28461), .Y(
        n28466) );
  sky130_fd_sc_hd__o21ai_1 U33038 ( .A1(n28590), .A2(n28463), .B1(n28462), .Y(
        n28465) );
  sky130_fd_sc_hd__a22o_1 U33040 ( .A1(n28466), .A2(n28465), .B1(n28464), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[26]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N66) );
  sky130_fd_sc_hd__a21oi_1 U33041 ( .A1(n28467), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[27]), .B1(
        gpio_en_o[27]), .Y(n28468) );
  sky130_fd_sc_hd__nand2_1 U33042 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[27]), .B(n28468), .Y(
        n28469) );
  sky130_fd_sc_hd__a21oi_1 U33043 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[27]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[27]), .B1(n28469), .Y(
        n28474) );
  sky130_fd_sc_hd__o21ai_1 U33044 ( .A1(n28590), .A2(n28471), .B1(n28470), .Y(
        n28473) );
  sky130_fd_sc_hd__a22o_1 U33046 ( .A1(n28474), .A2(n28473), .B1(n28472), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[27]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N67) );
  sky130_fd_sc_hd__nor2_1 U33047 ( .A(n28590), .B(n28475), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N31) );
  sky130_fd_sc_hd__o21ai_1 U33048 ( .A1(n28477), .A2(n28476), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[28]), .Y(n28484) );
  sky130_fd_sc_hd__o21ai_1 U33049 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[28]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[28]), .B1(n12142), 
        .Y(n28478) );
  sky130_fd_sc_hd__a21oi_1 U33050 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[28]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[28]), .B1(n28478), .Y(
        n28482) );
  sky130_fd_sc_hd__nand2_1 U33051 ( .A(n28479), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[28]), .Y(n28481) );
  sky130_fd_sc_hd__nand4_1 U33052 ( .A(n28482), .B(n28481), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[28]), .D(n28480), .Y(
        n28483) );
  sky130_fd_sc_hd__nand2_1 U33053 ( .A(n28484), .B(n28483), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N68) );
  sky130_fd_sc_hd__a21oi_1 U33054 ( .A1(n28485), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[29]), .B1(
        gpio_en_o[29]), .Y(n28486) );
  sky130_fd_sc_hd__nand2_1 U33055 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[29]), .B(n28486), .Y(
        n28487) );
  sky130_fd_sc_hd__a21oi_1 U33056 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[29]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[29]), .B1(n28487), .Y(
        n28492) );
  sky130_fd_sc_hd__o21ai_1 U33057 ( .A1(n28590), .A2(n28489), .B1(n28488), .Y(
        n28491) );
  sky130_fd_sc_hd__a22o_1 U33059 ( .A1(n28492), .A2(n28491), .B1(n28490), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[29]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N69) );
  sky130_fd_sc_hd__a21oi_1 U33060 ( .A1(n28493), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[30]), .B1(
        gpio_en_o[30]), .Y(n28494) );
  sky130_fd_sc_hd__nand2_1 U33061 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[30]), .B(n28494), .Y(
        n28495) );
  sky130_fd_sc_hd__a21oi_1 U33062 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[30]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[30]), .B1(n28495), .Y(
        n28500) );
  sky130_fd_sc_hd__o21ai_1 U33063 ( .A1(n28590), .A2(n28497), .B1(n28496), .Y(
        n28499) );
  sky130_fd_sc_hd__o21ai_1 U33064 ( .A1(n28590), .A2(
        j202_soc_core_qspi_wb_wdat[30]), .B1(n28506), .Y(n28498) );
  sky130_fd_sc_hd__a22o_1 U33065 ( .A1(n28500), .A2(n28499), .B1(n28498), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[30]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N70) );
  sky130_fd_sc_hd__a21oi_1 U33066 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[31]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[31]), .B1(gpio_en_o[31]), 
        .Y(n28501) );
  sky130_fd_sc_hd__nand2_1 U33067 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[31]), .B(n28501), .Y(
        n28502) );
  sky130_fd_sc_hd__a21oi_1 U33068 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[31]), .A2(n28503), 
        .B1(n28502), .Y(n28509) );
  sky130_fd_sc_hd__o21ai_1 U33069 ( .A1(n28590), .A2(n28505), .B1(n28504), .Y(
        n28508) );
  sky130_fd_sc_hd__o21ai_1 U33070 ( .A1(n28590), .A2(
        j202_soc_core_qspi_wb_wdat[31]), .B1(n28506), .Y(n28507) );
  sky130_fd_sc_hd__a22o_1 U33071 ( .A1(n28509), .A2(n28508), .B1(n28507), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[31]), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N71) );
  sky130_fd_sc_hd__a22o_1 U33072 ( .A1(n28510), .A2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[4]), .B1(n12071), .B2(j202_soc_core_intr_vec__4_), .X(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N7) );
  sky130_fd_sc_hd__a22o_1 U33073 ( .A1(n28510), .A2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[6]), .B1(n12071), .B2(j202_soc_core_intr_vec__6_), .X(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N9) );
  sky130_fd_sc_hd__o22ai_1 U33074 ( .A1(n28518), .A2(n28512), .B1(n28511), 
        .B2(n28515), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N4) );
  sky130_fd_sc_hd__o22ai_1 U33075 ( .A1(n28518), .A2(n28514), .B1(n28513), 
        .B2(n28515), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N5) );
  sky130_fd_sc_hd__o22ai_1 U33076 ( .A1(n28518), .A2(n28517), .B1(n28516), 
        .B2(n28515), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N6) );
  sky130_fd_sc_hd__o22a_1 U33077 ( .A1(n28520), .A2(
        j202_soc_core_intc_core_00_rg_ipr[96]), .B1(n29086), .B2(n28519), .X(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U33078 ( .A1(n28614), .A2(n28526), .B1(n28521), 
        .B2(n28524), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U33079 ( .A1(n28614), .A2(n28538), .B1(n28522), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U33080 ( .A1(n28614), .A2(n28535), .B1(n28523), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U33081 ( .A1(n28610), .A2(n28526), .B1(n28525), 
        .B2(n28524), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U33082 ( .A1(n28544), .A2(n28610), .B1(n28527), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U33083 ( .A1(n28596), .A2(n28541), .B1(n28528), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U33084 ( .A1(n28598), .A2(n28541), .B1(n28529), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U33085 ( .A1(n28602), .A2(n28535), .B1(n28530), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U33086 ( .A1(n28605), .A2(n28547), .B1(n28531), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U33087 ( .A1(n28544), .A2(n28605), .B1(n28532), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U33088 ( .A1(n28605), .A2(n28535), .B1(n28534), 
        .B2(n28533), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U33089 ( .A1(n28605), .A2(n28538), .B1(n28537), 
        .B2(n28536), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U33090 ( .A1(n28605), .A2(n28541), .B1(n28540), 
        .B2(n28539), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U33091 ( .A1(n28544), .A2(n28600), .B1(n28543), 
        .B2(n28542), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U33092 ( .A1(n28600), .A2(n28547), .B1(n28546), 
        .B2(n28545), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__a21o_1 U33093 ( .A1(n28549), .A2(
        j202_soc_core_wbqspiflash_00_spi_out[1]), .B1(n28548), .X(
        j202_soc_core_wbqspiflash_00_N606) );
  sky130_fd_sc_hd__xnor2_1 U33095 ( .A(j202_soc_core_uart_TOP_rxd_s), .B(
        j202_soc_core_uart_TOP_rxd_r), .Y(n28553) );
  sky130_fd_sc_hd__nor2_1 U33096 ( .A(n28590), .B(n28553), .Y(
        j202_soc_core_uart_TOP_N102) );
  sky130_fd_sc_hd__nand3_1 U33097 ( .A(n28553), .B(n29593), .C(n28559), .Y(
        j202_soc_core_uart_TOP_N101) );
  sky130_fd_sc_hd__nand2_1 U33098 ( .A(n29087), .B(
        j202_soc_core_uart_TOP_change), .Y(n28555) );
  sky130_fd_sc_hd__nor2_1 U33099 ( .A(j202_soc_core_uart_TOP_change), .B(
        j202_soc_core_uart_TOP_dpll_state[0]), .Y(n28557) );
  sky130_fd_sc_hd__nand2_1 U33100 ( .A(n28557), .B(
        j202_soc_core_uart_sio_ce_x4), .Y(n28554) );
  sky130_fd_sc_hd__o211ai_1 U33101 ( .A1(j202_soc_core_uart_sio_ce_x4), .A2(
        n28556), .B1(n28555), .C1(n28554), .Y(n132) );
  sky130_fd_sc_hd__o21ai_1 U33102 ( .A1(n28559), .A2(n28557), .B1(
        j202_soc_core_uart_TOP_dpll_state[1]), .Y(n28558) );
  sky130_fd_sc_hd__nor2_1 U33104 ( .A(j202_soc_core_uart_TOP_shift_en), .B(
        j202_soc_core_uart_TOP_shift_en_r), .Y(n28561) );
  sky130_fd_sc_hd__nor2_1 U33105 ( .A(j202_soc_core_uart_TOP_hold_reg[0]), .B(
        n28561), .Y(n28563) );
  sky130_fd_sc_hd__xnor2_1 U33107 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[4]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[4]), .Y(n28568) );
  sky130_fd_sc_hd__xnor2_1 U33108 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[1]), .Y(n28567) );
  sky130_fd_sc_hd__xnor2_1 U33109 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[0]), .Y(n28566) );
  sky130_fd_sc_hd__xnor2_1 U33110 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[2]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[2]), .Y(n28565) );
  sky130_fd_sc_hd__nand4_1 U33111 ( .A(n28568), .B(n28567), .C(n28566), .D(
        n28565), .Y(n28579) );
  sky130_fd_sc_hd__xnor2_1 U33112 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[7]), .Y(n28572) );
  sky130_fd_sc_hd__xnor2_1 U33113 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[10]), .Y(n28571) );
  sky130_fd_sc_hd__xnor2_1 U33114 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[8]), .Y(n28570) );
  sky130_fd_sc_hd__xnor2_1 U33115 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[11]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[11]), .Y(n28569) );
  sky130_fd_sc_hd__nand4_1 U33116 ( .A(n28572), .B(n28571), .C(n28570), .D(
        n28569), .Y(n28578) );
  sky130_fd_sc_hd__xnor2_1 U33117 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[5]), .Y(n28576) );
  sky130_fd_sc_hd__xnor2_1 U33118 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[3]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[3]), .Y(n28575) );
  sky130_fd_sc_hd__xnor2_1 U33119 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[6]), .Y(n28574) );
  sky130_fd_sc_hd__xnor2_1 U33120 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]), .B(
        j202_soc_core_bldc_core_00_pwm_duty[9]), .Y(n28573) );
  sky130_fd_sc_hd__nand4_1 U33121 ( .A(n28576), .B(n28575), .C(n28574), .D(
        n28573), .Y(n28577) );
  sky130_fd_sc_hd__o31ai_1 U33122 ( .A1(n28579), .A2(n28578), .A3(n28577), 
        .B1(j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld), .Y(n28580) );
  sky130_fd_sc_hd__o31ai_1 U33123 ( .A1(n28582), .A2(n28581), .A3(io_in[25]), 
        .B1(n28580), .Y(n26) );
  sky130_fd_sc_hd__xnor2_1 U33124 ( .A(j202_soc_core_bldc_core_00_comm[1]), 
        .B(j202_soc_core_bldc_core_00_comm[0]), .Y(n28587) );
  sky130_fd_sc_hd__nor2_1 U33125 ( .A(n28585), .B(n28587), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posa) );
  sky130_fd_sc_hd__o21a_1 U33126 ( .A1(n29089), .A2(n29088), .B1(n28587), .X(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posb) );
  sky130_fd_sc_hd__or3_1 U33127 ( .A(j202_soc_core_bldc_core_00_comm[0]), .B(
        n28583), .C(n28588), .X(n28584) );
  sky130_fd_sc_hd__o31ai_1 U33128 ( .A1(j202_soc_core_bldc_core_00_comm[1]), 
        .A2(n28586), .A3(n28585), .B1(n28584), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_negb) );
  sky130_fd_sc_hd__nor2_1 U33129 ( .A(n28588), .B(n28587), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posc) );
  sky130_fd_sc_hd__nor2_1 U33130 ( .A(n28590), .B(n28589), .Y(n28739) );
  sky130_fd_sc_hd__or3_1 U33131 ( .A(n28637), .B(n28731), .C(n28743), .X(
        j202_soc_core_wbqspiflash_00_lldriver_N315) );
  sky130_fd_sc_hd__a22oi_1 U33132 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[27]), .B1(n28733), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[24]), .Y(n28592) );
  sky130_fd_sc_hd__a22oi_1 U33133 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[27]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[24]), .B2(n28734), .Y(n28591) );
  sky130_fd_sc_hd__o211ai_1 U33134 ( .A1(n28726), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B1(n28592), .C1(n28591), 
        .Y(j202_soc_core_wbqspiflash_00_lldriver_N419) );
  sky130_fd_sc_hd__a22oi_1 U33135 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[2]), .B1(n28719), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[2]), .Y(n28593) );
  sky130_fd_sc_hd__nand2_1 U33137 ( .A(n28595), .B(
        j202_soc_core_intc_core_00_bs_addr[7]), .Y(n28616) );
  sky130_fd_sc_hd__nor2_1 U33138 ( .A(n28596), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N14) );
  sky130_fd_sc_hd__nor2_1 U33139 ( .A(n28597), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N17) );
  sky130_fd_sc_hd__nor2_1 U33140 ( .A(n28598), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N16) );
  sky130_fd_sc_hd__nor2_1 U33141 ( .A(n28599), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N11) );
  sky130_fd_sc_hd__nor2_1 U33142 ( .A(n28600), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N22) );
  sky130_fd_sc_hd__nor2_1 U33143 ( .A(n28601), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N12) );
  sky130_fd_sc_hd__nor2_1 U33144 ( .A(n28602), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N20) );
  sky130_fd_sc_hd__nor2_1 U33145 ( .A(n28603), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N4) );
  sky130_fd_sc_hd__nor2_1 U33146 ( .A(n28604), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N23) );
  sky130_fd_sc_hd__nor2_1 U33147 ( .A(n28605), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N21) );
  sky130_fd_sc_hd__nor2_1 U33148 ( .A(n28606), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N19) );
  sky130_fd_sc_hd__nor2_1 U33149 ( .A(n28607), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N18) );
  sky130_fd_sc_hd__nor2_1 U33150 ( .A(n28608), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N15) );
  sky130_fd_sc_hd__nor2_1 U33151 ( .A(n28609), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N13) );
  sky130_fd_sc_hd__nor2_1 U33152 ( .A(n28610), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N10) );
  sky130_fd_sc_hd__nor2_1 U33153 ( .A(n28611), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N9) );
  sky130_fd_sc_hd__nor2_1 U33154 ( .A(n28612), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N8) );
  sky130_fd_sc_hd__nor2_1 U33155 ( .A(n28613), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N7) );
  sky130_fd_sc_hd__nor2_1 U33156 ( .A(n28614), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N6) );
  sky130_fd_sc_hd__nor2_1 U33157 ( .A(n28615), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N5) );
  sky130_fd_sc_hd__nor2_1 U33158 ( .A(n28881), .B(n28616), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N3) );
  sky130_fd_sc_hd__or3_1 U33159 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[0]), .C(n28901), .X(io_oeb[11]) );
  sky130_fd_sc_hd__nor3_1 U33160 ( .A(n28619), .B(n28618), .C(n28617), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt0_to1) );
  sky130_fd_sc_hd__nor2_1 U33161 ( .A(n28622), .B(n28621), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt1_to1) );
  sky130_fd_sc_hd__nor2b_1 U33162 ( .B_N(j202_soc_core_uart_TOP_rx_sio_ce_r1), 
        .A(j202_soc_core_uart_TOP_rx_sio_ce_r2), .Y(
        j202_soc_core_uart_TOP_N118) );
  sky130_fd_sc_hd__nor2_1 U33163 ( .A(j202_soc_core_uart_TOP_shift_en), .B(
        j202_soc_core_uart_TOP_txf_empty_r), .Y(j202_soc_core_uart_TOP_N137)
         );
  sky130_fd_sc_hd__nand3_1 U33164 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[1]), 
        .B(n28624), .C(n28623), .Y(j202_soc_core_uart_TOP_N128) );
  sky130_fd_sc_hd__nand4b_1 U33165 ( .A_N(j202_soc_core_uart_TOP_tx_bit_cnt[1]), .B(j202_soc_core_uart_TOP_tx_bit_cnt[0]), .C(
        j202_soc_core_uart_TOP_tx_bit_cnt[3]), .D(n28625), .Y(
        j202_soc_core_uart_TOP_N123) );
  sky130_fd_sc_hd__nor2b_1 U33166 ( .B_N(n29090), .A(
        j202_soc_core_uart_BRG_sio_ce_r), .Y(j202_soc_core_uart_BRG_N59) );
  sky130_fd_sc_hd__o21ai_1 U33167 ( .A1(j202_soc_core_uart_BRG_ps[7]), .A2(
        n28628), .B1(n28626), .Y(n28627) );
  sky130_fd_sc_hd__a21oi_1 U33168 ( .A1(j202_soc_core_uart_BRG_ps[7]), .A2(
        n28628), .B1(n28627), .Y(j202_soc_core_uart_BRG_N19) );
  sky130_fd_sc_hd__o21ai_1 U33169 ( .A1(j202_soc_core_uart_BRG_br_cnt[7]), 
        .A2(n28632), .B1(n28630), .Y(n28631) );
  sky130_fd_sc_hd__a21oi_1 U33170 ( .A1(j202_soc_core_uart_BRG_br_cnt[7]), 
        .A2(n28632), .B1(n28631), .Y(j202_soc_core_uart_BRG_N42) );
  sky130_fd_sc_hd__a31oi_1 U33171 ( .A1(n29092), .A2(wbs_we_i), .A3(
        wbs_sel_i[0]), .B1(wb_rst_i), .Y(n28633) );
  sky130_fd_sc_hd__nand2_1 U33172 ( .A(start_n_reg[1]), .B(n28633), .Y(n10) );
  sky130_fd_sc_hd__nand2_1 U33173 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .B(
        j202_soc_core_wbqspiflash_00_alt_ctrl), .Y(n28634) );
  sky130_fd_sc_hd__o21ai_0 U33174 ( .A1(n28635), .A2(
        j202_soc_core_wbqspiflash_00_spif_override), .B1(n28634), .Y(io_out[9]) );
  sky130_fd_sc_hd__a22o_1 U33175 ( .A1(n28636), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_dir), .B1(n28734), .B2(
        j202_soc_core_wbqspiflash_00_spi_dir), .X(
        j202_soc_core_wbqspiflash_00_lldriver_N355) );
  sky130_fd_sc_hd__nand2b_1 U33176 ( .A_N(n28636), .B(n28723), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N356) );
  sky130_fd_sc_hd__or3_1 U33177 ( .A(n28647), .B(n28637), .C(n28646), .X(
        j202_soc_core_wbqspiflash_00_lldriver_N354) );
  sky130_fd_sc_hd__nand2_1 U33178 ( .A(n28638), .B(
        j202_soc_core_wbqspiflash_00_spi_wr), .Y(n28639) );
  sky130_fd_sc_hd__a21o_1 U33179 ( .A1(n28642), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .B1(n28641), .X(
        n28643) );
  sky130_fd_sc_hd__or4_1 U33180 ( .A(n28645), .B(n28644), .C(n28643), .D(
        n29091), .X(j202_soc_core_wbqspiflash_00_lldriver_N321) );
  sky130_fd_sc_hd__nor2_1 U33181 ( .A(n28647), .B(n28646), .Y(n28648) );
  sky130_fd_sc_hd__nand2_1 U33182 ( .A(n28649), .B(n28648), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N313) );
  sky130_fd_sc_hd__a22oi_1 U33183 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[3]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[0]), .B2(n28733), .Y(
        n28651) );
  sky130_fd_sc_hd__a22oi_1 U33184 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[3]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[4]), .Y(n28650) );
  sky130_fd_sc_hd__o211ai_1 U33185 ( .A1(n28652), .A2(n28723), .B1(n28651), 
        .C1(n28650), .Y(j202_soc_core_wbqspiflash_00_lldriver_N395) );
  sky130_fd_sc_hd__a22oi_1 U33186 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[4]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[1]), .B2(n28733), .Y(
        n28654) );
  sky130_fd_sc_hd__a22oi_1 U33187 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[4]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[5]), .Y(n28653) );
  sky130_fd_sc_hd__o211ai_1 U33188 ( .A1(n28655), .A2(n28723), .B1(n28654), 
        .C1(n28653), .Y(j202_soc_core_wbqspiflash_00_lldriver_N396) );
  sky130_fd_sc_hd__a22oi_1 U33189 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[5]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[2]), .B2(n28733), .Y(
        n28657) );
  sky130_fd_sc_hd__a22oi_1 U33190 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[5]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[6]), .Y(n28656) );
  sky130_fd_sc_hd__o211ai_1 U33191 ( .A1(n28658), .A2(n28723), .B1(n28657), 
        .C1(n28656), .Y(j202_soc_core_wbqspiflash_00_lldriver_N397) );
  sky130_fd_sc_hd__a22oi_1 U33192 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[6]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[3]), .B2(n28733), .Y(
        n28660) );
  sky130_fd_sc_hd__a22oi_1 U33193 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[6]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[7]), .Y(n28659) );
  sky130_fd_sc_hd__o211ai_1 U33194 ( .A1(n28661), .A2(n28723), .B1(n28660), 
        .C1(n28659), .Y(j202_soc_core_wbqspiflash_00_lldriver_N398) );
  sky130_fd_sc_hd__a22oi_1 U33195 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[7]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[4]), .B2(n28733), .Y(
        n28663) );
  sky130_fd_sc_hd__a22oi_1 U33196 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[7]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[8]), .Y(n28662) );
  sky130_fd_sc_hd__o211ai_1 U33197 ( .A1(n28723), .A2(n28664), .B1(n28663), 
        .C1(n28662), .Y(j202_soc_core_wbqspiflash_00_lldriver_N399) );
  sky130_fd_sc_hd__a22oi_1 U33198 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[8]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[5]), .B2(n28733), .Y(
        n28666) );
  sky130_fd_sc_hd__a22oi_1 U33199 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[8]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[9]), .Y(n28665) );
  sky130_fd_sc_hd__o211ai_1 U33200 ( .A1(n28723), .A2(n28667), .B1(n28666), 
        .C1(n28665), .Y(j202_soc_core_wbqspiflash_00_lldriver_N400) );
  sky130_fd_sc_hd__a22oi_1 U33201 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[9]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[6]), .B2(n28733), .Y(
        n28669) );
  sky130_fd_sc_hd__a22oi_1 U33202 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[9]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[10]), .Y(n28668) );
  sky130_fd_sc_hd__o211ai_1 U33203 ( .A1(n28723), .A2(n28670), .B1(n28669), 
        .C1(n28668), .Y(j202_soc_core_wbqspiflash_00_lldriver_N401) );
  sky130_fd_sc_hd__a22oi_1 U33204 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[10]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[7]), .B2(n28733), .Y(
        n28672) );
  sky130_fd_sc_hd__a22oi_1 U33205 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[10]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[11]), .Y(n28671) );
  sky130_fd_sc_hd__o211ai_1 U33206 ( .A1(n28723), .A2(n28673), .B1(n28672), 
        .C1(n28671), .Y(j202_soc_core_wbqspiflash_00_lldriver_N402) );
  sky130_fd_sc_hd__a22oi_1 U33207 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[11]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[8]), .B2(n28733), .Y(
        n28675) );
  sky130_fd_sc_hd__a22oi_1 U33208 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[11]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[12]), .Y(n28674) );
  sky130_fd_sc_hd__o211ai_1 U33209 ( .A1(n28723), .A2(n28676), .B1(n28675), 
        .C1(n28674), .Y(j202_soc_core_wbqspiflash_00_lldriver_N403) );
  sky130_fd_sc_hd__a22oi_1 U33210 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[12]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[9]), .B2(n28733), .Y(
        n28678) );
  sky130_fd_sc_hd__a22oi_1 U33211 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[12]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[13]), .Y(n28677) );
  sky130_fd_sc_hd__o211ai_1 U33212 ( .A1(n28723), .A2(n28679), .B1(n28678), 
        .C1(n28677), .Y(j202_soc_core_wbqspiflash_00_lldriver_N404) );
  sky130_fd_sc_hd__a22oi_1 U33213 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[13]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[10]), .B2(n28733), .Y(
        n28681) );
  sky130_fd_sc_hd__a22oi_1 U33214 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[13]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[14]), .Y(n28680) );
  sky130_fd_sc_hd__o211ai_1 U33215 ( .A1(n28723), .A2(n28682), .B1(n28681), 
        .C1(n28680), .Y(j202_soc_core_wbqspiflash_00_lldriver_N405) );
  sky130_fd_sc_hd__a22oi_1 U33216 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[14]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[11]), .B2(n28733), .Y(
        n28684) );
  sky130_fd_sc_hd__a22oi_1 U33217 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[14]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[15]), .Y(n28683) );
  sky130_fd_sc_hd__o211ai_1 U33218 ( .A1(n28723), .A2(n28685), .B1(n28684), 
        .C1(n28683), .Y(j202_soc_core_wbqspiflash_00_lldriver_N406) );
  sky130_fd_sc_hd__a22oi_1 U33219 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[15]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[12]), .B2(n28733), .Y(
        n28687) );
  sky130_fd_sc_hd__a22oi_1 U33220 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[15]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[16]), .Y(n28686) );
  sky130_fd_sc_hd__o211ai_1 U33221 ( .A1(n28723), .A2(n28688), .B1(n28687), 
        .C1(n28686), .Y(j202_soc_core_wbqspiflash_00_lldriver_N407) );
  sky130_fd_sc_hd__a22oi_1 U33222 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[16]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[13]), .B2(n28733), .Y(
        n28690) );
  sky130_fd_sc_hd__a22oi_1 U33223 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[16]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[17]), .Y(n28689) );
  sky130_fd_sc_hd__o211ai_1 U33224 ( .A1(n28723), .A2(n28691), .B1(n28690), 
        .C1(n28689), .Y(j202_soc_core_wbqspiflash_00_lldriver_N408) );
  sky130_fd_sc_hd__a22oi_1 U33225 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[17]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[14]), .B2(n28733), .Y(
        n28693) );
  sky130_fd_sc_hd__a22oi_1 U33226 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[17]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[18]), .Y(n28692) );
  sky130_fd_sc_hd__o211ai_1 U33227 ( .A1(n28723), .A2(n28694), .B1(n28693), 
        .C1(n28692), .Y(j202_soc_core_wbqspiflash_00_lldriver_N409) );
  sky130_fd_sc_hd__a22oi_1 U33228 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[18]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[15]), .B2(n28733), .Y(
        n28696) );
  sky130_fd_sc_hd__a22oi_1 U33229 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[18]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[19]), .Y(n28695) );
  sky130_fd_sc_hd__o211ai_1 U33230 ( .A1(n28723), .A2(n28697), .B1(n28696), 
        .C1(n28695), .Y(j202_soc_core_wbqspiflash_00_lldriver_N410) );
  sky130_fd_sc_hd__a22oi_1 U33231 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[19]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[16]), .B2(n28733), .Y(
        n28699) );
  sky130_fd_sc_hd__a22oi_1 U33232 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[19]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[20]), .Y(n28698) );
  sky130_fd_sc_hd__o211ai_1 U33233 ( .A1(n28723), .A2(n28700), .B1(n28699), 
        .C1(n28698), .Y(j202_soc_core_wbqspiflash_00_lldriver_N411) );
  sky130_fd_sc_hd__a22oi_1 U33234 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[20]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[17]), .B2(n28733), .Y(
        n28702) );
  sky130_fd_sc_hd__a22oi_1 U33235 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[20]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[21]), .Y(n28701) );
  sky130_fd_sc_hd__o211ai_1 U33236 ( .A1(n28723), .A2(n28703), .B1(n28702), 
        .C1(n28701), .Y(j202_soc_core_wbqspiflash_00_lldriver_N412) );
  sky130_fd_sc_hd__a22oi_1 U33237 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[21]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[18]), .B2(n28733), .Y(
        n28705) );
  sky130_fd_sc_hd__a22oi_1 U33238 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[21]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[22]), .Y(n28704) );
  sky130_fd_sc_hd__o211ai_1 U33239 ( .A1(n28723), .A2(n28706), .B1(n28705), 
        .C1(n28704), .Y(j202_soc_core_wbqspiflash_00_lldriver_N413) );
  sky130_fd_sc_hd__a22oi_1 U33240 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[22]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[19]), .B2(n28733), .Y(
        n28708) );
  sky130_fd_sc_hd__a22oi_1 U33241 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[22]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[23]), .Y(n28707) );
  sky130_fd_sc_hd__o211ai_1 U33242 ( .A1(n28723), .A2(n28709), .B1(n28708), 
        .C1(n28707), .Y(j202_soc_core_wbqspiflash_00_lldriver_N414) );
  sky130_fd_sc_hd__a22oi_1 U33243 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[23]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[20]), .B2(n28733), .Y(
        n28711) );
  sky130_fd_sc_hd__a22oi_1 U33244 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[23]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[24]), .Y(n28710) );
  sky130_fd_sc_hd__o211ai_1 U33245 ( .A1(n28723), .A2(n28712), .B1(n28711), 
        .C1(n28710), .Y(j202_soc_core_wbqspiflash_00_lldriver_N415) );
  sky130_fd_sc_hd__a22oi_1 U33246 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[24]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[21]), .B2(n28733), .Y(
        n28714) );
  sky130_fd_sc_hd__a22oi_1 U33247 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[24]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[25]), .Y(n28713) );
  sky130_fd_sc_hd__o211ai_1 U33248 ( .A1(n28723), .A2(n28715), .B1(n28714), 
        .C1(n28713), .Y(j202_soc_core_wbqspiflash_00_lldriver_N416) );
  sky130_fd_sc_hd__a22oi_1 U33249 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[25]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[22]), .B2(n28733), .Y(
        n28717) );
  sky130_fd_sc_hd__a22oi_1 U33250 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[25]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[26]), .Y(n28716) );
  sky130_fd_sc_hd__o211ai_1 U33251 ( .A1(n28723), .A2(n28718), .B1(n28717), 
        .C1(n28716), .Y(j202_soc_core_wbqspiflash_00_lldriver_N417) );
  sky130_fd_sc_hd__a22oi_1 U33252 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[26]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[23]), .B2(n28733), .Y(
        n28721) );
  sky130_fd_sc_hd__a22oi_1 U33253 ( .A1(n28719), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[26]), .B1(n28727), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[27]), .Y(n28720) );
  sky130_fd_sc_hd__o211ai_1 U33254 ( .A1(n28723), .A2(n28722), .B1(n28721), 
        .C1(n28720), .Y(j202_soc_core_wbqspiflash_00_lldriver_N418) );
  sky130_fd_sc_hd__a22oi_1 U33255 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[28]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[25]), .B2(n28733), .Y(
        n28725) );
  sky130_fd_sc_hd__a22oi_1 U33256 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_in[25]), .A2(n28734), .B1(n28727), 
        .B2(j202_soc_core_wbqspiflash_00_spi_in[29]), .Y(n28724) );
  sky130_fd_sc_hd__o211ai_1 U33257 ( .A1(n28740), .A2(n28726), .B1(n28725), 
        .C1(n28724), .Y(j202_soc_core_wbqspiflash_00_lldriver_N420) );
  sky130_fd_sc_hd__a22oi_1 U33258 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[29]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[26]), .B2(n28733), .Y(
        n28729) );
  sky130_fd_sc_hd__a22oi_1 U33259 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_in[26]), .A2(n28734), .B1(n28727), 
        .B2(j202_soc_core_wbqspiflash_00_spi_in[30]), .Y(n28728) );
  sky130_fd_sc_hd__o211ai_1 U33260 ( .A1(n28740), .A2(n28730), .B1(n28729), 
        .C1(n28728), .Y(j202_soc_core_wbqspiflash_00_lldriver_N421) );
  sky130_fd_sc_hd__nand2_1 U33261 ( .A(j202_soc_core_wbqspiflash_00_spi_in[31]), .B(n28737), .Y(n28745) );
  sky130_fd_sc_hd__a21oi_1 U33262 ( .A1(n28732), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[31]), .B1(n28731), .Y(
        n28736) );
  sky130_fd_sc_hd__a22oi_1 U33263 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_in[28]), .A2(n28734), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[28]), .B2(n28733), .Y(
        n28735) );
  sky130_fd_sc_hd__o211ai_1 U33264 ( .A1(j202_soc_core_wbqspiflash_00_spi_spd), 
        .A2(n28745), .B1(n28736), .C1(n28735), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N316) );
  sky130_fd_sc_hd__nand2_1 U33265 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[30]), .B(n28743), .Y(
        n28742) );
  sky130_fd_sc_hd__nand2_1 U33266 ( .A(j202_soc_core_wbqspiflash_00_spi_in[30]), .B(n28737), .Y(n28741) );
  sky130_fd_sc_hd__and3_1 U33267 ( .A(n28740), .B(n28739), .C(n28738), .X(
        n28744) );
  sky130_fd_sc_hd__nand3_1 U33268 ( .A(n28742), .B(n28741), .C(n28744), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N318) );
  sky130_fd_sc_hd__nand2_1 U33269 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[31]), .B(n28743), .Y(
        n28746) );
  sky130_fd_sc_hd__nand3_1 U33270 ( .A(n28746), .B(n28745), .C(n28744), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N319) );
  sky130_fd_sc_hd__nand2_1 U33271 ( .A(n28748), .B(n28747), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N310) );
  sky130_fd_sc_hd__a21oi_1 U33272 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[0]), .A2(
        j202_soc_core_wbqspiflash_00_reset_counter[1]), .B1(n28749), .Y(n28750) );
  sky130_fd_sc_hd__nor2_1 U33273 ( .A(n28751), .B(n28750), .Y(
        j202_soc_core_wbqspiflash_00_N615) );
  sky130_fd_sc_hd__nor2_1 U33274 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[0]), 
        .B(j202_soc_core_uart_TOP_tx_fifo_rp[1]), .Y(n28778) );
  sky130_fd_sc_hd__a22oi_1 U33275 ( .A1(n28777), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[0]), .B1(n28778), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[24]), .Y(n28755) );
  sky130_fd_sc_hd__nor2_1 U33276 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[0]), 
        .B(n28752), .Y(n28780) );
  sky130_fd_sc_hd__nor2_1 U33277 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[1]), 
        .B(n28753), .Y(n28779) );
  sky130_fd_sc_hd__a22oi_1 U33278 ( .A1(n28780), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[8]), .B1(n28779), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[16]), .Y(n28754) );
  sky130_fd_sc_hd__a21oi_1 U33279 ( .A1(n28755), .A2(n28754), .B1(n28776), .Y(
        n28756) );
  sky130_fd_sc_hd__a21o_1 U33280 ( .A1(j202_soc_core_uart_TOP_hold_reg[2]), 
        .A2(n28775), .B1(n28756), .X(j202_soc_core_uart_TOP_N26) );
  sky130_fd_sc_hd__a22oi_1 U33281 ( .A1(n28779), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[17]), .B1(n28778), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[25]), .Y(n28758) );
  sky130_fd_sc_hd__a22oi_1 U33282 ( .A1(n28780), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[9]), .B1(n28777), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[1]), .Y(n28757) );
  sky130_fd_sc_hd__a21oi_1 U33283 ( .A1(n28758), .A2(n28757), .B1(n28776), .Y(
        n28759) );
  sky130_fd_sc_hd__a21o_1 U33284 ( .A1(j202_soc_core_uart_TOP_hold_reg[3]), 
        .A2(n28775), .B1(n28759), .X(j202_soc_core_uart_TOP_N27) );
  sky130_fd_sc_hd__a22oi_1 U33285 ( .A1(n28777), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[2]), .B1(n28778), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[26]), .Y(n28761) );
  sky130_fd_sc_hd__a22oi_1 U33286 ( .A1(n28780), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[10]), .B1(n28779), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[18]), .Y(n28760) );
  sky130_fd_sc_hd__a21oi_1 U33287 ( .A1(n28761), .A2(n28760), .B1(n28776), .Y(
        n28762) );
  sky130_fd_sc_hd__a21o_1 U33288 ( .A1(j202_soc_core_uart_TOP_hold_reg[4]), 
        .A2(n28775), .B1(n28762), .X(j202_soc_core_uart_TOP_N28) );
  sky130_fd_sc_hd__a22oi_1 U33289 ( .A1(n28780), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[11]), .B1(n28778), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[27]), .Y(n28764) );
  sky130_fd_sc_hd__a22oi_1 U33290 ( .A1(n28779), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[19]), .B1(n28777), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[3]), .Y(n28763) );
  sky130_fd_sc_hd__a21oi_1 U33291 ( .A1(n28764), .A2(n28763), .B1(n28776), .Y(
        n28765) );
  sky130_fd_sc_hd__a21o_1 U33292 ( .A1(j202_soc_core_uart_TOP_hold_reg[5]), 
        .A2(n28775), .B1(n28765), .X(j202_soc_core_uart_TOP_N29) );
  sky130_fd_sc_hd__a22oi_1 U33293 ( .A1(n28780), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[12]), .B1(n28779), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[20]), .Y(n28767) );
  sky130_fd_sc_hd__a22oi_1 U33294 ( .A1(n28777), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[4]), .B1(n28778), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[28]), .Y(n28766) );
  sky130_fd_sc_hd__a21oi_1 U33295 ( .A1(n28767), .A2(n28766), .B1(n28776), .Y(
        n28768) );
  sky130_fd_sc_hd__a21o_1 U33296 ( .A1(j202_soc_core_uart_TOP_hold_reg[6]), 
        .A2(n28775), .B1(n28768), .X(j202_soc_core_uart_TOP_N30) );
  sky130_fd_sc_hd__a22oi_1 U33297 ( .A1(n28779), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[21]), .B1(n28778), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[29]), .Y(n28770) );
  sky130_fd_sc_hd__a22oi_1 U33298 ( .A1(n28780), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[13]), .B1(n28777), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[5]), .Y(n28769) );
  sky130_fd_sc_hd__a21oi_1 U33299 ( .A1(n28770), .A2(n28769), .B1(n28776), .Y(
        n28771) );
  sky130_fd_sc_hd__a21o_1 U33300 ( .A1(j202_soc_core_uart_TOP_hold_reg[7]), 
        .A2(n28775), .B1(n28771), .X(j202_soc_core_uart_TOP_N31) );
  sky130_fd_sc_hd__a22oi_1 U33301 ( .A1(n28779), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[22]), .B1(n28778), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[30]), .Y(n28773) );
  sky130_fd_sc_hd__a22oi_1 U33302 ( .A1(n28780), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[14]), .B1(n28777), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[6]), .Y(n28772) );
  sky130_fd_sc_hd__a21oi_1 U33303 ( .A1(n28773), .A2(n28772), .B1(n28776), .Y(
        n28774) );
  sky130_fd_sc_hd__a21o_1 U33304 ( .A1(j202_soc_core_uart_TOP_hold_reg[8]), 
        .A2(n28775), .B1(n28774), .X(j202_soc_core_uart_TOP_N32) );
  sky130_fd_sc_hd__a21oi_1 U33305 ( .A1(n28777), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[7]), .B1(n28776), .Y(n28784) );
  sky130_fd_sc_hd__a22oi_1 U33306 ( .A1(n28779), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[23]), .B1(n28778), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[31]), .Y(n28783) );
  sky130_fd_sc_hd__nand2_1 U33307 ( .A(n28780), .B(
        j202_soc_core_uart_TOP_tx_fifo_mem[15]), .Y(n28782) );
  sky130_fd_sc_hd__a31oi_1 U33308 ( .A1(n28784), .A2(n28783), .A3(n28782), 
        .B1(n28781), .Y(j202_soc_core_uart_TOP_N33) );
  sky130_fd_sc_hd__a22oi_1 U33309 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[2]), .A2(n28874), .B1(
        n28869), .B2(la_data_out[2]), .Y(n28787) );
  sky130_fd_sc_hd__a22oi_1 U33310 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[2]), .A2(n28873), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_ier[2]), .B2(n13289), .Y(
        n28786) );
  sky130_fd_sc_hd__a22oi_1 U33311 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[2]), .A2(n28875), .B1(
        gpio_en_o[2]), .B2(n28876), .Y(n28785) );
  sky130_fd_sc_hd__nand3_1 U33312 ( .A(n28787), .B(n28786), .C(n28785), .Y(
        j202_soc_core_ahb2apb_02_N130) );
  sky130_fd_sc_hd__a22oi_1 U33313 ( .A1(n28876), .A2(gpio_en_o[3]), .B1(n13289), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_ier[3]), .Y(n28790) );
  sky130_fd_sc_hd__a22oi_1 U33314 ( .A1(n28873), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]), .B1(n28869), 
        .B2(la_data_out[3]), .Y(n28789) );
  sky130_fd_sc_hd__a22oi_1 U33315 ( .A1(n28875), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[3]), .B1(n28874), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[3]), .Y(n28788) );
  sky130_fd_sc_hd__nand3_1 U33316 ( .A(n28790), .B(n28789), .C(n28788), .Y(
        j202_soc_core_ahb2apb_02_N131) );
  sky130_fd_sc_hd__a22oi_1 U33317 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[4]), .A2(n28873), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_dtr[4]), .B2(n28874), .Y(
        n28793) );
  sky130_fd_sc_hd__a22oi_1 U33318 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[4]), .A2(n28875), .B1(
        gpio_en_o[4]), .B2(n28876), .Y(n28792) );
  sky130_fd_sc_hd__a22oi_1 U33319 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[4]), .A2(n13289), .B1(
        n28869), .B2(la_data_out[4]), .Y(n28791) );
  sky130_fd_sc_hd__nand3_1 U33320 ( .A(n28793), .B(n28792), .C(n28791), .Y(
        j202_soc_core_ahb2apb_02_N132) );
  sky130_fd_sc_hd__a22oi_1 U33321 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[5]), .A2(n28874), .B1(
        gpio_en_o[5]), .B2(n28876), .Y(n28796) );
  sky130_fd_sc_hd__a22oi_1 U33322 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[5]), .A2(n28875), .B1(
        n28869), .B2(la_data_out[5]), .Y(n28795) );
  sky130_fd_sc_hd__a22oi_1 U33323 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]), .A2(n28873), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_ier[5]), .B2(n13289), .Y(
        n28794) );
  sky130_fd_sc_hd__nand3_1 U33324 ( .A(n28796), .B(n28795), .C(n28794), .Y(
        j202_soc_core_ahb2apb_02_N133) );
  sky130_fd_sc_hd__a22oi_1 U33325 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[6]), .A2(n28874), .B1(
        n28869), .B2(la_data_out[6]), .Y(n28799) );
  sky130_fd_sc_hd__a22oi_1 U33326 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[6]), .A2(n13289), .B1(
        gpio_en_o[6]), .B2(n28876), .Y(n28798) );
  sky130_fd_sc_hd__a22oi_1 U33327 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[6]), .A2(n28875), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]), .B2(n28873), 
        .Y(n28797) );
  sky130_fd_sc_hd__nand3_1 U33328 ( .A(n28799), .B(n28798), .C(n28797), .Y(
        j202_soc_core_ahb2apb_02_N134) );
  sky130_fd_sc_hd__a22oi_1 U33329 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[7]), .A2(n28875), .B1(
        n28869), .B2(la_data_out[7]), .Y(n28802) );
  sky130_fd_sc_hd__a22oi_1 U33330 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[7]), .A2(n28874), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]), .B2(n28873), 
        .Y(n28801) );
  sky130_fd_sc_hd__a22oi_1 U33331 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[7]), .A2(n13289), .B1(
        gpio_en_o[7]), .B2(n28876), .Y(n28800) );
  sky130_fd_sc_hd__nand3_1 U33332 ( .A(n28802), .B(n28801), .C(n28800), .Y(
        j202_soc_core_ahb2apb_02_N135) );
  sky130_fd_sc_hd__a22oi_1 U33333 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]), .A2(n28873), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_ier[8]), .B2(n13289), .Y(
        n28805) );
  sky130_fd_sc_hd__a22oi_1 U33334 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[8]), .A2(n28874), .B1(
        n28869), .B2(la_data_out[8]), .Y(n28804) );
  sky130_fd_sc_hd__a22oi_1 U33335 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[8]), .A2(n28875), .B1(
        gpio_en_o[8]), .B2(n28876), .Y(n28803) );
  sky130_fd_sc_hd__nand3_1 U33336 ( .A(n28805), .B(n28804), .C(n28803), .Y(
        j202_soc_core_ahb2apb_02_N136) );
  sky130_fd_sc_hd__a22oi_1 U33337 ( .A1(n28875), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[9]), .B1(n28869), .B2(
        la_data_out[9]), .Y(n28808) );
  sky130_fd_sc_hd__a22oi_1 U33338 ( .A1(n28873), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[9]), .B1(n28876), 
        .B2(gpio_en_o[9]), .Y(n28807) );
  sky130_fd_sc_hd__a22oi_1 U33339 ( .A1(n28874), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[9]), .B1(n13289), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[9]), .Y(n28806) );
  sky130_fd_sc_hd__nand3_1 U33340 ( .A(n28808), .B(n28807), .C(n28806), .Y(
        j202_soc_core_ahb2apb_02_N137) );
  sky130_fd_sc_hd__a22oi_1 U33341 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[10]), .A2(n28875), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[10]), .B2(n13289), .Y(
        n28811) );
  sky130_fd_sc_hd__a22oi_1 U33342 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[10]), .A2(n28873), 
        .B1(gpio_en_o[10]), .B2(n28876), .Y(n28810) );
  sky130_fd_sc_hd__a22oi_1 U33343 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[10]), .A2(n28874), .B1(
        n28869), .B2(la_data_out[10]), .Y(n28809) );
  sky130_fd_sc_hd__nand3_1 U33344 ( .A(n28811), .B(n28810), .C(n28809), .Y(
        j202_soc_core_ahb2apb_02_N138) );
  sky130_fd_sc_hd__a22oi_1 U33345 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[11]), .A2(n28873), 
        .B1(gpio_en_o[11]), .B2(n28876), .Y(n28814) );
  sky130_fd_sc_hd__a22oi_1 U33346 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[11]), .A2(n28875), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[11]), .B2(n13289), .Y(
        n28813) );
  sky130_fd_sc_hd__a22oi_1 U33347 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[11]), .A2(n28874), .B1(
        n28869), .B2(la_data_out[11]), .Y(n28812) );
  sky130_fd_sc_hd__nand3_1 U33348 ( .A(n28814), .B(n28813), .C(n28812), .Y(
        j202_soc_core_ahb2apb_02_N139) );
  sky130_fd_sc_hd__a22oi_1 U33349 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[12]), .A2(n28873), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_dtr[12]), .B2(n28874), .Y(
        n28817) );
  sky130_fd_sc_hd__a22oi_1 U33350 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[12]), .A2(n13289), .B1(
        n28869), .B2(la_data_out[12]), .Y(n28816) );
  sky130_fd_sc_hd__a22oi_1 U33351 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[12]), .A2(n28875), .B1(
        gpio_en_o[12]), .B2(n28876), .Y(n28815) );
  sky130_fd_sc_hd__nand3_1 U33352 ( .A(n28817), .B(n28816), .C(n28815), .Y(
        j202_soc_core_ahb2apb_02_N140) );
  sky130_fd_sc_hd__a22oi_1 U33353 ( .A1(n28876), .A2(gpio_en_o[13]), .B1(
        n28874), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_dtr[13]), .Y(
        n28820) );
  sky130_fd_sc_hd__a22oi_1 U33354 ( .A1(n28875), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[13]), .B1(n13289), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[13]), .Y(n28819) );
  sky130_fd_sc_hd__a22oi_1 U33355 ( .A1(n28873), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13]), .B1(n28869), 
        .B2(la_data_out[13]), .Y(n28818) );
  sky130_fd_sc_hd__nand3_1 U33356 ( .A(n28820), .B(n28819), .C(n28818), .Y(
        j202_soc_core_ahb2apb_02_N141) );
  sky130_fd_sc_hd__a22oi_1 U33357 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[14]), .A2(n28875), .B1(
        n28869), .B2(la_data_out[14]), .Y(n28823) );
  sky130_fd_sc_hd__a22oi_1 U33358 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[14]), .A2(n13289), .B1(
        gpio_en_o[14]), .B2(n28876), .Y(n28822) );
  sky130_fd_sc_hd__a22oi_1 U33359 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[14]), .A2(n28874), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14]), .B2(n28873), 
        .Y(n28821) );
  sky130_fd_sc_hd__nand3_1 U33360 ( .A(n28823), .B(n28822), .C(n28821), .Y(
        j202_soc_core_ahb2apb_02_N142) );
  sky130_fd_sc_hd__a22oi_1 U33361 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15]), .A2(n28873), 
        .B1(gpio_en_o[15]), .B2(n28876), .Y(n28826) );
  sky130_fd_sc_hd__a22oi_1 U33362 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[15]), .A2(n28875), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[15]), .B2(n28874), .Y(
        n28825) );
  sky130_fd_sc_hd__a22oi_1 U33363 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[15]), .A2(n13289), .B1(
        n28869), .B2(la_data_out[15]), .Y(n28824) );
  sky130_fd_sc_hd__nand3_1 U33364 ( .A(n28826), .B(n28825), .C(n28824), .Y(
        j202_soc_core_ahb2apb_02_N143) );
  sky130_fd_sc_hd__a22oi_1 U33365 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[16]), .A2(n28875), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[16]), .B2(n28874), .Y(
        n28829) );
  sky130_fd_sc_hd__a22oi_1 U33366 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[16]), .A2(n13289), .B1(
        n28869), .B2(la_data_out[16]), .Y(n28828) );
  sky130_fd_sc_hd__a22oi_1 U33367 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16]), .A2(n28873), 
        .B1(gpio_en_o[16]), .B2(n28876), .Y(n28827) );
  sky130_fd_sc_hd__nand3_1 U33368 ( .A(n28829), .B(n28828), .C(n28827), .Y(
        j202_soc_core_ahb2apb_02_N144) );
  sky130_fd_sc_hd__a22oi_1 U33369 ( .A1(n28873), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[17]), .B1(n28875), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_isr[17]), .Y(n28832) );
  sky130_fd_sc_hd__a22oi_1 U33370 ( .A1(n28876), .A2(gpio_en_o[17]), .B1(
        n28869), .B2(la_data_out[17]), .Y(n28831) );
  sky130_fd_sc_hd__a22oi_1 U33371 ( .A1(n28874), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[17]), .B1(n13289), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[17]), .Y(n28830) );
  sky130_fd_sc_hd__nand3_1 U33372 ( .A(n28832), .B(n28831), .C(n28830), .Y(
        j202_soc_core_ahb2apb_02_N145) );
  sky130_fd_sc_hd__a22oi_1 U33373 ( .A1(gpio_en_o[18]), .A2(n28876), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[18]), .B2(n13289), .Y(
        n28835) );
  sky130_fd_sc_hd__a22oi_1 U33374 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[18]), .A2(n28875), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[18]), .B2(n28874), .Y(
        n28834) );
  sky130_fd_sc_hd__a22oi_1 U33375 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[18]), .A2(n28873), 
        .B1(n28869), .B2(la_data_out[18]), .Y(n28833) );
  sky130_fd_sc_hd__nand3_1 U33376 ( .A(n28835), .B(n28834), .C(n28833), .Y(
        j202_soc_core_ahb2apb_02_N146) );
  sky130_fd_sc_hd__a22oi_1 U33377 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[19]), .A2(n28874), .B1(
        gpio_en_o[19]), .B2(n28876), .Y(n28838) );
  sky130_fd_sc_hd__a22oi_1 U33378 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[19]), .A2(n28875), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[19]), .B2(n28873), 
        .Y(n28837) );
  sky130_fd_sc_hd__a22oi_1 U33379 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[19]), .A2(n13289), .B1(
        n28869), .B2(la_data_out[19]), .Y(n28836) );
  sky130_fd_sc_hd__nand3_1 U33380 ( .A(n28838), .B(n28837), .C(n28836), .Y(
        j202_soc_core_ahb2apb_02_N147) );
  sky130_fd_sc_hd__a22oi_1 U33381 ( .A1(gpio_en_o[20]), .A2(n28876), .B1(
        n28869), .B2(la_data_out[20]), .Y(n28841) );
  sky130_fd_sc_hd__a22oi_1 U33382 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[20]), .A2(n28873), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_ier[20]), .B2(n13289), .Y(
        n28840) );
  sky130_fd_sc_hd__a22oi_1 U33383 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[20]), .A2(n28875), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[20]), .B2(n28874), .Y(
        n28839) );
  sky130_fd_sc_hd__nand3_1 U33384 ( .A(n28841), .B(n28840), .C(n28839), .Y(
        j202_soc_core_ahb2apb_02_N148) );
  sky130_fd_sc_hd__a22oi_1 U33385 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[21]), .A2(n13289), .B1(
        gpio_en_o[21]), .B2(n28876), .Y(n28844) );
  sky130_fd_sc_hd__a22oi_1 U33386 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[21]), .A2(n28875), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[21]), .B2(n28873), 
        .Y(n28843) );
  sky130_fd_sc_hd__a22oi_1 U33387 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[21]), .A2(n28874), .B1(
        n28869), .B2(la_data_out[21]), .Y(n28842) );
  sky130_fd_sc_hd__nand3_1 U33388 ( .A(n28844), .B(n28843), .C(n28842), .Y(
        j202_soc_core_ahb2apb_02_N149) );
  sky130_fd_sc_hd__a22oi_1 U33389 ( .A1(gpio_en_o[22]), .A2(n28876), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[22]), .B2(n13289), .Y(
        n28847) );
  sky130_fd_sc_hd__a22oi_1 U33390 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[22]), .A2(n28875), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[22]), .B2(n28874), .Y(
        n28846) );
  sky130_fd_sc_hd__a22oi_1 U33391 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[22]), .A2(n28873), 
        .B1(n28869), .B2(la_data_out[22]), .Y(n28845) );
  sky130_fd_sc_hd__nand3_1 U33392 ( .A(n28847), .B(n28846), .C(n28845), .Y(
        j202_soc_core_ahb2apb_02_N150) );
  sky130_fd_sc_hd__a22oi_1 U33393 ( .A1(n28873), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[23]), .B1(n28875), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_isr[23]), .Y(n28850) );
  sky130_fd_sc_hd__a22oi_1 U33394 ( .A1(n28876), .A2(gpio_en_o[23]), .B1(
        n28874), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_dtr[23]), .Y(
        n28849) );
  sky130_fd_sc_hd__a22oi_1 U33395 ( .A1(n28869), .A2(la_data_out[23]), .B1(
        n13289), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_ier[23]), .Y(
        n28848) );
  sky130_fd_sc_hd__nand3_1 U33396 ( .A(n28850), .B(n28849), .C(n28848), .Y(
        j202_soc_core_ahb2apb_02_N151) );
  sky130_fd_sc_hd__a22oi_1 U33397 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[24]), .A2(n28874), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[24]), .B2(n28873), 
        .Y(n28853) );
  sky130_fd_sc_hd__a22oi_1 U33398 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[24]), .A2(n13289), .B1(
        gpio_en_o[24]), .B2(n28876), .Y(n28852) );
  sky130_fd_sc_hd__a22oi_1 U33399 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[24]), .A2(n28875), .B1(
        n28869), .B2(la_data_out[24]), .Y(n28851) );
  sky130_fd_sc_hd__nand3_1 U33400 ( .A(n28853), .B(n28852), .C(n28851), .Y(
        j202_soc_core_ahb2apb_02_N152) );
  sky130_fd_sc_hd__a22oi_1 U33401 ( .A1(gpio_en_o[25]), .A2(n28876), .B1(
        n28869), .B2(la_data_out[25]), .Y(n28856) );
  sky130_fd_sc_hd__a22oi_1 U33402 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[25]), .A2(n28875), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[25]), .B2(n28874), .Y(
        n28855) );
  sky130_fd_sc_hd__a22oi_1 U33403 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[25]), .A2(n28873), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_ier[25]), .B2(n13289), .Y(
        n28854) );
  sky130_fd_sc_hd__nand3_1 U33404 ( .A(n28856), .B(n28855), .C(n28854), .Y(
        j202_soc_core_ahb2apb_02_N153) );
  sky130_fd_sc_hd__a22oi_1 U33405 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[26]), .A2(n28873), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_dtr[26]), .B2(n28874), .Y(
        n28859) );
  sky130_fd_sc_hd__a22oi_1 U33406 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[26]), .A2(n28875), .B1(
        n28869), .B2(la_data_out[26]), .Y(n28858) );
  sky130_fd_sc_hd__a22oi_1 U33407 ( .A1(gpio_en_o[26]), .A2(n28876), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[26]), .B2(n13289), .Y(
        n28857) );
  sky130_fd_sc_hd__nand3_1 U33408 ( .A(n28859), .B(n28858), .C(n28857), .Y(
        j202_soc_core_ahb2apb_02_N154) );
  sky130_fd_sc_hd__a22oi_1 U33409 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[27]), .A2(n28873), 
        .B1(j202_soc_core_gpio_core_00_gpio_regs_00_ier[27]), .B2(n13289), .Y(
        n28862) );
  sky130_fd_sc_hd__a22oi_1 U33410 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[27]), .A2(n28874), .B1(
        n28869), .B2(la_data_out[27]), .Y(n28861) );
  sky130_fd_sc_hd__a22oi_1 U33411 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[27]), .A2(n28875), .B1(
        gpio_en_o[27]), .B2(n28876), .Y(n28860) );
  sky130_fd_sc_hd__nand3_1 U33412 ( .A(n28862), .B(n28861), .C(n28860), .Y(
        j202_soc_core_ahb2apb_02_N155) );
  sky130_fd_sc_hd__a22oi_1 U33413 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[28]), .A2(n28875), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[28]), .B2(n13289), .Y(
        n28865) );
  sky130_fd_sc_hd__a22oi_1 U33414 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[28]), .A2(n28873), 
        .B1(gpio_en_o[28]), .B2(n28876), .Y(n28864) );
  sky130_fd_sc_hd__a22oi_1 U33415 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[28]), .A2(n28874), .B1(
        n28869), .B2(la_data_out[28]), .Y(n28863) );
  sky130_fd_sc_hd__nand3_1 U33416 ( .A(n28865), .B(n28864), .C(n28863), .Y(
        j202_soc_core_ahb2apb_02_N156) );
  sky130_fd_sc_hd__a22oi_1 U33417 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[29]), .A2(n28874), .B1(
        gpio_en_o[29]), .B2(n28876), .Y(n28868) );
  sky130_fd_sc_hd__a22oi_1 U33418 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[29]), .A2(n13289), .B1(
        n28869), .B2(la_data_out[29]), .Y(n28867) );
  sky130_fd_sc_hd__a22oi_1 U33419 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[29]), .A2(n28875), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[29]), .B2(n28873), 
        .Y(n28866) );
  sky130_fd_sc_hd__nand3_1 U33420 ( .A(n28868), .B(n28867), .C(n28866), .Y(
        j202_soc_core_ahb2apb_02_N157) );
  sky130_fd_sc_hd__a22oi_1 U33421 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[30]), .A2(n28873), 
        .B1(n28869), .B2(la_data_out[30]), .Y(n28872) );
  sky130_fd_sc_hd__a22oi_1 U33422 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[30]), .A2(n28875), .B1(
        gpio_en_o[30]), .B2(n28876), .Y(n28871) );
  sky130_fd_sc_hd__a22oi_1 U33423 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[30]), .A2(n28874), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[30]), .B2(n13289), .Y(
        n28870) );
  sky130_fd_sc_hd__nand3_1 U33424 ( .A(n28872), .B(n28871), .C(n28870), .Y(
        j202_soc_core_ahb2apb_02_N158) );
  sky130_fd_sc_hd__a22oi_1 U33425 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[31]), .A2(n28874), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[31]), .B2(n28873), 
        .Y(n28879) );
  sky130_fd_sc_hd__a22oi_1 U33426 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[31]), .A2(n28875), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[31]), .B2(n13289), .Y(
        n28878) );
  sky130_fd_sc_hd__a22oi_1 U33427 ( .A1(gpio_en_o[31]), .A2(n28876), .B1(
        n28869), .B2(la_data_out[31]), .Y(n28877) );
  sky130_fd_sc_hd__nand3_1 U33428 ( .A(n28879), .B(n28878), .C(n28877), .Y(
        j202_soc_core_ahb2apb_02_N159) );
  sky130_fd_sc_hd__nor3_1 U33429 ( .A(n28882), .B(n28881), .C(n28880), .Y(
        n28887) );
  sky130_fd_sc_hd__nand3_1 U33430 ( .A(n28887), .B(
        j202_soc_core_intc_core_00_bs_addr[3]), .C(
        j202_soc_core_intc_core_00_bs_addr[2]), .Y(n28896) );
  sky130_fd_sc_hd__nor2_1 U33431 ( .A(n28884), .B(n28883), .Y(n28895) );
  sky130_fd_sc_hd__nand3_1 U33432 ( .A(n28895), .B(
        j202_soc_core_intc_core_00_bs_addr[5]), .C(
        j202_soc_core_intc_core_00_bs_addr[4]), .Y(n28889) );
  sky130_fd_sc_hd__nor2_1 U33433 ( .A(n28896), .B(n28889), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_15__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand2_1 U33434 ( .A(n28885), .B(n28887), .Y(n28897) );
  sky130_fd_sc_hd__nor2_1 U33435 ( .A(n28889), .B(n28897), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_14__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand3_1 U33436 ( .A(n28887), .B(
        j202_soc_core_intc_core_00_bs_addr[2]), .C(n28886), .Y(n28898) );
  sky130_fd_sc_hd__nor2_1 U33437 ( .A(n28889), .B(n28898), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_13__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand2_1 U33438 ( .A(n28888), .B(n28887), .Y(n28900) );
  sky130_fd_sc_hd__nor2_1 U33439 ( .A(n28889), .B(n28900), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_12__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand3_1 U33440 ( .A(n28895), .B(
        j202_soc_core_intc_core_00_bs_addr[5]), .C(n28890), .Y(n28891) );
  sky130_fd_sc_hd__nor2_1 U33441 ( .A(n28896), .B(n28891), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_11__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33442 ( .A(n28897), .B(n28891), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_10__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33443 ( .A(n28898), .B(n28891), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_9__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33444 ( .A(n28900), .B(n28891), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_8__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand3_1 U33445 ( .A(n28895), .B(
        j202_soc_core_intc_core_00_bs_addr[4]), .C(n28892), .Y(n28893) );
  sky130_fd_sc_hd__nor2_1 U33446 ( .A(n28896), .B(n28893), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_7__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33447 ( .A(n28897), .B(n28893), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_6__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33448 ( .A(n28898), .B(n28893), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_5__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33449 ( .A(n28900), .B(n28893), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_4__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand2_1 U33450 ( .A(n28895), .B(n28894), .Y(n28899) );
  sky130_fd_sc_hd__nor2_1 U33451 ( .A(n28896), .B(n28899), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_3__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33452 ( .A(n28897), .B(n28899), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_2__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33453 ( .A(n28898), .B(n28899), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_1__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U33454 ( .A(n28900), .B(n28899), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_0__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__or3_1 U33455 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[2]), .C(n28901), .X(io_out[12]) );
  sky130_fd_sc_hd__or3_1 U33456 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[3]), .C(n28901), .X(io_out[13]) );
  sky130_fd_sc_hd__nand2_1 U33457 ( .A(n29092), .B(wbs_dat_i[0]), .Y(n28902)
         );
  sky130_fd_sc_hd__nand2_1 U33458 ( .A(n470), .B(n28902), .Y(n11) );
  sky130_fd_sc_hd__xnor2_1 U33459 ( .A(j202_soc_core_uart_div0[1]), .B(
        j202_soc_core_uart_BRG_ps[1]), .Y(n28904) );
  sky130_fd_sc_hd__xnor2_1 U33460 ( .A(j202_soc_core_uart_div0[5]), .B(
        j202_soc_core_uart_BRG_ps[5]), .Y(n28903) );
  sky130_fd_sc_hd__xor2_1 U33461 ( .A(j202_soc_core_uart_BRG_ps[6]), .B(
        j202_soc_core_uart_div0[6]), .X(n28906) );
  sky130_fd_sc_hd__xor2_1 U33462 ( .A(j202_soc_core_uart_BRG_ps[3]), .B(
        j202_soc_core_uart_div0[3]), .X(n28905) );
  sky130_fd_sc_hd__nor2_1 U33463 ( .A(n28906), .B(n28905), .Y(n28913) );
  sky130_fd_sc_hd__xor2_1 U33464 ( .A(j202_soc_core_uart_BRG_ps[2]), .B(
        j202_soc_core_uart_div0[2]), .X(n28908) );
  sky130_fd_sc_hd__xor2_1 U33465 ( .A(j202_soc_core_uart_BRG_ps[7]), .B(
        j202_soc_core_uart_div0[7]), .X(n28907) );
  sky130_fd_sc_hd__nor2_1 U33466 ( .A(n28908), .B(n28907), .Y(n28912) );
  sky130_fd_sc_hd__xor2_1 U33467 ( .A(j202_soc_core_uart_BRG_ps[4]), .B(
        j202_soc_core_uart_div0[4]), .X(n28910) );
  sky130_fd_sc_hd__xor2_1 U33468 ( .A(j202_soc_core_uart_BRG_ps[0]), .B(
        j202_soc_core_uart_div0[0]), .X(n28909) );
  sky130_fd_sc_hd__nor2_1 U33469 ( .A(n28910), .B(n28909), .Y(n28911) );
  sky130_fd_sc_hd__and4_1 U33470 ( .A(n28914), .B(n28913), .C(n28912), .D(
        n28911), .X(j202_soc_core_uart_BRG_N21) );
  sky130_fd_sc_hd__nand2_2 U20531 ( .A(n12350), .B(
        j202_soc_core_j22_cpu_regop_Rb__1_), .Y(n13702) );
  sky130_fd_sc_hd__o21a_4 U18044 ( .A1(n23822), .A2(n12876), .B1(n27980), .X(
        j202_soc_core_j22_cpu_id_idec_N857) );
  sky130_fd_sc_hd__nand3_2 U19008 ( .A(n12326), .B(n12875), .C(n24256), .Y(
        n12876) );
  sky130_fd_sc_hd__nand3_2 U17584 ( .A(n23145), .B(n23146), .C(n27564), .Y(
        n12485) );
  sky130_fd_sc_hd__nor3_2 U17467 ( .A(n23962), .B(n24420), .C(n23961), .Y(
        n23963) );
  sky130_fd_sc_hd__nand3_1 U18176 ( .A(n12555), .B(n27174), .C(n12557), .Y(
        n12560) );
  sky130_fd_sc_hd__nand2_1 U19232 ( .A(n24423), .B(n13180), .Y(n27174) );
  sky130_fd_sc_hd__clkbuf_1 U13920 ( .A(n27890), .X(n12581) );
  sky130_fd_sc_hd__inv_1 U17720 ( .A(n11901), .Y(n12880) );
  sky130_fd_sc_hd__a21oi_1 U18379 ( .A1(n22944), .A2(n21975), .B1(n21974), .Y(
        n21976) );
  sky130_fd_sc_hd__a21oi_2 U14620 ( .A1(n18824), .A2(n21791), .B1(n18823), .Y(
        n18825) );
  sky130_fd_sc_hd__nand2_2 U13482 ( .A(n26529), .B(n22581), .Y(n11723) );
  sky130_fd_sc_hd__nand3_1 U18200 ( .A(n12732), .B(n27298), .C(n12150), .Y(
        n27550) );
  sky130_fd_sc_hd__inv_1 U15315 ( .A(n12663), .Y(n12661) );
  sky130_fd_sc_hd__nand2_2 U13638 ( .A(n17396), .B(n17688), .Y(n17397) );
  sky130_fd_sc_hd__o21ai_2 U13397 ( .A1(n21499), .A2(n18872), .B1(n18873), .Y(
        n22754) );
  sky130_fd_sc_hd__o21ai_2 U16963 ( .A1(n21495), .A2(n22912), .B1(n21494), .Y(
        n21496) );
  sky130_fd_sc_hd__nand3_2 U28334 ( .A(n12757), .B(n23149), .C(n12735), .Y(
        n23802) );
  sky130_fd_sc_hd__nand2_1 U17594 ( .A(n27551), .B(n11816), .Y(n27686) );
  sky130_fd_sc_hd__nor2_1 U13553 ( .A(n10974), .B(n12501), .Y(n10973) );
  sky130_fd_sc_hd__nor2_2 U19227 ( .A(n23211), .B(n27890), .Y(n23961) );
  sky130_fd_sc_hd__nand2_2 U19219 ( .A(n23602), .B(n24336), .Y(n24420) );
  sky130_fd_sc_hd__nand3_2 U19123 ( .A(n13191), .B(n13192), .C(n13190), .Y(
        n12439) );
  sky130_fd_sc_hd__inv_1 U13722 ( .A(n19473), .Y(n21447) );
  sky130_fd_sc_hd__o22ai_2 U17065 ( .A1(n11514), .A2(n18342), .B1(n18719), 
        .B2(n18374), .Y(n18361) );
  sky130_fd_sc_hd__o21a_2 U13333 ( .A1(n26352), .A2(n11573), .B1(n11571), .X(
        n25711) );
  sky130_fd_sc_hd__inv_4 U13910 ( .A(n12353), .Y(n11521) );
  sky130_fd_sc_hd__nand2_2 U13317 ( .A(n12124), .B(n11790), .Y(n12644) );
  sky130_fd_sc_hd__inv_1 U13981 ( .A(n12983), .Y(n12013) );
  sky130_fd_sc_hd__inv_2 U17645 ( .A(n11846), .Y(n13191) );
  sky130_fd_sc_hd__nand2_2 U13483 ( .A(n26529), .B(n21776), .Y(n21783) );
  sky130_fd_sc_hd__inv_2 U13921 ( .A(n23157), .Y(n22282) );
  sky130_fd_sc_hd__nand2_2 U13861 ( .A(n20974), .B(n12182), .Y(n12460) );
  sky130_fd_sc_hd__inv_2 U17601 ( .A(n11820), .Y(n12646) );
  sky130_fd_sc_hd__nand3_1 U13365 ( .A(n23607), .B(n24266), .C(n13179), .Y(
        n23566) );
  sky130_fd_sc_hd__inv_1 U17873 ( .A(n23162), .Y(n12022) );
  sky130_fd_sc_hd__nand2_1 U17562 ( .A(n23607), .B(n24266), .Y(n27791) );
  sky130_fd_sc_hd__nor2_4 U16823 ( .A(n12692), .B(n29546), .Y(n27898) );
  sky130_fd_sc_hd__inv_1 U16780 ( .A(n19942), .Y(n11313) );
  sky130_fd_sc_hd__inv_1 U16806 ( .A(n12804), .Y(n11326) );
  sky130_fd_sc_hd__inv_1 U17566 ( .A(n13156), .Y(n13155) );
  sky130_fd_sc_hd__inv_2 U13721 ( .A(n12374), .Y(n12371) );
  sky130_fd_sc_hd__nor2_1 U17651 ( .A(n11106), .B(n11874), .Y(n11849) );
  sky130_fd_sc_hd__nand2_1 U13361 ( .A(n11533), .B(n23138), .Y(n24446) );
  sky130_fd_sc_hd__nand2_2 U13370 ( .A(n11132), .B(n29077), .Y(n23602) );
  sky130_fd_sc_hd__o22ai_1 U30930 ( .A1(n27575), .A2(n27464), .B1(n27574), 
        .B2(n27463), .Y(j202_soc_core_j22_cpu_rf_N3097) );
  sky130_fd_sc_hd__nand2_1 U14548 ( .A(n11811), .B(n13052), .Y(n11820) );
  sky130_fd_sc_hd__inv_2 U17520 ( .A(n12353), .Y(n11769) );
  sky130_fd_sc_hd__nand2_2 U13362 ( .A(n12036), .B(n23950), .Y(n27232) );
  sky130_fd_sc_hd__inv_2 U17329 ( .A(n24123), .Y(n22669) );
  sky130_fd_sc_hd__clkinv_1 U17253 ( .A(n13054), .Y(n12558) );
  sky130_fd_sc_hd__nand2_2 U13414 ( .A(n11918), .B(n11917), .Y(n12200) );
  sky130_fd_sc_hd__nor2_1 U20496 ( .A(j202_soc_core_ahb2apb_00_state[1]), .B(
        j202_soc_core_ahb2apb_00_state[0]), .Y(n24815) );
  sky130_fd_sc_hd__bufinv_8 U17256 ( .A(n27928), .Y(n27980) );
  sky130_fd_sc_hd__inv_2 U17602 ( .A(n11821), .Y(n13053) );
  sky130_fd_sc_hd__nand2_2 U13390 ( .A(n12470), .B(n13180), .Y(n12621) );
  sky130_fd_sc_hd__nand2_1 U16869 ( .A(n24350), .B(n29546), .Y(n11903) );
  sky130_fd_sc_hd__nor2_1 U16801 ( .A(n11106), .B(n11325), .Y(n12804) );
  sky130_fd_sc_hd__a22oi_2 U13799 ( .A1(j202_soc_core_memory0_ram_dout0[99]), 
        .A2(n21591), .B1(n21592), .B2(j202_soc_core_memory0_ram_dout0[131]), 
        .Y(n19937) );
  sky130_fd_sc_hd__inv_4 U19344 ( .A(n12621), .Y(n24350) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__1_ ( .D(
        j202_soc_core_j22_cpu_ml_N153), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]) );
  sky130_fd_sc_hd__buf_4 U13648 ( .A(n18112), .X(n18344) );
  sky130_fd_sc_hd__clkbuf_1 U14314 ( .A(n17406), .X(n18469) );
  sky130_fd_sc_hd__buf_2 U14289 ( .A(n18366), .X(n18711) );
  sky130_fd_sc_hd__nand2_1 U20290 ( .A(n25881), .B(n28562), .Y(n10539) );
  sky130_fd_sc_hd__fa_1 U13417 ( .A(n18326), .B(n18325), .CIN(n18324), .COUT(
        n18355), .SUM(n18577) );
  sky130_fd_sc_hd__or2b_1 U20511 ( .A(n13529), .B_N(
        j202_soc_core_j22_cpu_regop_We__3_), .X(n23172) );
  sky130_fd_sc_hd__fa_1 U18011 ( .A(n18755), .B(n18754), .CIN(n18753), .COUT(
        n18768), .SUM(n18758) );
  sky130_fd_sc_hd__fa_1 U13407 ( .A(n17680), .B(n17679), .CIN(n17678), .COUT(
        n17905), .SUM(n17705) );
  sky130_fd_sc_hd__nor2_1 U14171 ( .A(n17890), .B(n17891), .Y(n21889) );
  sky130_fd_sc_hd__nor2_2 U13779 ( .A(n13374), .B(n13496), .Y(n21734) );
  sky130_fd_sc_hd__nor2_1 U17079 ( .A(n18821), .B(n18822), .Y(n21785) );
  sky130_fd_sc_hd__nor2_1 U13994 ( .A(n21785), .B(n19159), .Y(n11515) );
  sky130_fd_sc_hd__nand2_2 U16786 ( .A(n22277), .B(n22278), .Y(n11377) );
  sky130_fd_sc_hd__and2_1 U18840 ( .A(n13163), .B(n20144), .X(n12175) );
  sky130_fd_sc_hd__nand2_2 U17558 ( .A(n20836), .B(n20835), .Y(n29015) );
  sky130_fd_sc_hd__nand2_1 U13495 ( .A(n23731), .B(n22581), .Y(n11395) );
  sky130_fd_sc_hd__inv_2 U16871 ( .A(n11377), .Y(n27556) );
  sky130_fd_sc_hd__nand3_1 U18049 ( .A(n21817), .B(n21816), .C(n21815), .Y(
        n12449) );
  sky130_fd_sc_hd__a2bb2oi_1 U14918 ( .B1(n23940), .B2(n25871), .A1_N(n26423), 
        .A2_N(n27392), .Y(n23836) );
  sky130_fd_sc_hd__nand2b_1 U26839 ( .A_N(n26536), .B(n22581), .Y(n21005) );
  sky130_fd_sc_hd__inv_2 U14497 ( .A(n12692), .Y(n23586) );
  sky130_fd_sc_hd__a2bb2oi_1 U14894 ( .B1(n26085), .B2(n25137), .A1_N(n26423), 
        .A2_N(n25122), .Y(n25124) );
  sky130_fd_sc_hd__nand2_1 U14097 ( .A(n11769), .B(n26548), .Y(n13214) );
  sky130_fd_sc_hd__nand2_1 U17009 ( .A(n11519), .B(n12152), .Y(n27340) );
  sky130_fd_sc_hd__clkbuf_1 U17565 ( .A(n27260), .X(n11798) );
  sky130_fd_sc_hd__nand4_1 U17532 ( .A(n22282), .B(n23154), .C(n23156), .D(
        n23155), .Y(n12438) );
  sky130_fd_sc_hd__a2bb2oi_1 U19376 ( .B1(n23955), .B2(n23954), .A1_N(n23952), 
        .A2_N(n23953), .Y(n27779) );
  sky130_fd_sc_hd__nand2_1 U13372 ( .A(n11769), .B(n11768), .Y(n26550) );
  sky130_fd_sc_hd__nand2_1 U17093 ( .A(n11521), .B(n26524), .Y(n11574) );
  sky130_fd_sc_hd__nor2_2 U14133 ( .A(n23559), .B(n23558), .Y(n26948) );
  sky130_fd_sc_hd__nand3_1 U27657 ( .A(n22228), .B(n26398), .C(n22227), .Y(
        n25545) );
  sky130_fd_sc_hd__nand3_1 U14405 ( .A(n22109), .B(n12310), .C(n12309), .Y(
        n26068) );
  sky130_fd_sc_hd__o21ai_1 U14088 ( .A1(n26443), .A2(n27044), .B1(n12724), .Y(
        n23981) );
  sky130_fd_sc_hd__nand2_1 U14455 ( .A(n24163), .B(n24157), .Y(n11773) );
  sky130_fd_sc_hd__nor2_1 U13881 ( .A(n27897), .B(n27896), .Y(n12393) );
  sky130_fd_sc_hd__inv_2 U16917 ( .A(n11410), .Y(n27467) );
  sky130_fd_sc_hd__nand2_1 U17156 ( .A(n13214), .B(n11574), .Y(n24633) );
  sky130_fd_sc_hd__clkinv_2 U13349 ( .A(n27182), .Y(n27414) );
  sky130_fd_sc_hd__nand2_1 U19235 ( .A(n11127), .B(n29010), .Y(n23815) );
  sky130_fd_sc_hd__nor2_2 U14134 ( .A(n23170), .B(n23169), .Y(n27333) );
  sky130_fd_sc_hd__nor2_2 U14135 ( .A(n23099), .B(n23169), .Y(n27221) );
  sky130_fd_sc_hd__nor2_2 U17472 ( .A(n23105), .B(n23169), .Y(n27213) );
  sky130_fd_sc_hd__nand2_1 U13510 ( .A(n24210), .B(n29012), .Y(n23552) );
  sky130_fd_sc_hd__clkinv_1 U14434 ( .A(n25269), .Y(n11131) );
  sky130_fd_sc_hd__nor2_2 U17525 ( .A(n23090), .B(n23169), .Y(n27466) );
  sky130_fd_sc_hd__nand3_1 U13325 ( .A(n11694), .B(n11051), .C(n11697), .Y(
        n11586) );
  sky130_fd_sc_hd__o21ai_1 U18835 ( .A1(n23563), .A2(n23562), .B1(n11127), .Y(
        n12168) );
  sky130_fd_sc_hd__inv_1 U13328 ( .A(n23815), .Y(n12534) );
  sky130_fd_sc_hd__clkbuf_1 U17524 ( .A(n27044), .X(n11764) );
  sky130_fd_sc_hd__nand2_2 U13913 ( .A(n25156), .B(n25152), .Y(n25158) );
  sky130_fd_sc_hd__nand2_2 U18273 ( .A(n13072), .B(n13240), .Y(n27300) );
  sky130_fd_sc_hd__buf_8 U19177 ( .A(n23812), .X(n12479) );
  sky130_fd_sc_hd__nor2_1 U17334 ( .A(n24118), .B(n25107), .Y(n12458) );
  sky130_fd_sc_hd__inv_2 U18278 ( .A(n24213), .Y(n24214) );
  sky130_fd_sc_hd__buf_2 U14052 ( .A(n25661), .X(n12474) );
  sky130_fd_sc_hd__and2_0 U13905 ( .A(n28985), .B(n11129), .X(n11083) );
  sky130_fd_sc_hd__inv_2 U19163 ( .A(n25705), .Y(n25707) );
  sky130_fd_sc_hd__o22ai_1 U31570 ( .A1(n27575), .A2(n27370), .B1(n27574), 
        .B2(n26469), .Y(j202_soc_core_j22_cpu_rf_N3117) );
  sky130_fd_sc_hd__nand2_2 U13284 ( .A(n12464), .B(n29595), .Y(
        j202_soc_core_ahb2apb_00_N22) );
  sky130_fd_sc_hd__inv_2 U19985 ( .A(n23173), .Y(n23168) );
  sky130_fd_sc_hd__nand3_2 U13502 ( .A(n11948), .B(n12214), .C(n11064), .Y(
        n26710) );
  sky130_fd_sc_hd__fa_2 U13408 ( .A(n18725), .B(n18724), .CIN(n18723), .COUT(
        n18756), .SUM(n18746) );
  sky130_fd_sc_hd__nor2_2 U17304 ( .A(j202_soc_core_memory0_ram_dout0_sel[14]), 
        .B(n13498), .Y(n21598) );
  sky130_fd_sc_hd__nor2_1 U13406 ( .A(n14128), .B(n14127), .Y(n21526) );
  sky130_fd_sc_hd__nand2_1 U13461 ( .A(n21007), .B(n21006), .Y(n26524) );
  sky130_fd_sc_hd__nand2_1 U16796 ( .A(n20988), .B(n11706), .Y(n11323) );
  sky130_fd_sc_hd__clkbuf_1 U25640 ( .A(n19223), .X(n19483) );
  sky130_fd_sc_hd__clkbuf_1 U19225 ( .A(n12415), .X(n12727) );
  sky130_fd_sc_hd__nand2_1 U13393 ( .A(n11135), .B(n22581), .Y(n11394) );
  sky130_fd_sc_hd__nand2_2 U13467 ( .A(n12732), .B(n23139), .Y(n27877) );
  sky130_fd_sc_hd__nand2_1 U17630 ( .A(n11072), .B(n12395), .Y(n13072) );
  sky130_fd_sc_hd__buf_2 U13898 ( .A(n23561), .X(n11126) );
  sky130_fd_sc_hd__inv_4 U19073 ( .A(n12644), .Y(n12383) );
  sky130_fd_sc_hd__nand2_1 U13289 ( .A(n25557), .B(n25559), .Y(n24733) );
  sky130_fd_sc_hd__nand2_1 U13302 ( .A(n11769), .B(n12643), .Y(n27044) );
  sky130_fd_sc_hd__nand3_1 U13303 ( .A(n11933), .B(n11067), .C(n11079), .Y(
        n11932) );
  sky130_fd_sc_hd__clkbuf_1 U13305 ( .A(n17139), .X(n10934) );
  sky130_fd_sc_hd__inv_2 U13309 ( .A(n11970), .Y(n11974) );
  sky130_fd_sc_hd__nand2_2 U13321 ( .A(n11723), .B(n29504), .Y(n28918) );
  sky130_fd_sc_hd__nand3_1 U13323 ( .A(n19251), .B(n22581), .C(n19250), .Y(
        n16664) );
  sky130_fd_sc_hd__inv_4 U13326 ( .A(n24733), .Y(n25639) );
  sky130_fd_sc_hd__clkinv_2 U13327 ( .A(n12167), .Y(n27063) );
  sky130_fd_sc_hd__inv_8 U13334 ( .A(n29507), .Y(n29249) );
  sky130_fd_sc_hd__and2_1 U13342 ( .A(n28993), .B(n11127), .X(n12193) );
  sky130_fd_sc_hd__inv_8 U13345 ( .A(n11126), .Y(n12538) );
  sky130_fd_sc_hd__nand2_2 U13346 ( .A(n12627), .B(n29492), .Y(n12042) );
  sky130_fd_sc_hd__clkbuf_1 U13351 ( .A(n27182), .X(n29549) );
  sky130_fd_sc_hd__nor2_4 U13353 ( .A(n12416), .B(n29508), .Y(n29507) );
  sky130_fd_sc_hd__nand2_1 U13355 ( .A(n11797), .B(n27898), .Y(n24266) );
  sky130_fd_sc_hd__and2_1 U13356 ( .A(n17130), .B(n17129), .X(n11933) );
  sky130_fd_sc_hd__nor2_1 U13360 ( .A(n11899), .B(n29560), .Y(n11898) );
  sky130_fd_sc_hd__buf_2 U13366 ( .A(n11377), .X(n29546) );
  sky130_fd_sc_hd__nand2_1 U13388 ( .A(n13008), .B(n12250), .Y(n11324) );
  sky130_fd_sc_hd__nor3_1 U13392 ( .A(n14962), .B(n15816), .C(n15819), .Y(
        n17077) );
  sky130_fd_sc_hd__o21ai_0 U13395 ( .A1(n22177), .A2(n22795), .B1(n22178), .Y(
        n22081) );
  sky130_fd_sc_hd__o21ai_0 U13404 ( .A1(n18388), .A2(n18389), .B1(n18387), .Y(
        n11599) );
  sky130_fd_sc_hd__o21ai_0 U13451 ( .A1(n16076), .A2(n16075), .B1(n17273), .Y(
        n16084) );
  sky130_fd_sc_hd__clkinv_1 U13452 ( .A(n18432), .Y(n29555) );
  sky130_fd_sc_hd__o21ai_0 U13454 ( .A1(n15423), .A2(n15846), .B1(n16058), .Y(
        n14906) );
  sky130_fd_sc_hd__o21ai_0 U13458 ( .A1(n17550), .A2(n17551), .B1(n17549), .Y(
        n11637) );
  sky130_fd_sc_hd__o21ai_0 U13459 ( .A1(n18394), .A2(n18395), .B1(n18393), .Y(
        n11741) );
  sky130_fd_sc_hd__o21ai_0 U13462 ( .A1(n22085), .A2(n22183), .B1(n22084), .Y(
        n22161) );
  sky130_fd_sc_hd__clkinv_1 U13464 ( .A(n17453), .Y(n12584) );
  sky130_fd_sc_hd__o21ai_0 U13466 ( .A1(n18491), .A2(n18492), .B1(n18490), .Y(
        n18494) );
  sky130_fd_sc_hd__o21ai_0 U13468 ( .A1(n18434), .A2(n18435), .B1(n18433), .Y(
        n12703) );
  sky130_fd_sc_hd__o21ai_0 U13470 ( .A1(n18432), .A2(n29556), .B1(n18430), .Y(
        n29553) );
  sky130_fd_sc_hd__o21ai_0 U13471 ( .A1(n17059), .A2(n13436), .B1(n15324), .Y(
        n15561) );
  sky130_fd_sc_hd__clkinv_1 U13472 ( .A(n14936), .Y(n14874) );
  sky130_fd_sc_hd__o21ai_0 U13474 ( .A1(n15673), .A2(n15703), .B1(n15672), .Y(
        n15732) );
  sky130_fd_sc_hd__or2_0 U13475 ( .A(n18043), .B(n18042), .X(n18117) );
  sky130_fd_sc_hd__o21ai_0 U13476 ( .A1(n18166), .A2(n18170), .B1(n18167), .Y(
        n18165) );
  sky130_fd_sc_hd__clkinv_1 U13477 ( .A(n18401), .Y(n11743) );
  sky130_fd_sc_hd__o21ai_0 U13479 ( .A1(n17486), .A2(n17485), .B1(n17484), .Y(
        n11375) );
  sky130_fd_sc_hd__o21ai_0 U13481 ( .A1(n18476), .A2(n18475), .B1(n18474), .Y(
        n12923) );
  sky130_fd_sc_hd__o21ai_0 U13484 ( .A1(n16755), .A2(n16878), .B1(n16945), .Y(
        n16756) );
  sky130_fd_sc_hd__o21ai_0 U13485 ( .A1(n13423), .A2(n13422), .B1(n15584), .Y(
        n13424) );
  sky130_fd_sc_hd__clkinv_1 U13503 ( .A(n20603), .Y(n20674) );
  sky130_fd_sc_hd__o21ai_0 U13504 ( .A1(n15846), .A2(n15845), .B1(n15844), .Y(
        n15848) );
  sky130_fd_sc_hd__clkinv_1 U13505 ( .A(n14928), .Y(n15871) );
  sky130_fd_sc_hd__o21ai_0 U13506 ( .A1(n14937), .A2(n14936), .B1(n14942), .Y(
        n14938) );
  sky130_fd_sc_hd__o21ai_0 U13507 ( .A1(n14907), .A2(n17034), .B1(n13388), .Y(
        n14908) );
  sky130_fd_sc_hd__o21ai_0 U13513 ( .A1(n19873), .A2(n17164), .B1(n20920), .Y(
        n20355) );
  sky130_fd_sc_hd__o21ai_0 U13521 ( .A1(n16611), .A2(n16913), .B1(n16585), .Y(
        n16586) );
  sky130_fd_sc_hd__clkinv_1 U13526 ( .A(n17059), .Y(n15308) );
  sky130_fd_sc_hd__o21ai_0 U13530 ( .A1(n17615), .A2(n12756), .B1(n17614), .Y(
        n12754) );
  sky130_fd_sc_hd__o21ai_0 U13533 ( .A1(n19468), .A2(n18844), .B1(n18843), .Y(
        n18845) );
  sky130_fd_sc_hd__o21ai_0 U13535 ( .A1(n18246), .A2(n18247), .B1(n18245), .Y(
        n13203) );
  sky130_fd_sc_hd__o21ai_0 U13536 ( .A1(n18026), .A2(n18027), .B1(n18025), .Y(
        n18029) );
  sky130_fd_sc_hd__o21ai_0 U13541 ( .A1(n18677), .A2(n11428), .B1(n18676), .Y(
        n11426) );
  sky130_fd_sc_hd__o21ai_0 U13558 ( .A1(n18801), .A2(n18802), .B1(n18800), .Y(
        n12778) );
  sky130_fd_sc_hd__o21ai_0 U13565 ( .A1(n17523), .A2(n17522), .B1(n17521), .Y(
        n12571) );
  sky130_fd_sc_hd__clkinv_1 U13588 ( .A(n26419), .Y(n24483) );
  sky130_fd_sc_hd__o21ai_0 U13590 ( .A1(n18604), .A2(n18603), .B1(n12057), .Y(
        n12054) );
  sky130_fd_sc_hd__o21ai_0 U13595 ( .A1(n16215), .A2(n16214), .B1(n16945), .Y(
        n16224) );
  sky130_fd_sc_hd__o21ai_0 U13596 ( .A1(n15597), .A2(n15596), .B1(n15630), .Y(
        n15598) );
  sky130_fd_sc_hd__o21ai_0 U13597 ( .A1(n20790), .A2(n20789), .B1(n21631), .Y(
        n21717) );
  sky130_fd_sc_hd__clkinv_1 U13625 ( .A(n21614), .Y(n21046) );
  sky130_fd_sc_hd__clkinv_1 U13626 ( .A(n20473), .Y(n20491) );
  sky130_fd_sc_hd__and2_0 U13643 ( .A(n20632), .B(n16171), .X(n15716) );
  sky130_fd_sc_hd__o21ai_0 U13651 ( .A1(n17011), .A2(n17046), .B1(n17273), .Y(
        n17019) );
  sky130_fd_sc_hd__o21ai_0 U13652 ( .A1(n17009), .A2(n17008), .B1(n13387), .Y(
        n17020) );
  sky130_fd_sc_hd__o21ai_0 U13663 ( .A1(n15352), .A2(n15351), .B1(n16090), .Y(
        n15353) );
  sky130_fd_sc_hd__o21ai_0 U13666 ( .A1(n15330), .A2(n15547), .B1(n15584), .Y(
        n15336) );
  sky130_fd_sc_hd__and2_0 U13675 ( .A(n20350), .B(n20325), .X(n13279) );
  sky130_fd_sc_hd__inv_2 U13678 ( .A(n21117), .Y(n18961) );
  sky130_fd_sc_hd__o21ai_0 U13680 ( .A1(j202_soc_core_intc_core_00_rg_ipr[65]), 
        .A2(n26900), .B1(j202_soc_core_intc_core_00_rg_ipr[64]), .Y(n19505) );
  sky130_fd_sc_hd__o21ai_0 U13683 ( .A1(n16595), .A2(n16594), .B1(n16919), .Y(
        n16603) );
  sky130_fd_sc_hd__o21ai_0 U13685 ( .A1(n16878), .A2(n16877), .B1(n16919), .Y(
        n16899) );
  sky130_fd_sc_hd__and2_0 U13687 ( .A(n24350), .B(n12595), .X(n13317) );
  sky130_fd_sc_hd__clkinv_1 U13689 ( .A(n18719), .Y(n11162) );
  sky130_fd_sc_hd__clkinv_1 U13693 ( .A(n11419), .Y(n18595) );
  sky130_fd_sc_hd__o21ai_0 U13694 ( .A1(n18594), .A2(n18595), .B1(n18593), .Y(
        n13205) );
  sky130_fd_sc_hd__o21ai_0 U13698 ( .A1(n25302), .A2(n25301), .B1(n26329), .Y(
        n25303) );
  sky130_fd_sc_hd__o21ai_0 U13703 ( .A1(n19470), .A2(n19469), .B1(n19468), .Y(
        n19471) );
  sky130_fd_sc_hd__o21ai_0 U13713 ( .A1(n17735), .A2(n17734), .B1(n17733), .Y(
        n11622) );
  sky130_fd_sc_hd__o21ai_0 U13718 ( .A1(n18790), .A2(n18791), .B1(n18789), .Y(
        n18793) );
  sky130_fd_sc_hd__o21ai_0 U13724 ( .A1(n23920), .A2(n23919), .B1(n23918), .Y(
        n23921) );
  sky130_fd_sc_hd__a21boi_0 U13727 ( .A1(n22102), .A2(n11476), .B1_N(n11474), 
        .Y(n22618) );
  sky130_fd_sc_hd__o21ai_0 U13728 ( .A1(n18400), .A2(n18401), .B1(n18399), .Y(
        n11745) );
  sky130_fd_sc_hd__o21ai_0 U13731 ( .A1(n18088), .A2(n18089), .B1(n18087), .Y(
        n13002) );
  sky130_fd_sc_hd__o21ai_0 U13732 ( .A1(n18545), .A2(n18546), .B1(n18544), .Y(
        n18548) );
  sky130_fd_sc_hd__o21ai_0 U13733 ( .A1(n18550), .A2(n18551), .B1(n18549), .Y(
        n12920) );
  sky130_fd_sc_hd__o21ai_0 U13737 ( .A1(n15572), .A2(n15571), .B1(n16090), .Y(
        n15573) );
  sky130_fd_sc_hd__o21ai_0 U13742 ( .A1(n21695), .A2(n21705), .B1(n21694), .Y(
        n21696) );
  sky130_fd_sc_hd__o21ai_0 U13745 ( .A1(n20866), .A2(n20865), .B1(n20864), .Y(
        n20867) );
  sky130_fd_sc_hd__o21ai_0 U13746 ( .A1(n18438), .A2(n18439), .B1(n18437), .Y(
        n18441) );
  sky130_fd_sc_hd__clkinv_1 U13752 ( .A(n20736), .Y(n21643) );
  sky130_fd_sc_hd__o21ai_0 U13753 ( .A1(n21189), .A2(n21188), .B1(n21235), .Y(
        n21195) );
  sky130_fd_sc_hd__o21ai_0 U13771 ( .A1(n16694), .A2(n16906), .B1(n16945), .Y(
        n16695) );
  sky130_fd_sc_hd__o21ai_0 U13776 ( .A1(n20787), .A2(n17057), .B1(n11670), .Y(
        n17058) );
  sky130_fd_sc_hd__o21ai_0 U13781 ( .A1(n17055), .A2(n14959), .B1(n14958), .Y(
        n14964) );
  sky130_fd_sc_hd__clkinv_1 U13792 ( .A(n21256), .Y(n21226) );
  sky130_fd_sc_hd__o21ai_0 U13798 ( .A1(n20810), .A2(n19259), .B1(n21251), .Y(
        n19262) );
  sky130_fd_sc_hd__clkinv_1 U13800 ( .A(n20202), .Y(n19848) );
  sky130_fd_sc_hd__o21ai_0 U13810 ( .A1(n15556), .A2(n15243), .B1(n15584), .Y(
        n15244) );
  sky130_fd_sc_hd__o21ai_0 U13816 ( .A1(n15224), .A2(n15547), .B1(n15584), .Y(
        n15233) );
  sky130_fd_sc_hd__o21ai_0 U13826 ( .A1(n18265), .A2(n18267), .B1(n18264), .Y(
        n18260) );
  sky130_fd_sc_hd__clkinv_1 U13827 ( .A(n22680), .Y(n22400) );
  sky130_fd_sc_hd__o21ai_0 U13829 ( .A1(n17760), .A2(n17759), .B1(n17758), .Y(
        n11501) );
  sky130_fd_sc_hd__o21ai_0 U13830 ( .A1(n22361), .A2(n22360), .B1(n22359), .Y(
        n22362) );
  sky130_fd_sc_hd__or2_0 U13831 ( .A(n26791), .B(n19026), .X(n26333) );
  sky130_fd_sc_hd__and2_0 U13833 ( .A(n17781), .B(n11499), .X(n11041) );
  sky130_fd_sc_hd__o21ai_0 U13834 ( .A1(n22893), .A2(n22892), .B1(n22891), .Y(
        n22894) );
  sky130_fd_sc_hd__clkinv_1 U13835 ( .A(n26424), .Y(n25063) );
  sky130_fd_sc_hd__o21ai_0 U13839 ( .A1(n22620), .A2(n22619), .B1(n22618), .Y(
        n22621) );
  sky130_fd_sc_hd__o21ai_0 U13840 ( .A1(n22937), .A2(n22941), .B1(n22938), .Y(
        n22166) );
  sky130_fd_sc_hd__clkinv_1 U13846 ( .A(n22360), .Y(n22132) );
  sky130_fd_sc_hd__o21ai_0 U13848 ( .A1(n26705), .A2(n26432), .B1(n26431), .Y(
        n26433) );
  sky130_fd_sc_hd__clkinv_1 U13849 ( .A(n13612), .Y(n13611) );
  sky130_fd_sc_hd__o21ai_0 U13856 ( .A1(n16551), .A2(n17109), .B1(n16550), .Y(
        n16552) );
  sky130_fd_sc_hd__o21ai_0 U13865 ( .A1(n21794), .A2(n21793), .B1(n21792), .Y(
        n21795) );
  sky130_fd_sc_hd__o21ai_0 U13867 ( .A1(n19368), .A2(n19367), .B1(n20908), .Y(
        n19375) );
  sky130_fd_sc_hd__clkinv_1 U13876 ( .A(n21649), .Y(n19257) );
  sky130_fd_sc_hd__o21ai_0 U13883 ( .A1(n15540), .A2(n15539), .B1(n15630), .Y(
        n15541) );
  sky130_fd_sc_hd__o21ai_0 U13885 ( .A1(n15536), .A2(n15544), .B1(n16090), .Y(
        n15542) );
  sky130_fd_sc_hd__clkinv_1 U13886 ( .A(n14742), .Y(n11146) );
  sky130_fd_sc_hd__o21ai_0 U13891 ( .A1(n13478), .A2(n13477), .B1(n15630), .Y(
        n13482) );
  sky130_fd_sc_hd__clkinv_1 U13892 ( .A(n16988), .Y(n16810) );
  sky130_fd_sc_hd__o21ai_0 U13893 ( .A1(n17278), .A2(n15878), .B1(n15877), .Y(
        n15884) );
  sky130_fd_sc_hd__o21ai_0 U13894 ( .A1(n18938), .A2(n21044), .B1(n21636), .Y(
        n18939) );
  sky130_fd_sc_hd__nand2_1 U13895 ( .A(n19388), .B(n20788), .Y(n21256) );
  sky130_fd_sc_hd__o21ai_0 U13900 ( .A1(n21200), .A2(n19285), .B1(n21235), .Y(
        n19289) );
  sky130_fd_sc_hd__clkinv_1 U13907 ( .A(n20872), .Y(n20073) );
  sky130_fd_sc_hd__clkinv_1 U13908 ( .A(n19971), .Y(n20046) );
  sky130_fd_sc_hd__o21ai_0 U13909 ( .A1(n19126), .A2(n19998), .B1(n20912), .Y(
        n19127) );
  sky130_fd_sc_hd__clkinv_1 U13916 ( .A(n18925), .Y(n21710) );
  sky130_fd_sc_hd__clkinv_1 U13922 ( .A(n21628), .Y(n21126) );
  sky130_fd_sc_hd__clkinv_1 U13923 ( .A(n20904), .Y(n19135) );
  sky130_fd_sc_hd__o21ai_0 U13924 ( .A1(n19876), .A2(n20323), .B1(n20892), .Y(
        n17196) );
  sky130_fd_sc_hd__clkinv_1 U13925 ( .A(n19994), .Y(n19905) );
  sky130_fd_sc_hd__clkinv_1 U13927 ( .A(n20298), .Y(n20313) );
  sky130_fd_sc_hd__clkinv_1 U13928 ( .A(n19767), .Y(n19757) );
  sky130_fd_sc_hd__o21ai_0 U13930 ( .A1(n27380), .A2(n22592), .B1(n16031), .Y(
        n16032) );
  sky130_fd_sc_hd__and2_0 U13937 ( .A(n13268), .B(n13271), .X(n12286) );
  sky130_fd_sc_hd__o21ai_0 U13941 ( .A1(n18806), .A2(n11605), .B1(n18805), .Y(
        n11603) );
  sky130_fd_sc_hd__o21ai_0 U13943 ( .A1(n21345), .A2(n21332), .B1(n21333), .Y(
        n14566) );
  sky130_fd_sc_hd__and2_0 U13956 ( .A(n12926), .B(n22681), .X(n11053) );
  sky130_fd_sc_hd__o21ai_0 U13960 ( .A1(n26352), .A2(n26726), .B1(n26351), .Y(
        n24157) );
  sky130_fd_sc_hd__o21ai_0 U13972 ( .A1(n23919), .A2(n26714), .B1(n23047), .Y(
        n23048) );
  sky130_fd_sc_hd__o21ai_0 U13997 ( .A1(n16536), .A2(n16535), .B1(n16534), .Y(
        n16537) );
  sky130_fd_sc_hd__o21ai_0 U14031 ( .A1(n14742), .A2(n25122), .B1(n15950), .Y(
        n15955) );
  sky130_fd_sc_hd__o21ai_0 U14034 ( .A1(n15664), .A2(n15418), .B1(n15419), .Y(
        n15199) );
  sky130_fd_sc_hd__clkinv_1 U14046 ( .A(n27964), .Y(n24445) );
  sky130_fd_sc_hd__o21ai_0 U14051 ( .A1(n18916), .A2(n22312), .B1(n19193), .Y(
        n19194) );
  sky130_fd_sc_hd__o21ai_0 U14054 ( .A1(n22794), .A2(n22798), .B1(n22795), .Y(
        n22190) );
  sky130_fd_sc_hd__clkinv_1 U14056 ( .A(n14466), .Y(n14393) );
  sky130_fd_sc_hd__clkinv_1 U14061 ( .A(n21785), .Y(n21787) );
  sky130_fd_sc_hd__o21ai_0 U14062 ( .A1(n21071), .A2(n19376), .B1(n13275), .Y(
        n19377) );
  sky130_fd_sc_hd__clkinv_1 U14068 ( .A(n19352), .Y(n17284) );
  sky130_fd_sc_hd__o21ai_0 U14099 ( .A1(j202_soc_core_intc_core_00_rg_ipr[74]), 
        .A2(n26850), .B1(n19520), .Y(n19536) );
  sky130_fd_sc_hd__and2_0 U14101 ( .A(n18981), .B(n22714), .X(n11710) );
  sky130_fd_sc_hd__clkinv_1 U14111 ( .A(n21418), .Y(n11139) );
  sky130_fd_sc_hd__o21ai_0 U14116 ( .A1(j202_soc_core_j22_cpu_exuop_EXU_[5]), 
        .A2(n26745), .B1(n26744), .Y(n26752) );
  sky130_fd_sc_hd__o21ai_0 U14142 ( .A1(n21290), .A2(n21289), .B1(n21288), .Y(
        n21291) );
  sky130_fd_sc_hd__o21ai_0 U14144 ( .A1(n15773), .A2(n15194), .B1(n15193), .Y(
        n15414) );
  sky130_fd_sc_hd__o21ai_0 U14180 ( .A1(j202_soc_core_qspi_wb_addr[2]), .A2(
        n26029), .B1(n28225), .Y(n23460) );
  sky130_fd_sc_hd__clkinv_1 U14181 ( .A(n26716), .Y(n26578) );
  sky130_fd_sc_hd__clkinv_1 U14277 ( .A(n19926), .Y(n29538) );
  sky130_fd_sc_hd__clkinv_1 U14288 ( .A(n20925), .Y(n20335) );
  sky130_fd_sc_hd__o21ai_0 U14315 ( .A1(n18940), .A2(n21720), .B1(n18939), .Y(
        n18941) );
  sky130_fd_sc_hd__o21ai_0 U14332 ( .A1(n20122), .A2(n20121), .B1(n20892), .Y(
        n20123) );
  sky130_fd_sc_hd__clkinv_1 U14343 ( .A(n20326), .Y(n20916) );
  sky130_fd_sc_hd__o21ai_0 U14344 ( .A1(n20873), .A2(n17210), .B1(n17209), .Y(
        n17214) );
  sky130_fd_sc_hd__o21ai_0 U14355 ( .A1(j202_soc_core_j22_cpu_rfuo_sr__i__1_), 
        .A2(n16041), .B1(n16040), .Y(n16044) );
  sky130_fd_sc_hd__o21ai_0 U14362 ( .A1(n19887), .A2(n19886), .B1(n20864), .Y(
        n19888) );
  sky130_fd_sc_hd__o21ai_0 U14366 ( .A1(n12505), .A2(n13547), .B1(
        j202_soc_core_j22_cpu_regop_Rs__0_), .Y(n13548) );
  sky130_fd_sc_hd__o21ai_0 U14371 ( .A1(n21015), .A2(n15512), .B1(n15513), .Y(
        n14834) );
  sky130_fd_sc_hd__clkinv_1 U14374 ( .A(n11874), .Y(n11866) );
  sky130_fd_sc_hd__inv_2 U14375 ( .A(n23241), .Y(n12349) );
  sky130_fd_sc_hd__o2bb2ai_1 U14381 ( .B1(j202_soc_core_j22_cpu_regop_Rs__1_), 
        .B2(n13530), .A1_N(n16513), .A2_N(n12350), .Y(n13553) );
  sky130_fd_sc_hd__clkinv_1 U14386 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[3]), 
        .Y(n26744) );
  sky130_fd_sc_hd__and2_0 U14403 ( .A(n27602), .B(n17137), .X(n12279) );
  sky130_fd_sc_hd__o21ai_0 U14411 ( .A1(n14742), .A2(n27372), .B1(n14307), .Y(
        n14561) );
  sky130_fd_sc_hd__o21ai_0 U14418 ( .A1(n19486), .A2(n22837), .B1(n19485), .Y(
        n19487) );
  sky130_fd_sc_hd__o21ai_0 U14425 ( .A1(n22402), .A2(n22897), .B1(n22401), .Y(
        n22403) );
  sky130_fd_sc_hd__clkinv_1 U14437 ( .A(n22828), .Y(n22830) );
  sky130_fd_sc_hd__o21ai_0 U14439 ( .A1(n21982), .A2(n22837), .B1(n21981), .Y(
        n21983) );
  sky130_fd_sc_hd__clkinv_1 U14440 ( .A(n21428), .Y(n11142) );
  sky130_fd_sc_hd__o21ai_0 U14441 ( .A1(n14742), .A2(n27383), .B1(n14516), .Y(
        n14555) );
  sky130_fd_sc_hd__o21ai_0 U14461 ( .A1(n26352), .A2(n26722), .B1(n26351), .Y(
        n25043) );
  sky130_fd_sc_hd__o21ai_0 U14472 ( .A1(n14742), .A2(n27405), .B1(n15163), .Y(
        n15198) );
  sky130_fd_sc_hd__o21ai_0 U14480 ( .A1(n22802), .A2(n22897), .B1(n22801), .Y(
        n22803) );
  sky130_fd_sc_hd__clkinv_1 U14484 ( .A(n23249), .Y(n23224) );
  sky130_fd_sc_hd__clkinv_1 U14502 ( .A(n11669), .Y(n23789) );
  sky130_fd_sc_hd__and2_0 U14505 ( .A(n13159), .B(n27772), .X(n11076) );
  sky130_fd_sc_hd__o21ai_0 U14527 ( .A1(n24772), .A2(n23926), .B1(n23925), .Y(
        n23938) );
  sky130_fd_sc_hd__o21ai_0 U14532 ( .A1(n26352), .A2(n26600), .B1(n26351), .Y(
        n21550) );
  sky130_fd_sc_hd__and2_0 U14556 ( .A(n13159), .B(n24336), .X(n11077) );
  sky130_fd_sc_hd__o21ai_0 U14590 ( .A1(n21805), .A2(n21804), .B1(n21803), .Y(
        n21806) );
  sky130_fd_sc_hd__o21ai_0 U14598 ( .A1(n27313), .A2(n26846), .B1(n19530), .Y(
        n19540) );
  sky130_fd_sc_hd__o21ai_0 U14626 ( .A1(n18916), .A2(n24492), .B1(n24491), .Y(
        n24493) );
  sky130_fd_sc_hd__o21ai_0 U14640 ( .A1(n26413), .A2(n26412), .B1(n26411), .Y(
        n26438) );
  sky130_fd_sc_hd__o21ai_0 U14654 ( .A1(n18916), .A2(n22305), .B1(n21944), .Y(
        n21945) );
  sky130_fd_sc_hd__clkinv_1 U14658 ( .A(n12556), .Y(n12437) );
  sky130_fd_sc_hd__clkinv_1 U14687 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .Y(n13398) );
  sky130_fd_sc_hd__clkinv_1 U14694 ( .A(n21756), .Y(n21758) );
  sky130_fd_sc_hd__o21ai_0 U14717 ( .A1(n14742), .A2(n24613), .B1(n14797), .Y(
        n14831) );
  sky130_fd_sc_hd__clkinv_1 U14772 ( .A(n13635), .Y(n13641) );
  sky130_fd_sc_hd__o21ai_0 U14786 ( .A1(n20925), .A2(n20895), .B1(n20894), .Y(
        n20910) );
  sky130_fd_sc_hd__o21ai_0 U14797 ( .A1(n23012), .A2(n26604), .B1(n23011), .Y(
        n21384) );
  sky130_fd_sc_hd__o21ai_0 U14864 ( .A1(n14742), .A2(n27361), .B1(n14203), .Y(
        n14565) );
  sky130_fd_sc_hd__o21ai_0 U14869 ( .A1(n21705), .A2(n21292), .B1(n21291), .Y(
        n21293) );
  sky130_fd_sc_hd__o21ai_0 U14892 ( .A1(n14742), .A2(n27412), .B1(n15192), .Y(
        n15196) );
  sky130_fd_sc_hd__o21ai_0 U14905 ( .A1(n26012), .A2(n25972), .B1(n25886), .Y(
        n23462) );
  sky130_fd_sc_hd__o21ai_0 U14910 ( .A1(n14742), .A2(n27357), .B1(n16530), .Y(
        n16547) );
  sky130_fd_sc_hd__and2_0 U14923 ( .A(n18981), .B(n21776), .X(n29586) );
  sky130_fd_sc_hd__clkinv_1 U15021 ( .A(n16012), .Y(n11095) );
  sky130_fd_sc_hd__nand2_1 U15093 ( .A(j202_soc_core_memory0_ram_dout0[320]), 
        .B(n21593), .Y(n11382) );
  sky130_fd_sc_hd__o21ai_0 U15204 ( .A1(n20101), .A2(n20238), .B1(n20892), .Y(
        n20102) );
  sky130_fd_sc_hd__o21ai_0 U15225 ( .A1(n20002), .A2(n20001), .B1(n13481), .Y(
        n20025) );
  sky130_fd_sc_hd__o21ai_0 U15253 ( .A1(n14742), .A2(n27419), .B1(n14840), .Y(
        n14842) );
  sky130_fd_sc_hd__clkinv_1 U15298 ( .A(n23599), .Y(n23180) );
  sky130_fd_sc_hd__clkinv_1 U15350 ( .A(n17259), .Y(n17261) );
  sky130_fd_sc_hd__clkinv_1 U15436 ( .A(n17137), .Y(n17155) );
  sky130_fd_sc_hd__clkinv_1 U15498 ( .A(n27168), .Y(n12765) );
  sky130_fd_sc_hd__o21ai_0 U15517 ( .A1(j202_soc_core_cmt_core_00_cks1[0]), 
        .A2(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[3]), .B1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[7]), .Y(n23678) );
  sky130_fd_sc_hd__o21ai_0 U15529 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[5]), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[9]), .B1(n24846), .Y(
        n23652) );
  sky130_fd_sc_hd__clkinv_1 U15536 ( .A(n22759), .Y(n22761) );
  sky130_fd_sc_hd__clkinv_1 U15538 ( .A(n27865), .Y(n27758) );
  sky130_fd_sc_hd__clkinv_1 U15544 ( .A(n22582), .Y(n22584) );
  sky130_fd_sc_hd__o21ai_0 U15656 ( .A1(n25993), .A2(n25886), .B1(n25885), .Y(
        n25887) );
  sky130_fd_sc_hd__o21ai_0 U15754 ( .A1(n23296), .A2(n22452), .B1(n22451), .Y(
        n22453) );
  sky130_fd_sc_hd__clkinv_1 U15783 ( .A(n19240), .Y(n21460) );
  sky130_fd_sc_hd__o21ai_0 U15789 ( .A1(n19481), .A2(n22837), .B1(n19483), .Y(
        n19224) );
  sky130_fd_sc_hd__clkinv_1 U15790 ( .A(n17897), .Y(n18889) );
  sky130_fd_sc_hd__nand2_1 U15806 ( .A(n11773), .B(n11772), .Y(n25269) );
  sky130_fd_sc_hd__o21ai_0 U15818 ( .A1(n26352), .A2(n26725), .B1(n26351), .Y(
        n25319) );
  sky130_fd_sc_hd__clkinv_1 U15915 ( .A(j202_soc_core_j22_cpu_regop_Rb__1_), 
        .Y(n13700) );
  sky130_fd_sc_hd__o21ai_0 U16630 ( .A1(n22859), .A2(n11095), .B1(n14540), .Y(
        n14543) );
  sky130_fd_sc_hd__clkinv_1 U16631 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[5]), 
        .Y(n27910) );
  sky130_fd_sc_hd__o21ai_0 U16632 ( .A1(n18916), .A2(n25178), .B1(n25177), .Y(
        n25179) );
  sky130_fd_sc_hd__o21ai_0 U16633 ( .A1(n21951), .A2(n11095), .B1(n14054), .Y(
        n14056) );
  sky130_fd_sc_hd__clkinv_1 U16634 ( .A(n25159), .Y(n26406) );
  sky130_fd_sc_hd__clkinv_1 U16635 ( .A(n26537), .Y(n23735) );
  sky130_fd_sc_hd__nand2_1 U16636 ( .A(n27925), .B(n27553), .Y(n24357) );
  sky130_fd_sc_hd__clkinv_1 U16637 ( .A(n22029), .Y(n17975) );
  sky130_fd_sc_hd__clkinv_1 U16638 ( .A(n13043), .Y(n11803) );
  sky130_fd_sc_hd__a21boi_0 U16639 ( .A1(n26970), .A2(n12688), .B1_N(n24045), 
        .Y(n24047) );
  sky130_fd_sc_hd__o21ai_0 U16640 ( .A1(n15899), .A2(n17110), .B1(n15953), .Y(
        n15205) );
  sky130_fd_sc_hd__clkinv_1 U16641 ( .A(n27780), .Y(n27255) );
  sky130_fd_sc_hd__clkinv_1 U16642 ( .A(n13266), .Y(n13265) );
  sky130_fd_sc_hd__clkinv_1 U16643 ( .A(n21014), .Y(n21016) );
  sky130_fd_sc_hd__clkinv_1 U16644 ( .A(n15413), .Y(n15770) );
  sky130_fd_sc_hd__o21ai_0 U16645 ( .A1(n26684), .A2(n26685), .B1(n26683), .Y(
        n11729) );
  sky130_fd_sc_hd__and2_0 U16646 ( .A(n12888), .B(n12887), .X(n11052) );
  sky130_fd_sc_hd__o21ai_0 U16647 ( .A1(j202_soc_core_wbqspiflash_00_state[3]), 
        .A2(n28067), .B1(n26251), .Y(n26118) );
  sky130_fd_sc_hd__clkinv_1 U16648 ( .A(io_in[15]), .Y(n17154) );
  sky130_fd_sc_hd__and2_0 U16649 ( .A(n20973), .B(n21750), .X(n12182) );
  sky130_fd_sc_hd__a21boi_0 U16650 ( .A1(n17354), .A2(n17355), .B1_N(n17353), 
        .Y(n28916) );
  sky130_fd_sc_hd__clkinv_1 U16651 ( .A(n11644), .Y(n11643) );
  sky130_fd_sc_hd__o21ai_0 U16652 ( .A1(n20320), .A2(n20927), .B1(n20319), .Y(
        n20321) );
  sky130_fd_sc_hd__o21ai_0 U16653 ( .A1(n20212), .A2(n20906), .B1(n20211), .Y(
        n20213) );
  sky130_fd_sc_hd__o21ai_0 U16654 ( .A1(n15413), .A2(n15772), .B1(n15773), .Y(
        n14838) );
  sky130_fd_sc_hd__o21ai_0 U16655 ( .A1(n20275), .A2(n20279), .B1(n20276), .Y(
        n17263) );
  sky130_fd_sc_hd__nor2_1 U16656 ( .A(n24437), .B(n27772), .Y(n24328) );
  sky130_fd_sc_hd__nand2_1 U16657 ( .A(n21752), .B(n21751), .Y(n26530) );
  sky130_fd_sc_hd__o21ai_0 U16658 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[13]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[13]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13]), .Y(n28362) );
  sky130_fd_sc_hd__o21ai_0 U16659 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[3]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[3]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]), .Y(n28293) );
  sky130_fd_sc_hd__o21ai_0 U16660 ( .A1(n26352), .A2(n27183), .B1(n26407), .Y(
        n25419) );
  sky130_fd_sc_hd__o21ai_0 U16661 ( .A1(n24692), .A2(n23236), .B1(n22922), .Y(
        n22928) );
  sky130_fd_sc_hd__o21ai_0 U16662 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[8]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[8]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]), .Y(n28328) );
  sky130_fd_sc_hd__o21ai_0 U16663 ( .A1(n28415), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[20]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[20]), .Y(n28413) );
  sky130_fd_sc_hd__nor2_1 U16664 ( .A(n29030), .B(n11972), .Y(n11971) );
  sky130_fd_sc_hd__o21ai_0 U16665 ( .A1(n22587), .A2(n22586), .B1(n22585), .Y(
        n22588) );
  sky130_fd_sc_hd__o21ai_0 U16666 ( .A1(n25906), .A2(n25986), .B1(n28249), .Y(
        n25892) );
  sky130_fd_sc_hd__o21ai_0 U16667 ( .A1(n22545), .A2(n22352), .B1(n22351), .Y(
        n22354) );
  sky130_fd_sc_hd__clkinv_1 U16668 ( .A(n25273), .Y(n11590) );
  sky130_fd_sc_hd__and2_0 U16669 ( .A(n25703), .B(n26802), .X(n11050) );
  sky130_fd_sc_hd__o21ai_0 U16670 ( .A1(n22847), .A2(n22846), .B1(n22845), .Y(
        n22848) );
  sky130_fd_sc_hd__clkinv_1 U16671 ( .A(n23012), .Y(n26691) );
  sky130_fd_sc_hd__nand2_1 U16672 ( .A(n24417), .B(n11042), .Y(n24388) );
  sky130_fd_sc_hd__or2_0 U16673 ( .A(n13664), .B(n13684), .X(n12171) );
  sky130_fd_sc_hd__and2_0 U16674 ( .A(n22492), .B(n22491), .X(n11045) );
  sky130_fd_sc_hd__clkinv_1 U16675 ( .A(n25337), .Y(n12313) );
  sky130_fd_sc_hd__clkinv_1 U16676 ( .A(n24094), .Y(n24436) );
  sky130_fd_sc_hd__o21ai_0 U16677 ( .A1(n22546), .A2(n23292), .B1(n21964), .Y(
        n21965) );
  sky130_fd_sc_hd__clkinv_1 U16678 ( .A(n23563), .Y(n23306) );
  sky130_fd_sc_hd__o21ai_0 U16679 ( .A1(n21482), .A2(n22586), .B1(n21481), .Y(
        n22328) );
  sky130_fd_sc_hd__o21ai_0 U16680 ( .A1(n24654), .A2(n11774), .B1(n21458), .Y(
        n21465) );
  sky130_fd_sc_hd__and2_0 U16681 ( .A(n21164), .B(n21776), .X(n12281) );
  sky130_fd_sc_hd__o21ai_0 U16682 ( .A1(n26127), .A2(n26054), .B1(n26053), .Y(
        n26055) );
  sky130_fd_sc_hd__o21ai_0 U16683 ( .A1(n26009), .A2(n26051), .B1(n26008), .Y(
        n26010) );
  sky130_fd_sc_hd__o21ai_0 U16684 ( .A1(n25938), .A2(n25937), .B1(n26155), .Y(
        n25939) );
  sky130_fd_sc_hd__o21ai_0 U16685 ( .A1(n28080), .A2(n25961), .B1(n26173), .Y(
        n25965) );
  sky130_fd_sc_hd__o21ai_0 U16686 ( .A1(n25920), .A2(n26254), .B1(n28126), .Y(
        n26122) );
  sky130_fd_sc_hd__and2_0 U16687 ( .A(n21520), .B(n21750), .X(n12235) );
  sky130_fd_sc_hd__and2_0 U16688 ( .A(n21006), .B(n21776), .X(n12282) );
  sky130_fd_sc_hd__o21ai_0 U16689 ( .A1(n20128), .A2(n20925), .B1(n20127), .Y(
        n20129) );
  sky130_fd_sc_hd__o21ai_0 U16690 ( .A1(n17336), .A2(n17335), .B1(n13481), .Y(
        n17349) );
  sky130_fd_sc_hd__clkinv_1 U16691 ( .A(n27256), .Y(n27257) );
  sky130_fd_sc_hd__o21a_1 U16692 ( .A1(n24117), .A2(n23580), .B1(n11129), .X(
        n12411) );
  sky130_fd_sc_hd__o21ai_0 U16693 ( .A1(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .A2(n24285), .B1(n17357), 
        .Y(n24286) );
  sky130_fd_sc_hd__clkinv_1 U16694 ( .A(n24660), .Y(n25815) );
  sky130_fd_sc_hd__o21ai_0 U16695 ( .A1(n24395), .A2(n27956), .B1(n27954), .Y(
        n24396) );
  sky130_fd_sc_hd__o21ai_0 U16696 ( .A1(n24282), .A2(n17357), .B1(n24285), .Y(
        n24283) );
  sky130_fd_sc_hd__o21ai_0 U16697 ( .A1(n28180), .A2(n28187), .B1(n28179), .Y(
        n28181) );
  sky130_fd_sc_hd__o21ai_0 U16698 ( .A1(n25692), .A2(n27764), .B1(n27865), .Y(
        n25693) );
  sky130_fd_sc_hd__o21ai_0 U16699 ( .A1(n25205), .A2(n27097), .B1(n25204), .Y(
        n25206) );
  sky130_fd_sc_hd__o21ai_0 U16700 ( .A1(n22978), .A2(n24624), .B1(n22820), .Y(
        n22821) );
  sky130_fd_sc_hd__o21ai_0 U16701 ( .A1(j202_soc_core_cmt_core_00_cnt1[2]), 
        .A2(n24939), .B1(j202_soc_core_cmt_core_00_cnt1[1]), .Y(n24940) );
  sky130_fd_sc_hd__o21ai_0 U16702 ( .A1(n23780), .A2(n21584), .B1(n21368), .Y(
        n21369) );
  sky130_fd_sc_hd__o21ai_0 U16703 ( .A1(n25860), .A2(n27097), .B1(n25859), .Y(
        n25861) );
  sky130_fd_sc_hd__o21ai_0 U16704 ( .A1(n27540), .A2(n27760), .B1(n27539), .Y(
        n27541) );
  sky130_fd_sc_hd__o21ai_0 U16705 ( .A1(n28590), .A2(n28415), .B1(n28414), .Y(
        n28416) );
  sky130_fd_sc_hd__o21ai_0 U16706 ( .A1(n28438), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[23]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[23]), .Y(n28439) );
  sky130_fd_sc_hd__clkinv_1 U16707 ( .A(n24127), .Y(n11891) );
  sky130_fd_sc_hd__o21ai_0 U16708 ( .A1(n22614), .A2(n22613), .B1(n22612), .Y(
        n22634) );
  sky130_fd_sc_hd__o21ai_0 U16709 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), 
        .A2(n28063), .B1(n26248), .Y(n23688) );
  sky130_fd_sc_hd__o21ai_0 U16710 ( .A1(n25990), .A2(n25993), .B1(n25989), .Y(
        n26004) );
  sky130_fd_sc_hd__o21ai_0 U16711 ( .A1(n22456), .A2(n24380), .B1(n22455), .Y(
        n22457) );
  sky130_fd_sc_hd__nand3_1 U16712 ( .A(n13820), .B(n13324), .C(n12218), .Y(
        n27429) );
  sky130_fd_sc_hd__inv_2 U16713 ( .A(n12918), .Y(n13000) );
  sky130_fd_sc_hd__nor2_1 U16714 ( .A(n22997), .B(n14849), .Y(n23177) );
  sky130_fd_sc_hd__o21ai_0 U16715 ( .A1(n18916), .A2(n26513), .B1(n26512), .Y(
        n26518) );
  sky130_fd_sc_hd__clkinv_1 U16716 ( .A(n11293), .Y(n12556) );
  sky130_fd_sc_hd__o21ai_0 U16717 ( .A1(n24437), .A2(n24436), .B1(n24435), .Y(
        n24439) );
  sky130_fd_sc_hd__buf_1 U16718 ( .A(n27428), .X(n12120) );
  sky130_fd_sc_hd__o21ai_0 U16719 ( .A1(n26301), .A2(n26297), .B1(n26300), .Y(
        n26293) );
  sky130_fd_sc_hd__o21ai_0 U16720 ( .A1(n26808), .A2(n26807), .B1(n26806), .Y(
        n26809) );
  sky130_fd_sc_hd__o21ai_0 U16721 ( .A1(n25953), .A2(n23636), .B1(n28079), .Y(
        n23637) );
  sky130_fd_sc_hd__o21ai_0 U16722 ( .A1(n26018), .A2(n28250), .B1(n28083), .Y(
        n28238) );
  sky130_fd_sc_hd__o21ai_0 U16723 ( .A1(n28229), .A2(n28243), .B1(n26252), .Y(
        n26253) );
  sky130_fd_sc_hd__o21ai_0 U16724 ( .A1(j202_soc_core_wbqspiflash_00_spi_wr), 
        .A2(n26244), .B1(n26243), .Y(n26245) );
  sky130_fd_sc_hd__o21ai_0 U16725 ( .A1(n26152), .A2(n26151), .B1(n26150), .Y(
        n26157) );
  sky130_fd_sc_hd__o211a_2 U16726 ( .A1(n26417), .A2(n11143), .B1(n13723), 
        .C1(n13722), .X(n12197) );
  sky130_fd_sc_hd__buf_1 U16727 ( .A(n26519), .X(n11771) );
  sky130_fd_sc_hd__nor2_1 U16728 ( .A(n13209), .B(n13206), .Y(n17354) );
  sky130_fd_sc_hd__clkinv_1 U16729 ( .A(n23770), .Y(n24534) );
  sky130_fd_sc_hd__clkinv_1 U16730 ( .A(n13055), .Y(n24423) );
  sky130_fd_sc_hd__o21ai_0 U16731 ( .A1(n27930), .A2(n29593), .B1(n27950), .Y(
        n27922) );
  sky130_fd_sc_hd__inv_2 U16732 ( .A(n23812), .Y(n23813) );
  sky130_fd_sc_hd__and2_0 U16733 ( .A(n28743), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd), .X(n28733) );
  sky130_fd_sc_hd__o21ai_0 U16734 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[7]), .A2(n27829), .B1(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_0_), .Y(
        n27322) );
  sky130_fd_sc_hd__o21ai_0 U16735 ( .A1(n27014), .A2(n27013), .B1(n27012), .Y(
        n27017) );
  sky130_fd_sc_hd__and2_0 U16736 ( .A(n15306), .B(n12216), .X(n12247) );
  sky130_fd_sc_hd__o21ai_0 U16737 ( .A1(n25506), .A2(n27013), .B1(n25497), .Y(
        n25500) );
  sky130_fd_sc_hd__o21ai_0 U16738 ( .A1(j202_soc_core_uart_BRG_br_cnt[5]), 
        .A2(n28041), .B1(n28037), .Y(n28038) );
  sky130_fd_sc_hd__o21ai_0 U16739 ( .A1(j202_soc_core_uart_TOP_tx_bit_cnt[0]), 
        .A2(j202_soc_core_uart_TOP_tx_bit_cnt[1]), .B1(n28007), .Y(n28002) );
  sky130_fd_sc_hd__o21ai_0 U16740 ( .A1(n25515), .A2(n25514), .B1(n25513), .Y(
        n25518) );
  sky130_fd_sc_hd__o21ai_0 U16741 ( .A1(n25475), .A2(n25514), .B1(n25474), .Y(
        n25478) );
  sky130_fd_sc_hd__o21ai_0 U16742 ( .A1(n28590), .A2(
        j202_soc_core_qspi_wb_wdat[19]), .B1(n28506), .Y(n28409) );
  sky130_fd_sc_hd__o21ai_0 U16743 ( .A1(n27014), .A2(n25514), .B1(n25468), .Y(
        n25471) );
  sky130_fd_sc_hd__o21ai_0 U16744 ( .A1(n27479), .A2(n27478), .B1(
        j202_soc_core_cmt_core_00_cnt0[15]), .Y(n27485) );
  sky130_fd_sc_hd__o21ai_0 U16745 ( .A1(n28619), .A2(n26277), .B1(n25583), .Y(
        n25586) );
  sky130_fd_sc_hd__o21ai_0 U16746 ( .A1(n28619), .A2(n25573), .B1(n25583), .Y(
        n26916) );
  sky130_fd_sc_hd__o21ai_0 U16747 ( .A1(n28619), .A2(n25568), .B1(n25583), .Y(
        n25560) );
  sky130_fd_sc_hd__o21ai_0 U16748 ( .A1(n28590), .A2(
        j202_soc_core_qspi_wb_wdat[25]), .B1(n28506), .Y(n28456) );
  sky130_fd_sc_hd__o21ai_0 U16749 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[2]), .A2(n24887), .B1(
        n24890), .Y(n24888) );
  sky130_fd_sc_hd__o21ai_0 U16750 ( .A1(n26301), .A2(n25593), .B1(n25592), .Y(
        n25594) );
  sky130_fd_sc_hd__o21ai_0 U16751 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[2]), .A2(n24825), .B1(
        n24828), .Y(n24826) );
  sky130_fd_sc_hd__clkinv_1 U16752 ( .A(j202_soc_core_intc_core_00_rg_ipr[44]), 
        .Y(n25461) );
  sky130_fd_sc_hd__clkinv_1 U16753 ( .A(j202_soc_core_intc_core_00_rg_ipr[69]), 
        .Y(n26900) );
  sky130_fd_sc_hd__o21ai_0 U16754 ( .A1(n25515), .A2(n27013), .B1(n25488), .Y(
        n25491) );
  sky130_fd_sc_hd__o21ai_0 U16755 ( .A1(n28590), .A2(
        j202_soc_core_qspi_wb_wdat[27]), .B1(n28506), .Y(n28472) );
  sky130_fd_sc_hd__o21ai_0 U16764 ( .A1(j202_soc_core_uart_BRG_ps[3]), .A2(
        n28019), .B1(n28021), .Y(n28020) );
  sky130_fd_sc_hd__or2_0 U16768 ( .A(n28948), .B(n22676), .X(n12162) );
  sky130_fd_sc_hd__o21ai_0 U16781 ( .A1(n27755), .A2(n28476), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[0]), .Y(n27744) );
  sky130_fd_sc_hd__o21ai_0 U16783 ( .A1(n28300), .A2(n28476), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[4]), .Y(n28301) );
  sky130_fd_sc_hd__o21ai_0 U16787 ( .A1(n28326), .A2(n28476), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[8]), .Y(n28331) );
  sky130_fd_sc_hd__o21ai_0 U16790 ( .A1(n28355), .A2(n28476), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[12]), .Y(n28356) );
  sky130_fd_sc_hd__o21ai_0 U16794 ( .A1(n28590), .A2(
        j202_soc_core_qspi_wb_wdat[18]), .B1(n28506), .Y(n28401) );
  sky130_fd_sc_hd__o21ai_0 U16803 ( .A1(n28590), .A2(
        j202_soc_core_qspi_wb_wdat[22]), .B1(n28506), .Y(n28434) );
  sky130_fd_sc_hd__o21ai_0 U16829 ( .A1(n28590), .A2(
        j202_soc_core_qspi_wb_wdat[26]), .B1(n28506), .Y(n28464) );
  sky130_fd_sc_hd__o21ai_0 U16831 ( .A1(n28590), .A2(
        j202_soc_core_qspi_wb_wdat[29]), .B1(n28506), .Y(n28490) );
  sky130_fd_sc_hd__nor2_1 U16835 ( .A(n23179), .B(n24127), .Y(n11895) );
  sky130_fd_sc_hd__o21ai_0 U16843 ( .A1(n25787), .A2(n23235), .B1(n25786), .Y(
        n25845) );
  sky130_fd_sc_hd__and4_2 U16858 ( .A(n24796), .B(n24794), .C(n11372), .D(
        n11370), .X(n12433) );
  sky130_fd_sc_hd__o21ai_0 U16865 ( .A1(n28230), .A2(n23440), .B1(n28067), .Y(
        n24996) );
  sky130_fd_sc_hd__clkinv_1 U16879 ( .A(n24163), .Y(n25276) );
  sky130_fd_sc_hd__clkinv_1 U16887 ( .A(n27395), .Y(n27524) );
  sky130_fd_sc_hd__clkinv_1 U16892 ( .A(n26393), .Y(n26382) );
  sky130_fd_sc_hd__clkinv_1 U16895 ( .A(n23079), .Y(n26379) );
  sky130_fd_sc_hd__clkinv_1 U16914 ( .A(n24629), .Y(n11103) );
  sky130_fd_sc_hd__nor2_1 U16927 ( .A(n24053), .B(n27356), .Y(n27441) );
  sky130_fd_sc_hd__and2_0 U16940 ( .A(n27273), .B(n12783), .X(n12276) );
  sky130_fd_sc_hd__and2_0 U17035 ( .A(n27273), .B(n12781), .X(n12275) );
  sky130_fd_sc_hd__nor2_1 U17041 ( .A(n24118), .B(n25107), .Y(n12459) );
  sky130_fd_sc_hd__o21ai_0 U17082 ( .A1(n29523), .A2(n12712), .B1(n27980), .Y(
        n24415) );
  sky130_fd_sc_hd__clkinv_1 U17083 ( .A(n27333), .Y(n11137) );
  sky130_fd_sc_hd__clkinv_1 U17094 ( .A(n27417), .Y(n12504) );
  sky130_fd_sc_hd__o21ai_0 U17110 ( .A1(n26518), .A2(n26517), .B1(n26516), .Y(
        n26522) );
  sky130_fd_sc_hd__a21o_1 U17150 ( .A1(n13526), .A2(n13527), .B1(n12200), .X(
        n24113) );
  sky130_fd_sc_hd__o21ai_0 U17176 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[7]), .A2(n27831), .B1(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_0_), .Y(
        n27324) );
  sky130_fd_sc_hd__o21ai_0 U17177 ( .A1(n24426), .A2(n24438), .B1(n27980), .Y(
        n24427) );
  sky130_fd_sc_hd__o21ai_0 U17188 ( .A1(n29523), .A2(n12556), .B1(n27980), .Y(
        n27981) );
  sky130_fd_sc_hd__o21ai_0 U17193 ( .A1(n26800), .A2(n26799), .B1(n26798), .Y(
        n26811) );
  sky130_fd_sc_hd__and2_0 U17205 ( .A(n15777), .B(n12199), .X(n11046) );
  sky130_fd_sc_hd__o21ai_0 U17225 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), 
        .A2(n26257), .B1(n26256), .Y(n26258) );
  sky130_fd_sc_hd__a2bb2oi_1 U17230 ( .B1(n23563), .B2(n24119), .A1_N(n23304), 
        .A2_N(n12085), .Y(n25111) );
  sky130_fd_sc_hd__a21oi_1 U17233 ( .A1(j202_soc_core_memory0_ram_dout0[481]), 
        .A2(n21771), .B1(n19913), .Y(n20562) );
  sky130_fd_sc_hd__o21ai_0 U17244 ( .A1(n25506), .A2(n25514), .B1(n25505), .Y(
        n25509) );
  sky130_fd_sc_hd__and2_0 U17254 ( .A(n27961), .B(n27969), .X(n13303) );
  sky130_fd_sc_hd__and2_0 U17262 ( .A(n19244), .B(n19245), .X(n11060) );
  sky130_fd_sc_hd__clkinv_1 U17263 ( .A(n29066), .Y(n27619) );
  sky130_fd_sc_hd__o21ai_0 U17265 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[3]), .A2(n24232), .B1(
        n24236), .Y(n24234) );
  sky130_fd_sc_hd__and2_0 U17266 ( .A(n28998), .B(n24210), .X(n11080) );
  sky130_fd_sc_hd__o21ai_0 U17283 ( .A1(n24288), .A2(n27272), .B1(n24287), .Y(
        j202_soc_core_j22_cpu_ml_N153) );
  sky130_fd_sc_hd__o21ai_0 U17284 ( .A1(n28063), .A2(n25025), .B1(n12142), .Y(
        j202_soc_core_wbqspiflash_00_N742) );
  sky130_fd_sc_hd__o21ai_0 U17298 ( .A1(n26398), .A2(n27272), .B1(n24284), .Y(
        j202_soc_core_j22_cpu_ml_N152) );
  sky130_fd_sc_hd__o21ai_0 U17299 ( .A1(n28661), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B1(n28593), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N394) );
  sky130_fd_sc_hd__o21ai_0 U17300 ( .A1(n26231), .A2(n26216), .B1(n26215), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N428) );
  sky130_fd_sc_hd__o21ai_0 U17301 ( .A1(n28352), .A2(n28351), .B1(n28350), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N51) );
  sky130_fd_sc_hd__o21ai_0 U17302 ( .A1(n27501), .A2(n27500), .B1(n27499), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[15]) );
  sky130_fd_sc_hd__o21ai_0 U17303 ( .A1(n28564), .A2(n28563), .B1(n12142), .Y(
        j202_soc_core_uart_TOP_N43) );
  sky130_fd_sc_hd__o21ai_0 U17314 ( .A1(j202_soc_core_uart_TOP_tx_bit_cnt[0]), 
        .A2(n28003), .B1(n12142), .Y(j202_soc_core_uart_TOP_N58) );
  sky130_fd_sc_hd__o21ai_0 U17318 ( .A1(n28560), .A2(n28559), .B1(n28558), .Y(
        n24) );
  sky130_fd_sc_hd__o21ai_0 U17333 ( .A1(n25699), .A2(n27593), .B1(n25698), .Y(
        n25) );
  sky130_fd_sc_hd__and2_0 U17335 ( .A(n27190), .B(n26450), .X(n12269) );
  sky130_fd_sc_hd__o21ai_0 U17338 ( .A1(n27192), .A2(n27414), .B1(n27191), .Y(
        j202_soc_core_j22_cpu_rf_N3294) );
  sky130_fd_sc_hd__o21ai_0 U17350 ( .A1(n27799), .A2(n27473), .B1(n27472), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[13]) );
  sky130_fd_sc_hd__o21ai_0 U17365 ( .A1(j202_soc_core_cmt_core_00_cnt0[7]), 
        .A2(n25589), .B1(n25580), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[7]) );
  sky130_fd_sc_hd__o21ai_0 U17419 ( .A1(n25562), .A2(n25560), .B1(n24879), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[2]) );
  sky130_fd_sc_hd__o21ai_0 U17420 ( .A1(n25742), .A2(n27983), .B1(n25741), .Y(
        n31) );
  sky130_fd_sc_hd__o21ai_0 U17422 ( .A1(n27647), .A2(n27646), .B1(n27645), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N41) );
  sky130_fd_sc_hd__o21ai_0 U17425 ( .A1(n24938), .A2(n24943), .B1(n24937), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[1]) );
  sky130_fd_sc_hd__o21ai_0 U17439 ( .A1(n25604), .A2(n25603), .B1(n25602), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[6]) );
  sky130_fd_sc_hd__o21ai_0 U17442 ( .A1(n27611), .A2(n27829), .B1(n24847), .Y(
        n33) );
  sky130_fd_sc_hd__and2_0 U17443 ( .A(n29067), .B(n29062), .X(n13315) );
  sky130_fd_sc_hd__and2_0 U17445 ( .A(n29067), .B(n29010), .X(n12243) );
  sky130_fd_sc_hd__o21ai_0 U17447 ( .A1(n28289), .A2(n28288), .B1(n28287), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N42) );
  sky130_fd_sc_hd__o21ai_0 U17448 ( .A1(n28387), .A2(n28386), .B1(n28385), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N56) );
  sky130_fd_sc_hd__o21ai_0 U17451 ( .A1(n28380), .A2(n28379), .B1(n28378), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N55) );
  sky130_fd_sc_hd__and2_0 U17453 ( .A(n12899), .B(n27620), .X(n29590) );
  sky130_fd_sc_hd__and2_0 U17459 ( .A(n12435), .B(n26450), .X(n13344) );
  sky130_fd_sc_hd__o21ai_0 U17466 ( .A1(n27109), .A2(n27108), .B1(n27107), .Y(
        n43) );
  sky130_fd_sc_hd__o21ai_0 U17468 ( .A1(n27741), .A2(n27728), .B1(n27727), .Y(
        n47) );
  sky130_fd_sc_hd__o21ai_0 U17476 ( .A1(n27984), .A2(n27983), .B1(n27982), .Y(
        n58) );
  sky130_fd_sc_hd__o21ai_0 U17477 ( .A1(n25870), .A2(n27108), .B1(n25869), .Y(
        n69) );
  sky130_fd_sc_hd__o21ai_0 U17478 ( .A1(n27460), .A2(n12433), .B1(n25260), .Y(
        j202_soc_core_j22_cpu_rf_N3290) );
  sky130_fd_sc_hd__o21ai_0 U17481 ( .A1(n28552), .A2(n28551), .B1(n28550), .Y(
        j202_soc_core_wbqspiflash_00_N608) );
  sky130_fd_sc_hd__o21ai_0 U17483 ( .A1(n10959), .A2(n26130), .B1(n26251), .Y(
        j202_soc_core_wbqspiflash_00_N663) );
  sky130_fd_sc_hd__o21ai_0 U17498 ( .A1(n26478), .A2(n28096), .B1(n26477), .Y(
        j202_soc_core_wbqspiflash_00_N740) );
  sky130_fd_sc_hd__o21ai_0 U17503 ( .A1(n26187), .A2(n26252), .B1(n26186), .Y(
        j202_soc_core_wbqspiflash_00_N592) );
  sky130_fd_sc_hd__o21ai_0 U17510 ( .A1(n27043), .A2(n27042), .B1(n27041), .Y(
        n71) );
  sky130_fd_sc_hd__o21ai_0 U17511 ( .A1(n26981), .A2(n24513), .B1(n24512), .Y(
        j202_soc_core_j22_cpu_ml_maclj[30]) );
  sky130_fd_sc_hd__o21ai_0 U17515 ( .A1(n25114), .A2(n27108), .B1(n25113), .Y(
        n73) );
  sky130_fd_sc_hd__and2_0 U17518 ( .A(n12644), .B(n26450), .X(n13331) );
  sky130_fd_sc_hd__o21ai_0 U17521 ( .A1(n27192), .A2(n27451), .B1(n24747), .Y(
        j202_soc_core_j22_cpu_rf_N3288) );
  sky130_fd_sc_hd__o21ai_0 U17523 ( .A1(n27275), .A2(n27274), .B1(n27273), .Y(
        j202_soc_core_j22_cpu_ml_machj[10]) );
  sky130_fd_sc_hd__o21ai_0 U17533 ( .A1(n25335), .A2(n27275), .B1(n25055), .Y(
        j202_soc_core_j22_cpu_rf_N3356) );
  sky130_fd_sc_hd__and2_0 U17539 ( .A(n25878), .B(n26450), .X(n29115) );
  sky130_fd_sc_hd__o21ai_0 U17560 ( .A1(n26951), .A2(n25853), .B1(n25852), .Y(
        j202_soc_core_j22_cpu_rf_N3372) );
  sky130_fd_sc_hd__o21ai_0 U17561 ( .A1(n27192), .A2(n27407), .B1(n26104), .Y(
        j202_soc_core_j22_cpu_rf_N3295) );
  sky130_fd_sc_hd__o21ai_0 U17563 ( .A1(n27460), .A2(n27127), .B1(n27126), .Y(
        j202_soc_core_j22_cpu_rf_N3286) );
  sky130_fd_sc_hd__o21ai_0 U17579 ( .A1(n27217), .A2(n26395), .B1(n26366), .Y(
        j202_soc_core_j22_cpu_rf_N2839) );
  sky130_fd_sc_hd__o21ai_0 U17586 ( .A1(n25335), .A2(n24691), .B1(n24690), .Y(
        j202_soc_core_j22_cpu_rf_N3357) );
  sky130_fd_sc_hd__and2_0 U17591 ( .A(n12385), .B(n26450), .X(n12270) );
  sky130_fd_sc_hd__o21ai_0 U17592 ( .A1(n27209), .A2(n25157), .B1(n23040), .Y(
        j202_soc_core_j22_cpu_rf_N2745) );
  sky130_fd_sc_hd__o21ai_0 U17597 ( .A1(n27460), .A2(n12473), .B1(n25660), .Y(
        j202_soc_core_j22_cpu_rf_N3291) );
  sky130_fd_sc_hd__o21ai_0 U17611 ( .A1(n27418), .A2(n27417), .B1(n27416), .Y(
        j202_soc_core_j22_cpu_ml_N417) );
  sky130_fd_sc_hd__and2_0 U17612 ( .A(n29242), .B(n24112), .X(n29119) );
  sky130_fd_sc_hd__o21ai_0 U17653 ( .A1(n24948), .A2(n27829), .B1(n24881), .Y(
        n75) );
  sky130_fd_sc_hd__o21ai_0 U17668 ( .A1(n27731), .A2(n24883), .B1(n24821), .Y(
        n80) );
  sky130_fd_sc_hd__o21ai_0 U17669 ( .A1(n24278), .A2(n27337), .B1(n27336), .Y(
        j202_soc_core_j22_cpu_ml_N194) );
  sky130_fd_sc_hd__o21ai_0 U17674 ( .A1(n14849), .A2(n25554), .B1(n26814), .Y(
        j202_soc_core_j22_cpu_rf_N2639) );
  sky130_fd_sc_hd__o21ai_0 U17676 ( .A1(n27192), .A2(n25640), .B1(n24734), .Y(
        j202_soc_core_j22_cpu_rf_N3280) );
  sky130_fd_sc_hd__o21ai_0 U17684 ( .A1(n26951), .A2(n25559), .B1(n25558), .Y(
        j202_soc_core_j22_cpu_rf_N3355) );
  sky130_fd_sc_hd__o21ai_0 U17685 ( .A1(n27460), .A2(n26066), .B1(n26065), .Y(
        j202_soc_core_j22_cpu_rf_N3296) );
  sky130_fd_sc_hd__o21ai_0 U17708 ( .A1(n28318), .A2(n28281), .B1(n28280), .Y(
        n88) );
  sky130_fd_sc_hd__o21ai_0 U17709 ( .A1(n28291), .A2(n28281), .B1(n28275), .Y(
        n92) );
  sky130_fd_sc_hd__o21ai_0 U17710 ( .A1(n27928), .A2(n24256), .B1(n24259), .Y(
        n10589) );
  sky130_fd_sc_hd__o21ai_0 U17712 ( .A1(n27226), .A2(n27359), .B1(n13032), .Y(
        j202_soc_core_j22_cpu_rf_N3156) );
  sky130_fd_sc_hd__o21ai_2 U17714 ( .A1(n23543), .A2(n23541), .B1(n27574), .Y(
        j202_soc_core_j22_cpu_rf_N3116) );
  sky130_fd_sc_hd__o21ai_0 U17740 ( .A1(n27215), .A2(n27461), .B1(n24555), .Y(
        j202_soc_core_j22_cpu_rf_N2914) );
  sky130_fd_sc_hd__o21ai_0 U17764 ( .A1(n27460), .A2(n25223), .B1(n25076), .Y(
        j202_soc_core_j22_cpu_rf_N3299) );
  sky130_fd_sc_hd__o21ai_0 U17765 ( .A1(n26986), .A2(n27827), .B1(n26982), .Y(
        n97) );
  sky130_fd_sc_hd__o21ai_0 U17766 ( .A1(n27326), .A2(n27833), .B1(n27325), .Y(
        n107) );
  sky130_fd_sc_hd__o21ai_0 U17767 ( .A1(n27722), .A2(n27721), .B1(n27720), .Y(
        j202_soc_core_j22_cpu_ma_N53) );
  sky130_fd_sc_hd__o21ai_0 U17768 ( .A1(n12397), .A2(n27928), .B1(n24314), .Y(
        n10603) );
  sky130_fd_sc_hd__o21ai_0 U17808 ( .A1(n27834), .A2(n27833), .B1(n27832), .Y(
        n115) );
  sky130_fd_sc_hd__o21ai_0 U17824 ( .A1(n27237), .A2(n27833), .B1(n27236), .Y(
        n120) );
  sky130_fd_sc_hd__o21ai_0 U17827 ( .A1(n27138), .A2(n27135), .B1(n27132), .Y(
        n131) );
  sky130_fd_sc_hd__o21ai_0 U17828 ( .A1(n28389), .A2(n27593), .B1(n25739), .Y(
        n133) );
  sky130_fd_sc_hd__o21ai_0 U17829 ( .A1(n27527), .A2(n27829), .B1(n25762), .Y(
        n134) );
  sky130_fd_sc_hd__o21ai_0 U17830 ( .A1(n25012), .A2(n25011), .B1(n25010), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N314) );
  sky130_fd_sc_hd__o21ai_0 U17832 ( .A1(n24293), .A2(n27337), .B1(n24289), .Y(
        j202_soc_core_j22_cpu_ml_N195) );
  sky130_fd_sc_hd__o21ai_0 U17842 ( .A1(n29076), .A2(n27607), .B1(n27606), .Y(
        n136) );
  sky130_fd_sc_hd__clkinv_1 U17843 ( .A(n29027), .Y(n10543) );
  sky130_fd_sc_hd__clkinv_1 U17847 ( .A(n29024), .Y(n10549) );
  sky130_fd_sc_hd__clkinv_1 U17857 ( .A(n29022), .Y(n10553) );
  sky130_fd_sc_hd__conb_1 U17867 ( .LO(n29363), .HI(
        j202_soc_core_ahb2aqu_00_N127) );
  sky130_fd_sc_hd__clkinv_1 U17875 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        user_irq[0]) );
  sky130_fd_sc_hd__clkinv_1 U17900 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        user_irq[1]) );
  sky130_fd_sc_hd__clkinv_1 U17908 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        user_irq[2]) );
  sky130_fd_sc_hd__clkinv_1 U17920 ( .A(n29363), .Y(io_oeb[5]) );
  sky130_fd_sc_hd__clkinv_1 U17927 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[6]) );
  sky130_fd_sc_hd__clkinv_1 U17956 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[8]) );
  sky130_fd_sc_hd__clkinv_1 U17977 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[9]) );
  sky130_fd_sc_hd__clkinv_1 U17983 ( .A(n29363), .Y(io_oeb[14]) );
  sky130_fd_sc_hd__clkinv_1 U17998 ( .A(n29363), .Y(io_oeb[15]) );
  sky130_fd_sc_hd__clkinv_1 U17999 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[16]) );
  sky130_fd_sc_hd__clkinv_1 U18000 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[17]) );
  sky130_fd_sc_hd__clkinv_1 U18001 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[18]) );
  sky130_fd_sc_hd__clkinv_1 U18023 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[19]) );
  sky130_fd_sc_hd__clkinv_1 U18033 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[20]) );
  sky130_fd_sc_hd__clkinv_1 U18045 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[21]) );
  sky130_fd_sc_hd__clkinv_1 U18052 ( .A(n29363), .Y(io_oeb[22]) );
  sky130_fd_sc_hd__clkinv_1 U18054 ( .A(n29363), .Y(io_oeb[23]) );
  sky130_fd_sc_hd__clkinv_1 U18062 ( .A(n29363), .Y(io_oeb[24]) );
  sky130_fd_sc_hd__clkinv_1 U18067 ( .A(n29363), .Y(io_oeb[25]) );
  sky130_fd_sc_hd__clkinv_1 U18074 ( .A(n29363), .Y(io_oeb[37]) );
  sky130_fd_sc_hd__clkinv_1 U18082 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[5]) );
  sky130_fd_sc_hd__clkinv_1 U18083 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[14]) );
  sky130_fd_sc_hd__clkinv_1 U18084 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[15]) );
  sky130_fd_sc_hd__clkinv_1 U18091 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[22]) );
  sky130_fd_sc_hd__clkinv_1 U18114 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[23]) );
  sky130_fd_sc_hd__clkinv_1 U18130 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[24]) );
  sky130_fd_sc_hd__clkinv_1 U18140 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[25]) );
  sky130_fd_sc_hd__clkinv_1 U18161 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[37]) );
  sky130_fd_sc_hd__clkinv_1 U18166 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[32]) );
  sky130_fd_sc_hd__clkinv_1 U18169 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[33]) );
  sky130_fd_sc_hd__clkinv_1 U18180 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[34]) );
  sky130_fd_sc_hd__clkinv_1 U18185 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[35]) );
  sky130_fd_sc_hd__clkinv_1 U18189 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[36]) );
  sky130_fd_sc_hd__clkinv_1 U18209 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[37]) );
  sky130_fd_sc_hd__clkinv_1 U18268 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[38]) );
  sky130_fd_sc_hd__clkinv_1 U18327 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[39]) );
  sky130_fd_sc_hd__clkinv_1 U18337 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[40]) );
  sky130_fd_sc_hd__clkinv_1 U18338 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[41]) );
  sky130_fd_sc_hd__clkinv_1 U18372 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[42]) );
  sky130_fd_sc_hd__clkinv_1 U18402 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[43]) );
  sky130_fd_sc_hd__clkinv_1 U18417 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[44]) );
  sky130_fd_sc_hd__clkinv_1 U18418 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[45]) );
  sky130_fd_sc_hd__clkinv_1 U18465 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[46]) );
  sky130_fd_sc_hd__clkinv_1 U18477 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[47]) );
  sky130_fd_sc_hd__clkinv_1 U18492 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[48]) );
  sky130_fd_sc_hd__clkinv_1 U18494 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[49]) );
  sky130_fd_sc_hd__clkinv_1 U18526 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[50]) );
  sky130_fd_sc_hd__clkinv_1 U18536 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[51]) );
  sky130_fd_sc_hd__clkinv_1 U18568 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[52]) );
  sky130_fd_sc_hd__clkinv_1 U18601 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[53]) );
  sky130_fd_sc_hd__clkinv_1 U18629 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[54]) );
  sky130_fd_sc_hd__clkinv_1 U18655 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[55]) );
  sky130_fd_sc_hd__clkinv_1 U18664 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[56]) );
  sky130_fd_sc_hd__clkinv_1 U18736 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[57]) );
  sky130_fd_sc_hd__clkinv_1 U18817 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[58]) );
  sky130_fd_sc_hd__clkinv_1 U18819 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[59]) );
  sky130_fd_sc_hd__clkinv_1 U18828 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[60]) );
  sky130_fd_sc_hd__clkinv_1 U18829 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[61]) );
  sky130_fd_sc_hd__clkinv_1 U18837 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[62]) );
  sky130_fd_sc_hd__clkinv_1 U18845 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[63]) );
  sky130_fd_sc_hd__clkinv_1 U18859 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[64]) );
  sky130_fd_sc_hd__clkinv_1 U18865 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[65]) );
  sky130_fd_sc_hd__clkinv_1 U18890 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[66]) );
  sky130_fd_sc_hd__clkinv_1 U18907 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[67]) );
  sky130_fd_sc_hd__clkinv_1 U18908 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[68]) );
  sky130_fd_sc_hd__clkinv_1 U18915 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[69]) );
  sky130_fd_sc_hd__clkinv_1 U18918 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[70]) );
  sky130_fd_sc_hd__clkinv_1 U18932 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[71]) );
  sky130_fd_sc_hd__clkinv_1 U18941 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[72]) );
  sky130_fd_sc_hd__clkinv_1 U19045 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[73]) );
  sky130_fd_sc_hd__clkinv_1 U19053 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[74]) );
  sky130_fd_sc_hd__clkinv_1 U19058 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[75]) );
  sky130_fd_sc_hd__clkinv_1 U19077 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[76]) );
  sky130_fd_sc_hd__clkinv_1 U19082 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[77]) );
  sky130_fd_sc_hd__clkinv_1 U19085 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[78]) );
  sky130_fd_sc_hd__clkinv_1 U19088 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[79]) );
  sky130_fd_sc_hd__clkinv_1 U19108 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[80]) );
  sky130_fd_sc_hd__clkinv_1 U19135 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[81]) );
  sky130_fd_sc_hd__clkinv_1 U19146 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[82]) );
  sky130_fd_sc_hd__clkinv_1 U19154 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[83]) );
  sky130_fd_sc_hd__clkinv_1 U19157 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[84]) );
  sky130_fd_sc_hd__clkinv_1 U19172 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[85]) );
  sky130_fd_sc_hd__clkinv_1 U19258 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[86]) );
  sky130_fd_sc_hd__clkinv_1 U19275 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[87]) );
  sky130_fd_sc_hd__clkinv_1 U19284 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[88]) );
  sky130_fd_sc_hd__clkinv_1 U19300 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[89]) );
  sky130_fd_sc_hd__clkinv_1 U19338 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[90]) );
  sky130_fd_sc_hd__clkinv_1 U19383 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[91]) );
  sky130_fd_sc_hd__clkinv_1 U19397 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[92]) );
  sky130_fd_sc_hd__clkinv_1 U19406 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[93]) );
  sky130_fd_sc_hd__clkinv_1 U19415 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[94]) );
  sky130_fd_sc_hd__clkinv_1 U19433 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[95]) );
  sky130_fd_sc_hd__clkinv_1 U19435 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[96]) );
  sky130_fd_sc_hd__clkinv_1 U19438 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[97]) );
  sky130_fd_sc_hd__clkinv_1 U19461 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[98]) );
  sky130_fd_sc_hd__clkinv_1 U19467 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[99]) );
  sky130_fd_sc_hd__clkinv_1 U19484 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[100]) );
  sky130_fd_sc_hd__clkinv_1 U19498 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[101]) );
  sky130_fd_sc_hd__clkinv_1 U19508 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[102]) );
  sky130_fd_sc_hd__clkinv_1 U19614 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[103]) );
  sky130_fd_sc_hd__clkinv_1 U19615 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[104]) );
  sky130_fd_sc_hd__clkinv_1 U19617 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[105]) );
  sky130_fd_sc_hd__clkinv_1 U19618 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[106]) );
  sky130_fd_sc_hd__clkinv_1 U19619 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[107]) );
  sky130_fd_sc_hd__clkinv_1 U19620 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[108]) );
  sky130_fd_sc_hd__clkinv_1 U19621 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[109]) );
  sky130_fd_sc_hd__clkinv_1 U19622 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[110]) );
  sky130_fd_sc_hd__clkinv_1 U19623 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[111]) );
  sky130_fd_sc_hd__clkinv_1 U19624 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[112]) );
  sky130_fd_sc_hd__clkinv_1 U19625 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[113]) );
  sky130_fd_sc_hd__clkinv_1 U19626 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[114]) );
  sky130_fd_sc_hd__clkinv_1 U19627 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[115]) );
  sky130_fd_sc_hd__clkinv_1 U19628 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[116]) );
  sky130_fd_sc_hd__clkinv_1 U19629 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[117]) );
  sky130_fd_sc_hd__clkinv_1 U19630 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[118]) );
  sky130_fd_sc_hd__clkinv_1 U19631 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[119]) );
  sky130_fd_sc_hd__clkinv_1 U19637 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[120]) );
  sky130_fd_sc_hd__clkinv_1 U19641 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[121]) );
  sky130_fd_sc_hd__clkinv_1 U19684 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[122]) );
  sky130_fd_sc_hd__clkinv_1 U19718 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[123]) );
  sky130_fd_sc_hd__clkinv_1 U19726 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[124]) );
  sky130_fd_sc_hd__clkinv_1 U19739 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[125]) );
  sky130_fd_sc_hd__clkinv_1 U19742 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[126]) );
  sky130_fd_sc_hd__clkinv_1 U19743 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[127]) );
  sky130_fd_sc_hd__and2_4 U19755 ( .A(n11129), .B(n29013), .X(n29488) );
  sky130_fd_sc_hd__buf_2 U19759 ( .A(n28562), .X(n12142) );
  sky130_fd_sc_hd__clkinv_1 U19787 ( .A(n28590), .Y(n29595) );
  sky130_fd_sc_hd__clkinv_1 U19788 ( .A(n26802), .Y(n29535) );
  sky130_fd_sc_hd__clkinv_1 U19791 ( .A(n12480), .Y(n27948) );
  sky130_fd_sc_hd__and2_0 U19826 ( .A(n12902), .B(n12899), .X(n29489) );
  sky130_fd_sc_hd__and2_0 U19827 ( .A(n29516), .B(n27948), .X(n29490) );
  sky130_fd_sc_hd__or2_0 U19829 ( .A(n27775), .B(n27774), .X(n29491) );
  sky130_fd_sc_hd__and2_0 U19831 ( .A(n17159), .B(n12237), .X(n29492) );
  sky130_fd_sc_hd__or2_0 U19853 ( .A(n11536), .B(n11537), .X(n29493) );
  sky130_fd_sc_hd__and2_4 U19854 ( .A(n11129), .B(n23578), .X(n29494) );
  sky130_fd_sc_hd__nand2_1 U19855 ( .A(n11895), .B(n24565), .Y(n12464) );
  sky130_fd_sc_hd__inv_2 U19872 ( .A(n11892), .Y(n11894) );
  sky130_fd_sc_hd__clkinv_1 U19874 ( .A(n27561), .Y(n24338) );
  sky130_fd_sc_hd__clkinv_1 U19910 ( .A(n29009), .Y(n27523) );
  sky130_fd_sc_hd__or2_0 U19919 ( .A(n25144), .B(n23015), .X(n29495) );
  sky130_fd_sc_hd__and2_0 U19925 ( .A(n26399), .B(n12294), .X(n29496) );
  sky130_fd_sc_hd__and2_0 U19937 ( .A(n11567), .B(n11582), .X(n29497) );
  sky130_fd_sc_hd__and3_1 U19947 ( .A(n24535), .B(n24537), .C(n29550), .X(
        n29498) );
  sky130_fd_sc_hd__nand2_1 U19965 ( .A(n29498), .B(n24540), .Y(n12435) );
  sky130_fd_sc_hd__nand2b_1 U19981 ( .A_N(n24737), .B(n12123), .Y(n12151) );
  sky130_fd_sc_hd__and2_4 U20015 ( .A(n24210), .B(n29063), .X(n29499) );
  sky130_fd_sc_hd__and4_1 U20055 ( .A(n15283), .B(n15280), .C(n15282), .D(
        n15281), .X(n29500) );
  sky130_fd_sc_hd__and2_4 U20091 ( .A(n24210), .B(n29034), .X(n29501) );
  sky130_fd_sc_hd__clkinv_1 U20134 ( .A(n29033), .Y(n29559) );
  sky130_fd_sc_hd__and2_2 U20135 ( .A(n20720), .B(n20722), .X(n29502) );
  sky130_fd_sc_hd__nand2_1 U20138 ( .A(n11317), .B(n11314), .Y(n29530) );
  sky130_fd_sc_hd__inv_2 U20153 ( .A(n29530), .Y(n29529) );
  sky130_fd_sc_hd__clkinv_1 U20195 ( .A(j202_soc_core_j22_cpu_regop_Rn__0_), 
        .Y(n10964) );
  sky130_fd_sc_hd__clkinv_1 U20215 ( .A(n12656), .Y(n29524) );
  sky130_fd_sc_hd__and2_0 U20417 ( .A(n16155), .B(n16156), .X(n29503) );
  sky130_fd_sc_hd__and2_0 U20428 ( .A(n14848), .B(n12197), .X(n29504) );
  sky130_fd_sc_hd__a21boi_2 U20479 ( .A1(n19423), .A2(n19425), .B1_N(n19424), 
        .Y(n21824) );
  sky130_fd_sc_hd__inv_1 U20513 ( .A(n11036), .Y(n11038) );
  sky130_fd_sc_hd__nor2_2 U20534 ( .A(n12042), .B(n29066), .Y(n29505) );
  sky130_fd_sc_hd__nor2_2 U20606 ( .A(n12042), .B(n29066), .Y(n29506) );
  sky130_fd_sc_hd__nor2_2 U20661 ( .A(n12042), .B(n29066), .Y(n17160) );
  sky130_fd_sc_hd__nor2_4 U20712 ( .A(n11129), .B(n17143), .Y(n29066) );
  sky130_fd_sc_hd__nand2_1 U20871 ( .A(n12122), .B(n27823), .Y(n25107) );
  sky130_fd_sc_hd__inv_2 U21116 ( .A(n12122), .Y(n12627) );
  sky130_fd_sc_hd__nand2_2 U21263 ( .A(n17145), .B(n12416), .Y(n12122) );
  sky130_fd_sc_hd__bufinv_8 U21376 ( .A(n12416), .Y(n24225) );
  sky130_fd_sc_hd__and4bb_1 U21598 ( .C(n17150), .D(n21026), .A_N(n28920), 
        .B_N(n28919), .X(n17153) );
  sky130_fd_sc_hd__clkinv_1 U21627 ( .A(n12626), .Y(n17131) );
  sky130_fd_sc_hd__inv_2 U21649 ( .A(n29064), .Y(n29508) );
  sky130_fd_sc_hd__inv_1 U21883 ( .A(n27429), .Y(n26792) );
  sky130_fd_sc_hd__inv_1 U21924 ( .A(n12416), .Y(n24210) );
  sky130_fd_sc_hd__inv_1 U21926 ( .A(n12416), .Y(n27824) );
  sky130_fd_sc_hd__nor2_2 U21930 ( .A(n13497), .B(n13496), .Y(n21592) );
  sky130_fd_sc_hd__nand3_2 U22092 ( .A(n13487), .B(n13486), .C(n13371), .Y(
        n13496) );
  sky130_fd_sc_hd__inv_1 U22096 ( .A(n13487), .Y(n13499) );
  sky130_fd_sc_hd__bufinv_8 U22123 ( .A(n29249), .Y(n29509) );
  sky130_fd_sc_hd__bufinv_8 U22138 ( .A(n29249), .Y(n29510) );
  sky130_fd_sc_hd__bufinv_8 U22141 ( .A(n29249), .Y(n29511) );
  sky130_fd_sc_hd__bufinv_8 U22352 ( .A(n29249), .Y(n29512) );
  sky130_fd_sc_hd__buf_2 U22385 ( .A(n29070), .X(n11767) );
  sky130_fd_sc_hd__nand2_2 U22391 ( .A(n17107), .B(n13314), .Y(n29513) );
  sky130_fd_sc_hd__nand2_1 U22394 ( .A(n17107), .B(n13314), .Y(n26525) );
  sky130_fd_sc_hd__clkinv_1 U22399 ( .A(n28963), .Y(n11107) );
  sky130_fd_sc_hd__nand3_2 U22418 ( .A(n13053), .B(n12448), .C(n12646), .Y(
        n11650) );
  sky130_fd_sc_hd__nand3_2 U22443 ( .A(n11656), .B(n12062), .C(n29576), .Y(
        n23967) );
  sky130_fd_sc_hd__and2_1 U22514 ( .A(n12064), .B(n12060), .X(n11078) );
  sky130_fd_sc_hd__inv_1 U22528 ( .A(n26311), .Y(n23727) );
  sky130_fd_sc_hd__buf_1 U22589 ( .A(n24420), .X(n29514) );
  sky130_fd_sc_hd__o21a_2 U22753 ( .A1(n24297), .A2(n13045), .B1(n27949), .X(
        n29322) );
  sky130_fd_sc_hd__nand2_1 U22755 ( .A(n23603), .B(n27260), .Y(n23161) );
  sky130_fd_sc_hd__nand2_1 U22766 ( .A(n23603), .B(n27556), .Y(n23150) );
  sky130_fd_sc_hd__and2_1 U22781 ( .A(n23603), .B(n29071), .X(n11042) );
  sky130_fd_sc_hd__nor2_1 U22821 ( .A(n21023), .B(n28919), .Y(n29515) );
  sky130_fd_sc_hd__clkinv_4 U22943 ( .A(n25878), .Y(n25853) );
  sky130_fd_sc_hd__nand2_1 U22958 ( .A(n23045), .B(n23001), .Y(n23758) );
  sky130_fd_sc_hd__buf_6 U23026 ( .A(n12193), .X(n29283) );
  sky130_fd_sc_hd__nand3_1 U23096 ( .A(n27558), .B(n23144), .C(n12021), .Y(
        n23145) );
  sky130_fd_sc_hd__inv_1 U23106 ( .A(n11390), .Y(n11717) );
  sky130_fd_sc_hd__nand2_2 U23132 ( .A(j202_soc_core_memory0_ram_dout0[188]), 
        .B(n21590), .Y(n16633) );
  sky130_fd_sc_hd__nor2_2 U23305 ( .A(n11767), .B(n12012), .Y(n13056) );
  sky130_fd_sc_hd__inv_1 U23610 ( .A(n24455), .Y(n27924) );
  sky130_fd_sc_hd__nor2_1 U23617 ( .A(n12023), .B(n27174), .Y(n23611) );
  sky130_fd_sc_hd__nor2_1 U23626 ( .A(n12712), .B(n24092), .Y(n29516) );
  sky130_fd_sc_hd__nor2_1 U23667 ( .A(n12712), .B(n24092), .Y(n24656) );
  sky130_fd_sc_hd__buf_1 U23673 ( .A(n11135), .X(n29517) );
  sky130_fd_sc_hd__nand2_1 U23700 ( .A(n20146), .B(n20145), .Y(n12024) );
  sky130_fd_sc_hd__nand2_1 U23743 ( .A(n11393), .B(n29503), .Y(n29518) );
  sky130_fd_sc_hd__nand2_1 U23775 ( .A(n12743), .B(n22581), .Y(n11393) );
  sky130_fd_sc_hd__nand2_1 U23849 ( .A(n11393), .B(n29503), .Y(n17146) );
  sky130_fd_sc_hd__nand2_1 U23907 ( .A(n12884), .B(n29534), .Y(n29519) );
  sky130_fd_sc_hd__buf_6 U23908 ( .A(n12193), .X(n29284) );
  sky130_fd_sc_hd__nand3_1 U23958 ( .A(n27684), .B(n11996), .C(n13152), .Y(
        n24705) );
  sky130_fd_sc_hd__nor2_2 U23965 ( .A(n23148), .B(n12502), .Y(n27684) );
  sky130_fd_sc_hd__nand3_1 U23987 ( .A(n29585), .B(n22274), .C(n12462), .Y(
        n23140) );
  sky130_fd_sc_hd__nand3_1 U24078 ( .A(n22274), .B(n12735), .C(n12462), .Y(
        n12714) );
  sky130_fd_sc_hd__nand2_1 U24100 ( .A(n22274), .B(n12735), .Y(n23157) );
  sky130_fd_sc_hd__nor2_1 U24149 ( .A(n11802), .B(n12128), .Y(n29520) );
  sky130_fd_sc_hd__nor2_1 U24281 ( .A(n11802), .B(n12128), .Y(n12386) );
  sky130_fd_sc_hd__nand2_2 U24579 ( .A(n22827), .B(n22826), .Y(n11686) );
  sky130_fd_sc_hd__bufinv_8 U24605 ( .A(n29249), .Y(n12520) );
  sky130_fd_sc_hd__nand2_1 U24721 ( .A(n26315), .B(n26543), .Y(n27388) );
  sky130_fd_sc_hd__nor2_1 U24724 ( .A(n20715), .B(n20716), .Y(n29521) );
  sky130_fd_sc_hd__nor2_1 U24813 ( .A(n10975), .B(n12501), .Y(n29522) );
  sky130_fd_sc_hd__nand2_2 U24896 ( .A(n11873), .B(n10970), .Y(n23165) );
  sky130_fd_sc_hd__nand3_4 U24958 ( .A(n16664), .B(n16663), .C(n16662), .Y(
        n24123) );
  sky130_fd_sc_hd__a22oi_2 U25026 ( .A1(n21676), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[27]), .B1(n17099), .B2(
        n17098), .Y(n17104) );
  sky130_fd_sc_hd__nand3_2 U25073 ( .A(n11316), .B(n11066), .C(n11052), .Y(
        n20715) );
  sky130_fd_sc_hd__nand2_2 U25107 ( .A(n12656), .B(n28972), .Y(n23148) );
  sky130_fd_sc_hd__clkbuf_1 U25139 ( .A(n11875), .X(n29523) );
  sky130_fd_sc_hd__nand2_1 U25231 ( .A(n27776), .B(n27779), .Y(n11875) );
  sky130_fd_sc_hd__clkbuf_2 U25255 ( .A(n12743), .X(n11669) );
  sky130_fd_sc_hd__nand2_1 U25333 ( .A(n11669), .B(n22714), .Y(n12989) );
  sky130_fd_sc_hd__nand2_1 U25334 ( .A(n24417), .B(n24257), .Y(n24105) );
  sky130_fd_sc_hd__nand2b_1 U25361 ( .A_N(n27566), .B(n27298), .Y(n12476) );
  sky130_fd_sc_hd__clkbuf_1 U25566 ( .A(n27878), .X(n12655) );
  sky130_fd_sc_hd__inv_2 U25619 ( .A(n28957), .Y(n17152) );
  sky130_fd_sc_hd__clkinv_2 U25672 ( .A(n22019), .Y(n12656) );
  sky130_fd_sc_hd__nor2_2 U25707 ( .A(n27556), .B(n12512), .Y(n11848) );
  sky130_fd_sc_hd__inv_1 U25770 ( .A(n21022), .Y(n22672) );
  sky130_fd_sc_hd__nand2_2 U25778 ( .A(n12502), .B(n11107), .Y(n11845) );
  sky130_fd_sc_hd__nand2_1 U25857 ( .A(n12595), .B(n13152), .Y(n13269) );
  sky130_fd_sc_hd__nand3_1 U25864 ( .A(n23153), .B(n23152), .C(n23187), .Y(
        n23585) );
  sky130_fd_sc_hd__inv_1 U25920 ( .A(n12005), .Y(n22023) );
  sky130_fd_sc_hd__nand2_1 U25930 ( .A(n22020), .B(n12595), .Y(n27780) );
  sky130_fd_sc_hd__inv_2 U25946 ( .A(n11997), .Y(n11996) );
  sky130_fd_sc_hd__nand3_1 U26191 ( .A(n12734), .B(n12716), .C(n21166), .Y(
        n28963) );
  sky130_fd_sc_hd__nand2_2 U26284 ( .A(n21164), .B(n21165), .Y(n26538) );
  sky130_fd_sc_hd__inv_2 U26353 ( .A(n12010), .Y(n24417) );
  sky130_fd_sc_hd__nand3_4 U26367 ( .A(n13053), .B(n12646), .C(n12448), .Y(
        n12745) );
  sky130_fd_sc_hd__nand2_1 U26370 ( .A(n12088), .B(n12087), .Y(n21165) );
  sky130_fd_sc_hd__nor2_1 U26416 ( .A(n27790), .B(n23165), .Y(n24262) );
  sky130_fd_sc_hd__nand2_1 U26476 ( .A(n21165), .B(n12281), .Y(n12716) );
  sky130_fd_sc_hd__bufinv_8 U26735 ( .A(n29249), .Y(n12521) );
  sky130_fd_sc_hd__bufinv_8 U26781 ( .A(n29249), .Y(n12518) );
  sky130_fd_sc_hd__inv_8 U26794 ( .A(n23816), .Y(n29527) );
  sky130_fd_sc_hd__bufinv_8 U26968 ( .A(n23816), .Y(n29525) );
  sky130_fd_sc_hd__bufinv_8 U27020 ( .A(n23816), .Y(n29526) );
  sky130_fd_sc_hd__nand2_4 U27021 ( .A(n11127), .B(n29035), .Y(n23816) );
  sky130_fd_sc_hd__inv_4 U27060 ( .A(n12538), .Y(n11012) );
  sky130_fd_sc_hd__inv_16 U27074 ( .A(n12538), .Y(n11119) );
  sky130_fd_sc_hd__inv_16 U27131 ( .A(n12538), .Y(n11013) );
  sky130_fd_sc_hd__inv_4 U27149 ( .A(n29249), .Y(n29528) );
  sky130_fd_sc_hd__buf_4 U27212 ( .A(n10951), .X(n12408) );
  sky130_fd_sc_hd__clkinv_8 U27285 ( .A(n10940), .Y(n10951) );
  sky130_fd_sc_hd__buf_2 U27327 ( .A(n12692), .X(n29532) );
  sky130_fd_sc_hd__nand2_1 U27331 ( .A(n24310), .B(n12475), .Y(n24264) );
  sky130_fd_sc_hd__nand4_1 U27434 ( .A(n11921), .B(n11922), .C(n11923), .D(
        n11924), .Y(n11928) );
  sky130_fd_sc_hd__inv_2 U27451 ( .A(n24712), .Y(n22766) );
  sky130_fd_sc_hd__nand3_2 U27464 ( .A(n11662), .B(n22745), .C(n22746), .Y(
        n24712) );
  sky130_fd_sc_hd__nand4_1 U27552 ( .A(n19927), .B(n19929), .C(n10933), .D(
        n19930), .Y(n13158) );
  sky130_fd_sc_hd__nand2_1 U27554 ( .A(n12001), .B(n29520), .Y(n29531) );
  sky130_fd_sc_hd__nor2_1 U27616 ( .A(n10938), .B(n12006), .Y(n12001) );
  sky130_fd_sc_hd__nand2_1 U27630 ( .A(n27878), .B(n23950), .Y(n11815) );
  sky130_fd_sc_hd__nand3_2 U27725 ( .A(n13115), .B(n11392), .C(n25048), .Y(
        n27878) );
  sky130_fd_sc_hd__nand2b_1 U27733 ( .A_N(n23959), .B(n27551), .Y(n11656) );
  sky130_fd_sc_hd__nor2_4 U27764 ( .A(n13180), .B(n29070), .Y(n23603) );
  sky130_fd_sc_hd__nand3_4 U27809 ( .A(n29529), .B(n20721), .C(n29502), .Y(
        n29070) );
  sky130_fd_sc_hd__nand3_1 U27811 ( .A(n29529), .B(n29502), .C(n20721), .Y(
        n11763) );
  sky130_fd_sc_hd__nand2_1 U27910 ( .A(n29531), .B(n23968), .Y(n12622) );
  sky130_fd_sc_hd__nand2_1 U27928 ( .A(n29533), .B(n11297), .Y(n20710) );
  sky130_fd_sc_hd__nor2_1 U27932 ( .A(n11301), .B(n11302), .Y(n29533) );
  sky130_fd_sc_hd__nor2_1 U28074 ( .A(n13241), .B(n13242), .Y(n20964) );
  sky130_fd_sc_hd__buf_2 U28118 ( .A(n11698), .X(n29534) );
  sky130_fd_sc_hd__nand4_1 U28122 ( .A(n29493), .B(n13595), .C(n13593), .D(
        n13594), .Y(n11535) );
  sky130_fd_sc_hd__nand2_1 U28131 ( .A(n11568), .B(n29497), .Y(n11566) );
  sky130_fd_sc_hd__nor2_2 U28156 ( .A(n17919), .B(n17918), .Y(n22759) );
  sky130_fd_sc_hd__o21ai_2 U28171 ( .A1(n24691), .A2(n29535), .B1(n24689), .Y(
        n24686) );
  sky130_fd_sc_hd__nor2_1 U28256 ( .A(n29536), .B(n11346), .Y(n11345) );
  sky130_fd_sc_hd__nand4_1 U28260 ( .A(n29541), .B(n11352), .C(n11357), .D(
        n11353), .Y(n29536) );
  sky130_fd_sc_hd__nand2_1 U28325 ( .A(n29537), .B(n12974), .Y(n21007) );
  sky130_fd_sc_hd__nor2_1 U28374 ( .A(n11522), .B(n11527), .Y(n29537) );
  sky130_fd_sc_hd__nand3_1 U28444 ( .A(n29539), .B(n20708), .C(n29538), .Y(
        n11644) );
  sky130_fd_sc_hd__nand2_1 U28584 ( .A(j202_soc_core_memory0_ram_dout0[321]), 
        .B(n21593), .Y(n29539) );
  sky130_fd_sc_hd__nand3_1 U28615 ( .A(n12017), .B(n12018), .C(n12395), .Y(
        n12020) );
  sky130_fd_sc_hd__nor2_1 U28618 ( .A(n29540), .B(n11987), .Y(n12000) );
  sky130_fd_sc_hd__nand4_1 U28737 ( .A(n21145), .B(n21031), .C(n21034), .D(
        n11989), .Y(n29540) );
  sky130_fd_sc_hd__a21oi_2 U28824 ( .A1(n24682), .A2(n26720), .B1(n24681), .Y(
        n24689) );
  sky130_fd_sc_hd__nand2_1 U28848 ( .A(j202_soc_core_memory0_ram_dout0[368]), 
        .B(n21596), .Y(n29541) );
  sky130_fd_sc_hd__nor2_1 U28887 ( .A(n29542), .B(n13030), .Y(n12770) );
  sky130_fd_sc_hd__nand4_1 U28907 ( .A(n13219), .B(n13218), .C(n13216), .D(
        n13215), .Y(n29542) );
  sky130_fd_sc_hd__nand3_2 U29043 ( .A(n12150), .B(n10973), .C(n23143), .Y(
        n23163) );
  sky130_fd_sc_hd__nand3_2 U29080 ( .A(n11322), .B(n11318), .C(n29543), .Y(
        n22277) );
  sky130_fd_sc_hd__nand2_1 U29085 ( .A(n11320), .B(n11321), .Y(n29543) );
  sky130_fd_sc_hd__nand3_2 U29128 ( .A(n11134), .B(n11392), .C(n29544), .Y(
        n27261) );
  sky130_fd_sc_hd__inv_2 U29181 ( .A(n29545), .Y(n29544) );
  sky130_fd_sc_hd__nand2_1 U29262 ( .A(n27523), .B(n25048), .Y(n29545) );
  sky130_fd_sc_hd__nand3_1 U29357 ( .A(n12716), .B(n12734), .C(n21166), .Y(
        n11997) );
  sky130_fd_sc_hd__nand2_1 U29408 ( .A(n11965), .B(n23803), .Y(n11817) );
  sky130_fd_sc_hd__nand2_2 U29425 ( .A(n11818), .B(n12641), .Y(n11965) );
  sky130_fd_sc_hd__nand2_1 U29426 ( .A(n12001), .B(n12386), .Y(n11964) );
  sky130_fd_sc_hd__nor2_1 U29454 ( .A(n12480), .B(n12558), .Y(n12557) );
  sky130_fd_sc_hd__buf_2 U29455 ( .A(n27790), .X(n29548) );
  sky130_fd_sc_hd__nand2_1 U29468 ( .A(n28974), .B(n24225), .Y(n23973) );
  sky130_fd_sc_hd__nand3_2 U29491 ( .A(n22935), .B(n22934), .C(n22933), .Y(
        n28974) );
  sky130_fd_sc_hd__and2_0 U29506 ( .A(n24536), .B(n24539), .X(n29550) );
  sky130_fd_sc_hd__nor2_1 U29513 ( .A(n29551), .B(n12975), .Y(n12974) );
  sky130_fd_sc_hd__nand4_1 U29515 ( .A(n20565), .B(n20564), .C(n20563), .D(
        n12977), .Y(n29551) );
  sky130_fd_sc_hd__a21boi_1 U29516 ( .A1(n17354), .A2(n17355), .B1_N(n17353), 
        .Y(n12415) );
  sky130_fd_sc_hd__nor2_2 U29518 ( .A(n21909), .B(n22747), .Y(n18816) );
  sky130_fd_sc_hd__nor2_2 U29519 ( .A(n18814), .B(n18813), .Y(n22747) );
  sky130_fd_sc_hd__nand2_1 U29538 ( .A(n29553), .B(n29552), .Y(n18460) );
  sky130_fd_sc_hd__nand2_1 U29555 ( .A(n29556), .B(n18432), .Y(n29552) );
  sky130_fd_sc_hd__xor2_1 U29592 ( .A(n18430), .B(n29554), .X(n18418) );
  sky130_fd_sc_hd__xnor2_1 U29612 ( .A(n29556), .B(n29555), .Y(n29554) );
  sky130_fd_sc_hd__nand2_1 U29621 ( .A(n18352), .B(n22071), .Y(n29556) );
  sky130_fd_sc_hd__nand2_4 U29658 ( .A(n11717), .B(n20977), .Y(n12502) );
  sky130_fd_sc_hd__nand4_1 U29672 ( .A(n13100), .B(n29561), .C(n13101), .D(
        n29557), .Y(n13098) );
  sky130_fd_sc_hd__nand2_1 U29721 ( .A(j202_soc_core_memory0_ram_dout0[84]), 
        .B(n21734), .Y(n29557) );
  sky130_fd_sc_hd__nand2_1 U29727 ( .A(n29558), .B(n24709), .Y(n10502) );
  sky130_fd_sc_hd__nand2_1 U29732 ( .A(n24707), .B(n27980), .Y(n29558) );
  sky130_fd_sc_hd__nor2b_1 U29869 ( .B_N(n29067), .A(n29559), .Y(n12264) );
  sky130_fd_sc_hd__nand2_1 U29878 ( .A(n12640), .B(n23209), .Y(n27888) );
  sky130_fd_sc_hd__nand2_1 U29909 ( .A(n12883), .B(n24414), .Y(n12640) );
  sky130_fd_sc_hd__nand4_1 U29910 ( .A(n28918), .B(n29518), .C(n27602), .D(
        n24123), .Y(n29560) );
  sky130_fd_sc_hd__nand2_1 U29950 ( .A(j202_soc_core_memory0_ram_dout0[20]), 
        .B(n21733), .Y(n29561) );
  sky130_fd_sc_hd__nand2_1 U29961 ( .A(n23963), .B(n23965), .Y(n12128) );
  sky130_fd_sc_hd__inv_2 U29981 ( .A(n24161), .Y(n24163) );
  sky130_fd_sc_hd__o21a_1 U30056 ( .A1(n22759), .A2(n22762), .B1(n22760), .X(
        n29562) );
  sky130_fd_sc_hd__nor2_4 U30061 ( .A(n13702), .B(n19053), .Y(n29563) );
  sky130_fd_sc_hd__nor2_4 U30065 ( .A(n13638), .B(n23445), .Y(n29564) );
  sky130_fd_sc_hd__nor2_2 U30081 ( .A(n12137), .B(n11994), .Y(n13387) );
  sky130_fd_sc_hd__a21oi_4 U30111 ( .A1(n25744), .A2(n26802), .B1(n12591), .Y(
        n29565) );
  sky130_fd_sc_hd__nand2_4 U30115 ( .A(n24225), .B(n29356), .Y(n23581) );
  sky130_fd_sc_hd__nor2_4 U30120 ( .A(n13658), .B(n13675), .Y(n29566) );
  sky130_fd_sc_hd__nor2_4 U30126 ( .A(n13702), .B(n19050), .Y(n29567) );
  sky130_fd_sc_hd__or2_0 U30167 ( .A(n13638), .B(n23513), .X(n12169) );
  sky130_fd_sc_hd__or2_1 U30169 ( .A(n13678), .B(n13687), .X(n29568) );
  sky130_fd_sc_hd__and2_4 U30226 ( .A(n24350), .B(n24265), .X(n29569) );
  sky130_fd_sc_hd__and2_4 U30238 ( .A(n29006), .B(n24225), .X(n29570) );
  sky130_fd_sc_hd__and2_4 U30253 ( .A(n28987), .B(n11127), .X(n29571) );
  sky130_fd_sc_hd__and2_0 U30268 ( .A(n20714), .B(n21776), .X(n29572) );
  sky130_fd_sc_hd__clkinv_1 U30285 ( .A(n29077), .Y(n27553) );
  sky130_fd_sc_hd__or2_0 U30308 ( .A(n17772), .B(n18353), .X(n29573) );
  sky130_fd_sc_hd__clkinv_1 U30325 ( .A(n17302), .Y(n17055) );
  sky130_fd_sc_hd__or2_0 U30359 ( .A(n22763), .B(n22759), .X(n29574) );
  sky130_fd_sc_hd__inv_2 U30418 ( .A(n11661), .Y(n12740) );
  sky130_fd_sc_hd__inv_2 U30454 ( .A(n11692), .Y(n12743) );
  sky130_fd_sc_hd__and2_1 U30509 ( .A(n12899), .B(n29033), .X(n29575) );
  sky130_fd_sc_hd__and2_0 U30553 ( .A(n23960), .B(n23958), .X(n29576) );
  sky130_fd_sc_hd__inv_1 U30565 ( .A(n13686), .Y(n23118) );
  sky130_fd_sc_hd__or2_0 U30674 ( .A(n23206), .B(n24325), .X(n29577) );
  sky130_fd_sc_hd__and2_1 U30757 ( .A(n12899), .B(n27621), .X(n29578) );
  sky130_fd_sc_hd__and2_1 U30763 ( .A(n12899), .B(n29010), .X(n29579) );
  sky130_fd_sc_hd__and2_1 U30777 ( .A(n12899), .B(n29012), .X(n29580) );
  sky130_fd_sc_hd__and2_1 U30785 ( .A(n12899), .B(n29061), .X(n29581) );
  sky130_fd_sc_hd__and2_1 U30793 ( .A(n12899), .B(n29034), .X(n29582) );
  sky130_fd_sc_hd__and2_1 U30800 ( .A(n12899), .B(n29013), .X(n29583) );
  sky130_fd_sc_hd__and2_1 U30842 ( .A(n12899), .B(n29011), .X(n29584) );
  sky130_fd_sc_hd__inv_1 U30844 ( .A(n11867), .Y(n24385) );
  sky130_fd_sc_hd__and2_1 U30853 ( .A(n10974), .B(n13103), .X(n29585) );
  sky130_fd_sc_hd__and2_0 U30863 ( .A(n24134), .B(n21434), .X(n29587) );
  sky130_fd_sc_hd__and2_0 U30866 ( .A(n29065), .B(n24567), .X(n29588) );
  sky130_fd_sc_hd__or2_0 U30876 ( .A(n24562), .B(n12457), .X(n29589) );
  sky130_fd_sc_hd__inv_1 U30888 ( .A(n27791), .Y(n23608) );
  sky130_fd_sc_hd__clkinv_1 U30898 ( .A(n10939), .Y(n21026) );
  sky130_fd_sc_hd__clkinv_1 U30963 ( .A(n26443), .Y(n26352) );
  sky130_fd_sc_hd__inv_2 U30992 ( .A(n27409), .Y(n11977) );
  sky130_fd_sc_hd__clkinv_1 U30998 ( .A(n26085), .Y(n26422) );
  sky130_fd_sc_hd__clkinv_2 U31040 ( .A(n28590), .Y(n29592) );
  sky130_fd_sc_hd__clkinv_2 U31044 ( .A(n28590), .Y(n29593) );
  sky130_fd_sc_hd__clkinv_1 U31062 ( .A(n28590), .Y(n29591) );
  sky130_fd_sc_hd__clkinv_2 U31123 ( .A(n28590), .Y(n29594) );
endmodule

