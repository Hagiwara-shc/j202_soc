magic
tech sky130A
magscale 1 2
timestamp 1670651684
<< metal1 >>
rect 186498 702992 186504 703044
rect 186556 703032 186562 703044
rect 188430 703032 188436 703044
rect 186556 703004 188436 703032
rect 186556 702992 186562 703004
rect 188430 702992 188436 703004
rect 188488 702992 188494 703044
rect 235166 702992 235172 703044
rect 235224 703032 235230 703044
rect 236178 703032 236184 703044
rect 235224 703004 236184 703032
rect 235224 702992 235230 703004
rect 236178 702992 236184 703004
rect 236236 702992 236242 703044
rect 522758 702992 522764 703044
rect 522816 703032 522822 703044
rect 527082 703032 527088 703044
rect 522816 703004 527088 703032
rect 522816 702992 522822 703004
rect 527082 702992 527088 703004
rect 527140 702992 527146 703044
rect 570506 702992 570512 703044
rect 570564 703032 570570 703044
rect 575842 703032 575848 703044
rect 570564 703004 575848 703032
rect 570564 702992 570570 703004
rect 575842 702992 575848 703004
rect 575900 702992 575906 703044
rect 490926 702720 490932 702772
rect 490984 702760 490990 702772
rect 494790 702760 494796 702772
rect 490984 702732 494796 702760
rect 490984 702720 490990 702732
rect 494790 702720 494796 702732
rect 494848 702720 494854 702772
rect 538674 702720 538680 702772
rect 538732 702760 538738 702772
rect 543458 702760 543464 702772
rect 538732 702732 543464 702760
rect 538732 702720 538738 702732
rect 543458 702720 543464 702732
rect 543516 702720 543522 702772
rect 24302 702448 24308 702500
rect 24360 702488 24366 702500
rect 29270 702488 29276 702500
rect 24360 702460 29276 702488
rect 24360 702448 24366 702460
rect 29270 702448 29276 702460
rect 29328 702448 29334 702500
rect 218974 702448 218980 702500
rect 219032 702488 219038 702500
rect 220262 702488 220268 702500
rect 219032 702460 220268 702488
rect 219032 702448 219038 702460
rect 220262 702448 220268 702460
rect 220320 702448 220326 702500
rect 459094 702448 459100 702500
rect 459152 702488 459158 702500
rect 462314 702488 462320 702500
rect 459152 702460 462320 702488
rect 459152 702448 459158 702460
rect 462314 702448 462320 702460
rect 462372 702448 462378 702500
rect 506842 702448 506848 702500
rect 506900 702488 506906 702500
rect 510982 702488 510988 702500
rect 506900 702460 510988 702488
rect 506900 702448 506906 702460
rect 510982 702448 510988 702460
rect 511040 702448 511046 702500
rect 554590 702448 554596 702500
rect 554648 702488 554654 702500
rect 559650 702488 559656 702500
rect 554648 702460 559656 702488
rect 554648 702448 554654 702460
rect 559650 702448 559656 702460
rect 559708 702448 559714 702500
rect 8110 700952 8116 701004
rect 8168 700992 8174 701004
rect 13078 700992 13084 701004
rect 8168 700964 13084 700992
rect 8168 700952 8174 700964
rect 13078 700952 13084 700964
rect 13136 700952 13142 701004
rect 40494 700952 40500 701004
rect 40552 700992 40558 701004
rect 44910 700992 44916 701004
rect 40552 700964 44916 700992
rect 40552 700952 40558 700964
rect 44910 700952 44916 700964
rect 44968 700952 44974 701004
rect 56778 700952 56784 701004
rect 56836 700992 56842 701004
rect 60734 700992 60740 701004
rect 56836 700964 60740 700992
rect 56836 700952 56842 700964
rect 60734 700952 60740 700964
rect 60792 700952 60798 701004
rect 72970 700952 72976 701004
rect 73028 700992 73034 701004
rect 76742 700992 76748 701004
rect 73028 700964 76748 700992
rect 73028 700952 73034 700964
rect 76742 700952 76748 700964
rect 76800 700952 76806 701004
rect 89162 700952 89168 701004
rect 89220 700992 89226 701004
rect 92566 700992 92572 701004
rect 89220 700964 92572 700992
rect 89220 700952 89226 700964
rect 92566 700952 92572 700964
rect 92624 700952 92630 701004
rect 105446 700952 105452 701004
rect 105504 700992 105510 701004
rect 108574 700992 108580 701004
rect 105504 700964 108580 700992
rect 105504 700952 105510 700964
rect 108574 700952 108580 700964
rect 108632 700952 108638 701004
rect 121638 700952 121644 701004
rect 121696 700992 121702 701004
rect 124398 700992 124404 701004
rect 121696 700964 124404 700992
rect 121696 700952 121702 700964
rect 124398 700952 124404 700964
rect 124456 700952 124462 701004
rect 137830 700952 137836 701004
rect 137888 700992 137894 701004
rect 140406 700992 140412 701004
rect 137888 700964 140412 700992
rect 137888 700952 137894 700964
rect 140406 700952 140412 700964
rect 140464 700952 140470 701004
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 156230 700992 156236 701004
rect 154172 700964 156236 700992
rect 154172 700952 154178 700964
rect 156230 700952 156236 700964
rect 156288 700952 156294 701004
rect 170306 700952 170312 701004
rect 170364 700992 170370 701004
rect 172422 700992 172428 701004
rect 170364 700964 172428 700992
rect 170364 700952 170370 700964
rect 172422 700952 172428 700964
rect 172480 700952 172486 701004
rect 202782 700952 202788 701004
rect 202840 700992 202846 701004
rect 204254 700992 204260 701004
rect 202840 700964 204260 700992
rect 202840 700952 202846 700964
rect 204254 700952 204260 700964
rect 204312 700952 204318 701004
rect 348050 700952 348056 701004
rect 348108 700992 348114 701004
rect 348786 700992 348792 701004
rect 348108 700964 348792 700992
rect 348108 700952 348114 700964
rect 348786 700952 348792 700964
rect 348844 700952 348850 701004
rect 363874 700952 363880 701004
rect 363932 700992 363938 701004
rect 364978 700992 364984 701004
rect 363932 700964 364984 700992
rect 363932 700952 363938 700964
rect 364978 700952 364984 700964
rect 365036 700952 365042 701004
rect 379330 700952 379336 701004
rect 379388 700992 379394 701004
rect 381170 700992 381176 701004
rect 379388 700964 381176 700992
rect 379388 700952 379394 700964
rect 381170 700952 381176 700964
rect 381228 700952 381234 701004
rect 395706 700952 395712 701004
rect 395764 700992 395770 701004
rect 397454 700992 397460 701004
rect 395764 700964 397460 700992
rect 395764 700952 395770 700964
rect 397454 700952 397460 700964
rect 397512 700952 397518 701004
rect 411714 700952 411720 701004
rect 411772 700992 411778 701004
rect 413646 700992 413652 701004
rect 411772 700964 413652 700992
rect 411772 700952 411778 700964
rect 413646 700952 413652 700964
rect 413704 700952 413710 701004
rect 427538 700952 427544 701004
rect 427596 700992 427602 701004
rect 429838 700992 429844 701004
rect 427596 700964 429844 700992
rect 427596 700952 427602 700964
rect 429838 700952 429844 700964
rect 429896 700952 429902 701004
rect 443546 700952 443552 701004
rect 443604 700992 443610 701004
rect 446122 700992 446128 701004
rect 443604 700964 446128 700992
rect 443604 700952 443610 700964
rect 446122 700952 446128 700964
rect 446180 700952 446186 701004
rect 475378 700952 475384 701004
rect 475436 700992 475442 701004
rect 478506 700992 478512 701004
rect 475436 700964 478512 700992
rect 475436 700952 475442 700964
rect 478506 700952 478512 700964
rect 478564 700952 478570 701004
rect 73522 3952 73528 4004
rect 73580 3992 73586 4004
rect 87966 3992 87972 4004
rect 73580 3964 87972 3992
rect 73580 3952 73586 3964
rect 87966 3952 87972 3964
rect 88024 3952 88030 4004
rect 64322 3884 64328 3936
rect 64380 3924 64386 3936
rect 79134 3924 79140 3936
rect 64380 3896 79140 3924
rect 64380 3884 64386 3896
rect 79134 3884 79140 3896
rect 79192 3884 79198 3936
rect 70118 3816 70124 3868
rect 70176 3856 70182 3868
rect 84654 3856 84660 3868
rect 70176 3828 84660 3856
rect 70176 3816 70182 3828
rect 84654 3816 84660 3828
rect 84712 3816 84718 3868
rect 99834 3816 99840 3868
rect 99892 3856 99898 3868
rect 112254 3856 112260 3868
rect 99892 3828 112260 3856
rect 99892 3816 99898 3828
rect 112254 3816 112260 3828
rect 112312 3816 112318 3868
rect 58802 3748 58808 3800
rect 58860 3788 58866 3800
rect 73614 3788 73620 3800
rect 58860 3760 73620 3788
rect 58860 3748 58866 3760
rect 73614 3748 73620 3760
rect 73672 3748 73678 3800
rect 77386 3748 77392 3800
rect 77444 3788 77450 3800
rect 91278 3788 91284 3800
rect 77444 3760 91284 3788
rect 77444 3748 77450 3760
rect 91278 3748 91284 3760
rect 91336 3748 91342 3800
rect 105722 3748 105728 3800
rect 105780 3788 105786 3800
rect 117774 3788 117780 3800
rect 105780 3760 117780 3788
rect 105780 3748 105786 3760
rect 117774 3748 117780 3760
rect 117832 3748 117838 3800
rect 125962 3748 125968 3800
rect 126020 3788 126026 3800
rect 136634 3788 136640 3800
rect 126020 3760 136640 3788
rect 126020 3748 126026 3760
rect 136634 3748 136640 3760
rect 136692 3748 136698 3800
rect 63218 3680 63224 3732
rect 63276 3720 63282 3732
rect 78030 3720 78036 3732
rect 63276 3692 78036 3720
rect 63276 3680 63282 3692
rect 78030 3680 78036 3692
rect 78088 3680 78094 3732
rect 83274 3680 83280 3732
rect 83332 3720 83338 3732
rect 96798 3720 96804 3732
rect 83332 3692 96804 3720
rect 83332 3680 83338 3692
rect 96798 3680 96804 3692
rect 96856 3680 96862 3732
rect 98914 3680 98920 3732
rect 98972 3720 98978 3732
rect 103422 3720 103428 3732
rect 98972 3692 103428 3720
rect 98972 3680 98978 3692
rect 103422 3680 103428 3692
rect 103480 3680 103486 3732
rect 118786 3680 118792 3732
rect 118844 3720 118850 3732
rect 129918 3720 129924 3732
rect 118844 3692 129924 3720
rect 118844 3680 118850 3692
rect 129918 3680 129924 3692
rect 129976 3680 129982 3732
rect 60826 3612 60832 3664
rect 60884 3652 60890 3664
rect 75822 3652 75828 3664
rect 60884 3624 75828 3652
rect 60884 3612 60890 3624
rect 75822 3612 75828 3624
rect 75880 3612 75886 3664
rect 79686 3612 79692 3664
rect 79744 3652 79750 3664
rect 93486 3652 93492 3664
rect 79744 3624 93492 3652
rect 79744 3612 79750 3624
rect 93486 3612 93492 3624
rect 93544 3612 93550 3664
rect 95142 3612 95148 3664
rect 95200 3652 95206 3664
rect 107838 3652 107844 3664
rect 95200 3624 107844 3652
rect 95200 3612 95206 3624
rect 107838 3612 107844 3624
rect 107896 3612 107902 3664
rect 117590 3612 117596 3664
rect 117648 3652 117654 3664
rect 128814 3652 128820 3664
rect 117648 3624 128820 3652
rect 117648 3612 117654 3624
rect 128814 3612 128820 3624
rect 128872 3612 128878 3664
rect 144730 3612 144736 3664
rect 144788 3652 144794 3664
rect 154206 3652 154212 3664
rect 144788 3624 154212 3652
rect 144788 3612 144794 3624
rect 154206 3612 154212 3624
rect 154264 3612 154270 3664
rect 56962 3544 56968 3596
rect 57020 3584 57026 3596
rect 72510 3584 72516 3596
rect 57020 3556 72516 3584
rect 57020 3544 57026 3556
rect 72510 3544 72516 3556
rect 72568 3544 72574 3596
rect 72602 3544 72608 3596
rect 72660 3584 72666 3596
rect 86862 3584 86868 3596
rect 72660 3556 86868 3584
rect 72660 3544 72666 3556
rect 86862 3544 86868 3556
rect 86920 3544 86926 3596
rect 89530 3544 89536 3596
rect 89588 3584 89594 3596
rect 102318 3584 102324 3596
rect 89588 3556 102324 3584
rect 89588 3544 89594 3556
rect 102318 3544 102324 3556
rect 102376 3544 102382 3596
rect 103330 3544 103336 3596
rect 103388 3584 103394 3596
rect 115566 3584 115572 3596
rect 103388 3556 115572 3584
rect 103388 3544 103394 3556
rect 115566 3544 115572 3556
rect 115624 3544 115630 3596
rect 120902 3544 120908 3596
rect 120960 3584 120966 3596
rect 132126 3584 132132 3596
rect 120960 3556 132132 3584
rect 120960 3544 120966 3556
rect 132126 3544 132132 3556
rect 132184 3544 132190 3596
rect 132954 3544 132960 3596
rect 133012 3584 133018 3596
rect 143166 3584 143172 3596
rect 133012 3556 143172 3584
rect 133012 3544 133018 3556
rect 143166 3544 143172 3556
rect 143224 3544 143230 3596
rect 148318 3544 148324 3596
rect 148376 3584 148382 3596
rect 157518 3584 157524 3596
rect 148376 3556 157524 3584
rect 148376 3544 148382 3556
rect 157518 3544 157524 3556
rect 157576 3544 157582 3596
rect 71314 3476 71320 3528
rect 71372 3516 71378 3528
rect 85758 3516 85764 3528
rect 71372 3488 85764 3516
rect 71372 3476 71378 3488
rect 85758 3476 85764 3488
rect 85816 3476 85822 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 111150 3516 111156 3528
rect 98696 3488 111156 3516
rect 98696 3476 98702 3488
rect 111150 3476 111156 3488
rect 111208 3476 111214 3528
rect 129366 3476 129372 3528
rect 129424 3516 129430 3528
rect 139854 3516 139860 3528
rect 129424 3488 139860 3516
rect 129424 3476 129430 3488
rect 139854 3476 139860 3488
rect 139912 3476 139918 3528
rect 142522 3476 142528 3528
rect 142580 3516 142586 3528
rect 151998 3516 152004 3528
rect 142580 3488 152004 3516
rect 142580 3476 142586 3488
rect 151998 3476 152004 3488
rect 152056 3476 152062 3528
rect 163682 3476 163688 3528
rect 163740 3516 163746 3528
rect 171870 3516 171876 3528
rect 163740 3488 171876 3516
rect 163740 3476 163746 3488
rect 171870 3476 171876 3488
rect 171928 3476 171934 3528
rect 59722 3408 59728 3460
rect 59780 3448 59786 3460
rect 74442 3448 74448 3460
rect 59780 3420 74448 3448
rect 59780 3408 59786 3420
rect 74442 3408 74448 3420
rect 74500 3408 74506 3460
rect 75362 3408 75368 3460
rect 75420 3448 75426 3460
rect 89070 3448 89076 3460
rect 75420 3420 89076 3448
rect 75420 3408 75426 3420
rect 89070 3408 89076 3420
rect 89128 3408 89134 3460
rect 93946 3408 93952 3460
rect 94004 3448 94010 3460
rect 100754 3448 100760 3460
rect 94004 3420 100760 3448
rect 94004 3408 94010 3420
rect 100754 3408 100760 3420
rect 100812 3408 100818 3460
rect 109034 3448 109040 3460
rect 100956 3420 109040 3448
rect 52546 3340 52552 3392
rect 52604 3380 52610 3392
rect 68094 3380 68100 3392
rect 52604 3352 68100 3380
rect 52604 3340 52610 3352
rect 68094 3340 68100 3352
rect 68152 3340 68158 3392
rect 68554 3340 68560 3392
rect 68612 3380 68618 3392
rect 82446 3380 82452 3392
rect 68612 3352 82452 3380
rect 68612 3340 68618 3352
rect 82446 3340 82452 3352
rect 82504 3340 82510 3392
rect 90082 3340 90088 3392
rect 90140 3380 90146 3392
rect 98914 3380 98920 3392
rect 90140 3352 98920 3380
rect 90140 3340 90146 3352
rect 98914 3340 98920 3352
rect 98972 3340 98978 3392
rect 48958 3272 48964 3324
rect 49016 3312 49022 3324
rect 49016 3284 60044 3312
rect 49016 3272 49022 3284
rect 40402 3204 40408 3256
rect 40460 3244 40466 3256
rect 57054 3244 57060 3256
rect 40460 3216 57060 3244
rect 40460 3204 40466 3216
rect 57054 3204 57060 3216
rect 57112 3204 57118 3256
rect 60016 3244 60044 3284
rect 62022 3272 62028 3324
rect 62080 3312 62086 3324
rect 76926 3312 76932 3324
rect 62080 3284 76932 3312
rect 62080 3272 62086 3284
rect 76926 3272 76932 3284
rect 76984 3272 76990 3324
rect 85666 3272 85672 3324
rect 85724 3312 85730 3324
rect 99006 3312 99012 3324
rect 85724 3284 99012 3312
rect 85724 3272 85730 3284
rect 99006 3272 99012 3284
rect 99064 3272 99070 3324
rect 64690 3244 64696 3256
rect 60016 3216 64696 3244
rect 64690 3204 64696 3216
rect 64748 3204 64754 3256
rect 66714 3204 66720 3256
rect 66772 3244 66778 3256
rect 66772 3216 74534 3244
rect 66772 3204 66778 3216
rect 51350 3136 51356 3188
rect 51408 3176 51414 3188
rect 66990 3176 66996 3188
rect 51408 3148 66996 3176
rect 51408 3136 51414 3148
rect 66990 3136 66996 3148
rect 67048 3136 67054 3188
rect 74506 3176 74534 3216
rect 80882 3204 80888 3256
rect 80940 3244 80946 3256
rect 94590 3244 94596 3256
rect 80940 3216 94596 3244
rect 80940 3204 80946 3216
rect 94590 3204 94596 3216
rect 94648 3204 94654 3256
rect 96246 3204 96252 3256
rect 96304 3244 96310 3256
rect 100956 3244 100984 3420
rect 109034 3408 109040 3420
rect 109092 3408 109098 3460
rect 116394 3408 116400 3460
rect 116452 3448 116458 3460
rect 127710 3448 127716 3460
rect 116452 3420 127716 3448
rect 116452 3408 116458 3420
rect 127710 3408 127716 3420
rect 127768 3408 127774 3460
rect 137462 3408 137468 3460
rect 137520 3448 137526 3460
rect 137520 3420 137784 3448
rect 137520 3408 137526 3420
rect 101030 3340 101036 3392
rect 101088 3380 101094 3392
rect 101088 3352 104296 3380
rect 101088 3340 101094 3352
rect 96304 3216 100984 3244
rect 104268 3244 104296 3352
rect 114002 3340 114008 3392
rect 114060 3380 114066 3392
rect 125594 3380 125600 3392
rect 114060 3352 125600 3380
rect 114060 3340 114066 3352
rect 125594 3340 125600 3352
rect 125652 3340 125658 3392
rect 127066 3340 127072 3392
rect 127124 3380 127130 3392
rect 137646 3380 137652 3392
rect 127124 3352 137652 3380
rect 127124 3340 127130 3352
rect 137646 3340 137652 3352
rect 137704 3340 137710 3392
rect 137756 3380 137784 3420
rect 153010 3408 153016 3460
rect 153068 3448 153074 3460
rect 161934 3448 161940 3460
rect 153068 3420 161940 3448
rect 153068 3408 153074 3420
rect 161934 3408 161940 3420
rect 161992 3408 161998 3460
rect 169570 3408 169576 3460
rect 169628 3448 169634 3460
rect 177390 3448 177396 3460
rect 169628 3420 177396 3448
rect 169628 3408 169634 3420
rect 177390 3408 177396 3420
rect 177448 3408 177454 3460
rect 183738 3408 183744 3460
rect 183796 3448 183802 3460
rect 190638 3448 190644 3460
rect 183796 3420 190644 3448
rect 183796 3408 183802 3420
rect 190638 3408 190644 3420
rect 190696 3408 190702 3460
rect 147674 3380 147680 3392
rect 137756 3352 147680 3380
rect 147674 3340 147680 3352
rect 147732 3340 147738 3392
rect 155402 3340 155408 3392
rect 155460 3380 155466 3392
rect 164234 3380 164240 3392
rect 155460 3352 164240 3380
rect 155460 3340 155466 3352
rect 164234 3340 164240 3352
rect 164292 3340 164298 3392
rect 167178 3340 167184 3392
rect 167236 3380 167242 3392
rect 175274 3380 175280 3392
rect 167236 3352 175280 3380
rect 167236 3340 167242 3352
rect 175274 3340 175280 3352
rect 175332 3340 175338 3392
rect 180242 3340 180248 3392
rect 180300 3380 180306 3392
rect 187326 3380 187332 3392
rect 180300 3352 187332 3380
rect 180300 3340 180306 3352
rect 187326 3340 187332 3352
rect 187384 3340 187390 3392
rect 109402 3272 109408 3324
rect 109460 3312 109466 3324
rect 121086 3312 121092 3324
rect 109460 3284 121092 3312
rect 109460 3272 109466 3284
rect 121086 3272 121092 3284
rect 121144 3272 121150 3324
rect 130562 3272 130568 3324
rect 130620 3312 130626 3324
rect 140958 3312 140964 3324
rect 130620 3284 140964 3312
rect 130620 3272 130626 3284
rect 140958 3272 140964 3284
rect 141016 3272 141022 3324
rect 143626 3272 143632 3324
rect 143684 3312 143690 3324
rect 153194 3312 153200 3324
rect 143684 3284 153200 3312
rect 143684 3272 143690 3284
rect 153194 3272 153200 3284
rect 153252 3272 153258 3324
rect 154206 3272 154212 3324
rect 154264 3312 154270 3324
rect 163038 3312 163044 3324
rect 154264 3284 163044 3312
rect 154264 3272 154270 3284
rect 163038 3272 163044 3284
rect 163096 3272 163102 3324
rect 164878 3272 164884 3324
rect 164936 3312 164942 3324
rect 172974 3312 172980 3324
rect 164936 3284 172980 3312
rect 164936 3272 164942 3284
rect 172974 3272 172980 3284
rect 173032 3272 173038 3324
rect 174262 3272 174268 3324
rect 174320 3312 174326 3324
rect 181806 3312 181812 3324
rect 174320 3284 181812 3312
rect 174320 3272 174326 3284
rect 181806 3272 181812 3284
rect 181864 3272 181870 3324
rect 189718 3272 189724 3324
rect 189776 3312 189782 3324
rect 196158 3312 196164 3324
rect 189776 3284 196164 3312
rect 189776 3272 189782 3284
rect 196158 3272 196164 3284
rect 196216 3272 196222 3324
rect 560018 3272 560024 3324
rect 560076 3312 560082 3324
rect 578602 3312 578608 3324
rect 560076 3284 578608 3312
rect 560076 3272 560082 3284
rect 578602 3272 578608 3284
rect 578660 3272 578666 3324
rect 113082 3244 113088 3256
rect 104268 3216 113088 3244
rect 96304 3204 96310 3216
rect 113082 3204 113088 3216
rect 113140 3204 113146 3256
rect 122282 3204 122288 3256
rect 122340 3244 122346 3256
rect 133230 3244 133236 3256
rect 122340 3216 133236 3244
rect 122340 3204 122346 3216
rect 133230 3204 133236 3216
rect 133288 3204 133294 3256
rect 139210 3204 139216 3256
rect 139268 3244 139274 3256
rect 148686 3244 148692 3256
rect 139268 3216 148692 3244
rect 139268 3204 139274 3216
rect 148686 3204 148692 3216
rect 148744 3204 148750 3256
rect 150618 3204 150624 3256
rect 150676 3244 150682 3256
rect 159726 3244 159732 3256
rect 150676 3216 159732 3244
rect 150676 3204 150682 3216
rect 159726 3204 159732 3216
rect 159784 3204 159790 3256
rect 161290 3204 161296 3256
rect 161348 3244 161354 3256
rect 169754 3244 169760 3256
rect 161348 3216 169760 3244
rect 161348 3204 161354 3216
rect 169754 3204 169760 3216
rect 169812 3204 169818 3256
rect 173158 3204 173164 3256
rect 173216 3244 173222 3256
rect 180886 3244 180892 3256
rect 173216 3216 180892 3244
rect 173216 3204 173222 3216
rect 180886 3204 180892 3216
rect 180944 3204 180950 3256
rect 182542 3204 182548 3256
rect 182600 3244 182606 3256
rect 189534 3244 189540 3256
rect 182600 3216 189540 3244
rect 182600 3204 182606 3216
rect 189534 3204 189540 3216
rect 189592 3204 189598 3256
rect 190822 3204 190828 3256
rect 190880 3244 190886 3256
rect 197354 3244 197360 3256
rect 190880 3216 197360 3244
rect 190880 3204 190886 3216
rect 197354 3204 197360 3216
rect 197412 3204 197418 3256
rect 200298 3204 200304 3256
rect 200356 3244 200362 3256
rect 206094 3244 206100 3256
rect 200356 3216 206100 3244
rect 200356 3204 200362 3216
rect 206094 3204 206100 3216
rect 206152 3204 206158 3256
rect 553302 3204 553308 3256
rect 553360 3244 553366 3256
rect 571518 3244 571524 3256
rect 553360 3216 571524 3244
rect 553360 3204 553366 3216
rect 571518 3204 571524 3216
rect 571576 3204 571582 3256
rect 81342 3176 81348 3188
rect 74506 3148 81348 3176
rect 81342 3136 81348 3148
rect 81400 3136 81406 3188
rect 82078 3136 82084 3188
rect 82136 3176 82142 3188
rect 95694 3176 95700 3188
rect 82136 3148 95700 3176
rect 82136 3136 82142 3148
rect 95694 3136 95700 3148
rect 95752 3136 95758 3188
rect 97442 3136 97448 3188
rect 97500 3176 97506 3188
rect 110046 3176 110052 3188
rect 97500 3148 110052 3176
rect 97500 3136 97506 3148
rect 110046 3136 110052 3148
rect 110104 3136 110110 3188
rect 110874 3136 110880 3188
rect 110932 3176 110938 3188
rect 122190 3176 122196 3188
rect 110932 3148 122196 3176
rect 110932 3136 110938 3148
rect 122190 3136 122196 3148
rect 122248 3136 122254 3188
rect 135254 3136 135260 3188
rect 135312 3176 135318 3188
rect 145374 3176 145380 3188
rect 135312 3148 145380 3176
rect 135312 3136 135318 3148
rect 145374 3136 145380 3148
rect 145432 3136 145438 3188
rect 147122 3136 147128 3188
rect 147180 3176 147186 3188
rect 156414 3176 156420 3188
rect 147180 3148 156420 3176
rect 147180 3136 147186 3148
rect 156414 3136 156420 3148
rect 156472 3136 156478 3188
rect 162486 3136 162492 3188
rect 162544 3176 162550 3188
rect 162544 3148 168696 3176
rect 162544 3136 162550 3148
rect 56042 3068 56048 3120
rect 56100 3108 56106 3120
rect 71406 3108 71412 3120
rect 56100 3080 71412 3108
rect 56100 3068 56106 3080
rect 71406 3068 71412 3080
rect 71464 3068 71470 3120
rect 87966 3068 87972 3120
rect 88024 3108 88030 3120
rect 101214 3108 101220 3120
rect 88024 3080 101220 3108
rect 88024 3068 88030 3080
rect 101214 3068 101220 3080
rect 101272 3068 101278 3120
rect 102226 3068 102232 3120
rect 102284 3108 102290 3120
rect 114554 3108 114560 3120
rect 102284 3080 114560 3108
rect 102284 3068 102290 3080
rect 114554 3068 114560 3080
rect 114612 3068 114618 3120
rect 115198 3068 115204 3120
rect 115256 3108 115262 3120
rect 126606 3108 126612 3120
rect 115256 3080 126612 3108
rect 115256 3068 115262 3080
rect 126606 3068 126612 3080
rect 126664 3068 126670 3120
rect 134150 3068 134156 3120
rect 134208 3108 134214 3120
rect 144270 3108 144276 3120
rect 134208 3080 144276 3108
rect 134208 3068 134214 3080
rect 144270 3068 144276 3080
rect 144328 3068 144334 3120
rect 151814 3068 151820 3120
rect 151872 3108 151878 3120
rect 160830 3108 160836 3120
rect 151872 3080 160836 3108
rect 151872 3068 151878 3080
rect 160830 3068 160836 3080
rect 160888 3068 160894 3120
rect 164234 3068 164240 3120
rect 164292 3108 164298 3120
rect 168558 3108 168564 3120
rect 164292 3080 168564 3108
rect 164292 3068 164298 3080
rect 168558 3068 168564 3080
rect 168616 3068 168622 3120
rect 168668 3108 168696 3148
rect 170766 3136 170772 3188
rect 170824 3176 170830 3188
rect 178494 3176 178500 3188
rect 170824 3148 178500 3176
rect 170824 3136 170830 3148
rect 178494 3136 178500 3148
rect 178552 3136 178558 3188
rect 179046 3136 179052 3188
rect 179104 3176 179110 3188
rect 186314 3176 186320 3188
rect 179104 3148 186320 3176
rect 179104 3136 179110 3148
rect 186314 3136 186320 3148
rect 186372 3136 186378 3188
rect 192386 3136 192392 3188
rect 192444 3176 192450 3188
rect 198366 3176 198372 3188
rect 192444 3148 198372 3176
rect 192444 3136 192450 3148
rect 198366 3136 198372 3148
rect 198424 3136 198430 3188
rect 201494 3136 201500 3188
rect 201552 3176 201558 3188
rect 206922 3176 206928 3188
rect 201552 3148 206928 3176
rect 201552 3136 201558 3148
rect 206922 3136 206928 3148
rect 206980 3136 206986 3188
rect 214466 3136 214472 3188
rect 214524 3176 214530 3188
rect 219342 3176 219348 3188
rect 214524 3148 219348 3176
rect 214524 3136 214530 3148
rect 219342 3136 219348 3148
rect 219400 3136 219406 3188
rect 220262 3136 220268 3188
rect 220320 3176 220326 3188
rect 224862 3176 224868 3188
rect 220320 3148 224868 3176
rect 220320 3136 220326 3148
rect 224862 3136 224868 3148
rect 224920 3136 224926 3188
rect 229830 3136 229836 3188
rect 229888 3176 229894 3188
rect 233694 3176 233700 3188
rect 229888 3148 233700 3176
rect 229888 3136 229894 3148
rect 233694 3136 233700 3148
rect 233752 3136 233758 3188
rect 556706 3136 556712 3188
rect 556764 3176 556770 3188
rect 575106 3176 575112 3188
rect 556764 3148 575112 3176
rect 556764 3136 556770 3148
rect 575106 3136 575112 3148
rect 575164 3136 575170 3188
rect 170858 3108 170864 3120
rect 168668 3080 170864 3108
rect 170858 3068 170864 3080
rect 170916 3068 170922 3120
rect 176746 3068 176752 3120
rect 176804 3108 176810 3120
rect 184014 3108 184020 3120
rect 176804 3080 184020 3108
rect 176804 3068 176810 3080
rect 184014 3068 184020 3080
rect 184072 3068 184078 3120
rect 196802 3068 196808 3120
rect 196860 3108 196866 3120
rect 202874 3108 202880 3120
rect 196860 3080 202880 3108
rect 196860 3068 196866 3080
rect 202874 3068 202880 3080
rect 202932 3068 202938 3120
rect 208946 3068 208952 3120
rect 209004 3108 209010 3120
rect 213822 3108 213828 3120
rect 209004 3080 213828 3108
rect 209004 3068 209010 3080
rect 213822 3068 213828 3080
rect 213880 3068 213886 3120
rect 215662 3068 215668 3120
rect 215720 3108 215726 3120
rect 220446 3108 220452 3120
rect 215720 3080 220452 3108
rect 215720 3068 215726 3080
rect 220446 3068 220452 3080
rect 220504 3068 220510 3120
rect 221550 3068 221556 3120
rect 221608 3108 221614 3120
rect 225966 3108 225972 3120
rect 221608 3080 225972 3108
rect 221608 3068 221614 3080
rect 225966 3068 225972 3080
rect 226024 3068 226030 3120
rect 231026 3068 231032 3120
rect 231084 3108 231090 3120
rect 234798 3108 234804 3120
rect 231084 3080 234804 3108
rect 231084 3068 231090 3080
rect 234798 3068 234804 3080
rect 234856 3068 234862 3120
rect 530026 3068 530032 3120
rect 530084 3108 530090 3120
rect 546678 3108 546684 3120
rect 530084 3080 546684 3108
rect 530084 3068 530090 3080
rect 546678 3068 546684 3080
rect 546736 3068 546742 3120
rect 564342 3068 564348 3120
rect 564400 3108 564406 3120
rect 583386 3108 583392 3120
rect 564400 3080 583392 3108
rect 564400 3068 564406 3080
rect 583386 3068 583392 3080
rect 583444 3068 583450 3120
rect 47854 3000 47860 3052
rect 47912 3040 47918 3052
rect 63678 3040 63684 3052
rect 47912 3012 63684 3040
rect 47912 3000 47918 3012
rect 63678 3000 63684 3012
rect 63736 3000 63742 3052
rect 70302 3040 70308 3052
rect 64846 3012 70308 3040
rect 33594 2932 33600 2984
rect 33652 2972 33658 2984
rect 50430 2972 50436 2984
rect 33652 2944 50436 2972
rect 33652 2932 33658 2944
rect 50430 2932 50436 2944
rect 50488 2932 50494 2984
rect 54938 2932 54944 2984
rect 54996 2972 55002 2984
rect 64846 2972 64874 3012
rect 70302 3000 70308 3012
rect 70360 3000 70366 3052
rect 76282 3000 76288 3052
rect 76340 3040 76346 3052
rect 90174 3040 90180 3052
rect 76340 3012 90180 3040
rect 76340 3000 76346 3012
rect 90174 3000 90180 3012
rect 90232 3000 90238 3052
rect 91922 3000 91928 3052
rect 91980 3040 91986 3052
rect 104526 3040 104532 3052
rect 91980 3012 104532 3040
rect 91980 3000 91986 3012
rect 104526 3000 104532 3012
rect 104584 3000 104590 3052
rect 108482 3000 108488 3052
rect 108540 3040 108546 3052
rect 119982 3040 119988 3052
rect 108540 3012 119988 3040
rect 108540 3000 108546 3012
rect 119982 3000 119988 3012
rect 120040 3000 120046 3052
rect 128170 3000 128176 3052
rect 128228 3040 128234 3052
rect 138750 3040 138756 3052
rect 128228 3012 138756 3040
rect 128228 3000 128234 3012
rect 138750 3000 138756 3012
rect 138808 3000 138814 3052
rect 140038 3000 140044 3052
rect 140096 3040 140102 3052
rect 149790 3040 149796 3052
rect 140096 3012 149796 3040
rect 140096 3000 140102 3012
rect 149790 3000 149796 3012
rect 149848 3000 149854 3052
rect 156598 3000 156604 3052
rect 156656 3040 156662 3052
rect 165246 3040 165252 3052
rect 156656 3012 165252 3040
rect 156656 3000 156662 3012
rect 165246 3000 165252 3012
rect 165304 3000 165310 3052
rect 171962 3000 171968 3052
rect 172020 3040 172026 3052
rect 179598 3040 179604 3052
rect 172020 3012 179604 3040
rect 172020 3000 172026 3012
rect 179598 3000 179604 3012
rect 179656 3000 179662 3052
rect 187326 3000 187332 3052
rect 187384 3040 187390 3052
rect 193950 3040 193956 3052
rect 187384 3012 193956 3040
rect 187384 3000 187390 3012
rect 193950 3000 193956 3012
rect 194008 3000 194014 3052
rect 194410 3000 194416 3052
rect 194468 3040 194474 3052
rect 200574 3040 200580 3052
rect 194468 3012 200580 3040
rect 194468 3000 194474 3012
rect 200574 3000 200580 3012
rect 200632 3000 200638 3052
rect 202690 3000 202696 3052
rect 202748 3040 202754 3052
rect 208394 3040 208400 3052
rect 202748 3012 208400 3040
rect 202748 3000 202754 3012
rect 208394 3000 208400 3012
rect 208452 3000 208458 3052
rect 214926 3040 214932 3052
rect 209792 3012 214932 3040
rect 209792 2984 209820 3012
rect 214926 3000 214932 3012
rect 214984 3000 214990 3052
rect 218054 3000 218060 3052
rect 218112 3040 218118 3052
rect 222654 3040 222660 3052
rect 218112 3012 222660 3040
rect 218112 3000 218118 3012
rect 222654 3000 222660 3012
rect 222712 3000 222718 3052
rect 225506 3000 225512 3052
rect 225564 3040 225570 3052
rect 229278 3040 229284 3052
rect 225564 3012 229284 3040
rect 225564 3000 225570 3012
rect 229278 3000 229284 3012
rect 229336 3000 229342 3052
rect 233418 3000 233424 3052
rect 233476 3040 233482 3052
rect 237006 3040 237012 3052
rect 233476 3012 237012 3040
rect 233476 3000 233482 3012
rect 237006 3000 237012 3012
rect 237064 3000 237070 3052
rect 238110 3000 238116 3052
rect 238168 3040 238174 3052
rect 241514 3040 241520 3052
rect 238168 3012 241520 3040
rect 238168 3000 238174 3012
rect 241514 3000 241520 3012
rect 241572 3000 241578 3052
rect 248782 3000 248788 3052
rect 248840 3040 248846 3052
rect 251358 3040 251364 3052
rect 248840 3012 251364 3040
rect 248840 3000 248846 3012
rect 251358 3000 251364 3012
rect 251416 3000 251422 3052
rect 331306 3000 331312 3052
rect 331364 3040 331370 3052
rect 333882 3040 333888 3052
rect 331364 3012 333888 3040
rect 331364 3000 331370 3012
rect 333882 3000 333888 3012
rect 333940 3000 333946 3052
rect 334802 3000 334808 3052
rect 334860 3040 334866 3052
rect 337470 3040 337476 3052
rect 334860 3012 337476 3040
rect 334860 3000 334866 3012
rect 337470 3000 337476 3012
rect 337528 3000 337534 3052
rect 543458 3000 543464 3052
rect 543516 3040 543522 3052
rect 560478 3040 560484 3052
rect 543516 3012 560484 3040
rect 543516 3000 543522 3012
rect 560478 3000 560484 3012
rect 560536 3000 560542 3052
rect 562226 3000 562232 3052
rect 562284 3040 562290 3052
rect 580994 3040 581000 3052
rect 562284 3012 581000 3040
rect 562284 3000 562290 3012
rect 580994 3000 581000 3012
rect 581052 3000 581058 3052
rect 54996 2944 64874 2972
rect 54996 2932 55002 2944
rect 69106 2932 69112 2984
rect 69164 2972 69170 2984
rect 83826 2972 83832 2984
rect 69164 2944 83832 2972
rect 69164 2932 69170 2944
rect 83826 2932 83832 2944
rect 83884 2932 83890 2984
rect 84470 2932 84476 2984
rect 84528 2972 84534 2984
rect 98178 2972 98184 2984
rect 84528 2944 98184 2972
rect 84528 2932 84534 2944
rect 98178 2932 98184 2944
rect 98236 2932 98242 2984
rect 106918 2932 106924 2984
rect 106976 2972 106982 2984
rect 119154 2972 119160 2984
rect 106976 2944 119160 2972
rect 106976 2932 106982 2944
rect 119154 2932 119160 2944
rect 119212 2932 119218 2984
rect 119890 2932 119896 2984
rect 119948 2972 119954 2984
rect 131298 2972 131304 2984
rect 119948 2944 131304 2972
rect 119948 2932 119954 2944
rect 131298 2932 131304 2944
rect 131356 2932 131362 2984
rect 131758 2932 131764 2984
rect 131816 2972 131822 2984
rect 142338 2972 142344 2984
rect 131816 2944 142344 2972
rect 131816 2932 131822 2944
rect 142338 2932 142344 2944
rect 142396 2932 142402 2984
rect 145926 2932 145932 2984
rect 145984 2972 145990 2984
rect 155586 2972 155592 2984
rect 145984 2944 155592 2972
rect 145984 2932 145990 2944
rect 155586 2932 155592 2944
rect 155644 2932 155650 2984
rect 157794 2932 157800 2984
rect 157852 2972 157858 2984
rect 166626 2972 166632 2984
rect 157852 2944 166632 2972
rect 157852 2932 157858 2944
rect 166626 2932 166632 2944
rect 166684 2932 166690 2984
rect 174354 2972 174360 2984
rect 166736 2944 174360 2972
rect 26602 2864 26608 2916
rect 26660 2904 26666 2916
rect 43806 2904 43812 2916
rect 26660 2876 43812 2904
rect 26660 2864 26666 2876
rect 43806 2864 43812 2876
rect 43864 2864 43870 2916
rect 44266 2864 44272 2916
rect 44324 2904 44330 2916
rect 60366 2904 60372 2916
rect 44324 2876 60372 2904
rect 44324 2864 44330 2876
rect 60366 2864 60372 2876
rect 60424 2864 60430 2916
rect 65518 2864 65524 2916
rect 65576 2904 65582 2916
rect 65576 2876 74534 2904
rect 65576 2864 65582 2876
rect 27706 2796 27712 2848
rect 27764 2836 27770 2848
rect 44910 2836 44916 2848
rect 27764 2808 44916 2836
rect 27764 2796 27770 2808
rect 44910 2796 44916 2808
rect 44968 2796 44974 2848
rect 50154 2796 50160 2848
rect 50212 2836 50218 2848
rect 65886 2836 65892 2848
rect 50212 2808 65892 2836
rect 50212 2796 50218 2808
rect 65886 2796 65892 2808
rect 65944 2796 65950 2848
rect 67910 2796 67916 2848
rect 67968 2836 67974 2848
rect 68554 2836 68560 2848
rect 67968 2808 68560 2836
rect 67968 2796 67974 2808
rect 68554 2796 68560 2808
rect 68612 2796 68618 2848
rect 74506 2836 74534 2876
rect 78582 2864 78588 2916
rect 78640 2904 78646 2916
rect 92474 2904 92480 2916
rect 78640 2876 92480 2904
rect 78640 2864 78646 2876
rect 92474 2864 92480 2876
rect 92532 2864 92538 2916
rect 92750 2864 92756 2916
rect 92808 2904 92814 2916
rect 105906 2904 105912 2916
rect 92808 2876 105912 2904
rect 92808 2864 92814 2876
rect 105906 2864 105912 2876
rect 105964 2864 105970 2916
rect 112806 2864 112812 2916
rect 112864 2904 112870 2916
rect 124674 2904 124680 2916
rect 112864 2876 124680 2904
rect 112864 2864 112870 2876
rect 124674 2864 124680 2876
rect 124732 2864 124738 2916
rect 125042 2864 125048 2916
rect 125100 2904 125106 2916
rect 135714 2904 135720 2916
rect 125100 2876 135720 2904
rect 125100 2864 125106 2876
rect 135714 2864 135720 2876
rect 135772 2864 135778 2916
rect 141234 2864 141240 2916
rect 141292 2904 141298 2916
rect 151170 2904 151176 2916
rect 141292 2876 151176 2904
rect 141292 2864 141298 2876
rect 151170 2864 151176 2876
rect 151228 2864 151234 2916
rect 158898 2864 158904 2916
rect 158956 2904 158962 2916
rect 158956 2876 164372 2904
rect 158956 2864 158962 2876
rect 79962 2836 79968 2848
rect 74506 2808 79968 2836
rect 79962 2796 79968 2808
rect 80020 2796 80026 2848
rect 86862 2796 86868 2848
rect 86920 2836 86926 2848
rect 100386 2836 100392 2848
rect 86920 2808 100392 2836
rect 86920 2796 86926 2808
rect 100386 2796 100392 2808
rect 100444 2796 100450 2848
rect 104526 2796 104532 2848
rect 104584 2836 104590 2848
rect 110506 2836 110512 2848
rect 104584 2808 110512 2836
rect 104584 2796 104590 2808
rect 110506 2796 110512 2808
rect 110564 2796 110570 2848
rect 111610 2796 111616 2848
rect 111668 2836 111674 2848
rect 123570 2836 123576 2848
rect 111668 2808 123576 2836
rect 111668 2796 111674 2808
rect 123570 2796 123576 2808
rect 123628 2796 123634 2848
rect 134610 2836 134616 2848
rect 123680 2808 134616 2836
rect 123478 2728 123484 2780
rect 123536 2768 123542 2780
rect 123680 2768 123708 2808
rect 134610 2796 134616 2808
rect 134668 2796 134674 2848
rect 136450 2796 136456 2848
rect 136508 2836 136514 2848
rect 146754 2836 146760 2848
rect 136508 2808 146760 2836
rect 136508 2796 136514 2808
rect 146754 2796 146760 2808
rect 146812 2796 146818 2848
rect 149514 2796 149520 2848
rect 149572 2836 149578 2848
rect 158714 2836 158720 2848
rect 149572 2808 158720 2836
rect 149572 2796 149578 2808
rect 158714 2796 158720 2808
rect 158772 2796 158778 2848
rect 160094 2796 160100 2848
rect 160152 2836 160158 2848
rect 164234 2836 164240 2848
rect 160152 2808 164240 2836
rect 160152 2796 160158 2808
rect 164234 2796 164240 2808
rect 164292 2796 164298 2848
rect 164344 2836 164372 2876
rect 166074 2864 166080 2916
rect 166132 2904 166138 2916
rect 166736 2904 166764 2944
rect 174354 2932 174360 2944
rect 174412 2932 174418 2984
rect 177850 2932 177856 2984
rect 177908 2972 177914 2984
rect 185394 2972 185400 2984
rect 177908 2944 185400 2972
rect 177908 2932 177914 2944
rect 185394 2932 185400 2944
rect 185452 2932 185458 2984
rect 186130 2932 186136 2984
rect 186188 2972 186194 2984
rect 193122 2972 193128 2984
rect 186188 2944 193128 2972
rect 186188 2932 186194 2944
rect 193122 2932 193128 2944
rect 193180 2932 193186 2984
rect 195606 2932 195612 2984
rect 195664 2972 195670 2984
rect 201954 2972 201960 2984
rect 195664 2944 201960 2972
rect 195664 2932 195670 2944
rect 201954 2932 201960 2944
rect 202012 2932 202018 2984
rect 203886 2932 203892 2984
rect 203944 2972 203950 2984
rect 209406 2972 209412 2984
rect 203944 2944 209412 2972
rect 203944 2932 203950 2944
rect 209406 2932 209412 2944
rect 209464 2932 209470 2984
rect 209774 2932 209780 2984
rect 209832 2932 209838 2984
rect 212166 2932 212172 2984
rect 212224 2972 212230 2984
rect 217134 2972 217140 2984
rect 212224 2944 217140 2972
rect 212224 2932 212230 2944
rect 217134 2932 217140 2944
rect 217192 2932 217198 2984
rect 222746 2932 222752 2984
rect 222804 2972 222810 2984
rect 227346 2972 227352 2984
rect 222804 2944 227352 2972
rect 222804 2932 222810 2944
rect 227346 2932 227352 2944
rect 227404 2932 227410 2984
rect 227530 2932 227536 2984
rect 227588 2972 227594 2984
rect 231762 2972 231768 2984
rect 227588 2944 231768 2972
rect 227588 2932 227594 2944
rect 231762 2932 231768 2944
rect 231820 2932 231826 2984
rect 234614 2932 234620 2984
rect 234672 2972 234678 2984
rect 238386 2972 238392 2984
rect 234672 2944 238392 2972
rect 234672 2932 234678 2944
rect 238386 2932 238392 2944
rect 238444 2932 238450 2984
rect 239306 2932 239312 2984
rect 239364 2972 239370 2984
rect 242802 2972 242808 2984
rect 239364 2944 242808 2972
rect 239364 2932 239370 2944
rect 242802 2932 242808 2944
rect 242860 2932 242866 2984
rect 242894 2932 242900 2984
rect 242952 2972 242958 2984
rect 246114 2972 246120 2984
rect 242952 2944 246120 2972
rect 242952 2932 242958 2944
rect 246114 2932 246120 2944
rect 246172 2932 246178 2984
rect 246390 2932 246396 2984
rect 246448 2972 246454 2984
rect 249426 2972 249432 2984
rect 246448 2944 249432 2972
rect 246448 2932 246454 2944
rect 249426 2932 249432 2944
rect 249484 2932 249490 2984
rect 253474 2932 253480 2984
rect 253532 2972 253538 2984
rect 256050 2972 256056 2984
rect 253532 2944 256056 2972
rect 253532 2932 253538 2944
rect 256050 2932 256056 2944
rect 256108 2932 256114 2984
rect 310238 2932 310244 2984
rect 310296 2972 310302 2984
rect 311434 2972 311440 2984
rect 310296 2944 311440 2972
rect 310296 2932 310302 2944
rect 311434 2932 311440 2944
rect 311492 2932 311498 2984
rect 325694 2932 325700 2984
rect 325752 2972 325758 2984
rect 327994 2972 328000 2984
rect 325752 2944 328000 2972
rect 325752 2932 325758 2944
rect 327994 2932 328000 2944
rect 328052 2932 328058 2984
rect 329006 2932 329012 2984
rect 329064 2972 329070 2984
rect 331582 2972 331588 2984
rect 329064 2944 331588 2972
rect 329064 2932 329070 2944
rect 331582 2932 331588 2944
rect 331640 2932 331646 2984
rect 332318 2932 332324 2984
rect 332376 2972 332382 2984
rect 335078 2972 335084 2984
rect 332376 2944 335084 2972
rect 332376 2932 332382 2944
rect 335078 2932 335084 2944
rect 335136 2932 335142 2984
rect 341150 2932 341156 2984
rect 341208 2972 341214 2984
rect 344554 2972 344560 2984
rect 341208 2944 344560 2972
rect 341208 2932 341214 2944
rect 344554 2932 344560 2944
rect 344612 2932 344618 2984
rect 536558 2932 536564 2984
rect 536616 2972 536622 2984
rect 553762 2972 553768 2984
rect 536616 2944 553768 2972
rect 536616 2932 536622 2944
rect 553762 2932 553768 2944
rect 553820 2932 553826 2984
rect 560846 2932 560852 2984
rect 560904 2972 560910 2984
rect 579798 2972 579804 2984
rect 560904 2944 579804 2972
rect 560904 2932 560910 2944
rect 579798 2932 579804 2944
rect 579856 2932 579862 2984
rect 166132 2876 166764 2904
rect 166132 2864 166138 2876
rect 168374 2864 168380 2916
rect 168432 2904 168438 2916
rect 176562 2904 176568 2916
rect 168432 2876 176568 2904
rect 168432 2864 168438 2876
rect 176562 2864 176568 2876
rect 176620 2864 176626 2916
rect 181438 2864 181444 2916
rect 181496 2904 181502 2916
rect 188430 2904 188436 2916
rect 181496 2876 188436 2904
rect 181496 2864 181502 2876
rect 188430 2864 188436 2876
rect 188488 2864 188494 2916
rect 188522 2864 188528 2916
rect 188580 2904 188586 2916
rect 195330 2904 195336 2916
rect 188580 2876 195336 2904
rect 188580 2864 188586 2876
rect 195330 2864 195336 2876
rect 195388 2864 195394 2916
rect 199102 2864 199108 2916
rect 199160 2904 199166 2916
rect 204990 2904 204996 2916
rect 199160 2876 204996 2904
rect 199160 2864 199166 2876
rect 204990 2864 204996 2876
rect 205048 2864 205054 2916
rect 206186 2864 206192 2916
rect 206244 2904 206250 2916
rect 211614 2904 211620 2916
rect 206244 2876 211620 2904
rect 206244 2864 206250 2876
rect 211614 2864 211620 2876
rect 211672 2864 211678 2916
rect 213362 2864 213368 2916
rect 213420 2904 213426 2916
rect 218238 2904 218244 2916
rect 213420 2876 218244 2904
rect 213420 2864 213426 2876
rect 218238 2864 218244 2876
rect 218296 2864 218302 2916
rect 219250 2864 219256 2916
rect 219308 2904 219314 2916
rect 223482 2904 223488 2916
rect 219308 2876 223488 2904
rect 219308 2864 219314 2876
rect 223482 2864 223488 2876
rect 223540 2864 223546 2916
rect 226334 2864 226340 2916
rect 226392 2904 226398 2916
rect 230658 2904 230664 2916
rect 226392 2876 230664 2904
rect 226392 2864 226398 2876
rect 230658 2864 230664 2876
rect 230716 2864 230722 2916
rect 232222 2864 232228 2916
rect 232280 2904 232286 2916
rect 236178 2904 236184 2916
rect 232280 2876 236184 2904
rect 232280 2864 232286 2876
rect 236178 2864 236184 2876
rect 236236 2864 236242 2916
rect 237006 2864 237012 2916
rect 237064 2904 237070 2916
rect 240594 2904 240600 2916
rect 237064 2876 240600 2904
rect 237064 2864 237070 2876
rect 240594 2864 240600 2876
rect 240652 2864 240658 2916
rect 242066 2864 242072 2916
rect 242124 2904 242130 2916
rect 245010 2904 245016 2916
rect 242124 2876 245016 2904
rect 242124 2864 242130 2876
rect 245010 2864 245016 2876
rect 245068 2864 245074 2916
rect 245194 2864 245200 2916
rect 245252 2904 245258 2916
rect 248322 2904 248328 2916
rect 245252 2876 248328 2904
rect 245252 2864 245258 2876
rect 248322 2864 248328 2876
rect 248380 2864 248386 2916
rect 249978 2864 249984 2916
rect 250036 2904 250042 2916
rect 252738 2904 252744 2916
rect 250036 2876 252744 2904
rect 250036 2864 250042 2876
rect 252738 2864 252744 2876
rect 252796 2864 252802 2916
rect 254670 2864 254676 2916
rect 254728 2904 254734 2916
rect 257154 2904 257160 2916
rect 254728 2876 257160 2904
rect 254728 2864 254734 2876
rect 257154 2864 257160 2876
rect 257212 2864 257218 2916
rect 261754 2864 261760 2916
rect 261812 2904 261818 2916
rect 263778 2904 263784 2916
rect 261812 2876 263784 2904
rect 261812 2864 261818 2876
rect 263778 2864 263784 2876
rect 263836 2864 263842 2916
rect 312446 2864 312452 2916
rect 312504 2904 312510 2916
rect 313826 2904 313832 2916
rect 312504 2876 313832 2904
rect 312504 2864 312510 2876
rect 313826 2864 313832 2876
rect 313884 2864 313890 2916
rect 314562 2864 314568 2916
rect 314620 2904 314626 2916
rect 316218 2904 316224 2916
rect 314620 2876 316224 2904
rect 314620 2864 314626 2876
rect 316218 2864 316224 2876
rect 316276 2864 316282 2916
rect 316862 2864 316868 2916
rect 316920 2904 316926 2916
rect 318518 2904 318524 2916
rect 316920 2876 318524 2904
rect 316920 2864 316926 2876
rect 318518 2864 318524 2876
rect 318576 2864 318582 2916
rect 319070 2864 319076 2916
rect 319128 2904 319134 2916
rect 320910 2904 320916 2916
rect 319128 2876 320916 2904
rect 319128 2864 319134 2876
rect 320910 2864 320916 2876
rect 320968 2864 320974 2916
rect 321278 2864 321284 2916
rect 321336 2904 321342 2916
rect 323302 2904 323308 2916
rect 321336 2876 323308 2904
rect 321336 2864 321342 2876
rect 323302 2864 323308 2876
rect 323360 2864 323366 2916
rect 323486 2864 323492 2916
rect 323544 2904 323550 2916
rect 325602 2904 325608 2916
rect 323544 2876 325608 2904
rect 323544 2864 323550 2876
rect 325602 2864 325608 2876
rect 325660 2864 325666 2916
rect 327902 2864 327908 2916
rect 327960 2904 327966 2916
rect 330386 2904 330392 2916
rect 327960 2876 330392 2904
rect 327960 2864 327966 2876
rect 330386 2864 330392 2876
rect 330444 2864 330450 2916
rect 333422 2864 333428 2916
rect 333480 2904 333486 2916
rect 336274 2904 336280 2916
rect 333480 2876 336280 2904
rect 333480 2864 333486 2876
rect 336274 2864 336280 2876
rect 336332 2864 336338 2916
rect 340046 2864 340052 2916
rect 340104 2904 340110 2916
rect 342990 2904 342996 2916
rect 340104 2876 342996 2904
rect 340104 2864 340110 2876
rect 342990 2864 342996 2876
rect 343048 2864 343054 2916
rect 526622 2864 526628 2916
rect 526680 2904 526686 2916
rect 542814 2904 542820 2916
rect 526680 2876 542820 2904
rect 526680 2864 526686 2876
rect 542814 2864 542820 2876
rect 542872 2864 542878 2916
rect 549806 2864 549812 2916
rect 549864 2904 549870 2916
rect 568022 2904 568028 2916
rect 549864 2876 568028 2904
rect 549864 2864 549870 2876
rect 568022 2864 568028 2876
rect 568080 2864 568086 2916
rect 167730 2836 167736 2848
rect 164344 2808 167736 2836
rect 167730 2796 167736 2808
rect 167788 2796 167794 2848
rect 175458 2796 175464 2848
rect 175516 2836 175522 2848
rect 183186 2836 183192 2848
rect 175516 2808 183192 2836
rect 175516 2796 175522 2808
rect 183186 2796 183192 2808
rect 183244 2796 183250 2848
rect 184934 2796 184940 2848
rect 184992 2836 184998 2848
rect 192018 2836 192024 2848
rect 184992 2808 192024 2836
rect 184992 2796 184998 2808
rect 192018 2796 192024 2808
rect 192076 2796 192082 2848
rect 199470 2836 199476 2848
rect 193232 2808 199476 2836
rect 193232 2780 193260 2808
rect 199470 2796 199476 2808
rect 199528 2796 199534 2848
rect 205082 2796 205088 2848
rect 205140 2836 205146 2848
rect 210510 2836 210516 2848
rect 205140 2808 210516 2836
rect 205140 2796 205146 2808
rect 210510 2796 210516 2808
rect 210568 2796 210574 2848
rect 210970 2796 210976 2848
rect 211028 2836 211034 2848
rect 216030 2836 216036 2848
rect 211028 2808 216036 2836
rect 211028 2796 211034 2808
rect 216030 2796 216036 2808
rect 216088 2796 216094 2848
rect 216858 2796 216864 2848
rect 216916 2836 216922 2848
rect 221826 2836 221832 2848
rect 216916 2808 221832 2836
rect 216916 2796 216922 2808
rect 221826 2796 221832 2808
rect 221884 2796 221890 2848
rect 223942 2796 223948 2848
rect 224000 2836 224006 2848
rect 228450 2836 228456 2848
rect 224000 2808 228456 2836
rect 224000 2796 224006 2808
rect 228450 2796 228456 2808
rect 228508 2796 228514 2848
rect 228726 2796 228732 2848
rect 228784 2836 228790 2848
rect 232866 2836 232872 2848
rect 228784 2808 232872 2836
rect 228784 2796 228790 2808
rect 232866 2796 232872 2808
rect 232924 2796 232930 2848
rect 235810 2796 235816 2848
rect 235868 2836 235874 2848
rect 239490 2836 239496 2848
rect 235868 2808 239496 2836
rect 235868 2796 235874 2808
rect 239490 2796 239496 2808
rect 239548 2796 239554 2848
rect 240502 2796 240508 2848
rect 240560 2836 240566 2848
rect 243906 2836 243912 2848
rect 240560 2808 243912 2836
rect 240560 2796 240566 2808
rect 243906 2796 243912 2808
rect 243964 2796 243970 2848
rect 244090 2796 244096 2848
rect 244148 2836 244154 2848
rect 247218 2836 247224 2848
rect 244148 2808 247224 2836
rect 244148 2796 244154 2808
rect 247218 2796 247224 2808
rect 247276 2796 247282 2848
rect 247586 2796 247592 2848
rect 247644 2836 247650 2848
rect 250530 2836 250536 2848
rect 247644 2808 250536 2836
rect 247644 2796 247650 2808
rect 250530 2796 250536 2808
rect 250588 2796 250594 2848
rect 252370 2796 252376 2848
rect 252428 2836 252434 2848
rect 254946 2836 254952 2848
rect 252428 2808 254952 2836
rect 252428 2796 252434 2808
rect 254946 2796 254952 2808
rect 255004 2796 255010 2848
rect 255866 2796 255872 2848
rect 255924 2836 255930 2848
rect 258258 2836 258264 2848
rect 255924 2808 258264 2836
rect 255924 2796 255930 2808
rect 258258 2796 258264 2808
rect 258316 2796 258322 2848
rect 260650 2796 260656 2848
rect 260708 2836 260714 2848
rect 262674 2836 262680 2848
rect 260708 2808 262680 2836
rect 260708 2796 260714 2808
rect 262674 2796 262680 2808
rect 262732 2796 262738 2848
rect 304718 2796 304724 2848
rect 304776 2836 304782 2848
rect 305546 2836 305552 2848
rect 304776 2808 305552 2836
rect 304776 2796 304782 2808
rect 305546 2796 305552 2808
rect 305604 2796 305610 2848
rect 306926 2796 306932 2848
rect 306984 2836 306990 2848
rect 307938 2836 307944 2848
rect 306984 2808 307944 2836
rect 306984 2796 306990 2808
rect 307938 2796 307944 2808
rect 307996 2796 308002 2848
rect 309134 2796 309140 2848
rect 309192 2836 309198 2848
rect 310238 2836 310244 2848
rect 309192 2808 310244 2836
rect 309192 2796 309198 2808
rect 310238 2796 310244 2808
rect 310296 2796 310302 2848
rect 311342 2796 311348 2848
rect 311400 2836 311406 2848
rect 312630 2836 312636 2848
rect 311400 2808 312636 2836
rect 311400 2796 311406 2808
rect 312630 2796 312636 2808
rect 312688 2796 312694 2848
rect 313550 2796 313556 2848
rect 313608 2836 313614 2848
rect 315022 2836 315028 2848
rect 313608 2808 315028 2836
rect 313608 2796 313614 2808
rect 315022 2796 315028 2808
rect 315080 2796 315086 2848
rect 315758 2796 315764 2848
rect 315816 2836 315822 2848
rect 317322 2836 317328 2848
rect 315816 2808 317328 2836
rect 315816 2796 315822 2808
rect 317322 2796 317328 2808
rect 317380 2796 317386 2848
rect 317966 2796 317972 2848
rect 318024 2836 318030 2848
rect 319714 2836 319720 2848
rect 318024 2808 319720 2836
rect 318024 2796 318030 2808
rect 319714 2796 319720 2808
rect 319772 2796 319778 2848
rect 320082 2796 320088 2848
rect 320140 2836 320146 2848
rect 322106 2836 322112 2848
rect 320140 2808 322112 2836
rect 320140 2796 320146 2808
rect 322106 2796 322112 2808
rect 322164 2796 322170 2848
rect 322382 2796 322388 2848
rect 322440 2836 322446 2848
rect 324406 2836 324412 2848
rect 322440 2808 324412 2836
rect 322440 2796 322446 2808
rect 324406 2796 324412 2808
rect 324464 2796 324470 2848
rect 324590 2796 324596 2848
rect 324648 2836 324654 2848
rect 326798 2836 326804 2848
rect 324648 2808 326804 2836
rect 324648 2796 324654 2808
rect 326798 2796 326804 2808
rect 326856 2796 326862 2848
rect 326982 2796 326988 2848
rect 327040 2836 327046 2848
rect 329190 2836 329196 2848
rect 327040 2808 329196 2836
rect 327040 2796 327046 2808
rect 329190 2796 329196 2808
rect 329248 2796 329254 2848
rect 330110 2796 330116 2848
rect 330168 2836 330174 2848
rect 332686 2836 332692 2848
rect 330168 2808 332692 2836
rect 330168 2796 330174 2808
rect 332686 2796 332692 2808
rect 332744 2796 332750 2848
rect 335630 2796 335636 2848
rect 335688 2836 335694 2848
rect 338666 2836 338672 2848
rect 335688 2808 338672 2836
rect 335688 2796 335694 2808
rect 338666 2796 338672 2808
rect 338724 2796 338730 2848
rect 338942 2796 338948 2848
rect 339000 2836 339006 2848
rect 342070 2836 342076 2848
rect 339000 2808 342076 2836
rect 339000 2796 339006 2808
rect 342070 2796 342076 2808
rect 342128 2796 342134 2848
rect 346670 2796 346676 2848
rect 346728 2836 346734 2848
rect 350442 2836 350448 2848
rect 346728 2808 350448 2836
rect 346728 2796 346734 2808
rect 350442 2796 350448 2808
rect 350500 2796 350506 2848
rect 353202 2796 353208 2848
rect 353260 2836 353266 2848
rect 357526 2836 357532 2848
rect 353260 2808 357532 2836
rect 353260 2796 353266 2808
rect 357526 2796 357532 2808
rect 357584 2796 357590 2848
rect 372338 2796 372344 2848
rect 372396 2836 372402 2848
rect 377674 2836 377680 2848
rect 372396 2808 377680 2836
rect 372396 2796 372402 2808
rect 377674 2796 377680 2808
rect 377732 2796 377738 2848
rect 546494 2796 546500 2848
rect 546552 2836 546558 2848
rect 557350 2836 557356 2848
rect 546552 2808 557356 2836
rect 546552 2796 546558 2808
rect 557350 2796 557356 2808
rect 557408 2796 557414 2848
rect 562962 2796 562968 2848
rect 563020 2836 563026 2848
rect 582190 2836 582196 2848
rect 563020 2808 582196 2836
rect 563020 2796 563026 2808
rect 582190 2796 582196 2808
rect 582248 2796 582254 2848
rect 123536 2740 123708 2768
rect 123536 2728 123542 2740
rect 193214 2728 193220 2780
rect 193272 2728 193278 2780
rect 198274 1300 198280 1352
rect 198332 1340 198338 1352
rect 204162 1340 204168 1352
rect 198332 1312 204168 1340
rect 198332 1300 198338 1312
rect 204162 1300 204168 1312
rect 204220 1300 204226 1352
rect 207382 1300 207388 1352
rect 207440 1340 207446 1352
rect 212994 1340 213000 1352
rect 207440 1312 213000 1340
rect 207440 1300 207446 1312
rect 212994 1300 213000 1312
rect 213052 1300 213058 1352
rect 257062 1300 257068 1352
rect 257120 1340 257126 1352
rect 259362 1340 259368 1352
rect 257120 1312 259368 1340
rect 257120 1300 257126 1312
rect 259362 1300 259368 1312
rect 259420 1300 259426 1352
rect 259454 1300 259460 1352
rect 259512 1340 259518 1352
rect 261570 1340 261576 1352
rect 259512 1312 261576 1340
rect 259512 1300 259518 1312
rect 261570 1300 261576 1312
rect 261628 1300 261634 1352
rect 262950 1300 262956 1352
rect 263008 1340 263014 1352
rect 264882 1340 264888 1352
rect 263008 1312 264888 1340
rect 263008 1300 263014 1312
rect 264882 1300 264888 1312
rect 264940 1300 264946 1352
rect 265342 1300 265348 1352
rect 265400 1340 265406 1352
rect 267090 1340 267096 1352
rect 265400 1312 267096 1340
rect 265400 1300 265406 1312
rect 267090 1300 267096 1312
rect 267148 1300 267154 1352
rect 267734 1300 267740 1352
rect 267792 1340 267798 1352
rect 269298 1340 269304 1352
rect 267792 1312 269304 1340
rect 267792 1300 267798 1312
rect 269298 1300 269304 1312
rect 269356 1300 269362 1352
rect 271230 1300 271236 1352
rect 271288 1340 271294 1352
rect 272610 1340 272616 1352
rect 271288 1312 272616 1340
rect 271288 1300 271294 1312
rect 272610 1300 272616 1312
rect 272668 1300 272674 1352
rect 273622 1300 273628 1352
rect 273680 1340 273686 1352
rect 274818 1340 274824 1352
rect 273680 1312 274824 1340
rect 273680 1300 273686 1312
rect 274818 1300 274824 1312
rect 274876 1300 274882 1352
rect 277118 1300 277124 1352
rect 277176 1340 277182 1352
rect 278130 1340 278136 1352
rect 277176 1312 278136 1340
rect 277176 1300 277182 1312
rect 278130 1300 278136 1312
rect 278188 1300 278194 1352
rect 279510 1300 279516 1352
rect 279568 1340 279574 1352
rect 280338 1340 280344 1352
rect 279568 1312 280344 1340
rect 279568 1300 279574 1312
rect 280338 1300 280344 1312
rect 280396 1300 280402 1352
rect 336642 1300 336648 1352
rect 336700 1340 336706 1352
rect 339862 1340 339868 1352
rect 336700 1312 339868 1340
rect 336700 1300 336706 1312
rect 339862 1300 339868 1312
rect 339920 1300 339926 1352
rect 342162 1300 342168 1352
rect 342220 1340 342226 1352
rect 345750 1340 345756 1352
rect 342220 1312 345756 1340
rect 342220 1300 342226 1312
rect 345750 1300 345756 1312
rect 345808 1300 345814 1352
rect 348878 1300 348884 1352
rect 348936 1340 348942 1352
rect 352834 1340 352840 1352
rect 348936 1312 352840 1340
rect 348936 1300 348942 1312
rect 352834 1300 352840 1312
rect 352892 1300 352898 1352
rect 356606 1300 356612 1352
rect 356664 1340 356670 1352
rect 361114 1340 361120 1352
rect 356664 1312 361120 1340
rect 356664 1300 356670 1312
rect 361114 1300 361120 1312
rect 361172 1300 361178 1352
rect 364242 1300 364248 1352
rect 364300 1340 364306 1352
rect 369394 1340 369400 1352
rect 364300 1312 369400 1340
rect 364300 1300 364306 1312
rect 369394 1300 369400 1312
rect 369452 1300 369458 1352
rect 369762 1300 369768 1352
rect 369820 1340 369826 1352
rect 375282 1340 375288 1352
rect 369820 1312 375288 1340
rect 369820 1300 369826 1312
rect 375282 1300 375288 1312
rect 375340 1300 375346 1352
rect 376478 1300 376484 1352
rect 376536 1340 376542 1352
rect 382366 1340 382372 1352
rect 376536 1312 382372 1340
rect 376536 1300 376542 1312
rect 382366 1300 382372 1312
rect 382424 1300 382430 1352
rect 384206 1300 384212 1352
rect 384264 1340 384270 1352
rect 390646 1340 390652 1352
rect 384264 1312 390652 1340
rect 384264 1300 384270 1312
rect 390646 1300 390652 1312
rect 390704 1300 390710 1352
rect 394142 1300 394148 1352
rect 394200 1340 394206 1352
rect 401318 1340 401324 1352
rect 394200 1312 401324 1340
rect 394200 1300 394206 1312
rect 401318 1300 401324 1312
rect 401376 1300 401382 1352
rect 406286 1300 406292 1352
rect 406344 1340 406350 1352
rect 414290 1340 414296 1352
rect 406344 1312 414296 1340
rect 406344 1300 406350 1312
rect 414290 1300 414296 1312
rect 414348 1300 414354 1352
rect 436002 1300 436008 1352
rect 436060 1340 436066 1352
rect 445846 1340 445852 1352
rect 436060 1312 445852 1340
rect 436060 1300 436066 1312
rect 445846 1300 445852 1312
rect 445904 1300 445910 1352
rect 450446 1300 450452 1352
rect 450504 1340 450510 1352
rect 461578 1340 461584 1352
rect 450504 1312 461584 1340
rect 450504 1300 450510 1312
rect 461578 1300 461584 1312
rect 461636 1300 461642 1352
rect 462590 1300 462596 1352
rect 462648 1340 462654 1352
rect 474182 1340 474188 1352
rect 462648 1312 474188 1340
rect 462648 1300 462654 1312
rect 474182 1300 474188 1312
rect 474240 1300 474246 1352
rect 475838 1300 475844 1352
rect 475896 1340 475902 1352
rect 488810 1340 488816 1352
rect 475896 1312 488816 1340
rect 475896 1300 475902 1312
rect 488810 1300 488816 1312
rect 488868 1300 488874 1352
rect 493502 1300 493508 1352
rect 493560 1340 493566 1352
rect 500034 1340 500040 1352
rect 493560 1312 500040 1340
rect 493560 1300 493566 1312
rect 500034 1300 500040 1312
rect 500092 1300 500098 1352
rect 500126 1300 500132 1352
rect 500184 1340 500190 1352
rect 507026 1340 507032 1352
rect 500184 1312 507032 1340
rect 500184 1300 500190 1312
rect 507026 1300 507032 1312
rect 507084 1300 507090 1352
rect 516686 1300 516692 1352
rect 516744 1340 516750 1352
rect 532050 1340 532056 1352
rect 516744 1312 532056 1340
rect 516744 1300 516750 1312
rect 532050 1300 532056 1312
rect 532108 1300 532114 1352
rect 539870 1300 539876 1352
rect 539928 1340 539934 1352
rect 546494 1340 546500 1352
rect 539928 1312 546500 1340
rect 539928 1300 539934 1312
rect 546494 1300 546500 1312
rect 546552 1300 546558 1352
rect 100754 1232 100760 1284
rect 100812 1272 100818 1284
rect 107010 1272 107016 1284
rect 100812 1244 107016 1272
rect 100812 1232 100818 1244
rect 107010 1232 107016 1244
rect 107068 1232 107074 1284
rect 110506 1232 110512 1284
rect 110564 1272 110570 1284
rect 116946 1272 116952 1284
rect 110564 1244 116952 1272
rect 110564 1232 110570 1244
rect 116946 1232 116952 1244
rect 117004 1232 117010 1284
rect 258258 1232 258264 1284
rect 258316 1272 258322 1284
rect 260466 1272 260472 1284
rect 258316 1244 260472 1272
rect 258316 1232 258322 1244
rect 260466 1232 260472 1244
rect 260524 1232 260530 1284
rect 264146 1232 264152 1284
rect 264204 1272 264210 1284
rect 265986 1272 265992 1284
rect 264204 1244 265992 1272
rect 264204 1232 264210 1244
rect 265986 1232 265992 1244
rect 266044 1232 266050 1284
rect 266538 1232 266544 1284
rect 266596 1272 266602 1284
rect 268194 1272 268200 1284
rect 266596 1244 268200 1272
rect 266596 1232 266602 1244
rect 268194 1232 268200 1244
rect 268252 1232 268258 1284
rect 270034 1232 270040 1284
rect 270092 1272 270098 1284
rect 271506 1272 271512 1284
rect 270092 1244 271512 1272
rect 270092 1232 270098 1244
rect 271506 1232 271512 1244
rect 271564 1232 271570 1284
rect 272426 1232 272432 1284
rect 272484 1272 272490 1284
rect 273714 1272 273720 1284
rect 272484 1244 273720 1272
rect 272484 1232 272490 1244
rect 273714 1232 273720 1244
rect 273772 1232 273778 1284
rect 343358 1232 343364 1284
rect 343416 1272 343422 1284
rect 346946 1272 346952 1284
rect 343416 1244 346952 1272
rect 343416 1232 343422 1244
rect 346946 1232 346952 1244
rect 347004 1232 347010 1284
rect 349982 1232 349988 1284
rect 350040 1272 350046 1284
rect 354030 1272 354036 1284
rect 350040 1244 354036 1272
rect 350040 1232 350046 1244
rect 354030 1232 354036 1244
rect 354088 1232 354094 1284
rect 357710 1232 357716 1284
rect 357768 1272 357774 1284
rect 362310 1272 362316 1284
rect 357768 1244 362316 1272
rect 357768 1232 357774 1244
rect 362310 1232 362316 1244
rect 362368 1232 362374 1284
rect 365438 1232 365444 1284
rect 365496 1272 365502 1284
rect 370222 1272 370228 1284
rect 365496 1244 370228 1272
rect 365496 1232 365502 1244
rect 370222 1232 370228 1244
rect 370280 1232 370286 1284
rect 370958 1232 370964 1284
rect 371016 1272 371022 1284
rect 376110 1272 376116 1284
rect 371016 1244 376116 1272
rect 371016 1232 371022 1244
rect 376110 1232 376116 1244
rect 376168 1232 376174 1284
rect 378686 1232 378692 1284
rect 378744 1272 378750 1284
rect 384390 1272 384396 1284
rect 378744 1244 384396 1272
rect 378744 1232 378750 1244
rect 384390 1232 384396 1244
rect 384448 1232 384454 1284
rect 387518 1232 387524 1284
rect 387576 1272 387582 1284
rect 394234 1272 394240 1284
rect 387576 1244 394240 1272
rect 387576 1232 387582 1244
rect 394234 1232 394240 1244
rect 394292 1232 394298 1284
rect 396350 1232 396356 1284
rect 396408 1272 396414 1284
rect 403618 1272 403624 1284
rect 396408 1244 403624 1272
rect 396408 1232 396414 1244
rect 403618 1232 403624 1244
rect 403676 1232 403682 1284
rect 404078 1232 404084 1284
rect 404136 1272 404142 1284
rect 411898 1272 411904 1284
rect 404136 1244 411904 1272
rect 404136 1232 404142 1244
rect 411898 1232 411904 1244
rect 411956 1232 411962 1284
rect 430482 1232 430488 1284
rect 430540 1272 430546 1284
rect 439958 1272 439964 1284
rect 430540 1244 439964 1272
rect 430540 1232 430546 1244
rect 439958 1232 439964 1244
rect 440016 1232 440022 1284
rect 447042 1232 447048 1284
rect 447100 1272 447106 1284
rect 456426 1272 456432 1284
rect 447100 1244 456432 1272
rect 447100 1232 447106 1244
rect 456426 1232 456432 1244
rect 456484 1232 456490 1284
rect 474642 1232 474648 1284
rect 474700 1272 474706 1284
rect 487246 1272 487252 1284
rect 474700 1244 487252 1272
rect 474700 1232 474706 1244
rect 487246 1232 487252 1244
rect 487304 1232 487310 1284
rect 499022 1232 499028 1284
rect 499080 1272 499086 1284
rect 499080 1244 509234 1272
rect 499080 1232 499086 1244
rect 268838 1164 268844 1216
rect 268896 1204 268902 1216
rect 270402 1204 270408 1216
rect 268896 1176 270408 1204
rect 268896 1164 268902 1176
rect 270402 1164 270408 1176
rect 270460 1164 270466 1216
rect 359918 1164 359924 1216
rect 359976 1204 359982 1216
rect 364610 1204 364616 1216
rect 359976 1176 364616 1204
rect 359976 1164 359982 1176
rect 364610 1164 364616 1176
rect 364668 1164 364674 1216
rect 368750 1164 368756 1216
rect 368808 1204 368814 1216
rect 373902 1204 373908 1216
rect 368808 1176 373908 1204
rect 368808 1164 368814 1176
rect 373902 1164 373908 1176
rect 373960 1164 373966 1216
rect 374270 1164 374276 1216
rect 374328 1204 374334 1216
rect 379606 1204 379612 1216
rect 374328 1176 379612 1204
rect 374328 1164 374334 1176
rect 379606 1164 379612 1176
rect 379664 1164 379670 1216
rect 379790 1164 379796 1216
rect 379848 1204 379854 1216
rect 385954 1204 385960 1216
rect 379848 1176 385960 1204
rect 379848 1164 379854 1176
rect 385954 1164 385960 1176
rect 386012 1164 386018 1216
rect 395246 1164 395252 1216
rect 395304 1204 395310 1216
rect 402514 1204 402520 1216
rect 395304 1176 402520 1204
rect 395304 1164 395310 1176
rect 402514 1164 402520 1176
rect 402572 1164 402578 1216
rect 443822 1164 443828 1216
rect 443880 1204 443886 1216
rect 454126 1204 454132 1216
rect 443880 1176 454132 1204
rect 443880 1164 443886 1176
rect 454126 1164 454132 1176
rect 454184 1164 454190 1216
rect 457070 1164 457076 1216
rect 457128 1204 457134 1216
rect 468294 1204 468300 1216
rect 457128 1176 468300 1204
rect 457128 1164 457134 1176
rect 468294 1164 468300 1176
rect 468352 1164 468358 1216
rect 469122 1164 469128 1216
rect 469180 1204 469186 1216
rect 481358 1204 481364 1216
rect 469180 1176 481364 1204
rect 469180 1164 469186 1176
rect 481358 1164 481364 1176
rect 481416 1164 481422 1216
rect 490190 1164 490196 1216
rect 490248 1204 490254 1216
rect 503806 1204 503812 1216
rect 490248 1176 503812 1204
rect 490248 1164 490254 1176
rect 503806 1164 503812 1176
rect 503864 1164 503870 1216
rect 509206 1204 509234 1244
rect 512270 1232 512276 1284
rect 512328 1272 512334 1284
rect 527818 1272 527824 1284
rect 512328 1244 527824 1272
rect 512328 1232 512334 1244
rect 527818 1232 527824 1244
rect 527876 1232 527882 1284
rect 513374 1204 513380 1216
rect 509206 1176 513380 1204
rect 513374 1164 513380 1176
rect 513432 1164 513438 1216
rect 517790 1164 517796 1216
rect 517848 1204 517854 1216
rect 533706 1204 533712 1216
rect 517848 1176 533712 1204
rect 517848 1164 517854 1176
rect 533706 1164 533712 1176
rect 533764 1164 533770 1216
rect 352190 1096 352196 1148
rect 352248 1136 352254 1148
rect 356330 1136 356336 1148
rect 352248 1108 356336 1136
rect 352248 1096 352254 1108
rect 356330 1096 356336 1108
rect 356388 1096 356394 1148
rect 361022 1096 361028 1148
rect 361080 1136 361086 1148
rect 365438 1136 365444 1148
rect 361080 1108 365444 1136
rect 361080 1096 361086 1108
rect 365438 1096 365444 1108
rect 365496 1096 365502 1148
rect 366542 1096 366548 1148
rect 366600 1136 366606 1148
rect 371326 1136 371332 1148
rect 366600 1108 371332 1136
rect 366600 1096 366606 1108
rect 371326 1096 371332 1108
rect 371384 1096 371390 1148
rect 375190 1096 375196 1148
rect 375248 1136 375254 1148
rect 381170 1136 381176 1148
rect 375248 1108 381176 1136
rect 375248 1096 375254 1108
rect 381170 1096 381176 1108
rect 381228 1096 381234 1148
rect 385310 1096 385316 1148
rect 385368 1136 385374 1148
rect 391842 1136 391848 1148
rect 385368 1108 391848 1136
rect 385368 1096 385374 1108
rect 391842 1096 391848 1108
rect 391900 1096 391906 1148
rect 397362 1096 397368 1148
rect 397420 1136 397426 1148
rect 404814 1136 404820 1148
rect 397420 1108 404820 1136
rect 397420 1096 397426 1108
rect 404814 1096 404820 1108
rect 404872 1096 404878 1148
rect 412910 1096 412916 1148
rect 412968 1136 412974 1148
rect 421374 1136 421380 1148
rect 412968 1108 421380 1136
rect 412968 1096 412974 1108
rect 421374 1096 421380 1108
rect 421432 1096 421438 1148
rect 437198 1096 437204 1148
rect 437256 1136 437262 1148
rect 447410 1136 447416 1148
rect 437256 1108 447416 1136
rect 437256 1096 437262 1108
rect 447410 1096 447416 1108
rect 447468 1096 447474 1148
rect 485682 1096 485688 1148
rect 485740 1136 485746 1148
rect 499022 1136 499028 1148
rect 485740 1108 499028 1136
rect 485740 1096 485746 1108
rect 499022 1096 499028 1108
rect 499080 1096 499086 1148
rect 500402 1096 500408 1148
rect 500460 1136 500466 1148
rect 500460 1108 510568 1136
rect 500460 1096 500466 1108
rect 355502 1028 355508 1080
rect 355560 1068 355566 1080
rect 359918 1068 359924 1080
rect 355560 1040 359924 1068
rect 355560 1028 355566 1040
rect 359918 1028 359924 1040
rect 359976 1028 359982 1080
rect 367646 1028 367652 1080
rect 367704 1068 367710 1080
rect 372890 1068 372896 1080
rect 367704 1040 372896 1068
rect 367704 1028 367710 1040
rect 372890 1028 372896 1040
rect 372948 1028 372954 1080
rect 377582 1028 377588 1080
rect 377640 1068 377646 1080
rect 383562 1068 383568 1080
rect 377640 1040 383568 1068
rect 377640 1028 377646 1040
rect 383562 1028 383568 1040
rect 383620 1028 383626 1080
rect 451550 1028 451556 1080
rect 451608 1068 451614 1080
rect 462406 1068 462412 1080
rect 451608 1040 462412 1068
rect 451608 1028 451614 1040
rect 462406 1028 462412 1040
rect 462464 1028 462470 1080
rect 489086 1028 489092 1080
rect 489144 1068 489150 1080
rect 502978 1068 502984 1080
rect 489144 1040 502984 1068
rect 489144 1028 489150 1040
rect 502978 1028 502984 1040
rect 503036 1028 503042 1080
rect 503438 1028 503444 1080
rect 503496 1068 503502 1080
rect 510540 1068 510568 1108
rect 511166 1096 511172 1148
rect 511224 1136 511230 1148
rect 526254 1136 526260 1148
rect 511224 1108 526260 1136
rect 511224 1096 511230 1108
rect 526254 1096 526260 1108
rect 526312 1096 526318 1148
rect 512086 1068 512092 1080
rect 503496 1040 510476 1068
rect 510540 1040 512092 1068
rect 503496 1028 503502 1040
rect 21818 960 21824 1012
rect 21876 1000 21882 1012
rect 39666 1000 39672 1012
rect 21876 972 39672 1000
rect 21876 960 21882 972
rect 39666 960 39672 972
rect 39724 960 39730 1012
rect 345566 960 345572 1012
rect 345624 1000 345630 1012
rect 349246 1000 349252 1012
rect 345624 972 349252 1000
rect 345624 960 345630 972
rect 349246 960 349252 972
rect 349304 960 349310 1012
rect 351086 960 351092 1012
rect 351144 1000 351150 1012
rect 355226 1000 355232 1012
rect 351144 972 355232 1000
rect 351144 960 351150 972
rect 355226 960 355232 972
rect 355284 960 355290 1012
rect 362126 960 362132 1012
rect 362184 1000 362190 1012
rect 367002 1000 367008 1012
rect 362184 972 367008 1000
rect 362184 960 362190 972
rect 367002 960 367008 972
rect 367060 960 367066 1012
rect 373166 960 373172 1012
rect 373224 1000 373230 1012
rect 378502 1000 378508 1012
rect 373224 972 378508 1000
rect 373224 960 373230 972
rect 378502 960 378508 972
rect 378560 960 378566 1012
rect 416222 960 416228 1012
rect 416280 1000 416286 1012
rect 424962 1000 424968 1012
rect 416280 972 424968 1000
rect 416280 960 416286 972
rect 424962 960 424968 972
rect 425020 960 425026 1012
rect 448238 960 448244 1012
rect 448296 1000 448302 1012
rect 459186 1000 459192 1012
rect 448296 972 459192 1000
rect 448296 960 448302 972
rect 459186 960 459192 972
rect 459244 960 459250 1012
rect 482462 960 482468 1012
rect 482520 1000 482526 1012
rect 495526 1000 495532 1012
rect 482520 972 495532 1000
rect 482520 960 482526 972
rect 495526 960 495532 972
rect 495584 960 495590 1012
rect 495710 960 495716 1012
rect 495768 1000 495774 1012
rect 509694 1000 509700 1012
rect 495768 972 509700 1000
rect 495768 960 495774 972
rect 509694 960 509700 972
rect 509752 960 509758 1012
rect 510448 1000 510476 1040
rect 512086 1028 512092 1040
rect 512144 1028 512150 1080
rect 517974 1000 517980 1012
rect 510448 972 517980 1000
rect 517974 960 517980 972
rect 518032 960 518038 1012
rect 534350 960 534356 1012
rect 534408 1000 534414 1012
rect 551462 1000 551468 1012
rect 534408 972 551468 1000
rect 534408 960 534414 972
rect 551462 960 551468 972
rect 551520 960 551526 1012
rect 19426 892 19432 944
rect 19484 932 19490 944
rect 37458 932 37464 944
rect 19484 904 37464 932
rect 19484 892 19490 904
rect 37458 892 37464 904
rect 37516 892 37522 944
rect 358722 892 358728 944
rect 358780 932 358786 944
rect 363506 932 363512 944
rect 358780 904 363512 932
rect 358780 892 358786 904
rect 363506 892 363512 904
rect 363564 892 363570 944
rect 444926 892 444932 944
rect 444984 932 444990 944
rect 455690 932 455696 944
rect 444984 904 455696 932
rect 444984 892 444990 904
rect 455690 892 455696 904
rect 455748 892 455754 944
rect 455966 892 455972 944
rect 456024 932 456030 944
rect 467466 932 467472 944
rect 456024 904 467472 932
rect 456024 892 456030 904
rect 467466 892 467472 904
rect 467524 892 467530 944
rect 480162 892 480168 944
rect 480220 932 480226 944
rect 493134 932 493140 944
rect 480220 904 493140 932
rect 480220 892 480226 904
rect 493134 892 493140 904
rect 493192 892 493198 944
rect 494606 892 494612 944
rect 494664 932 494670 944
rect 508866 932 508872 944
rect 494664 904 508872 932
rect 494664 892 494670 904
rect 508866 892 508872 904
rect 508924 892 508930 944
rect 510062 892 510068 944
rect 510120 932 510126 944
rect 525426 932 525432 944
rect 510120 904 525432 932
rect 510120 892 510126 904
rect 525426 892 525432 904
rect 525484 892 525490 944
rect 532142 892 532148 944
rect 532200 932 532206 944
rect 549070 932 549076 944
rect 532200 904 549076 932
rect 532200 892 532206 904
rect 549070 892 549076 904
rect 549128 892 549134 944
rect 11146 824 11152 876
rect 11204 864 11210 876
rect 29730 864 29736 876
rect 11204 836 29736 864
rect 11204 824 11210 836
rect 29730 824 29736 836
rect 29788 824 29794 876
rect 337838 824 337844 876
rect 337896 864 337902 876
rect 340966 864 340972 876
rect 337896 836 340972 864
rect 337896 824 337902 836
rect 340966 824 340972 836
rect 341024 824 341030 876
rect 347682 824 347688 876
rect 347740 864 347746 876
rect 351638 864 351644 876
rect 347740 836 351644 864
rect 347740 824 347746 836
rect 351638 824 351644 836
rect 351696 824 351702 876
rect 441522 824 441528 876
rect 441580 864 441586 876
rect 451734 864 451740 876
rect 441580 836 451740 864
rect 441580 824 441586 836
rect 451734 824 451740 836
rect 451792 824 451798 876
rect 454862 824 454868 876
rect 454920 864 454926 876
rect 465902 864 465908 876
rect 454920 836 465908 864
rect 454920 824 454926 836
rect 465902 824 465908 836
rect 465960 824 465966 876
rect 492398 824 492404 876
rect 492456 864 492462 876
rect 506474 864 506480 876
rect 492456 836 506480 864
rect 492456 824 492462 836
rect 506474 824 506480 836
rect 506532 824 506538 876
rect 508958 824 508964 876
rect 509016 864 509022 876
rect 523862 864 523868 876
rect 509016 836 523868 864
rect 509016 824 509022 836
rect 523862 824 523868 836
rect 523920 824 523926 876
rect 550910 824 550916 876
rect 550968 864 550974 876
rect 569126 864 569132 876
rect 550968 836 569132 864
rect 550968 824 550974 836
rect 569126 824 569132 836
rect 569184 824 569190 876
rect 20622 756 20628 808
rect 20680 796 20686 808
rect 38562 796 38568 808
rect 20680 768 38568 796
rect 20680 756 20686 768
rect 38562 756 38568 768
rect 38620 756 38626 808
rect 251174 756 251180 808
rect 251232 796 251238 808
rect 253842 796 253848 808
rect 251232 768 253848 796
rect 251232 756 251238 768
rect 253842 756 253848 768
rect 253900 756 253906 808
rect 438302 756 438308 808
rect 438360 796 438366 808
rect 448238 796 448244 808
rect 438360 768 448244 796
rect 438360 756 438366 768
rect 448238 756 448244 768
rect 448296 756 448302 808
rect 449342 756 449348 808
rect 449400 796 449406 808
rect 460014 796 460020 808
rect 449400 768 460020 796
rect 449400 756 449406 768
rect 460014 756 460020 768
rect 460072 756 460078 808
rect 483566 756 483572 808
rect 483624 796 483630 808
rect 497090 796 497096 808
rect 483624 768 497096 796
rect 483624 756 483630 768
rect 497090 756 497096 768
rect 497148 756 497154 808
rect 502242 756 502248 808
rect 502300 796 502306 808
rect 502300 768 506980 796
rect 502300 756 502306 768
rect 14734 688 14740 740
rect 14792 728 14798 740
rect 33042 728 33048 740
rect 14792 700 33048 728
rect 14792 688 14798 700
rect 33042 688 33048 700
rect 33100 688 33106 740
rect 36354 728 36360 740
rect 35866 700 36360 728
rect 18230 620 18236 672
rect 18288 660 18294 672
rect 35866 660 35894 700
rect 36354 688 36360 700
rect 36412 688 36418 740
rect 386322 688 386328 740
rect 386380 728 386386 740
rect 392670 728 392676 740
rect 386380 700 392676 728
rect 386380 688 386386 700
rect 392670 688 392676 700
rect 392728 688 392734 740
rect 408402 688 408408 740
rect 408460 728 408466 740
rect 416682 728 416688 740
rect 408460 700 416688 728
rect 408460 688 408466 700
rect 416682 688 416688 700
rect 416740 688 416746 740
rect 423950 688 423956 740
rect 424008 728 424014 740
rect 433242 728 433248 740
rect 424008 700 433248 728
rect 424008 688 424014 700
rect 433242 688 433248 700
rect 433300 688 433306 740
rect 446030 688 446036 740
rect 446088 728 446094 740
rect 456518 728 456524 740
rect 446088 700 456524 728
rect 446088 688 446094 700
rect 456518 688 456524 700
rect 456576 688 456582 740
rect 480530 728 480536 740
rect 470566 700 480536 728
rect 18288 632 35894 660
rect 18288 620 18294 632
rect 35986 620 35992 672
rect 36044 660 36050 672
rect 52914 660 52920 672
rect 36044 632 52920 660
rect 36044 620 36050 632
rect 52914 620 52920 632
rect 52972 620 52978 672
rect 393038 620 393044 672
rect 393096 660 393102 672
rect 400122 660 400128 672
rect 393096 632 400128 660
rect 393096 620 393102 632
rect 400122 620 400128 632
rect 400180 620 400186 672
rect 400766 620 400772 672
rect 400824 660 400830 672
rect 400824 632 408448 660
rect 400824 620 400830 632
rect 408420 604 408448 632
rect 409598 620 409604 672
rect 409656 660 409662 672
rect 417878 660 417884 672
rect 409656 632 417884 660
rect 409656 620 409662 632
rect 417878 620 417884 632
rect 417936 620 417942 672
rect 418430 620 418436 672
rect 418488 660 418494 672
rect 427262 660 427268 672
rect 418488 632 427268 660
rect 418488 620 418494 632
rect 427262 620 427268 632
rect 427320 620 427326 672
rect 442718 620 442724 672
rect 442776 660 442782 672
rect 453298 660 453304 672
rect 442776 632 453304 660
rect 442776 620 442782 632
rect 453298 620 453304 632
rect 453356 620 453362 672
rect 468110 620 468116 672
rect 468168 660 468174 672
rect 470566 660 470594 700
rect 480530 688 480536 700
rect 480588 688 480594 740
rect 487982 688 487988 740
rect 488040 728 488046 740
rect 501414 728 501420 740
rect 488040 700 501420 728
rect 488040 688 488046 700
rect 501414 688 501420 700
rect 501472 688 501478 740
rect 504542 688 504548 740
rect 504600 728 504606 740
rect 506952 728 506980 768
rect 507026 756 507032 808
rect 507084 796 507090 808
rect 514754 796 514760 808
rect 507084 768 514760 796
rect 507084 756 507090 768
rect 514754 756 514760 768
rect 514812 756 514818 808
rect 527726 756 527732 808
rect 527784 796 527790 808
rect 544378 796 544384 808
rect 527784 768 544384 796
rect 527784 756 527790 768
rect 544378 756 544384 768
rect 544436 756 544442 808
rect 547598 756 547604 808
rect 547656 796 547662 808
rect 565630 796 565636 808
rect 547656 768 565636 796
rect 547656 756 547662 768
rect 565630 756 565636 768
rect 565688 756 565694 808
rect 517146 728 517152 740
rect 504600 700 506888 728
rect 506952 700 517152 728
rect 504600 688 504606 700
rect 476942 660 476948 672
rect 468168 632 470594 660
rect 473372 632 476948 660
rect 468168 620 468174 632
rect 15930 552 15936 604
rect 15988 592 15994 604
rect 34146 592 34152 604
rect 15988 564 34152 592
rect 15988 552 15994 564
rect 34146 552 34152 564
rect 34204 552 34210 604
rect 34790 552 34796 604
rect 34848 592 34854 604
rect 51810 592 51816 604
rect 34848 564 51816 592
rect 34848 552 34854 564
rect 51810 552 51816 564
rect 51868 552 51874 604
rect 388622 552 388628 604
rect 388680 592 388686 604
rect 395338 592 395344 604
rect 388680 564 395344 592
rect 388680 552 388686 564
rect 395338 552 395344 564
rect 395396 552 395402 604
rect 408402 552 408408 604
rect 408460 552 408466 604
rect 426158 552 426164 604
rect 426216 592 426222 604
rect 435542 592 435548 604
rect 426216 564 435548 592
rect 426216 552 426222 564
rect 435542 552 435548 564
rect 435600 552 435606 604
rect 439130 552 439136 604
rect 439188 552 439194 604
rect 464798 552 464804 604
rect 464856 592 464862 604
rect 473372 592 473400 632
rect 476942 620 476948 632
rect 477000 620 477006 672
rect 481542 620 481548 672
rect 481600 660 481606 672
rect 494698 660 494704 672
rect 481600 632 494704 660
rect 481600 620 481606 632
rect 494698 620 494704 632
rect 494756 620 494762 672
rect 497918 620 497924 672
rect 497976 660 497982 672
rect 500402 660 500408 672
rect 497976 632 500408 660
rect 497976 620 497982 632
rect 500402 620 500408 632
rect 500460 620 500466 672
rect 505370 660 505376 672
rect 500512 632 505376 660
rect 464856 564 473400 592
rect 464856 552 464862 564
rect 473446 552 473452 604
rect 473504 552 473510 604
rect 486418 552 486424 604
rect 486476 552 486482 604
rect 491202 552 491208 604
rect 491260 592 491266 604
rect 500512 592 500540 632
rect 505370 620 505376 632
rect 505428 620 505434 672
rect 506860 660 506888 700
rect 517146 688 517152 700
rect 517204 688 517210 740
rect 524322 688 524328 740
rect 524380 728 524386 740
rect 540790 728 540796 740
rect 524380 700 540796 728
rect 524380 688 524386 700
rect 540790 688 540796 700
rect 540848 688 540854 740
rect 540882 688 540888 740
rect 540940 728 540946 740
rect 558546 728 558552 740
rect 540940 700 558552 728
rect 540940 688 540946 700
rect 558546 688 558552 700
rect 558604 688 558610 740
rect 506860 632 509234 660
rect 491260 564 500540 592
rect 491260 552 491266 564
rect 500586 552 500592 604
rect 500644 552 500650 604
rect 509206 592 509234 632
rect 525518 620 525524 672
rect 525576 660 525582 672
rect 541986 660 541992 672
rect 525576 632 541992 660
rect 525576 620 525582 632
rect 541986 620 541992 632
rect 542044 620 542050 672
rect 545390 620 545396 672
rect 545448 660 545454 672
rect 563238 660 563244 672
rect 545448 632 563244 660
rect 545448 620 545454 632
rect 563238 620 563244 632
rect 563296 620 563302 672
rect 519538 592 519544 604
rect 509206 564 519544 592
rect 519538 552 519544 564
rect 519596 552 519602 604
rect 522206 552 522212 604
rect 522264 592 522270 604
rect 538398 592 538404 604
rect 522264 564 538404 592
rect 522264 552 522270 564
rect 538398 552 538404 564
rect 538456 552 538462 604
rect 542078 552 542084 604
rect 542136 592 542142 604
rect 559742 592 559748 604
rect 542136 564 559748 592
rect 542136 552 542142 564
rect 559742 552 559748 564
rect 559800 552 559806 604
rect 562042 552 562048 604
rect 562100 552 562106 604
rect 3234 484 3240 536
rect 3292 524 3298 536
rect 22002 524 22008 536
rect 3292 496 22008 524
rect 3292 484 3298 496
rect 22002 484 22008 496
rect 22060 484 22066 536
rect 22830 484 22836 536
rect 22888 524 22894 536
rect 40494 524 40500 536
rect 22888 496 40500 524
rect 22888 484 22894 496
rect 40494 484 40500 496
rect 40552 484 40558 536
rect 45278 484 45284 536
rect 45336 524 45342 536
rect 61746 524 61752 536
rect 45336 496 61752 524
rect 45336 484 45342 496
rect 61746 484 61752 496
rect 61804 484 61810 536
rect 420638 484 420644 536
rect 420696 524 420702 536
rect 429286 524 429292 536
rect 420696 496 429292 524
rect 420696 484 420702 496
rect 429286 484 429292 496
rect 429344 484 429350 536
rect 429470 484 429476 536
rect 429528 524 429534 536
rect 439148 524 439176 552
rect 429528 496 439176 524
rect 429528 484 429534 496
rect 461762 484 461768 536
rect 461820 524 461826 536
rect 473464 524 473492 552
rect 461820 496 473492 524
rect 461820 484 461826 496
rect 473630 484 473636 536
rect 473688 524 473694 536
rect 486436 524 486464 552
rect 473688 496 486464 524
rect 473688 484 473694 496
rect 486878 484 486884 536
rect 486936 524 486942 536
rect 500604 524 500632 552
rect 486936 496 500632 524
rect 486936 484 486942 496
rect 501230 484 501236 536
rect 501288 524 501294 536
rect 515582 524 515588 536
rect 501288 496 515588 524
rect 501288 484 501294 496
rect 515582 484 515588 496
rect 515640 484 515646 536
rect 518802 484 518808 536
rect 518860 524 518866 536
rect 534534 524 534540 536
rect 518860 496 534540 524
rect 518860 484 518866 496
rect 534534 484 534540 496
rect 534592 484 534598 536
rect 544562 484 544568 536
rect 544620 524 544626 536
rect 562060 524 562088 552
rect 544620 496 562088 524
rect 544620 484 544626 496
rect 9122 416 9128 468
rect 9180 456 9186 468
rect 27522 456 27528 468
rect 9180 428 27528 456
rect 9180 416 9186 428
rect 27522 416 27528 428
rect 27580 416 27586 468
rect 32214 416 32220 468
rect 32272 456 32278 468
rect 49602 456 49608 468
rect 32272 428 49608 456
rect 32272 416 32278 428
rect 49602 416 49608 428
rect 49660 416 49666 468
rect 401870 416 401876 468
rect 401928 456 401934 468
rect 409230 456 409236 468
rect 401928 428 409236 456
rect 401928 416 401934 428
rect 409230 416 409236 428
rect 409288 416 409294 468
rect 424778 416 424784 468
rect 424836 456 424842 468
rect 434070 456 434076 468
rect 424836 428 434076 456
rect 424836 416 424842 428
rect 434070 416 434076 428
rect 434128 416 434134 468
rect 434990 416 434996 468
rect 435048 456 435054 468
rect 445202 456 445208 468
rect 435048 428 445208 456
rect 435048 416 435054 428
rect 445202 416 445208 428
rect 445260 416 445266 468
rect 457898 416 457904 468
rect 457956 456 457962 468
rect 470042 456 470048 468
rect 457956 428 470048 456
rect 457956 416 457962 428
rect 470042 416 470048 428
rect 470100 416 470106 468
rect 470318 416 470324 468
rect 470376 456 470382 468
rect 482462 456 482468 468
rect 470376 428 482468 456
rect 470376 416 470382 428
rect 482462 416 482468 428
rect 482520 416 482526 468
rect 500034 416 500040 468
rect 500092 456 500098 468
rect 507302 456 507308 468
rect 500092 428 507308 456
rect 500092 416 500098 428
rect 507302 416 507308 428
rect 507360 416 507366 468
rect 507854 416 507860 468
rect 507912 456 507918 468
rect 523218 456 523224 468
rect 507912 428 523224 456
rect 507912 416 507918 428
rect 523218 416 523224 428
rect 523276 416 523282 468
rect 528830 416 528836 468
rect 528888 456 528894 468
rect 545666 456 545672 468
rect 528888 428 545672 456
rect 528888 416 528894 428
rect 545666 416 545672 428
rect 545724 416 545730 468
rect 548702 416 548708 468
rect 548760 456 548766 468
rect 567010 456 567016 468
rect 548760 428 567016 456
rect 548760 416 548766 428
rect 567010 416 567016 428
rect 567068 416 567074 468
rect 9766 348 9772 400
rect 9824 388 9830 400
rect 28626 388 28632 400
rect 9824 360 28632 388
rect 9824 348 9830 360
rect 28626 348 28632 360
rect 28684 348 28690 400
rect 39390 348 39396 400
rect 39448 388 39454 400
rect 56226 388 56232 400
rect 39448 360 56232 388
rect 39448 348 39454 360
rect 56226 348 56232 360
rect 56284 348 56290 400
rect 407390 348 407396 400
rect 407448 388 407454 400
rect 415302 388 415308 400
rect 407448 360 415308 388
rect 407448 348 407454 360
rect 415302 348 415308 360
rect 415360 348 415366 400
rect 417326 348 417332 400
rect 417384 388 417390 400
rect 425790 388 425796 400
rect 417384 360 425796 388
rect 417384 348 417390 360
rect 425790 348 425796 360
rect 425848 348 425854 400
rect 428642 348 428648 400
rect 428700 388 428706 400
rect 437566 388 437572 400
rect 428700 360 437572 388
rect 428700 348 428706 360
rect 437566 348 437572 360
rect 437624 348 437630 400
rect 459462 348 459468 400
rect 459520 388 459526 400
rect 470778 388 470784 400
rect 459520 360 470784 388
rect 459520 348 459526 360
rect 470778 348 470784 360
rect 470836 348 470842 400
rect 472526 348 472532 400
rect 472584 388 472590 400
rect 484854 388 484860 400
rect 472584 360 484860 388
rect 472584 348 472590 360
rect 484854 348 484860 360
rect 484912 348 484918 400
rect 496722 348 496728 400
rect 496780 388 496786 400
rect 511442 388 511448 400
rect 496780 360 511448 388
rect 496780 348 496786 360
rect 511442 348 511448 360
rect 511500 348 511506 400
rect 514478 348 514484 400
rect 514536 388 514542 400
rect 529934 388 529940 400
rect 514536 360 529940 388
rect 514536 348 514542 360
rect 529934 348 529940 360
rect 529992 348 529998 400
rect 533246 348 533252 400
rect 533304 388 533310 400
rect 550450 388 550456 400
rect 533304 360 550456 388
rect 533304 348 533310 360
rect 550450 348 550456 360
rect 550508 348 550514 400
rect 555326 348 555332 400
rect 555384 388 555390 400
rect 573542 388 573548 400
rect 555384 360 573548 388
rect 555384 348 555390 360
rect 573542 348 573548 360
rect 573600 348 573606 400
rect 17402 280 17408 332
rect 17460 320 17466 332
rect 35250 320 35256 332
rect 17460 292 35256 320
rect 17460 280 17466 292
rect 35250 280 35256 292
rect 35308 280 35314 332
rect 38562 280 38568 332
rect 38620 320 38626 332
rect 55122 320 55128 332
rect 38620 292 55128 320
rect 38620 280 38626 292
rect 55122 280 55128 292
rect 55180 280 55186 332
rect 381998 280 382004 332
rect 382056 320 382062 332
rect 387886 320 387892 332
rect 382056 292 387892 320
rect 382056 280 382062 292
rect 387886 280 387892 292
rect 387944 280 387950 332
rect 389726 280 389732 332
rect 389784 320 389790 332
rect 396166 320 396172 332
rect 389784 292 396172 320
rect 389784 280 389790 292
rect 396166 280 396172 292
rect 396224 280 396230 332
rect 413922 280 413928 332
rect 413980 320 413986 332
rect 422754 320 422760 332
rect 413980 292 422760 320
rect 413980 280 413986 292
rect 422754 280 422760 292
rect 422812 280 422818 332
rect 427538 280 427544 332
rect 427596 320 427602 332
rect 436922 320 436928 332
rect 427596 292 436928 320
rect 427596 280 427602 292
rect 436922 280 436928 292
rect 436980 280 436986 332
rect 440510 280 440516 332
rect 440568 320 440574 332
rect 451090 320 451096 332
rect 440568 292 451096 320
rect 440568 280 440574 292
rect 451090 280 451096 292
rect 451148 280 451154 332
rect 467006 280 467012 332
rect 467064 320 467070 332
rect 478966 320 478972 332
rect 467064 292 478972 320
rect 467064 280 467070 292
rect 478966 280 478972 292
rect 479024 280 479030 332
rect 479518 280 479524 332
rect 479576 320 479582 332
rect 492490 320 492496 332
rect 479576 292 492496 320
rect 479576 280 479582 292
rect 492490 280 492496 292
rect 492548 280 492554 332
rect 505646 280 505652 332
rect 505704 320 505710 332
rect 520366 320 520372 332
rect 505704 292 520372 320
rect 505704 280 505710 292
rect 520366 280 520372 292
rect 520424 280 520430 332
rect 521102 280 521108 332
rect 521160 320 521166 332
rect 537386 320 537392 332
rect 521160 292 537392 320
rect 521160 280 521166 292
rect 537386 280 537392 292
rect 537444 280 537450 332
rect 538766 280 538772 332
rect 538824 320 538830 332
rect 556338 320 556344 332
rect 538824 292 556344 320
rect 538824 280 538830 292
rect 556338 280 556344 292
rect 556396 280 556402 332
rect 557166 280 557172 332
rect 557224 320 557230 332
rect 575934 320 575940 332
rect 557224 292 575940 320
rect 557224 280 557230 292
rect 575934 280 575940 292
rect 575992 280 575998 332
rect 3878 212 3884 264
rect 3936 252 3942 264
rect 23198 252 23204 264
rect 3936 224 23204 252
rect 3936 212 3942 224
rect 23198 212 23204 224
rect 23256 212 23262 264
rect 42242 212 42248 264
rect 42300 252 42306 264
rect 58158 252 58164 264
rect 42300 224 58164 252
rect 42300 212 42306 224
rect 58158 212 58164 224
rect 58216 212 58222 264
rect 390830 212 390836 264
rect 390888 252 390894 264
rect 397914 252 397920 264
rect 390888 224 397920 252
rect 390888 212 390894 224
rect 397914 212 397920 224
rect 397972 212 397978 264
rect 402882 212 402888 264
rect 402940 252 402946 264
rect 410978 252 410984 264
rect 402940 224 410984 252
rect 402940 212 402946 224
rect 410978 212 410984 224
rect 411036 212 411042 264
rect 415118 212 415124 264
rect 415176 252 415182 264
rect 423582 252 423588 264
rect 415176 224 423588 252
rect 415176 212 415182 224
rect 423582 212 423588 224
rect 423640 212 423646 264
rect 432782 212 432788 264
rect 432840 252 432846 264
rect 442810 252 442816 264
rect 432840 224 442816 252
rect 432840 212 432846 224
rect 442810 212 442816 224
rect 442868 212 442874 264
rect 456426 212 456432 264
rect 456484 252 456490 264
rect 458266 252 458272 264
rect 456484 224 458272 252
rect 456484 212 456490 224
rect 458266 212 458272 224
rect 458324 212 458330 264
rect 460566 212 460572 264
rect 460624 252 460630 264
rect 472434 252 472440 264
rect 460624 224 472440 252
rect 460624 212 460630 224
rect 472434 212 472440 224
rect 472492 212 472498 264
rect 478322 212 478328 264
rect 478380 252 478386 264
rect 490742 252 490748 264
rect 478380 224 490748 252
rect 478380 212 478386 224
rect 490742 212 490748 224
rect 490800 212 490806 264
rect 515490 212 515496 264
rect 515548 252 515554 264
rect 531498 252 531504 264
rect 515548 224 531504 252
rect 515548 212 515554 224
rect 531498 212 531504 224
rect 531556 212 531562 264
rect 535362 212 535368 264
rect 535420 252 535426 264
rect 552842 252 552848 264
rect 535420 224 552848 252
rect 535420 212 535426 224
rect 552842 212 552848 224
rect 552900 212 552906 264
rect 554222 212 554228 264
rect 554280 252 554286 264
rect 572898 252 572904 264
rect 554280 224 572904 252
rect 554280 212 554286 224
rect 572898 212 572904 224
rect 572956 212 572962 264
rect 1486 144 1492 196
rect 1544 184 1550 196
rect 20898 184 20904 196
rect 1544 156 20904 184
rect 1544 144 1550 156
rect 20898 144 20904 156
rect 20956 144 20962 196
rect 24578 144 24584 196
rect 24636 184 24642 196
rect 41598 184 41604 196
rect 24636 156 41604 184
rect 24636 144 24642 156
rect 41598 144 41604 156
rect 41656 144 41662 196
rect 42886 144 42892 196
rect 42944 184 42950 196
rect 59354 184 59360 196
rect 42944 156 59360 184
rect 42944 144 42950 156
rect 59354 144 59360 156
rect 59412 144 59418 196
rect 380802 144 380808 196
rect 380860 184 380866 196
rect 386782 184 386788 196
rect 380860 156 386788 184
rect 380860 144 380866 156
rect 386782 144 386788 156
rect 386840 144 386846 196
rect 391658 144 391664 196
rect 391716 184 391722 196
rect 398742 184 398748 196
rect 391716 156 398748 184
rect 391716 144 391722 156
rect 398742 144 398748 156
rect 398800 144 398806 196
rect 405182 144 405188 196
rect 405240 184 405246 196
rect 412818 184 412824 196
rect 405240 156 412824 184
rect 405240 144 405246 156
rect 412818 144 412824 156
rect 412876 144 412882 196
rect 419442 144 419448 196
rect 419500 184 419506 196
rect 428642 184 428648 196
rect 419500 156 428648 184
rect 419500 144 419506 156
rect 428642 144 428648 156
rect 428700 144 428706 196
rect 431678 144 431684 196
rect 431736 184 431742 196
rect 441246 184 441252 196
rect 431736 156 441252 184
rect 431736 144 431742 156
rect 441246 144 441252 156
rect 441304 144 441310 196
rect 453758 144 453764 196
rect 453816 184 453822 196
rect 464982 184 464988 196
rect 453816 156 464988 184
rect 453816 144 453822 156
rect 464982 144 464988 156
rect 465040 144 465046 196
rect 471422 144 471428 196
rect 471480 184 471486 196
rect 484210 184 484216 196
rect 471480 156 484216 184
rect 471480 144 471486 156
rect 484210 144 484216 156
rect 484268 144 484274 196
rect 519998 144 520004 196
rect 520056 184 520062 196
rect 536282 184 536288 196
rect 520056 156 536288 184
rect 520056 144 520062 156
rect 536282 144 536288 156
rect 536340 144 536346 196
rect 537662 144 537668 196
rect 537720 184 537726 196
rect 554774 184 554780 196
rect 537720 156 554780 184
rect 537720 144 537726 156
rect 554774 144 554780 156
rect 554832 144 554838 196
rect 558822 144 558828 196
rect 558880 184 558886 196
rect 577130 184 577136 196
rect 558880 156 577136 184
rect 558880 144 558886 156
rect 577130 144 577136 156
rect 577188 144 577194 196
rect 8018 76 8024 128
rect 8076 116 8082 128
rect 26326 116 26332 128
rect 8076 88 26332 116
rect 8076 76 8082 88
rect 26326 76 26332 88
rect 26384 76 26390 128
rect 31110 76 31116 128
rect 31168 116 31174 128
rect 48498 116 48504 128
rect 31168 88 48504 116
rect 31168 76 31174 88
rect 48498 76 48504 88
rect 48556 76 48562 128
rect 344738 76 344744 128
rect 344796 116 344802 128
rect 348234 116 348240 128
rect 344796 88 348240 116
rect 344796 76 344802 88
rect 348234 76 348240 88
rect 348292 76 348298 128
rect 354398 76 354404 128
rect 354456 116 354462 128
rect 358906 116 358912 128
rect 354456 88 358912 116
rect 354456 76 354462 88
rect 358906 76 358912 88
rect 358964 76 358970 128
rect 383102 76 383108 128
rect 383160 116 383166 128
rect 389634 116 389640 128
rect 383160 88 389640 116
rect 383160 76 383166 88
rect 389634 76 389640 88
rect 389692 76 389698 128
rect 398558 76 398564 128
rect 398616 116 398622 128
rect 406194 116 406200 128
rect 398616 88 406200 116
rect 398616 76 398622 88
rect 406194 76 406200 88
rect 406252 76 406258 128
rect 412082 76 412088 128
rect 412140 116 412146 128
rect 420362 116 420368 128
rect 412140 88 420368 116
rect 412140 76 412146 88
rect 420362 76 420368 88
rect 420420 76 420426 128
rect 422846 76 422852 128
rect 422904 116 422910 128
rect 431862 116 431868 128
rect 422904 88 431868 116
rect 422904 76 422910 88
rect 431862 76 431868 88
rect 431920 76 431926 128
rect 433886 76 433892 128
rect 433944 116 433950 128
rect 443454 116 443460 128
rect 433944 88 443460 116
rect 433944 76 433950 88
rect 443454 76 443460 88
rect 443512 76 443518 128
rect 463602 76 463608 128
rect 463660 116 463666 128
rect 475930 116 475936 128
rect 463660 88 475936 116
rect 463660 76 463666 88
rect 475930 76 475936 88
rect 475988 76 475994 128
rect 477218 76 477224 128
rect 477276 116 477282 128
rect 490098 116 490104 128
rect 477276 88 490104 116
rect 477276 76 477282 88
rect 490098 76 490104 88
rect 490156 76 490162 128
rect 513282 76 513288 128
rect 513340 116 513346 128
rect 528738 116 528744 128
rect 513340 88 528744 116
rect 513340 76 513346 88
rect 528738 76 528744 88
rect 528796 76 528802 128
rect 531038 76 531044 128
rect 531096 116 531102 128
rect 548058 116 548064 128
rect 531096 88 548064 116
rect 531096 76 531102 88
rect 548058 76 548064 88
rect 548116 76 548122 128
rect 551922 76 551928 128
rect 551980 116 551986 128
rect 570506 116 570512 128
rect 551980 88 570512 116
rect 551980 76 551986 88
rect 570506 76 570512 88
rect 570564 76 570570 128
rect 382 8 388 60
rect 440 48 446 60
rect 19794 48 19800 60
rect 440 20 19800 48
rect 440 8 446 20
rect 19794 8 19800 20
rect 19852 8 19858 60
rect 30282 8 30288 60
rect 30340 48 30346 60
rect 47394 48 47400 60
rect 30340 20 47400 48
rect 30340 8 30346 20
rect 47394 8 47400 20
rect 47452 8 47458 60
rect 53558 8 53564 60
rect 53616 48 53622 60
rect 69474 48 69480 60
rect 53616 20 69480 48
rect 53616 8 53622 20
rect 69474 8 69480 20
rect 69532 8 69538 60
rect 363230 8 363236 60
rect 363288 48 363294 60
rect 367830 48 367836 60
rect 363288 20 367836 48
rect 363288 8 363294 20
rect 367830 8 367836 20
rect 367888 8 367894 60
rect 399662 8 399668 60
rect 399720 48 399726 60
rect 407022 48 407028 60
rect 399720 20 407028 48
rect 399720 8 399726 20
rect 407022 8 407028 20
rect 407080 8 407086 60
rect 410610 8 410616 60
rect 410668 48 410674 60
rect 418614 48 418620 60
rect 410668 20 418620 48
rect 410668 8 410674 20
rect 418614 8 418620 20
rect 418672 8 418678 60
rect 421742 8 421748 60
rect 421800 48 421806 60
rect 431034 48 431040 60
rect 421800 20 431040 48
rect 421800 8 421806 20
rect 431034 8 431040 20
rect 431092 8 431098 60
rect 439406 8 439412 60
rect 439464 48 439470 60
rect 449986 48 449992 60
rect 439464 20 449992 48
rect 439464 8 439470 20
rect 449986 8 449992 20
rect 450044 8 450050 60
rect 452562 8 452568 60
rect 452620 48 452626 60
rect 464154 48 464160 60
rect 452620 20 464160 48
rect 452620 8 452626 20
rect 464154 8 464160 20
rect 464212 8 464218 60
rect 465810 8 465816 60
rect 465868 48 465874 60
rect 478322 48 478328 60
rect 465868 20 478328 48
rect 465868 8 465874 20
rect 478322 8 478328 20
rect 478380 8 478386 60
rect 484670 8 484676 60
rect 484728 48 484734 60
rect 498378 48 498384 60
rect 484728 20 498384 48
rect 484728 8 484734 20
rect 498378 8 498384 20
rect 498436 8 498442 60
rect 506750 8 506756 60
rect 506808 48 506814 60
rect 521654 48 521660 60
rect 506808 20 521660 48
rect 506808 8 506814 20
rect 521654 8 521660 20
rect 521712 8 521718 60
rect 523310 8 523316 60
rect 523368 48 523374 60
rect 539778 48 539784 60
rect 523368 20 539784 48
rect 523368 8 523374 20
rect 539778 8 539784 20
rect 539836 8 539842 60
rect 546402 8 546408 60
rect 546460 48 546466 60
rect 564618 48 564624 60
rect 546460 20 564624 48
rect 546460 8 546466 20
rect 564618 8 564624 20
rect 564676 8 564682 60
<< via1 >>
rect 186504 702992 186556 703044
rect 188436 702992 188488 703044
rect 235172 702992 235224 703044
rect 236184 702992 236236 703044
rect 522764 702992 522816 703044
rect 527088 702992 527140 703044
rect 570512 702992 570564 703044
rect 575848 702992 575900 703044
rect 490932 702720 490984 702772
rect 494796 702720 494848 702772
rect 538680 702720 538732 702772
rect 543464 702720 543516 702772
rect 24308 702448 24360 702500
rect 29276 702448 29328 702500
rect 218980 702448 219032 702500
rect 220268 702448 220320 702500
rect 459100 702448 459152 702500
rect 462320 702448 462372 702500
rect 506848 702448 506900 702500
rect 510988 702448 511040 702500
rect 554596 702448 554648 702500
rect 559656 702448 559708 702500
rect 8116 700952 8168 701004
rect 13084 700952 13136 701004
rect 40500 700952 40552 701004
rect 44916 700952 44968 701004
rect 56784 700952 56836 701004
rect 60740 700952 60792 701004
rect 72976 700952 73028 701004
rect 76748 700952 76800 701004
rect 89168 700952 89220 701004
rect 92572 700952 92624 701004
rect 105452 700952 105504 701004
rect 108580 700952 108632 701004
rect 121644 700952 121696 701004
rect 124404 700952 124456 701004
rect 137836 700952 137888 701004
rect 140412 700952 140464 701004
rect 154120 700952 154172 701004
rect 156236 700952 156288 701004
rect 170312 700952 170364 701004
rect 172428 700952 172480 701004
rect 202788 700952 202840 701004
rect 204260 700952 204312 701004
rect 348056 700952 348108 701004
rect 348792 700952 348844 701004
rect 363880 700952 363932 701004
rect 364984 700952 365036 701004
rect 379336 700952 379388 701004
rect 381176 700952 381228 701004
rect 395712 700952 395764 701004
rect 397460 700952 397512 701004
rect 411720 700952 411772 701004
rect 413652 700952 413704 701004
rect 427544 700952 427596 701004
rect 429844 700952 429896 701004
rect 443552 700952 443604 701004
rect 446128 700952 446180 701004
rect 475384 700952 475436 701004
rect 478512 700952 478564 701004
rect 73528 3952 73580 4004
rect 87972 3952 88024 4004
rect 64328 3884 64380 3936
rect 79140 3884 79192 3936
rect 70124 3816 70176 3868
rect 84660 3816 84712 3868
rect 99840 3816 99892 3868
rect 112260 3816 112312 3868
rect 58808 3748 58860 3800
rect 73620 3748 73672 3800
rect 77392 3748 77444 3800
rect 91284 3748 91336 3800
rect 105728 3748 105780 3800
rect 117780 3748 117832 3800
rect 125968 3748 126020 3800
rect 136640 3748 136692 3800
rect 63224 3680 63276 3732
rect 78036 3680 78088 3732
rect 83280 3680 83332 3732
rect 96804 3680 96856 3732
rect 98920 3680 98972 3732
rect 103428 3680 103480 3732
rect 118792 3680 118844 3732
rect 129924 3680 129976 3732
rect 60832 3612 60884 3664
rect 75828 3612 75880 3664
rect 79692 3612 79744 3664
rect 93492 3612 93544 3664
rect 95148 3612 95200 3664
rect 107844 3612 107896 3664
rect 117596 3612 117648 3664
rect 128820 3612 128872 3664
rect 144736 3612 144788 3664
rect 154212 3612 154264 3664
rect 56968 3544 57020 3596
rect 72516 3544 72568 3596
rect 72608 3544 72660 3596
rect 86868 3544 86920 3596
rect 89536 3544 89588 3596
rect 102324 3544 102376 3596
rect 103336 3544 103388 3596
rect 115572 3544 115624 3596
rect 120908 3544 120960 3596
rect 132132 3544 132184 3596
rect 132960 3544 133012 3596
rect 143172 3544 143224 3596
rect 148324 3544 148376 3596
rect 157524 3544 157576 3596
rect 71320 3476 71372 3528
rect 85764 3476 85816 3528
rect 98644 3476 98696 3528
rect 111156 3476 111208 3528
rect 129372 3476 129424 3528
rect 139860 3476 139912 3528
rect 142528 3476 142580 3528
rect 152004 3476 152056 3528
rect 163688 3476 163740 3528
rect 171876 3476 171928 3528
rect 59728 3408 59780 3460
rect 74448 3408 74500 3460
rect 75368 3408 75420 3460
rect 89076 3408 89128 3460
rect 93952 3408 94004 3460
rect 100760 3408 100812 3460
rect 52552 3340 52604 3392
rect 68100 3340 68152 3392
rect 68560 3340 68612 3392
rect 82452 3340 82504 3392
rect 90088 3340 90140 3392
rect 98920 3340 98972 3392
rect 48964 3272 49016 3324
rect 40408 3204 40460 3256
rect 57060 3204 57112 3256
rect 62028 3272 62080 3324
rect 76932 3272 76984 3324
rect 85672 3272 85724 3324
rect 99012 3272 99064 3324
rect 64696 3204 64748 3256
rect 66720 3204 66772 3256
rect 51356 3136 51408 3188
rect 66996 3136 67048 3188
rect 80888 3204 80940 3256
rect 94596 3204 94648 3256
rect 96252 3204 96304 3256
rect 109040 3408 109092 3460
rect 116400 3408 116452 3460
rect 127716 3408 127768 3460
rect 137468 3408 137520 3460
rect 101036 3340 101088 3392
rect 114008 3340 114060 3392
rect 125600 3340 125652 3392
rect 127072 3340 127124 3392
rect 137652 3340 137704 3392
rect 153016 3408 153068 3460
rect 161940 3408 161992 3460
rect 169576 3408 169628 3460
rect 177396 3408 177448 3460
rect 183744 3408 183796 3460
rect 190644 3408 190696 3460
rect 147680 3340 147732 3392
rect 155408 3340 155460 3392
rect 164240 3340 164292 3392
rect 167184 3340 167236 3392
rect 175280 3340 175332 3392
rect 180248 3340 180300 3392
rect 187332 3340 187384 3392
rect 109408 3272 109460 3324
rect 121092 3272 121144 3324
rect 130568 3272 130620 3324
rect 140964 3272 141016 3324
rect 143632 3272 143684 3324
rect 153200 3272 153252 3324
rect 154212 3272 154264 3324
rect 163044 3272 163096 3324
rect 164884 3272 164936 3324
rect 172980 3272 173032 3324
rect 174268 3272 174320 3324
rect 181812 3272 181864 3324
rect 189724 3272 189776 3324
rect 196164 3272 196216 3324
rect 560024 3272 560076 3324
rect 578608 3272 578660 3324
rect 113088 3204 113140 3256
rect 122288 3204 122340 3256
rect 133236 3204 133288 3256
rect 139216 3204 139268 3256
rect 148692 3204 148744 3256
rect 150624 3204 150676 3256
rect 159732 3204 159784 3256
rect 161296 3204 161348 3256
rect 169760 3204 169812 3256
rect 173164 3204 173216 3256
rect 180892 3204 180944 3256
rect 182548 3204 182600 3256
rect 189540 3204 189592 3256
rect 190828 3204 190880 3256
rect 197360 3204 197412 3256
rect 200304 3204 200356 3256
rect 206100 3204 206152 3256
rect 553308 3204 553360 3256
rect 571524 3204 571576 3256
rect 81348 3136 81400 3188
rect 82084 3136 82136 3188
rect 95700 3136 95752 3188
rect 97448 3136 97500 3188
rect 110052 3136 110104 3188
rect 110880 3136 110932 3188
rect 122196 3136 122248 3188
rect 135260 3136 135312 3188
rect 145380 3136 145432 3188
rect 147128 3136 147180 3188
rect 156420 3136 156472 3188
rect 162492 3136 162544 3188
rect 56048 3068 56100 3120
rect 71412 3068 71464 3120
rect 87972 3068 88024 3120
rect 101220 3068 101272 3120
rect 102232 3068 102284 3120
rect 114560 3068 114612 3120
rect 115204 3068 115256 3120
rect 126612 3068 126664 3120
rect 134156 3068 134208 3120
rect 144276 3068 144328 3120
rect 151820 3068 151872 3120
rect 160836 3068 160888 3120
rect 164240 3068 164292 3120
rect 168564 3068 168616 3120
rect 170772 3136 170824 3188
rect 178500 3136 178552 3188
rect 179052 3136 179104 3188
rect 186320 3136 186372 3188
rect 192392 3136 192444 3188
rect 198372 3136 198424 3188
rect 201500 3136 201552 3188
rect 206928 3136 206980 3188
rect 214472 3136 214524 3188
rect 219348 3136 219400 3188
rect 220268 3136 220320 3188
rect 224868 3136 224920 3188
rect 229836 3136 229888 3188
rect 233700 3136 233752 3188
rect 556712 3136 556764 3188
rect 575112 3136 575164 3188
rect 170864 3068 170916 3120
rect 176752 3068 176804 3120
rect 184020 3068 184072 3120
rect 196808 3068 196860 3120
rect 202880 3068 202932 3120
rect 208952 3068 209004 3120
rect 213828 3068 213880 3120
rect 215668 3068 215720 3120
rect 220452 3068 220504 3120
rect 221556 3068 221608 3120
rect 225972 3068 226024 3120
rect 231032 3068 231084 3120
rect 234804 3068 234856 3120
rect 530032 3068 530084 3120
rect 546684 3068 546736 3120
rect 564348 3068 564400 3120
rect 583392 3068 583444 3120
rect 47860 3000 47912 3052
rect 63684 3000 63736 3052
rect 33600 2932 33652 2984
rect 50436 2932 50488 2984
rect 54944 2932 54996 2984
rect 70308 3000 70360 3052
rect 76288 3000 76340 3052
rect 90180 3000 90232 3052
rect 91928 3000 91980 3052
rect 104532 3000 104584 3052
rect 108488 3000 108540 3052
rect 119988 3000 120040 3052
rect 128176 3000 128228 3052
rect 138756 3000 138808 3052
rect 140044 3000 140096 3052
rect 149796 3000 149848 3052
rect 156604 3000 156656 3052
rect 165252 3000 165304 3052
rect 171968 3000 172020 3052
rect 179604 3000 179656 3052
rect 187332 3000 187384 3052
rect 193956 3000 194008 3052
rect 194416 3000 194468 3052
rect 200580 3000 200632 3052
rect 202696 3000 202748 3052
rect 208400 3000 208452 3052
rect 214932 3000 214984 3052
rect 218060 3000 218112 3052
rect 222660 3000 222712 3052
rect 225512 3000 225564 3052
rect 229284 3000 229336 3052
rect 233424 3000 233476 3052
rect 237012 3000 237064 3052
rect 238116 3000 238168 3052
rect 241520 3000 241572 3052
rect 248788 3000 248840 3052
rect 251364 3000 251416 3052
rect 331312 3000 331364 3052
rect 333888 3000 333940 3052
rect 334808 3000 334860 3052
rect 337476 3000 337528 3052
rect 543464 3000 543516 3052
rect 560484 3000 560536 3052
rect 562232 3000 562284 3052
rect 581000 3000 581052 3052
rect 69112 2932 69164 2984
rect 83832 2932 83884 2984
rect 84476 2932 84528 2984
rect 98184 2932 98236 2984
rect 106924 2932 106976 2984
rect 119160 2932 119212 2984
rect 119896 2932 119948 2984
rect 131304 2932 131356 2984
rect 131764 2932 131816 2984
rect 142344 2932 142396 2984
rect 145932 2932 145984 2984
rect 155592 2932 155644 2984
rect 157800 2932 157852 2984
rect 166632 2932 166684 2984
rect 26608 2864 26660 2916
rect 43812 2864 43864 2916
rect 44272 2864 44324 2916
rect 60372 2864 60424 2916
rect 65524 2864 65576 2916
rect 27712 2796 27764 2848
rect 44916 2796 44968 2848
rect 50160 2796 50212 2848
rect 65892 2796 65944 2848
rect 67916 2796 67968 2848
rect 68560 2796 68612 2848
rect 78588 2864 78640 2916
rect 92480 2864 92532 2916
rect 92756 2864 92808 2916
rect 105912 2864 105964 2916
rect 112812 2864 112864 2916
rect 124680 2864 124732 2916
rect 125048 2864 125100 2916
rect 135720 2864 135772 2916
rect 141240 2864 141292 2916
rect 151176 2864 151228 2916
rect 158904 2864 158956 2916
rect 79968 2796 80020 2848
rect 86868 2796 86920 2848
rect 100392 2796 100444 2848
rect 104532 2796 104584 2848
rect 110512 2796 110564 2848
rect 111616 2796 111668 2848
rect 123576 2796 123628 2848
rect 123484 2728 123536 2780
rect 134616 2796 134668 2848
rect 136456 2796 136508 2848
rect 146760 2796 146812 2848
rect 149520 2796 149572 2848
rect 158720 2796 158772 2848
rect 160100 2796 160152 2848
rect 164240 2796 164292 2848
rect 166080 2864 166132 2916
rect 174360 2932 174412 2984
rect 177856 2932 177908 2984
rect 185400 2932 185452 2984
rect 186136 2932 186188 2984
rect 193128 2932 193180 2984
rect 195612 2932 195664 2984
rect 201960 2932 202012 2984
rect 203892 2932 203944 2984
rect 209412 2932 209464 2984
rect 209780 2932 209832 2984
rect 212172 2932 212224 2984
rect 217140 2932 217192 2984
rect 222752 2932 222804 2984
rect 227352 2932 227404 2984
rect 227536 2932 227588 2984
rect 231768 2932 231820 2984
rect 234620 2932 234672 2984
rect 238392 2932 238444 2984
rect 239312 2932 239364 2984
rect 242808 2932 242860 2984
rect 242900 2932 242952 2984
rect 246120 2932 246172 2984
rect 246396 2932 246448 2984
rect 249432 2932 249484 2984
rect 253480 2932 253532 2984
rect 256056 2932 256108 2984
rect 310244 2932 310296 2984
rect 311440 2932 311492 2984
rect 325700 2932 325752 2984
rect 328000 2932 328052 2984
rect 329012 2932 329064 2984
rect 331588 2932 331640 2984
rect 332324 2932 332376 2984
rect 335084 2932 335136 2984
rect 341156 2932 341208 2984
rect 344560 2932 344612 2984
rect 536564 2932 536616 2984
rect 553768 2932 553820 2984
rect 560852 2932 560904 2984
rect 579804 2932 579856 2984
rect 168380 2864 168432 2916
rect 176568 2864 176620 2916
rect 181444 2864 181496 2916
rect 188436 2864 188488 2916
rect 188528 2864 188580 2916
rect 195336 2864 195388 2916
rect 199108 2864 199160 2916
rect 204996 2864 205048 2916
rect 206192 2864 206244 2916
rect 211620 2864 211672 2916
rect 213368 2864 213420 2916
rect 218244 2864 218296 2916
rect 219256 2864 219308 2916
rect 223488 2864 223540 2916
rect 226340 2864 226392 2916
rect 230664 2864 230716 2916
rect 232228 2864 232280 2916
rect 236184 2864 236236 2916
rect 237012 2864 237064 2916
rect 240600 2864 240652 2916
rect 242072 2864 242124 2916
rect 245016 2864 245068 2916
rect 245200 2864 245252 2916
rect 248328 2864 248380 2916
rect 249984 2864 250036 2916
rect 252744 2864 252796 2916
rect 254676 2864 254728 2916
rect 257160 2864 257212 2916
rect 261760 2864 261812 2916
rect 263784 2864 263836 2916
rect 312452 2864 312504 2916
rect 313832 2864 313884 2916
rect 314568 2864 314620 2916
rect 316224 2864 316276 2916
rect 316868 2864 316920 2916
rect 318524 2864 318576 2916
rect 319076 2864 319128 2916
rect 320916 2864 320968 2916
rect 321284 2864 321336 2916
rect 323308 2864 323360 2916
rect 323492 2864 323544 2916
rect 325608 2864 325660 2916
rect 327908 2864 327960 2916
rect 330392 2864 330444 2916
rect 333428 2864 333480 2916
rect 336280 2864 336332 2916
rect 340052 2864 340104 2916
rect 342996 2864 343048 2916
rect 526628 2864 526680 2916
rect 542820 2864 542872 2916
rect 549812 2864 549864 2916
rect 568028 2864 568080 2916
rect 167736 2796 167788 2848
rect 175464 2796 175516 2848
rect 183192 2796 183244 2848
rect 184940 2796 184992 2848
rect 192024 2796 192076 2848
rect 199476 2796 199528 2848
rect 205088 2796 205140 2848
rect 210516 2796 210568 2848
rect 210976 2796 211028 2848
rect 216036 2796 216088 2848
rect 216864 2796 216916 2848
rect 221832 2796 221884 2848
rect 223948 2796 224000 2848
rect 228456 2796 228508 2848
rect 228732 2796 228784 2848
rect 232872 2796 232924 2848
rect 235816 2796 235868 2848
rect 239496 2796 239548 2848
rect 240508 2796 240560 2848
rect 243912 2796 243964 2848
rect 244096 2796 244148 2848
rect 247224 2796 247276 2848
rect 247592 2796 247644 2848
rect 250536 2796 250588 2848
rect 252376 2796 252428 2848
rect 254952 2796 255004 2848
rect 255872 2796 255924 2848
rect 258264 2796 258316 2848
rect 260656 2796 260708 2848
rect 262680 2796 262732 2848
rect 304724 2796 304776 2848
rect 305552 2796 305604 2848
rect 306932 2796 306984 2848
rect 307944 2796 307996 2848
rect 309140 2796 309192 2848
rect 310244 2796 310296 2848
rect 311348 2796 311400 2848
rect 312636 2796 312688 2848
rect 313556 2796 313608 2848
rect 315028 2796 315080 2848
rect 315764 2796 315816 2848
rect 317328 2796 317380 2848
rect 317972 2796 318024 2848
rect 319720 2796 319772 2848
rect 320088 2796 320140 2848
rect 322112 2796 322164 2848
rect 322388 2796 322440 2848
rect 324412 2796 324464 2848
rect 324596 2796 324648 2848
rect 326804 2796 326856 2848
rect 326988 2796 327040 2848
rect 329196 2796 329248 2848
rect 330116 2796 330168 2848
rect 332692 2796 332744 2848
rect 335636 2796 335688 2848
rect 338672 2796 338724 2848
rect 338948 2796 339000 2848
rect 342076 2796 342128 2848
rect 346676 2796 346728 2848
rect 350448 2796 350500 2848
rect 353208 2796 353260 2848
rect 357532 2796 357584 2848
rect 372344 2796 372396 2848
rect 377680 2796 377732 2848
rect 546500 2796 546552 2848
rect 557356 2796 557408 2848
rect 562968 2796 563020 2848
rect 582196 2796 582248 2848
rect 193220 2728 193272 2780
rect 198280 1300 198332 1352
rect 204168 1300 204220 1352
rect 207388 1300 207440 1352
rect 213000 1300 213052 1352
rect 257068 1300 257120 1352
rect 259368 1300 259420 1352
rect 259460 1300 259512 1352
rect 261576 1300 261628 1352
rect 262956 1300 263008 1352
rect 264888 1300 264940 1352
rect 265348 1300 265400 1352
rect 267096 1300 267148 1352
rect 267740 1300 267792 1352
rect 269304 1300 269356 1352
rect 271236 1300 271288 1352
rect 272616 1300 272668 1352
rect 273628 1300 273680 1352
rect 274824 1300 274876 1352
rect 277124 1300 277176 1352
rect 278136 1300 278188 1352
rect 279516 1300 279568 1352
rect 280344 1300 280396 1352
rect 336648 1300 336700 1352
rect 339868 1300 339920 1352
rect 342168 1300 342220 1352
rect 345756 1300 345808 1352
rect 348884 1300 348936 1352
rect 352840 1300 352892 1352
rect 356612 1300 356664 1352
rect 361120 1300 361172 1352
rect 364248 1300 364300 1352
rect 369400 1300 369452 1352
rect 369768 1300 369820 1352
rect 375288 1300 375340 1352
rect 376484 1300 376536 1352
rect 382372 1300 382424 1352
rect 384212 1300 384264 1352
rect 390652 1300 390704 1352
rect 394148 1300 394200 1352
rect 401324 1300 401376 1352
rect 406292 1300 406344 1352
rect 414296 1300 414348 1352
rect 436008 1300 436060 1352
rect 445852 1300 445904 1352
rect 450452 1300 450504 1352
rect 461584 1300 461636 1352
rect 462596 1300 462648 1352
rect 474188 1300 474240 1352
rect 475844 1300 475896 1352
rect 488816 1300 488868 1352
rect 493508 1300 493560 1352
rect 500040 1300 500092 1352
rect 500132 1300 500184 1352
rect 507032 1300 507084 1352
rect 516692 1300 516744 1352
rect 532056 1300 532108 1352
rect 539876 1300 539928 1352
rect 546500 1300 546552 1352
rect 100760 1232 100812 1284
rect 107016 1232 107068 1284
rect 110512 1232 110564 1284
rect 116952 1232 117004 1284
rect 258264 1232 258316 1284
rect 260472 1232 260524 1284
rect 264152 1232 264204 1284
rect 265992 1232 266044 1284
rect 266544 1232 266596 1284
rect 268200 1232 268252 1284
rect 270040 1232 270092 1284
rect 271512 1232 271564 1284
rect 272432 1232 272484 1284
rect 273720 1232 273772 1284
rect 343364 1232 343416 1284
rect 346952 1232 347004 1284
rect 349988 1232 350040 1284
rect 354036 1232 354088 1284
rect 357716 1232 357768 1284
rect 362316 1232 362368 1284
rect 365444 1232 365496 1284
rect 370228 1232 370280 1284
rect 370964 1232 371016 1284
rect 376116 1232 376168 1284
rect 378692 1232 378744 1284
rect 384396 1232 384448 1284
rect 387524 1232 387576 1284
rect 394240 1232 394292 1284
rect 396356 1232 396408 1284
rect 403624 1232 403676 1284
rect 404084 1232 404136 1284
rect 411904 1232 411956 1284
rect 430488 1232 430540 1284
rect 439964 1232 440016 1284
rect 447048 1232 447100 1284
rect 456432 1232 456484 1284
rect 474648 1232 474700 1284
rect 487252 1232 487304 1284
rect 499028 1232 499080 1284
rect 268844 1164 268896 1216
rect 270408 1164 270460 1216
rect 359924 1164 359976 1216
rect 364616 1164 364668 1216
rect 368756 1164 368808 1216
rect 373908 1164 373960 1216
rect 374276 1164 374328 1216
rect 379612 1164 379664 1216
rect 379796 1164 379848 1216
rect 385960 1164 386012 1216
rect 395252 1164 395304 1216
rect 402520 1164 402572 1216
rect 443828 1164 443880 1216
rect 454132 1164 454184 1216
rect 457076 1164 457128 1216
rect 468300 1164 468352 1216
rect 469128 1164 469180 1216
rect 481364 1164 481416 1216
rect 490196 1164 490248 1216
rect 503812 1164 503864 1216
rect 512276 1232 512328 1284
rect 527824 1232 527876 1284
rect 513380 1164 513432 1216
rect 517796 1164 517848 1216
rect 533712 1164 533764 1216
rect 352196 1096 352248 1148
rect 356336 1096 356388 1148
rect 361028 1096 361080 1148
rect 365444 1096 365496 1148
rect 366548 1096 366600 1148
rect 371332 1096 371384 1148
rect 375196 1096 375248 1148
rect 381176 1096 381228 1148
rect 385316 1096 385368 1148
rect 391848 1096 391900 1148
rect 397368 1096 397420 1148
rect 404820 1096 404872 1148
rect 412916 1096 412968 1148
rect 421380 1096 421432 1148
rect 437204 1096 437256 1148
rect 447416 1096 447468 1148
rect 485688 1096 485740 1148
rect 499028 1096 499080 1148
rect 500408 1096 500460 1148
rect 355508 1028 355560 1080
rect 359924 1028 359976 1080
rect 367652 1028 367704 1080
rect 372896 1028 372948 1080
rect 377588 1028 377640 1080
rect 383568 1028 383620 1080
rect 451556 1028 451608 1080
rect 462412 1028 462464 1080
rect 489092 1028 489144 1080
rect 502984 1028 503036 1080
rect 503444 1028 503496 1080
rect 511172 1096 511224 1148
rect 526260 1096 526312 1148
rect 21824 960 21876 1012
rect 39672 960 39724 1012
rect 345572 960 345624 1012
rect 349252 960 349304 1012
rect 351092 960 351144 1012
rect 355232 960 355284 1012
rect 362132 960 362184 1012
rect 367008 960 367060 1012
rect 373172 960 373224 1012
rect 378508 960 378560 1012
rect 416228 960 416280 1012
rect 424968 960 425020 1012
rect 448244 960 448296 1012
rect 459192 960 459244 1012
rect 482468 960 482520 1012
rect 495532 960 495584 1012
rect 495716 960 495768 1012
rect 509700 960 509752 1012
rect 512092 1028 512144 1080
rect 517980 960 518032 1012
rect 534356 960 534408 1012
rect 551468 960 551520 1012
rect 19432 892 19484 944
rect 37464 892 37516 944
rect 358728 892 358780 944
rect 363512 892 363564 944
rect 444932 892 444984 944
rect 455696 892 455748 944
rect 455972 892 456024 944
rect 467472 892 467524 944
rect 480168 892 480220 944
rect 493140 892 493192 944
rect 494612 892 494664 944
rect 508872 892 508924 944
rect 510068 892 510120 944
rect 525432 892 525484 944
rect 532148 892 532200 944
rect 549076 892 549128 944
rect 11152 824 11204 876
rect 29736 824 29788 876
rect 337844 824 337896 876
rect 340972 824 341024 876
rect 347688 824 347740 876
rect 351644 824 351696 876
rect 441528 824 441580 876
rect 451740 824 451792 876
rect 454868 824 454920 876
rect 465908 824 465960 876
rect 492404 824 492456 876
rect 506480 824 506532 876
rect 508964 824 509016 876
rect 523868 824 523920 876
rect 550916 824 550968 876
rect 569132 824 569184 876
rect 20628 756 20680 808
rect 38568 756 38620 808
rect 251180 756 251232 808
rect 253848 756 253900 808
rect 438308 756 438360 808
rect 448244 756 448296 808
rect 449348 756 449400 808
rect 460020 756 460072 808
rect 483572 756 483624 808
rect 497096 756 497148 808
rect 502248 756 502300 808
rect 14740 688 14792 740
rect 33048 688 33100 740
rect 18236 620 18288 672
rect 36360 688 36412 740
rect 386328 688 386380 740
rect 392676 688 392728 740
rect 408408 688 408460 740
rect 416688 688 416740 740
rect 423956 688 424008 740
rect 433248 688 433300 740
rect 446036 688 446088 740
rect 456524 688 456576 740
rect 35992 620 36044 672
rect 52920 620 52972 672
rect 393044 620 393096 672
rect 400128 620 400180 672
rect 400772 620 400824 672
rect 409604 620 409656 672
rect 417884 620 417936 672
rect 418436 620 418488 672
rect 427268 620 427320 672
rect 442724 620 442776 672
rect 453304 620 453356 672
rect 468116 620 468168 672
rect 480536 688 480588 740
rect 487988 688 488040 740
rect 501420 688 501472 740
rect 504548 688 504600 740
rect 507032 756 507084 808
rect 514760 756 514812 808
rect 527732 756 527784 808
rect 544384 756 544436 808
rect 547604 756 547656 808
rect 565636 756 565688 808
rect 15936 552 15988 604
rect 34152 552 34204 604
rect 34796 552 34848 604
rect 51816 552 51868 604
rect 388628 552 388680 604
rect 395344 552 395396 604
rect 408408 552 408460 604
rect 426164 552 426216 604
rect 435548 552 435600 604
rect 439136 552 439188 604
rect 464804 552 464856 604
rect 476948 620 477000 672
rect 481548 620 481600 672
rect 494704 620 494756 672
rect 497924 620 497976 672
rect 500408 620 500460 672
rect 473452 552 473504 604
rect 486424 552 486476 604
rect 491208 552 491260 604
rect 505376 620 505428 672
rect 517152 688 517204 740
rect 524328 688 524380 740
rect 540796 688 540848 740
rect 540888 688 540940 740
rect 558552 688 558604 740
rect 500592 552 500644 604
rect 525524 620 525576 672
rect 541992 620 542044 672
rect 545396 620 545448 672
rect 563244 620 563296 672
rect 519544 552 519596 604
rect 522212 552 522264 604
rect 538404 552 538456 604
rect 542084 552 542136 604
rect 559748 552 559800 604
rect 562048 552 562100 604
rect 3240 484 3292 536
rect 22008 484 22060 536
rect 22836 484 22888 536
rect 40500 484 40552 536
rect 45284 484 45336 536
rect 61752 484 61804 536
rect 420644 484 420696 536
rect 429292 484 429344 536
rect 429476 484 429528 536
rect 461768 484 461820 536
rect 473636 484 473688 536
rect 486884 484 486936 536
rect 501236 484 501288 536
rect 515588 484 515640 536
rect 518808 484 518860 536
rect 534540 484 534592 536
rect 544568 484 544620 536
rect 9128 416 9180 468
rect 27528 416 27580 468
rect 32220 416 32272 468
rect 49608 416 49660 468
rect 401876 416 401928 468
rect 409236 416 409288 468
rect 424784 416 424836 468
rect 434076 416 434128 468
rect 434996 416 435048 468
rect 445208 416 445260 468
rect 457904 416 457956 468
rect 470048 416 470100 468
rect 470324 416 470376 468
rect 482468 416 482520 468
rect 500040 416 500092 468
rect 507308 416 507360 468
rect 507860 416 507912 468
rect 523224 416 523276 468
rect 528836 416 528888 468
rect 545672 416 545724 468
rect 548708 416 548760 468
rect 567016 416 567068 468
rect 9772 348 9824 400
rect 28632 348 28684 400
rect 39396 348 39448 400
rect 56232 348 56284 400
rect 407396 348 407448 400
rect 415308 348 415360 400
rect 417332 348 417384 400
rect 425796 348 425848 400
rect 428648 348 428700 400
rect 437572 348 437624 400
rect 459468 348 459520 400
rect 470784 348 470836 400
rect 472532 348 472584 400
rect 484860 348 484912 400
rect 496728 348 496780 400
rect 511448 348 511500 400
rect 514484 348 514536 400
rect 529940 348 529992 400
rect 533252 348 533304 400
rect 550456 348 550508 400
rect 555332 348 555384 400
rect 573548 348 573600 400
rect 17408 280 17460 332
rect 35256 280 35308 332
rect 38568 280 38620 332
rect 55128 280 55180 332
rect 382004 280 382056 332
rect 387892 280 387944 332
rect 389732 280 389784 332
rect 396172 280 396224 332
rect 413928 280 413980 332
rect 422760 280 422812 332
rect 427544 280 427596 332
rect 436928 280 436980 332
rect 440516 280 440568 332
rect 451096 280 451148 332
rect 467012 280 467064 332
rect 478972 280 479024 332
rect 479524 280 479576 332
rect 492496 280 492548 332
rect 505652 280 505704 332
rect 520372 280 520424 332
rect 521108 280 521160 332
rect 537392 280 537444 332
rect 538772 280 538824 332
rect 556344 280 556396 332
rect 557172 280 557224 332
rect 575940 280 575992 332
rect 3884 212 3936 264
rect 23204 212 23256 264
rect 42248 212 42300 264
rect 58164 212 58216 264
rect 390836 212 390888 264
rect 397920 212 397972 264
rect 402888 212 402940 264
rect 410984 212 411036 264
rect 415124 212 415176 264
rect 423588 212 423640 264
rect 432788 212 432840 264
rect 442816 212 442868 264
rect 456432 212 456484 264
rect 458272 212 458324 264
rect 460572 212 460624 264
rect 472440 212 472492 264
rect 478328 212 478380 264
rect 490748 212 490800 264
rect 515496 212 515548 264
rect 531504 212 531556 264
rect 535368 212 535420 264
rect 552848 212 552900 264
rect 554228 212 554280 264
rect 572904 212 572956 264
rect 1492 144 1544 196
rect 20904 144 20956 196
rect 24584 144 24636 196
rect 41604 144 41656 196
rect 42892 144 42944 196
rect 59360 144 59412 196
rect 380808 144 380860 196
rect 386788 144 386840 196
rect 391664 144 391716 196
rect 398748 144 398800 196
rect 405188 144 405240 196
rect 412824 144 412876 196
rect 419448 144 419500 196
rect 428648 144 428700 196
rect 431684 144 431736 196
rect 441252 144 441304 196
rect 453764 144 453816 196
rect 464988 144 465040 196
rect 471428 144 471480 196
rect 484216 144 484268 196
rect 520004 144 520056 196
rect 536288 144 536340 196
rect 537668 144 537720 196
rect 554780 144 554832 196
rect 558828 144 558880 196
rect 577136 144 577188 196
rect 8024 76 8076 128
rect 26332 76 26384 128
rect 31116 76 31168 128
rect 48504 76 48556 128
rect 344744 76 344796 128
rect 348240 76 348292 128
rect 354404 76 354456 128
rect 358912 76 358964 128
rect 383108 76 383160 128
rect 389640 76 389692 128
rect 398564 76 398616 128
rect 406200 76 406252 128
rect 412088 76 412140 128
rect 420368 76 420420 128
rect 422852 76 422904 128
rect 431868 76 431920 128
rect 433892 76 433944 128
rect 443460 76 443512 128
rect 463608 76 463660 128
rect 475936 76 475988 128
rect 477224 76 477276 128
rect 490104 76 490156 128
rect 513288 76 513340 128
rect 528744 76 528796 128
rect 531044 76 531096 128
rect 548064 76 548116 128
rect 551928 76 551980 128
rect 570512 76 570564 128
rect 388 8 440 60
rect 19800 8 19852 60
rect 30288 8 30340 60
rect 47400 8 47452 60
rect 53564 8 53616 60
rect 69480 8 69532 60
rect 363236 8 363288 60
rect 367836 8 367888 60
rect 399668 8 399720 60
rect 407028 8 407080 60
rect 410616 8 410668 60
rect 418620 8 418672 60
rect 421748 8 421800 60
rect 431040 8 431092 60
rect 439412 8 439464 60
rect 449992 8 450044 60
rect 452568 8 452620 60
rect 464160 8 464212 60
rect 465816 8 465868 60
rect 478328 8 478380 60
rect 484676 8 484728 60
rect 498384 8 498436 60
rect 506756 8 506808 60
rect 521660 8 521712 60
rect 523316 8 523368 60
rect 539784 8 539836 60
rect 546408 8 546460 60
rect 564624 8 564676 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 251652 703582 251864 703610
rect 8128 701010 8156 703520
rect 24320 702506 24348 703520
rect 24308 702500 24360 702506
rect 24308 702442 24360 702448
rect 29276 702500 29328 702506
rect 29276 702442 29328 702448
rect 8116 701004 8168 701010
rect 8116 700946 8168 700952
rect 13084 701004 13136 701010
rect 13084 700946 13136 700952
rect 13096 700890 13124 700946
rect 13096 700862 13386 700890
rect 29288 700876 29316 702442
rect 40512 701010 40540 703520
rect 56796 701010 56824 703520
rect 72988 701010 73016 703520
rect 89180 701010 89208 703520
rect 105464 701010 105492 703520
rect 121656 701010 121684 703520
rect 137848 701010 137876 703520
rect 154132 701010 154160 703520
rect 170324 701010 170352 703520
rect 186516 703050 186544 703520
rect 186504 703044 186556 703050
rect 186504 702986 186556 702992
rect 188436 703044 188488 703050
rect 188436 702986 188488 702992
rect 40500 701004 40552 701010
rect 40500 700946 40552 700952
rect 44916 701004 44968 701010
rect 44916 700946 44968 700952
rect 56784 701004 56836 701010
rect 56784 700946 56836 700952
rect 60740 701004 60792 701010
rect 60740 700946 60792 700952
rect 72976 701004 73028 701010
rect 72976 700946 73028 700952
rect 76748 701004 76800 701010
rect 76748 700946 76800 700952
rect 89168 701004 89220 701010
rect 89168 700946 89220 700952
rect 92572 701004 92624 701010
rect 92572 700946 92624 700952
rect 105452 701004 105504 701010
rect 105452 700946 105504 700952
rect 108580 701004 108632 701010
rect 108580 700946 108632 700952
rect 121644 701004 121696 701010
rect 121644 700946 121696 700952
rect 124404 701004 124456 701010
rect 124404 700946 124456 700952
rect 137836 701004 137888 701010
rect 137836 700946 137888 700952
rect 140412 701004 140464 701010
rect 140412 700946 140464 700952
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 156236 701004 156288 701010
rect 156236 700946 156288 700952
rect 170312 701004 170364 701010
rect 170312 700946 170364 700952
rect 172428 701004 172480 701010
rect 172428 700946 172480 700952
rect 44928 700890 44956 700946
rect 60752 700890 60780 700946
rect 76760 700890 76788 700946
rect 92584 700890 92612 700946
rect 108592 700890 108620 700946
rect 124416 700890 124444 700946
rect 140424 700890 140452 700946
rect 156248 700890 156276 700946
rect 172440 700890 172468 700946
rect 44928 700862 45218 700890
rect 60752 700862 61134 700890
rect 76760 700862 77050 700890
rect 92584 700862 92966 700890
rect 108592 700862 108882 700890
rect 124416 700862 124798 700890
rect 140424 700862 140714 700890
rect 156248 700862 156630 700890
rect 172440 700862 172546 700890
rect 188448 700876 188476 702986
rect 202800 701010 202828 703520
rect 218992 702506 219020 703520
rect 235184 703050 235212 703520
rect 251468 703474 251496 703520
rect 251652 703474 251680 703582
rect 251468 703446 251680 703474
rect 235172 703044 235224 703050
rect 235172 702986 235224 702992
rect 236184 703044 236236 703050
rect 236184 702986 236236 702992
rect 218980 702500 219032 702506
rect 218980 702442 219032 702448
rect 220268 702500 220320 702506
rect 220268 702442 220320 702448
rect 202788 701004 202840 701010
rect 202788 700946 202840 700952
rect 204260 701004 204312 701010
rect 204260 700946 204312 700952
rect 204272 700890 204300 700946
rect 204272 700862 204378 700890
rect 220280 700876 220308 702442
rect 236196 700876 236224 702986
rect 251836 700890 251864 703582
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332152 703582 332364 703610
rect 267660 700890 267688 703520
rect 283852 700890 283880 703520
rect 300136 700890 300164 703520
rect 316328 702434 316356 703520
rect 316052 702406 316356 702434
rect 316052 700890 316080 702406
rect 332152 700890 332180 703582
rect 332336 703474 332364 703582
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 332520 703474 332548 703520
rect 332336 703446 332548 703474
rect 348804 701010 348832 703520
rect 364996 701010 365024 703520
rect 381188 701010 381216 703520
rect 397472 701010 397500 703520
rect 413664 701010 413692 703520
rect 429856 701010 429884 703520
rect 446140 701010 446168 703520
rect 462332 702506 462360 703520
rect 459100 702500 459152 702506
rect 459100 702442 459152 702448
rect 462320 702500 462372 702506
rect 462320 702442 462372 702448
rect 348056 701004 348108 701010
rect 348056 700946 348108 700952
rect 348792 701004 348844 701010
rect 348792 700946 348844 700952
rect 363880 701004 363932 701010
rect 363880 700946 363932 700952
rect 364984 701004 365036 701010
rect 364984 700946 365036 700952
rect 379336 701004 379388 701010
rect 379336 700946 379388 700952
rect 381176 701004 381228 701010
rect 381176 700946 381228 700952
rect 395712 701004 395764 701010
rect 395712 700946 395764 700952
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 411720 701004 411772 701010
rect 411720 700946 411772 700952
rect 413652 701004 413704 701010
rect 413652 700946 413704 700952
rect 427544 701004 427596 701010
rect 427544 700946 427596 700952
rect 429844 701004 429896 701010
rect 429844 700946 429896 700952
rect 443552 701004 443604 701010
rect 443552 700946 443604 700952
rect 446128 701004 446180 701010
rect 446128 700946 446180 700952
rect 348068 700890 348096 700946
rect 363892 700890 363920 700946
rect 251836 700862 252126 700890
rect 267660 700862 268042 700890
rect 283852 700862 283958 700890
rect 299966 700862 300164 700890
rect 315882 700862 316080 700890
rect 331798 700862 332180 700890
rect 347714 700862 348096 700890
rect 363630 700862 363920 700890
rect 379348 700890 379376 700946
rect 395724 700890 395752 700946
rect 411732 700890 411760 700946
rect 427556 700890 427584 700946
rect 443564 700890 443592 700946
rect 379348 700862 379454 700890
rect 395462 700862 395752 700890
rect 411378 700862 411760 700890
rect 427294 700862 427584 700890
rect 443210 700862 443592 700890
rect 459112 700876 459140 702442
rect 478524 701010 478552 703520
rect 494808 702778 494836 703520
rect 490932 702772 490984 702778
rect 490932 702714 490984 702720
rect 494796 702772 494848 702778
rect 494796 702714 494848 702720
rect 475384 701004 475436 701010
rect 475384 700946 475436 700952
rect 478512 701004 478564 701010
rect 478512 700946 478564 700952
rect 475396 700890 475424 700946
rect 475042 700862 475424 700890
rect 490944 700876 490972 702714
rect 511000 702506 511028 703520
rect 527192 703066 527220 703520
rect 527100 703050 527220 703066
rect 522764 703044 522816 703050
rect 522764 702986 522816 702992
rect 527088 703044 527220 703050
rect 527140 703038 527220 703044
rect 527088 702986 527140 702992
rect 506848 702500 506900 702506
rect 506848 702442 506900 702448
rect 510988 702500 511040 702506
rect 510988 702442 511040 702448
rect 506860 700876 506888 702442
rect 522776 700876 522804 702986
rect 543476 702778 543504 703520
rect 538680 702772 538732 702778
rect 538680 702714 538732 702720
rect 543464 702772 543516 702778
rect 543464 702714 543516 702720
rect 538692 700876 538720 702714
rect 559668 702506 559696 703520
rect 575860 703050 575888 703520
rect 570512 703044 570564 703050
rect 570512 702986 570564 702992
rect 575848 703044 575900 703050
rect 575848 702986 575900 702992
rect 554596 702500 554648 702506
rect 554596 702442 554648 702448
rect 559656 702500 559708 702506
rect 559656 702442 559708 702448
rect 554608 700876 554636 702442
rect 570524 700876 570552 702986
rect 2042 697368 2098 697377
rect 2042 697303 2098 697312
rect 2056 690849 2084 697303
rect 581642 697232 581698 697241
rect 581642 697167 581698 697176
rect 581656 691529 581684 697167
rect 581642 691520 581698 691529
rect 581642 691455 581698 691464
rect 2042 690840 2098 690849
rect 2042 690775 2098 690784
rect 1030 684312 1086 684321
rect 1030 684247 1086 684256
rect 1044 678065 1072 684247
rect 582378 683904 582434 683913
rect 582378 683839 582434 683848
rect 582392 678473 582420 683839
rect 582378 678464 582434 678473
rect 582378 678399 582434 678408
rect 1030 678056 1086 678065
rect 1030 677991 1086 678000
rect 1030 671256 1086 671265
rect 1030 671191 1086 671200
rect 1044 665281 1072 671191
rect 582378 670712 582434 670721
rect 582378 670647 582434 670656
rect 582392 665417 582420 670647
rect 582378 665408 582434 665417
rect 582378 665343 582434 665352
rect 1030 665272 1086 665281
rect 1030 665207 1086 665216
rect 18 657656 74 657665
rect 18 657591 74 657600
rect 32 652497 60 657591
rect 582378 657384 582434 657393
rect 582378 657319 582434 657328
rect 18 652488 74 652497
rect 18 652423 74 652432
rect 582392 652361 582420 657319
rect 582378 652352 582434 652361
rect 582378 652287 582434 652296
rect 1306 645144 1362 645153
rect 1306 645079 1362 645088
rect 1320 639713 1348 645079
rect 581642 644056 581698 644065
rect 581642 643991 581698 644000
rect 1306 639704 1362 639713
rect 1306 639639 1362 639648
rect 581656 639305 581684 643991
rect 581642 639296 581698 639305
rect 581642 639231 581698 639240
rect 1306 632088 1362 632097
rect 1306 632023 1362 632032
rect 1320 626929 1348 632023
rect 582378 630864 582434 630873
rect 582378 630799 582434 630808
rect 1306 626920 1362 626929
rect 1306 626855 1362 626864
rect 582392 626249 582420 630799
rect 582378 626240 582434 626249
rect 582378 626175 582434 626184
rect 18 618624 74 618633
rect 18 618559 74 618568
rect 32 614009 60 618559
rect 581642 617536 581698 617545
rect 581642 617471 581698 617480
rect 18 614000 74 614009
rect 18 613935 74 613944
rect 581656 613193 581684 617471
rect 581642 613184 581698 613193
rect 581642 613119 581698 613128
rect 846 606112 902 606121
rect 846 606047 902 606056
rect 860 601361 888 606047
rect 581642 604208 581698 604217
rect 581642 604143 581698 604152
rect 846 601352 902 601361
rect 846 601287 902 601296
rect 581656 600137 581684 604143
rect 581642 600128 581698 600137
rect 581642 600063 581698 600072
rect 2778 593056 2834 593065
rect 2778 592991 2834 593000
rect 2792 588577 2820 592991
rect 581642 591016 581698 591025
rect 581642 590951 581698 590960
rect 2778 588568 2834 588577
rect 2778 588503 2834 588512
rect 581656 587081 581684 590951
rect 581642 587072 581698 587081
rect 581642 587007 581698 587016
rect 2778 580000 2834 580009
rect 2778 579935 2834 579944
rect 2792 575793 2820 579935
rect 581642 577688 581698 577697
rect 581642 577623 581698 577632
rect 2778 575784 2834 575793
rect 2778 575719 2834 575728
rect 581656 574025 581684 577623
rect 581642 574016 581698 574025
rect 581642 573951 581698 573960
rect 2778 566944 2834 566953
rect 2778 566879 2834 566888
rect 2792 563009 2820 566879
rect 582378 564360 582434 564369
rect 582378 564295 582434 564304
rect 2778 563000 2834 563009
rect 2778 562935 2834 562944
rect 582392 560969 582420 564295
rect 582378 560960 582434 560969
rect 582378 560895 582434 560904
rect 2778 553888 2834 553897
rect 2778 553823 2834 553832
rect 2792 550225 2820 553823
rect 581642 551168 581698 551177
rect 581642 551103 581698 551112
rect 2778 550216 2834 550225
rect 2778 550151 2834 550160
rect 581656 547777 581684 551103
rect 581642 547768 581698 547777
rect 581642 547703 581698 547712
rect 1398 540832 1454 540841
rect 1398 540767 1454 540776
rect 1412 537441 1440 540767
rect 582378 537840 582434 537849
rect 582378 537775 582434 537784
rect 1398 537432 1454 537441
rect 1398 537367 1454 537376
rect 582392 534857 582420 537775
rect 582378 534848 582434 534857
rect 582378 534783 582434 534792
rect 1490 527912 1546 527921
rect 1490 527847 1546 527856
rect 1504 524657 1532 527847
rect 1490 524648 1546 524657
rect 1490 524583 1546 524592
rect 582378 524512 582434 524521
rect 582378 524447 582434 524456
rect 582392 521801 582420 524447
rect 582378 521792 582434 521801
rect 582378 521727 582434 521736
rect 2778 514856 2834 514865
rect 2778 514791 2834 514800
rect 2792 511873 2820 514791
rect 2778 511864 2834 511873
rect 2778 511799 2834 511808
rect 582378 511320 582434 511329
rect 582378 511255 582434 511264
rect 582392 508745 582420 511255
rect 582378 508736 582434 508745
rect 582378 508671 582434 508680
rect 1582 501800 1638 501809
rect 1582 501735 1638 501744
rect 1596 499089 1624 501735
rect 1582 499080 1638 499089
rect 1582 499015 1638 499024
rect 581642 497992 581698 498001
rect 581642 497927 581698 497936
rect 581656 495689 581684 497927
rect 581642 495680 581698 495689
rect 581642 495615 581698 495624
rect 1582 488744 1638 488753
rect 1582 488679 1638 488688
rect 1596 486305 1624 488679
rect 1582 486296 1638 486305
rect 1582 486231 1638 486240
rect 582378 484664 582434 484673
rect 582378 484599 582434 484608
rect 582392 482633 582420 484599
rect 582378 482624 582434 482633
rect 582378 482559 582434 482568
rect 2778 475688 2834 475697
rect 2778 475623 2834 475632
rect 2792 473521 2820 475623
rect 2778 473512 2834 473521
rect 2778 473447 2834 473456
rect 581642 471472 581698 471481
rect 581642 471407 581698 471416
rect 581656 469577 581684 471407
rect 581642 469568 581698 469577
rect 581642 469503 581698 469512
rect 1582 462632 1638 462641
rect 1582 462567 1638 462576
rect 1596 460737 1624 462567
rect 1582 460728 1638 460737
rect 1582 460663 1638 460672
rect 581642 458144 581698 458153
rect 581642 458079 581698 458088
rect 581656 456521 581684 458079
rect 581642 456512 581698 456521
rect 581642 456447 581698 456456
rect 2778 449576 2834 449585
rect 2778 449511 2834 449520
rect 2792 447953 2820 449511
rect 2778 447944 2834 447953
rect 2778 447879 2834 447888
rect 2778 436656 2834 436665
rect 2778 436591 2834 436600
rect 2792 435169 2820 436591
rect 2778 435160 2834 435169
rect 2778 435095 2834 435104
rect 2778 423600 2834 423609
rect 2778 423535 2834 423544
rect 2792 422385 2820 423535
rect 2778 422376 2834 422385
rect 2778 422311 2834 422320
rect 1306 294400 1362 294409
rect 1306 294335 1362 294344
rect 1320 293185 1348 294335
rect 1306 293176 1362 293185
rect 1306 293111 1362 293120
rect 2778 281616 2834 281625
rect 2778 281551 2834 281560
rect 2792 280129 2820 281551
rect 2778 280120 2834 280129
rect 2778 280055 2834 280064
rect 1306 268832 1362 268841
rect 1306 268767 1362 268776
rect 1320 267209 1348 268767
rect 1306 267200 1362 267209
rect 1306 267135 1362 267144
rect 582378 260536 582434 260545
rect 582378 260471 582434 260480
rect 582392 258913 582420 260471
rect 582378 258904 582434 258913
rect 582378 258839 582434 258848
rect 1306 256048 1362 256057
rect 1306 255983 1362 255992
rect 1320 254153 1348 255983
rect 1306 254144 1362 254153
rect 1306 254079 1362 254088
rect 580906 247072 580962 247081
rect 580906 247007 580962 247016
rect 580920 245585 580948 247007
rect 580906 245576 580962 245585
rect 580906 245511 580962 245520
rect 2778 243264 2834 243273
rect 2778 243199 2834 243208
rect 2792 241097 2820 243199
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 582378 234424 582434 234433
rect 582378 234359 582434 234368
rect 582392 232393 582420 234359
rect 582378 232384 582434 232393
rect 582378 232319 582434 232328
rect 2778 230616 2834 230625
rect 2778 230551 2834 230560
rect 2792 228041 2820 230551
rect 2778 228032 2834 228041
rect 2778 227967 2834 227976
rect 580906 220960 580962 220969
rect 580906 220895 580962 220904
rect 580920 219065 580948 220895
rect 580906 219056 580962 219065
rect 580906 218991 580962 219000
rect 2778 217696 2834 217705
rect 2778 217631 2834 217640
rect 2792 214985 2820 217631
rect 2778 214976 2834 214985
rect 2778 214911 2834 214920
rect 582378 208312 582434 208321
rect 582378 208247 582434 208256
rect 582392 205737 582420 208247
rect 582378 205728 582434 205737
rect 582378 205663 582434 205672
rect 2778 204912 2834 204921
rect 2778 204847 2834 204856
rect 2792 201929 2820 204847
rect 2778 201920 2834 201929
rect 2778 201855 2834 201864
rect 580906 194712 580962 194721
rect 580906 194647 580962 194656
rect 580920 192545 580948 194647
rect 580906 192536 580962 192545
rect 580906 192471 580962 192480
rect 1306 192128 1362 192137
rect 1306 192063 1362 192072
rect 1320 188873 1348 192063
rect 1306 188864 1362 188873
rect 1306 188799 1362 188808
rect 580906 182472 580962 182481
rect 580906 182407 580962 182416
rect 2778 179344 2834 179353
rect 2778 179279 2834 179288
rect 2792 175953 2820 179279
rect 580920 179217 580948 182407
rect 580906 179208 580962 179217
rect 580906 179143 580962 179152
rect 2778 175944 2834 175953
rect 2778 175879 2834 175888
rect 580906 168600 580962 168609
rect 580906 168535 580962 168544
rect 2778 166560 2834 166569
rect 2778 166495 2834 166504
rect 2792 162897 2820 166495
rect 580920 165889 580948 168535
rect 580906 165880 580962 165889
rect 580906 165815 580962 165824
rect 2778 162888 2834 162897
rect 2778 162823 2834 162832
rect 580906 156360 580962 156369
rect 580906 156295 580962 156304
rect 1306 153776 1362 153785
rect 1306 153711 1362 153720
rect 1320 149841 1348 153711
rect 580920 152697 580948 156295
rect 580906 152688 580962 152697
rect 580906 152623 580962 152632
rect 1306 149832 1362 149841
rect 1306 149767 1362 149776
rect 580906 142624 580962 142633
rect 580906 142559 580962 142568
rect 570 140992 626 141001
rect 570 140927 626 140936
rect 584 136785 612 140927
rect 580920 139369 580948 142559
rect 580906 139360 580962 139369
rect 580906 139295 580962 139304
rect 570 136776 626 136785
rect 570 136711 626 136720
rect 580906 130248 580962 130257
rect 580906 130183 580962 130192
rect 754 128208 810 128217
rect 754 128143 810 128152
rect 768 123729 796 128143
rect 580920 126041 580948 130183
rect 580906 126032 580962 126041
rect 580906 125967 580962 125976
rect 754 123720 810 123729
rect 754 123655 810 123664
rect 579894 116376 579950 116385
rect 579894 116311 579950 116320
rect 1306 115424 1362 115433
rect 1306 115359 1362 115368
rect 1320 110673 1348 115359
rect 579908 112849 579936 116311
rect 579894 112840 579950 112849
rect 579894 112775 579950 112784
rect 1306 110664 1362 110673
rect 1306 110599 1362 110608
rect 580906 103592 580962 103601
rect 580906 103527 580962 103536
rect 1582 102640 1638 102649
rect 1582 102575 1638 102584
rect 1596 97617 1624 102575
rect 580920 99521 580948 103527
rect 580906 99512 580962 99521
rect 580906 99447 580962 99456
rect 1582 97608 1638 97617
rect 1582 97543 1638 97552
rect 580906 90264 580962 90273
rect 580906 90199 580962 90208
rect 1582 89856 1638 89865
rect 1582 89791 1638 89800
rect 1596 84697 1624 89791
rect 580920 86193 580948 90199
rect 580906 86184 580962 86193
rect 580906 86119 580962 86128
rect 1582 84688 1638 84697
rect 1582 84623 1638 84632
rect 579894 77344 579950 77353
rect 579894 77279 579950 77288
rect 1582 77072 1638 77081
rect 1582 77007 1638 77016
rect 1596 71641 1624 77007
rect 579908 73001 579936 77279
rect 579894 72992 579950 73001
rect 579894 72927 579950 72936
rect 1582 71632 1638 71641
rect 1582 71567 1638 71576
rect 1490 64288 1546 64297
rect 1490 64223 1546 64232
rect 1504 58585 1532 64223
rect 580906 64152 580962 64161
rect 580906 64087 580962 64096
rect 580920 59673 580948 64087
rect 580906 59664 580962 59673
rect 580906 59599 580962 59608
rect 1490 58576 1546 58585
rect 1490 58511 1546 58520
rect 2778 51504 2834 51513
rect 2778 51439 2834 51448
rect 2792 45529 2820 51439
rect 580906 51096 580962 51105
rect 580906 51031 580962 51040
rect 580920 46345 580948 51031
rect 580906 46336 580962 46345
rect 580906 46271 580962 46280
rect 2778 45520 2834 45529
rect 2778 45455 2834 45464
rect 2778 38720 2834 38729
rect 2778 38655 2834 38664
rect 2792 32473 2820 38655
rect 580906 38040 580962 38049
rect 580906 37975 580962 37984
rect 580920 33153 580948 37975
rect 580906 33144 580962 33153
rect 580906 33079 580962 33088
rect 2778 32464 2834 32473
rect 2778 32399 2834 32408
rect 1490 25936 1546 25945
rect 1490 25871 1546 25880
rect 1504 19417 1532 25871
rect 580906 24984 580962 24993
rect 580906 24919 580962 24928
rect 580920 19825 580948 24919
rect 580906 19816 580962 19825
rect 580906 19751 580962 19760
rect 1490 19408 1546 19417
rect 1490 19343 1546 19352
rect 2778 13152 2834 13161
rect 2778 13087 2834 13096
rect 2792 6497 2820 13087
rect 579894 12744 579950 12753
rect 579894 12679 579950 12688
rect 579908 6633 579936 12679
rect 579894 6624 579950 6633
rect 579894 6559 579950 6568
rect 2778 6488 2834 6497
rect 2778 6423 2834 6432
rect 87984 4010 88274 4026
rect 73528 4004 73580 4010
rect 73528 3946 73580 3952
rect 87972 4004 88274 4010
rect 88024 3998 88274 4004
rect 87972 3946 88024 3952
rect 64328 3936 64380 3942
rect 64328 3878 64380 3884
rect 58808 3800 58860 3806
rect 58808 3742 58860 3748
rect 56968 3596 57020 3602
rect 56968 3538 57020 3544
rect 52552 3392 52604 3398
rect 52552 3334 52604 3340
rect 48964 3324 49016 3330
rect 48964 3266 49016 3272
rect 40408 3256 40460 3262
rect 40408 3198 40460 3204
rect 19432 944 19484 950
rect 19432 886 19484 892
rect 11152 876 11204 882
rect 11152 818 11204 824
rect 3240 536 3292 542
rect 542 82 654 480
rect 1646 218 1758 480
rect 1504 202 1758 218
rect 1492 196 1758 202
rect 1544 190 1758 196
rect 1492 138 1544 144
rect 400 66 654 82
rect 388 60 654 66
rect 440 54 654 60
rect 388 2 440 8
rect 542 -960 654 54
rect 1646 -960 1758 190
rect 2842 354 2954 480
rect 3240 478 3292 484
rect 11164 480 11192 818
rect 14740 740 14792 746
rect 14740 682 14792 688
rect 12162 504 12218 513
rect 3252 354 3280 478
rect 2842 326 3280 354
rect 2842 -960 2954 326
rect 3884 264 3936 270
rect 4038 218 4150 480
rect 3936 212 4150 218
rect 3884 206 4150 212
rect 3896 190 4150 206
rect 4038 -960 4150 190
rect 5234 218 5346 480
rect 5446 232 5502 241
rect 5234 190 5446 218
rect 5234 -960 5346 190
rect 5446 167 5502 176
rect 6274 96 6330 105
rect 6430 82 6542 480
rect 6330 54 6542 82
rect 6274 31 6330 40
rect 6430 -960 6542 54
rect 7626 82 7738 480
rect 8730 354 8842 480
rect 9128 468 9180 474
rect 9128 410 9180 416
rect 9140 354 9168 410
rect 8730 326 9168 354
rect 9772 400 9824 406
rect 9926 354 10038 480
rect 9824 348 10038 354
rect 9772 342 10038 348
rect 9784 326 10038 342
rect 8024 128 8076 134
rect 7626 76 8024 82
rect 7626 70 8076 76
rect 7626 54 8064 70
rect 7626 -960 7738 54
rect 8730 -960 8842 326
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 14752 480 14780 682
rect 18236 672 18288 678
rect 18236 614 18288 620
rect 15936 604 15988 610
rect 15936 546 15988 552
rect 15948 480 15976 546
rect 18248 480 18276 614
rect 19444 480 19472 886
rect 12162 439 12218 448
rect 12176 354 12204 439
rect 12318 354 12430 480
rect 12176 326 12430 354
rect 12318 -960 12430 326
rect 13514 354 13626 480
rect 13726 368 13782 377
rect 13514 326 13726 354
rect 13514 -960 13626 326
rect 13726 303 13782 312
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 354 17122 480
rect 17010 338 17448 354
rect 17010 332 17460 338
rect 17010 326 17408 332
rect 17010 -960 17122 326
rect 17408 274 17460 280
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 19812 66 19840 3060
rect 20628 808 20680 814
rect 20628 750 20680 756
rect 20640 480 20668 750
rect 19800 60 19852 66
rect 19800 2 19852 8
rect 20598 -960 20710 480
rect 20916 202 20944 3060
rect 21824 1012 21876 1018
rect 21824 954 21876 960
rect 21836 480 21864 954
rect 22020 542 22048 3060
rect 22008 536 22060 542
rect 20904 196 20956 202
rect 20904 138 20956 144
rect 21794 -960 21906 480
rect 22008 478 22060 484
rect 22836 536 22888 542
rect 22836 478 22888 484
rect 22848 354 22876 478
rect 22990 354 23102 480
rect 22848 326 23102 354
rect 22990 -960 23102 326
rect 23216 270 23244 3060
rect 23952 3046 24242 3074
rect 25056 3046 25346 3074
rect 26344 3046 26450 3074
rect 23204 264 23256 270
rect 23952 241 23980 3046
rect 23204 206 23256 212
rect 23938 232 23994 241
rect 23938 167 23994 176
rect 24186 218 24298 480
rect 24186 202 24624 218
rect 24186 196 24636 202
rect 24186 190 24584 196
rect 24186 -960 24298 190
rect 24584 138 24636 144
rect 25056 105 25084 3046
rect 25290 218 25402 480
rect 25686 232 25742 241
rect 25290 190 25686 218
rect 25042 96 25098 105
rect 25042 31 25098 40
rect 25290 -960 25402 190
rect 25686 167 25742 176
rect 26344 134 26372 3046
rect 26608 2916 26660 2922
rect 26608 2858 26660 2864
rect 26620 1442 26648 2858
rect 26528 1414 26648 1442
rect 26528 480 26556 1414
rect 26332 128 26384 134
rect 26332 70 26384 76
rect 26486 -960 26598 480
rect 27540 474 27568 3060
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 27724 480 27752 2790
rect 27528 468 27580 474
rect 27528 410 27580 416
rect 27682 -960 27794 480
rect 28644 406 28672 3060
rect 29748 882 29776 3060
rect 29736 876 29788 882
rect 29736 818 29788 824
rect 28906 640 28962 649
rect 28906 575 28962 584
rect 28920 480 28948 575
rect 30852 513 30880 3060
rect 30838 504 30894 513
rect 28632 400 28684 406
rect 28632 342 28684 348
rect 28878 -960 28990 480
rect 30074 82 30186 480
rect 30838 439 30894 448
rect 31116 128 31168 134
rect 30074 66 30328 82
rect 31270 82 31382 480
rect 31956 377 31984 3060
rect 33060 746 33088 3060
rect 33600 2984 33652 2990
rect 33600 2926 33652 2932
rect 33048 740 33100 746
rect 33048 682 33100 688
rect 33612 480 33640 2926
rect 34164 610 34192 3060
rect 34152 604 34204 610
rect 34152 546 34204 552
rect 34796 604 34848 610
rect 34796 546 34848 552
rect 34808 480 34836 546
rect 32220 468 32272 474
rect 32220 410 32272 416
rect 31942 368 31998 377
rect 32232 354 32260 410
rect 32374 354 32486 480
rect 32232 326 32486 354
rect 31942 303 31998 312
rect 31168 76 31382 82
rect 31116 70 31382 76
rect 30074 60 30340 66
rect 30074 54 30288 60
rect 30074 -960 30186 54
rect 31128 54 31382 70
rect 30288 2 30340 8
rect 31270 -960 31382 54
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35268 338 35296 3060
rect 36372 746 36400 3060
rect 37476 950 37504 3060
rect 37464 944 37516 950
rect 37464 886 37516 892
rect 38580 814 38608 3060
rect 39684 1018 39712 3060
rect 39672 1012 39724 1018
rect 39672 954 39724 960
rect 38568 808 38620 814
rect 38568 750 38620 756
rect 36360 740 36412 746
rect 36360 682 36412 688
rect 35992 672 36044 678
rect 35992 614 36044 620
rect 36004 480 36032 614
rect 35256 332 35308 338
rect 35256 274 35308 280
rect 35962 -960 36074 480
rect 37002 96 37058 105
rect 37158 82 37270 480
rect 37058 54 37270 82
rect 37002 31 37058 40
rect 37158 -960 37270 54
rect 38354 354 38466 480
rect 39396 400 39448 406
rect 38354 338 38608 354
rect 39550 354 39662 480
rect 39448 348 39662 354
rect 39396 342 39662 348
rect 38354 332 38620 338
rect 38354 326 38568 332
rect 38354 -960 38466 326
rect 39408 326 39662 342
rect 40420 354 40448 3198
rect 40512 3046 40802 3074
rect 41616 3046 41906 3074
rect 42812 3046 43010 3074
rect 43824 3046 44114 3074
rect 44928 3046 45218 3074
rect 40512 542 40540 3046
rect 40500 536 40552 542
rect 40500 478 40552 484
rect 40654 354 40766 480
rect 40420 326 40766 354
rect 38568 274 38620 280
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41616 202 41644 3046
rect 41850 218 41962 480
rect 42248 264 42300 270
rect 41850 212 42248 218
rect 41850 206 42300 212
rect 42706 232 42762 241
rect 41604 196 41656 202
rect 41604 138 41656 144
rect 41850 190 42288 206
rect 41850 -960 41962 190
rect 42812 218 42840 3046
rect 43824 2922 43852 3046
rect 43812 2916 43864 2922
rect 43812 2858 43864 2864
rect 44272 2916 44324 2922
rect 44272 2858 44324 2864
rect 44284 480 44312 2858
rect 44928 2854 44956 3046
rect 44916 2848 44968 2854
rect 44916 2790 44968 2796
rect 46308 649 46336 3060
rect 46294 640 46350 649
rect 46294 575 46350 584
rect 45284 536 45336 542
rect 43046 218 43158 480
rect 42762 190 42840 218
rect 42904 202 43158 218
rect 42892 196 43158 202
rect 42706 167 42762 176
rect 42944 190 43158 196
rect 42892 138 42944 144
rect 43046 -960 43158 190
rect 44242 -960 44354 480
rect 45284 478 45336 484
rect 45296 354 45324 478
rect 45438 354 45550 480
rect 45296 326 45550 354
rect 45438 -960 45550 326
rect 46634 218 46746 480
rect 46846 232 46902 241
rect 46634 190 46846 218
rect 46634 -960 46746 190
rect 46846 167 46902 176
rect 47412 66 47440 3060
rect 47860 3052 47912 3058
rect 47860 2994 47912 3000
rect 47872 480 47900 2994
rect 47400 60 47452 66
rect 47400 2 47452 8
rect 47830 -960 47942 480
rect 48516 134 48544 3060
rect 48976 480 49004 3266
rect 51356 3188 51408 3194
rect 51356 3130 51408 3136
rect 48504 128 48556 134
rect 48504 70 48556 76
rect 48934 -960 49046 480
rect 49620 474 49648 3060
rect 50448 3046 50738 3074
rect 50448 2990 50476 3046
rect 50436 2984 50488 2990
rect 50436 2926 50488 2932
rect 50160 2848 50212 2854
rect 50160 2790 50212 2796
rect 50172 480 50200 2790
rect 51368 480 51396 3130
rect 51828 610 51856 3060
rect 51816 604 51868 610
rect 51816 546 51868 552
rect 52564 480 52592 3334
rect 56048 3120 56100 3126
rect 56048 3062 56100 3068
rect 52932 678 52960 3060
rect 52920 672 52972 678
rect 52920 614 52972 620
rect 49608 468 49660 474
rect 49608 410 49660 416
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 82 53830 480
rect 54036 105 54064 3060
rect 54944 2984 54996 2990
rect 54944 2926 54996 2932
rect 54956 480 54984 2926
rect 53576 66 53830 82
rect 53564 60 53830 66
rect 53616 54 53830 60
rect 53564 2 53616 8
rect 53718 -960 53830 54
rect 54022 96 54078 105
rect 54022 31 54078 40
rect 54914 -960 55026 480
rect 55140 338 55168 3060
rect 56060 480 56088 3062
rect 55128 332 55180 338
rect 55128 274 55180 280
rect 56018 -960 56130 480
rect 56244 406 56272 3060
rect 56232 400 56284 406
rect 56232 342 56284 348
rect 56980 354 57008 3538
rect 57060 3256 57112 3262
rect 57112 3204 57362 3210
rect 57060 3198 57362 3204
rect 57072 3182 57362 3198
rect 58176 3046 58466 3074
rect 57214 354 57326 480
rect 56980 326 57326 354
rect 57214 -960 57326 326
rect 58176 270 58204 3046
rect 58410 354 58522 480
rect 58820 354 58848 3742
rect 63224 3732 63276 3738
rect 63224 3674 63276 3680
rect 60832 3664 60884 3670
rect 60832 3606 60884 3612
rect 59728 3460 59780 3466
rect 59728 3402 59780 3408
rect 58410 326 58848 354
rect 59372 3046 59570 3074
rect 58164 264 58216 270
rect 58164 206 58216 212
rect 58410 -960 58522 326
rect 59372 202 59400 3046
rect 59740 1714 59768 3402
rect 60384 3046 60674 3074
rect 60384 2922 60412 3046
rect 60372 2916 60424 2922
rect 60372 2858 60424 2864
rect 59648 1686 59768 1714
rect 59648 480 59676 1686
rect 60844 480 60872 3606
rect 62028 3324 62080 3330
rect 62028 3266 62080 3272
rect 61764 542 61792 3060
rect 61752 536 61804 542
rect 59360 196 59412 202
rect 59360 138 59412 144
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61752 478 61804 484
rect 62040 480 62068 3266
rect 61998 -960 62110 480
rect 62868 241 62896 3060
rect 63236 480 63264 3674
rect 63696 3058 63986 3074
rect 63684 3052 63986 3058
rect 63736 3046 63986 3052
rect 63684 2994 63736 3000
rect 64340 480 64368 3878
rect 70124 3868 70176 3874
rect 70124 3810 70176 3816
rect 68100 3392 68152 3398
rect 68560 3392 68612 3398
rect 68152 3340 68402 3346
rect 68100 3334 68402 3340
rect 68560 3334 68612 3340
rect 68112 3318 68402 3334
rect 64696 3256 64748 3262
rect 64696 3198 64748 3204
rect 66720 3256 66772 3262
rect 66720 3198 66772 3204
rect 64708 3074 64736 3198
rect 64708 3046 65090 3074
rect 65904 3046 66194 3074
rect 65524 2916 65576 2922
rect 65524 2858 65576 2864
rect 65536 480 65564 2858
rect 65904 2854 65932 3046
rect 65892 2848 65944 2854
rect 65892 2790 65944 2796
rect 66732 480 66760 3198
rect 67008 3194 67298 3210
rect 66996 3188 67298 3194
rect 67048 3182 67298 3188
rect 66996 3130 67048 3136
rect 68572 2854 68600 3334
rect 69112 2984 69164 2990
rect 69112 2926 69164 2932
rect 67916 2848 67968 2854
rect 67916 2790 67968 2796
rect 68560 2848 68612 2854
rect 68560 2790 68612 2796
rect 67928 480 67956 2790
rect 69124 480 69152 2926
rect 62854 232 62910 241
rect 62854 167 62910 176
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69492 66 69520 3060
rect 70136 218 70164 3810
rect 72528 3726 72818 3754
rect 72528 3602 72556 3726
rect 72516 3596 72568 3602
rect 72516 3538 72568 3544
rect 72608 3596 72660 3602
rect 72608 3538 72660 3544
rect 71320 3528 71372 3534
rect 71320 3470 71372 3476
rect 70320 3058 70610 3074
rect 70308 3052 70610 3058
rect 70360 3046 70610 3052
rect 70308 2994 70360 3000
rect 71332 1850 71360 3470
rect 71412 3120 71464 3126
rect 71464 3068 71714 3074
rect 71412 3062 71714 3068
rect 71424 3046 71714 3062
rect 71332 1822 71544 1850
rect 71516 480 71544 1822
rect 72620 480 72648 3538
rect 70278 218 70390 480
rect 70136 190 70390 218
rect 69480 60 69532 66
rect 69480 2 69532 8
rect 70278 -960 70390 190
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73540 354 73568 3946
rect 79140 3936 79192 3942
rect 79192 3884 79442 3890
rect 79140 3878 79442 3884
rect 79152 3862 79442 3878
rect 84672 3874 84962 3890
rect 112272 3874 112562 3890
rect 84660 3868 84962 3874
rect 84712 3862 84962 3868
rect 99840 3868 99892 3874
rect 84660 3810 84712 3816
rect 99840 3810 99892 3816
rect 112260 3868 112562 3874
rect 112312 3862 112562 3868
rect 112260 3810 112312 3816
rect 73620 3800 73672 3806
rect 77392 3800 77444 3806
rect 73672 3748 73922 3754
rect 73620 3742 73922 3748
rect 91284 3800 91336 3806
rect 77392 3742 77444 3748
rect 73632 3726 73922 3742
rect 75828 3664 75880 3670
rect 75880 3612 76130 3618
rect 75828 3606 76130 3612
rect 75840 3590 76130 3606
rect 74460 3466 75026 3482
rect 74448 3460 75026 3466
rect 74500 3454 75026 3460
rect 75368 3460 75420 3466
rect 74448 3402 74500 3408
rect 75368 3402 75420 3408
rect 73774 354 73886 480
rect 73540 326 73886 354
rect 73774 -960 73886 326
rect 74970 354 75082 480
rect 75380 354 75408 3402
rect 76944 3330 77234 3346
rect 76932 3324 77234 3330
rect 76984 3318 77234 3324
rect 76932 3266 76984 3272
rect 76288 3052 76340 3058
rect 76288 2994 76340 3000
rect 76300 1578 76328 2994
rect 76208 1550 76328 1578
rect 76208 480 76236 1550
rect 77404 480 77432 3742
rect 78048 3738 78338 3754
rect 91336 3748 91586 3754
rect 91284 3742 91586 3748
rect 78036 3732 78338 3738
rect 78088 3726 78338 3732
rect 83280 3732 83332 3738
rect 78036 3674 78088 3680
rect 91296 3726 91586 3742
rect 96816 3738 97106 3754
rect 96804 3732 97106 3738
rect 83280 3674 83332 3680
rect 96856 3726 97106 3732
rect 98920 3732 98972 3738
rect 96804 3674 96856 3680
rect 98920 3674 98972 3680
rect 79692 3664 79744 3670
rect 79692 3606 79744 3612
rect 78588 2916 78640 2922
rect 78588 2858 78640 2864
rect 78600 480 78628 2858
rect 79704 480 79732 3606
rect 82452 3392 82504 3398
rect 82504 3340 82754 3346
rect 82452 3334 82754 3340
rect 82464 3318 82754 3334
rect 80888 3256 80940 3262
rect 80888 3198 80940 3204
rect 79980 3046 80546 3074
rect 79980 2854 80008 3046
rect 79968 2848 80020 2854
rect 79968 2790 80020 2796
rect 80900 480 80928 3198
rect 81360 3194 81650 3210
rect 81348 3188 81650 3194
rect 81400 3182 81650 3188
rect 82084 3188 82136 3194
rect 81348 3130 81400 3136
rect 82084 3130 82136 3136
rect 82096 480 82124 3130
rect 83292 480 83320 3674
rect 93492 3664 93544 3670
rect 86880 3602 87170 3618
rect 95148 3664 95200 3670
rect 93544 3612 93794 3618
rect 93492 3606 93794 3612
rect 95148 3606 95200 3612
rect 86868 3596 87170 3602
rect 86920 3590 87170 3596
rect 89536 3596 89588 3602
rect 86868 3538 86920 3544
rect 93504 3590 93794 3606
rect 89536 3538 89588 3544
rect 85764 3528 85816 3534
rect 85816 3476 86066 3482
rect 85764 3470 86066 3476
rect 85776 3454 86066 3470
rect 89088 3466 89378 3482
rect 89076 3460 89378 3466
rect 89128 3454 89378 3460
rect 89076 3402 89128 3408
rect 85672 3324 85724 3330
rect 85672 3266 85724 3272
rect 83844 2990 83872 3060
rect 83832 2984 83884 2990
rect 83832 2926 83884 2932
rect 84476 2984 84528 2990
rect 84476 2926 84528 2932
rect 84488 480 84516 2926
rect 85684 480 85712 3266
rect 87972 3120 88024 3126
rect 87972 3062 88024 3068
rect 86868 2848 86920 2854
rect 86868 2790 86920 2796
rect 86880 480 86908 2790
rect 87984 480 88012 3062
rect 74970 326 75408 354
rect 74970 -960 75082 326
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 354 89250 480
rect 89548 354 89576 3538
rect 93952 3460 94004 3466
rect 93952 3402 94004 3408
rect 90088 3392 90140 3398
rect 90088 3334 90140 3340
rect 89138 326 89576 354
rect 90100 354 90128 3334
rect 90192 3058 90482 3074
rect 90180 3052 90482 3058
rect 90232 3046 90482 3052
rect 91928 3052 91980 3058
rect 90180 2994 90232 3000
rect 91928 2994 91980 3000
rect 92492 3046 92690 3074
rect 90334 354 90446 480
rect 90100 326 90446 354
rect 89138 -960 89250 326
rect 90334 -960 90446 326
rect 91530 354 91642 480
rect 91940 354 91968 2994
rect 92492 2922 92520 3046
rect 92480 2916 92532 2922
rect 92480 2858 92532 2864
rect 92756 2916 92808 2922
rect 92756 2858 92808 2864
rect 92768 480 92796 2858
rect 93964 480 93992 3402
rect 94596 3256 94648 3262
rect 94648 3204 94898 3210
rect 94596 3198 94898 3204
rect 94608 3182 94898 3198
rect 95160 480 95188 3606
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 96252 3256 96304 3262
rect 95712 3194 96002 3210
rect 96252 3198 96304 3204
rect 95700 3188 96002 3194
rect 95752 3182 96002 3188
rect 95700 3130 95752 3136
rect 96264 480 96292 3198
rect 97448 3188 97500 3194
rect 97448 3130 97500 3136
rect 97460 480 97488 3130
rect 98196 2990 98224 3060
rect 98184 2984 98236 2990
rect 98184 2926 98236 2932
rect 98656 480 98684 3470
rect 98932 3398 98960 3674
rect 98920 3392 98972 3398
rect 98920 3334 98972 3340
rect 99024 3330 99314 3346
rect 99012 3324 99314 3330
rect 99064 3318 99314 3324
rect 99012 3266 99064 3272
rect 99852 480 99880 3810
rect 105728 3800 105780 3806
rect 103440 3738 103730 3754
rect 105728 3742 105780 3748
rect 117780 3800 117832 3806
rect 125968 3800 126020 3806
rect 117832 3748 118082 3754
rect 117780 3742 118082 3748
rect 136640 3800 136692 3806
rect 125968 3742 126020 3748
rect 103428 3732 103730 3738
rect 103480 3726 103730 3732
rect 103428 3674 103480 3680
rect 102336 3602 102626 3618
rect 102324 3596 102626 3602
rect 102376 3590 102626 3596
rect 103336 3596 103388 3602
rect 102324 3538 102376 3544
rect 103336 3538 103388 3544
rect 100760 3460 100812 3466
rect 100760 3402 100812 3408
rect 100404 2854 100432 3060
rect 100392 2848 100444 2854
rect 100392 2790 100444 2796
rect 100772 1290 100800 3402
rect 101036 3392 101088 3398
rect 101036 3334 101088 3340
rect 100760 1284 100812 1290
rect 100760 1226 100812 1232
rect 101048 480 101076 3334
rect 101220 3120 101272 3126
rect 102232 3120 102284 3126
rect 101272 3068 101522 3074
rect 101220 3062 101522 3068
rect 102232 3062 102284 3068
rect 101232 3046 101522 3062
rect 102244 480 102272 3062
rect 103348 480 103376 3538
rect 104544 3058 104834 3074
rect 104532 3052 104834 3058
rect 104584 3046 104834 3052
rect 104532 2994 104584 3000
rect 104532 2848 104584 2854
rect 104532 2790 104584 2796
rect 104544 480 104572 2790
rect 105740 480 105768 3742
rect 117792 3726 118082 3742
rect 118792 3732 118844 3738
rect 118792 3674 118844 3680
rect 107844 3664 107896 3670
rect 117596 3664 117648 3670
rect 107896 3612 108146 3618
rect 107844 3606 108146 3612
rect 107856 3590 108146 3606
rect 115584 3602 115874 3618
rect 117596 3606 117648 3612
rect 115572 3596 115874 3602
rect 115624 3590 115874 3596
rect 115572 3538 115624 3544
rect 111156 3528 111208 3534
rect 109052 3466 109250 3482
rect 111208 3476 111458 3482
rect 111156 3470 111458 3476
rect 109040 3460 109250 3466
rect 109092 3454 109250 3460
rect 111168 3454 111458 3470
rect 116400 3460 116452 3466
rect 109040 3402 109092 3408
rect 116400 3402 116452 3408
rect 114008 3392 114060 3398
rect 114008 3334 114060 3340
rect 109408 3324 109460 3330
rect 109408 3266 109460 3272
rect 105924 2922 105952 3060
rect 106924 2984 106976 2990
rect 106924 2926 106976 2932
rect 105912 2916 105964 2922
rect 105912 2858 105964 2864
rect 106936 480 106964 2926
rect 107028 1290 107056 3060
rect 108488 3052 108540 3058
rect 108488 2994 108540 3000
rect 107016 1284 107068 1290
rect 107016 1226 107068 1232
rect 91530 326 91968 354
rect 91530 -960 91642 326
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 354 108202 480
rect 108500 354 108528 2994
rect 109420 1714 109448 3266
rect 113088 3256 113140 3262
rect 110064 3194 110354 3210
rect 113140 3204 113666 3210
rect 113088 3198 113666 3204
rect 110052 3188 110354 3194
rect 110104 3182 110354 3188
rect 110880 3188 110932 3194
rect 110052 3130 110104 3136
rect 113100 3182 113666 3198
rect 110880 3130 110932 3136
rect 110512 2848 110564 2854
rect 110512 2790 110564 2796
rect 109328 1686 109448 1714
rect 109328 480 109356 1686
rect 110524 1290 110552 2790
rect 110512 1284 110564 1290
rect 110512 1226 110564 1232
rect 108090 326 108528 354
rect 108090 -960 108202 326
rect 109286 -960 109398 480
rect 110482 218 110594 480
rect 110892 218 110920 3130
rect 112812 2916 112864 2922
rect 112812 2858 112864 2864
rect 111616 2848 111668 2854
rect 111616 2790 111668 2796
rect 111628 480 111656 2790
rect 112824 480 112852 2858
rect 114020 480 114048 3334
rect 114560 3120 114612 3126
rect 115204 3120 115256 3126
rect 114612 3068 114770 3074
rect 114560 3062 114770 3068
rect 115204 3062 115256 3068
rect 114572 3046 114770 3062
rect 115216 480 115244 3062
rect 116412 480 116440 3402
rect 116964 1290 116992 3060
rect 116952 1284 117004 1290
rect 116952 1226 117004 1232
rect 117608 480 117636 3606
rect 118804 480 118832 3674
rect 120908 3596 120960 3602
rect 120908 3538 120960 3544
rect 119172 2990 119200 3060
rect 120000 3058 120290 3074
rect 119988 3052 120290 3058
rect 120040 3046 120290 3052
rect 119988 2994 120040 3000
rect 119160 2984 119212 2990
rect 119160 2926 119212 2932
rect 119896 2984 119948 2990
rect 119896 2926 119948 2932
rect 119908 480 119936 2926
rect 110482 190 110920 218
rect 110482 -960 110594 190
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120920 218 120948 3538
rect 125600 3392 125652 3398
rect 121104 3330 121394 3346
rect 121092 3324 121394 3330
rect 121144 3318 121394 3324
rect 122208 3318 122498 3346
rect 125652 3340 125810 3346
rect 125600 3334 125810 3340
rect 125612 3318 125810 3334
rect 121092 3266 121144 3272
rect 122208 3194 122236 3318
rect 122288 3256 122340 3262
rect 122288 3198 122340 3204
rect 122196 3188 122248 3194
rect 122196 3130 122248 3136
rect 122300 480 122328 3198
rect 123588 2854 123616 3060
rect 124692 2922 124720 3060
rect 124680 2916 124732 2922
rect 124680 2858 124732 2864
rect 125048 2916 125100 2922
rect 125048 2858 125100 2864
rect 123576 2848 123628 2854
rect 123576 2790 123628 2796
rect 123484 2780 123536 2786
rect 123484 2722 123536 2728
rect 123496 480 123524 2722
rect 121062 218 121174 480
rect 120920 190 121174 218
rect 121062 -960 121174 190
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 354 124762 480
rect 125060 354 125088 2858
rect 125980 1986 126008 3742
rect 129936 3738 130226 3754
rect 136692 3748 136850 3754
rect 136640 3742 136850 3748
rect 129924 3732 130226 3738
rect 129976 3726 130226 3732
rect 136652 3726 136850 3742
rect 129924 3674 129976 3680
rect 128820 3664 128872 3670
rect 144736 3664 144788 3670
rect 128872 3612 129122 3618
rect 128820 3606 129122 3612
rect 128832 3590 129122 3606
rect 132144 3602 132434 3618
rect 143184 3602 143474 3618
rect 144736 3606 144788 3612
rect 154212 3664 154264 3670
rect 154264 3612 154514 3618
rect 154212 3606 154514 3612
rect 132132 3596 132434 3602
rect 132184 3590 132434 3596
rect 132960 3596 133012 3602
rect 132132 3538 132184 3544
rect 132960 3538 133012 3544
rect 143172 3596 143474 3602
rect 143224 3590 143474 3596
rect 143172 3538 143224 3544
rect 129372 3528 129424 3534
rect 127728 3466 128018 3482
rect 129372 3470 129424 3476
rect 127716 3460 128018 3466
rect 127768 3454 128018 3460
rect 127716 3402 127768 3408
rect 127072 3392 127124 3398
rect 127072 3334 127124 3340
rect 126612 3120 126664 3126
rect 126664 3068 126914 3074
rect 126612 3062 126914 3068
rect 126624 3046 126914 3062
rect 125888 1958 126008 1986
rect 125888 480 125916 1958
rect 127084 1714 127112 3334
rect 128176 3052 128228 3058
rect 128176 2994 128228 3000
rect 126992 1686 127112 1714
rect 126992 480 127020 1686
rect 128188 480 128216 2994
rect 129384 480 129412 3470
rect 130568 3324 130620 3330
rect 130568 3266 130620 3272
rect 130580 480 130608 3266
rect 131316 2990 131344 3060
rect 131304 2984 131356 2990
rect 131304 2926 131356 2932
rect 131764 2984 131816 2990
rect 131764 2926 131816 2932
rect 131776 480 131804 2926
rect 132972 480 133000 3538
rect 139860 3528 139912 3534
rect 142528 3528 142580 3534
rect 139912 3476 140162 3482
rect 139860 3470 140162 3476
rect 142528 3470 142580 3476
rect 137468 3460 137520 3466
rect 139872 3454 140162 3470
rect 137468 3402 137520 3408
rect 133236 3256 133288 3262
rect 133288 3204 133538 3210
rect 133236 3198 133538 3204
rect 133248 3182 133538 3198
rect 135260 3188 135312 3194
rect 135260 3130 135312 3136
rect 134156 3120 134208 3126
rect 134156 3062 134208 3068
rect 134168 480 134196 3062
rect 134628 2854 134656 3060
rect 134616 2848 134668 2854
rect 134616 2790 134668 2796
rect 135272 480 135300 3130
rect 135732 2922 135760 3060
rect 135720 2916 135772 2922
rect 135720 2858 135772 2864
rect 136456 2848 136508 2854
rect 136456 2790 136508 2796
rect 136468 480 136496 2790
rect 124650 326 125088 354
rect 124650 -960 124762 326
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137480 218 137508 3402
rect 137652 3392 137704 3398
rect 137704 3340 137954 3346
rect 137652 3334 137954 3340
rect 137664 3318 137954 3334
rect 140976 3330 141266 3346
rect 140964 3324 141266 3330
rect 141016 3318 141266 3324
rect 140964 3266 141016 3272
rect 139216 3256 139268 3262
rect 139216 3198 139268 3204
rect 138768 3058 139058 3074
rect 138756 3052 139058 3058
rect 138808 3046 139058 3052
rect 138756 2994 138808 3000
rect 137622 218 137734 480
rect 137480 190 137734 218
rect 137622 -960 137734 190
rect 138818 354 138930 480
rect 139228 354 139256 3198
rect 140044 3052 140096 3058
rect 140044 2994 140096 3000
rect 140056 480 140084 2994
rect 142356 2990 142384 3060
rect 142344 2984 142396 2990
rect 142344 2926 142396 2932
rect 141240 2916 141292 2922
rect 141240 2858 141292 2864
rect 141252 480 141280 2858
rect 142540 1850 142568 3470
rect 143632 3324 143684 3330
rect 143632 3266 143684 3272
rect 142448 1822 142568 1850
rect 142448 480 142476 1822
rect 143644 1714 143672 3266
rect 144276 3120 144328 3126
rect 144328 3068 144578 3074
rect 144276 3062 144578 3068
rect 144288 3046 144578 3062
rect 143552 1686 143672 1714
rect 143552 480 143580 1686
rect 144748 480 144776 3606
rect 148324 3596 148376 3602
rect 154224 3590 154514 3606
rect 157536 3602 157826 3618
rect 157524 3596 157826 3602
rect 148324 3538 148376 3544
rect 157576 3590 157826 3596
rect 157524 3538 157576 3544
rect 147680 3392 147732 3398
rect 147732 3340 147890 3346
rect 147680 3334 147890 3340
rect 147692 3318 147890 3334
rect 145392 3194 145682 3210
rect 145380 3188 145682 3194
rect 145432 3182 145682 3188
rect 147128 3188 147180 3194
rect 145380 3130 145432 3136
rect 147128 3130 147180 3136
rect 145932 2984 145984 2990
rect 145932 2926 145984 2932
rect 145944 480 145972 2926
rect 146772 2854 146800 3060
rect 146760 2848 146812 2854
rect 146760 2790 146812 2796
rect 147140 480 147168 3130
rect 148336 480 148364 3538
rect 152004 3528 152056 3534
rect 163688 3528 163740 3534
rect 152056 3476 152306 3482
rect 152004 3470 152306 3476
rect 152016 3454 152306 3470
rect 161952 3466 162242 3482
rect 163688 3470 163740 3476
rect 171876 3528 171928 3534
rect 171928 3476 172178 3482
rect 171876 3470 172178 3476
rect 153016 3460 153068 3466
rect 153016 3402 153068 3408
rect 161940 3460 162242 3466
rect 161992 3454 162242 3460
rect 161940 3402 161992 3408
rect 148692 3256 148744 3262
rect 150624 3256 150676 3262
rect 148744 3204 148994 3210
rect 148692 3198 148994 3204
rect 150624 3198 150676 3204
rect 148704 3182 148994 3198
rect 149808 3058 150098 3074
rect 149796 3052 150098 3058
rect 149848 3046 150098 3052
rect 149796 2994 149848 3000
rect 149520 2848 149572 2854
rect 149520 2790 149572 2796
rect 149532 480 149560 2790
rect 150636 480 150664 3198
rect 151820 3120 151872 3126
rect 151820 3062 151872 3068
rect 151188 2922 151216 3060
rect 151176 2916 151228 2922
rect 151176 2858 151228 2864
rect 151832 480 151860 3062
rect 153028 480 153056 3402
rect 155408 3392 155460 3398
rect 153212 3330 153410 3346
rect 155408 3334 155460 3340
rect 153200 3324 153410 3330
rect 153252 3318 153410 3324
rect 154212 3324 154264 3330
rect 153200 3266 153252 3272
rect 154212 3266 154264 3272
rect 154224 480 154252 3266
rect 155420 480 155448 3334
rect 163056 3330 163346 3346
rect 163044 3324 163346 3330
rect 163096 3318 163346 3324
rect 163044 3266 163096 3272
rect 159732 3256 159784 3262
rect 156432 3194 156722 3210
rect 161296 3256 161348 3262
rect 159784 3204 160034 3210
rect 159732 3198 160034 3204
rect 161296 3198 161348 3204
rect 156420 3188 156722 3194
rect 156472 3182 156722 3188
rect 159744 3182 160034 3198
rect 156420 3130 156472 3136
rect 160836 3120 160888 3126
rect 155604 2990 155632 3060
rect 156604 3052 156656 3058
rect 156604 2994 156656 3000
rect 158732 3046 158930 3074
rect 160888 3068 161138 3074
rect 160836 3062 161138 3068
rect 160848 3046 161138 3062
rect 155592 2984 155644 2990
rect 155592 2926 155644 2932
rect 156616 480 156644 2994
rect 157800 2984 157852 2990
rect 157800 2926 157852 2932
rect 157812 480 157840 2926
rect 158732 2854 158760 3046
rect 158904 2916 158956 2922
rect 158904 2858 158956 2864
rect 158720 2848 158772 2854
rect 158720 2790 158772 2796
rect 158916 480 158944 2858
rect 160100 2848 160152 2854
rect 160100 2790 160152 2796
rect 160112 480 160140 2790
rect 161308 480 161336 3198
rect 162492 3188 162544 3194
rect 162492 3130 162544 3136
rect 162504 480 162532 3130
rect 163700 480 163728 3470
rect 169576 3460 169628 3466
rect 171888 3454 172178 3470
rect 177408 3466 177698 3482
rect 177396 3460 177698 3466
rect 169576 3402 169628 3408
rect 177448 3454 177698 3460
rect 183744 3460 183796 3466
rect 177396 3402 177448 3408
rect 183744 3402 183796 3408
rect 189552 3454 189842 3482
rect 190656 3466 190946 3482
rect 190644 3460 190946 3466
rect 164240 3392 164292 3398
rect 167184 3392 167236 3398
rect 164292 3340 164450 3346
rect 164240 3334 164450 3340
rect 167184 3334 167236 3340
rect 164252 3318 164450 3334
rect 164884 3324 164936 3330
rect 164884 3266 164936 3272
rect 164240 3120 164292 3126
rect 164240 3062 164292 3068
rect 164252 2854 164280 3062
rect 164240 2848 164292 2854
rect 164240 2790 164292 2796
rect 164896 480 164924 3266
rect 165264 3058 165554 3074
rect 165252 3052 165554 3058
rect 165304 3046 165554 3052
rect 165252 2994 165304 3000
rect 166644 2990 166672 3060
rect 166632 2984 166684 2990
rect 166632 2926 166684 2932
rect 166080 2916 166132 2922
rect 166080 2858 166132 2864
rect 166092 480 166120 2858
rect 167196 480 167224 3334
rect 168564 3120 168616 3126
rect 168616 3068 168866 3074
rect 168564 3062 168866 3068
rect 167748 2854 167776 3060
rect 168576 3046 168866 3062
rect 168380 2916 168432 2922
rect 168380 2858 168432 2864
rect 167736 2848 167788 2854
rect 167736 2790 167788 2796
rect 168392 480 168420 2858
rect 169588 480 169616 3402
rect 175280 3392 175332 3398
rect 172992 3330 173282 3346
rect 180248 3392 180300 3398
rect 175332 3340 175490 3346
rect 175280 3334 175490 3340
rect 180248 3334 180300 3340
rect 172980 3324 173282 3330
rect 173032 3318 173282 3324
rect 174268 3324 174320 3330
rect 172980 3266 173032 3272
rect 175292 3318 175490 3334
rect 174268 3266 174320 3272
rect 169760 3256 169812 3262
rect 173164 3256 173216 3262
rect 169812 3204 169970 3210
rect 169760 3198 169970 3204
rect 173164 3198 173216 3204
rect 169772 3182 169970 3198
rect 170772 3188 170824 3194
rect 170772 3130 170824 3136
rect 170784 480 170812 3130
rect 170864 3120 170916 3126
rect 170916 3068 171074 3074
rect 170864 3062 171074 3068
rect 170876 3046 171074 3062
rect 171968 3052 172020 3058
rect 171968 2994 172020 3000
rect 171980 480 172008 2994
rect 173176 480 173204 3198
rect 174280 480 174308 3266
rect 178512 3194 178802 3210
rect 178500 3188 178802 3194
rect 178552 3182 178802 3188
rect 179052 3188 179104 3194
rect 178500 3130 178552 3136
rect 179052 3130 179104 3136
rect 176752 3120 176804 3126
rect 176752 3062 176804 3068
rect 174372 2990 174400 3060
rect 174360 2984 174412 2990
rect 174360 2926 174412 2932
rect 176580 2922 176608 3060
rect 176568 2916 176620 2922
rect 176568 2858 176620 2864
rect 175464 2848 175516 2854
rect 175464 2790 175516 2796
rect 175476 480 175504 2790
rect 176764 1578 176792 3062
rect 177856 2984 177908 2990
rect 177856 2926 177908 2932
rect 176672 1550 176792 1578
rect 176672 480 176700 1550
rect 177868 480 177896 2926
rect 179064 480 179092 3130
rect 179616 3058 179906 3074
rect 179604 3052 179906 3058
rect 179656 3046 179906 3052
rect 179604 2994 179656 3000
rect 180260 480 180288 3334
rect 181824 3330 182114 3346
rect 181812 3324 182114 3330
rect 181864 3318 182114 3324
rect 181812 3266 181864 3272
rect 180892 3256 180944 3262
rect 182548 3256 182600 3262
rect 180944 3204 181010 3210
rect 180892 3198 181010 3204
rect 182548 3198 182600 3204
rect 180904 3182 181010 3198
rect 181444 2916 181496 2922
rect 181444 2858 181496 2864
rect 181456 480 181484 2858
rect 182560 480 182588 3198
rect 183204 2854 183232 3060
rect 183192 2848 183244 2854
rect 183192 2790 183244 2796
rect 183756 480 183784 3402
rect 187332 3392 187384 3398
rect 187384 3340 187634 3346
rect 187332 3334 187634 3340
rect 187344 3318 187634 3334
rect 189552 3262 189580 3454
rect 190696 3454 190946 3460
rect 190644 3402 190696 3408
rect 196176 3330 196466 3346
rect 189724 3324 189776 3330
rect 189724 3266 189776 3272
rect 196164 3324 196466 3330
rect 196216 3318 196466 3324
rect 559774 3330 560064 3346
rect 559774 3324 560076 3330
rect 559774 3318 560024 3324
rect 196164 3266 196216 3272
rect 560024 3266 560076 3272
rect 578608 3324 578660 3330
rect 578608 3266 578660 3272
rect 189540 3256 189592 3262
rect 186332 3194 186530 3210
rect 189540 3198 189592 3204
rect 186320 3188 186530 3194
rect 186372 3182 186530 3188
rect 186320 3130 186372 3136
rect 184020 3120 184072 3126
rect 184072 3068 184322 3074
rect 184020 3062 184322 3068
rect 184032 3046 184322 3062
rect 185412 2990 185440 3060
rect 187332 3052 187384 3058
rect 187332 2994 187384 3000
rect 188448 3046 188738 3074
rect 185400 2984 185452 2990
rect 185400 2926 185452 2932
rect 186136 2984 186188 2990
rect 186136 2926 186188 2932
rect 184940 2848 184992 2854
rect 184940 2790 184992 2796
rect 184952 480 184980 2790
rect 186148 480 186176 2926
rect 187344 480 187372 2994
rect 188448 2922 188476 3046
rect 188436 2916 188488 2922
rect 188436 2858 188488 2864
rect 188528 2916 188580 2922
rect 188528 2858 188580 2864
rect 188540 480 188568 2858
rect 189736 480 189764 3266
rect 190828 3256 190880 3262
rect 190828 3198 190880 3204
rect 197360 3256 197412 3262
rect 200304 3256 200356 3262
rect 197412 3204 197570 3210
rect 197360 3198 197570 3204
rect 190840 480 190868 3198
rect 192392 3188 192444 3194
rect 197372 3182 197570 3198
rect 198384 3194 198674 3210
rect 200304 3198 200356 3204
rect 206100 3256 206152 3262
rect 553308 3256 553360 3262
rect 206152 3204 206402 3210
rect 206100 3198 206402 3204
rect 198372 3188 198674 3194
rect 192392 3130 192444 3136
rect 198424 3182 198674 3188
rect 198372 3130 198424 3136
rect 192036 2854 192064 3060
rect 192024 2848 192076 2854
rect 192024 2790 192076 2796
rect 138818 326 139256 354
rect 138818 -960 138930 326
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 354 192106 480
rect 192404 354 192432 3130
rect 196808 3120 196860 3126
rect 193140 2990 193168 3060
rect 193968 3058 194258 3074
rect 196808 3062 196860 3068
rect 193956 3052 194258 3058
rect 194008 3046 194258 3052
rect 194416 3052 194468 3058
rect 193956 2994 194008 3000
rect 194416 2994 194468 3000
rect 193128 2984 193180 2990
rect 193128 2926 193180 2932
rect 193220 2780 193272 2786
rect 193220 2722 193272 2728
rect 193232 480 193260 2722
rect 194428 480 194456 2994
rect 195348 2922 195376 3060
rect 195612 2984 195664 2990
rect 195612 2926 195664 2932
rect 195336 2916 195388 2922
rect 195336 2858 195388 2864
rect 195624 480 195652 2926
rect 196820 480 196848 3062
rect 199488 3046 199778 3074
rect 199108 2916 199160 2922
rect 199108 2858 199160 2864
rect 198280 1352 198332 1358
rect 198280 1294 198332 1300
rect 191994 326 192432 354
rect 191994 -960 192106 326
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 354 197994 480
rect 198292 354 198320 1294
rect 199120 480 199148 2858
rect 199488 2854 199516 3046
rect 199476 2848 199528 2854
rect 199476 2790 199528 2796
rect 200316 480 200344 3198
rect 201500 3188 201552 3194
rect 206112 3182 206402 3198
rect 206940 3194 207506 3210
rect 224880 3194 225170 3210
rect 233712 3194 234002 3210
rect 206928 3188 207506 3194
rect 201500 3130 201552 3136
rect 206980 3182 207506 3188
rect 214472 3188 214524 3194
rect 206928 3130 206980 3136
rect 214472 3130 214524 3136
rect 219348 3188 219400 3194
rect 219348 3130 219400 3136
rect 220268 3188 220320 3194
rect 220268 3130 220320 3136
rect 224868 3188 225170 3194
rect 224920 3182 225170 3188
rect 229836 3188 229888 3194
rect 224868 3130 224920 3136
rect 229836 3130 229888 3136
rect 233700 3188 234002 3194
rect 233752 3182 234002 3188
rect 553150 3204 553308 3210
rect 571524 3256 571576 3262
rect 553150 3198 553360 3204
rect 553150 3182 553348 3198
rect 556462 3194 556752 3210
rect 571524 3198 571576 3204
rect 556462 3188 556764 3194
rect 556462 3182 556712 3188
rect 233700 3130 233752 3136
rect 556712 3130 556764 3136
rect 200592 3058 200882 3074
rect 200580 3052 200882 3058
rect 200632 3046 200882 3052
rect 200580 2994 200632 3000
rect 201512 480 201540 3130
rect 202880 3120 202932 3126
rect 208952 3120 209004 3126
rect 202932 3068 203090 3074
rect 202880 3062 203090 3068
rect 201972 2990 202000 3060
rect 202696 3052 202748 3058
rect 202892 3046 203090 3062
rect 202696 2994 202748 3000
rect 201960 2984 202012 2990
rect 201960 2926 202012 2932
rect 202708 480 202736 2994
rect 203892 2984 203944 2990
rect 203892 2926 203944 2932
rect 203904 480 203932 2926
rect 204180 1358 204208 3060
rect 205008 3046 205298 3074
rect 208412 3058 208610 3074
rect 213828 3120 213880 3126
rect 208952 3062 209004 3068
rect 208400 3052 208610 3058
rect 205008 2922 205036 3046
rect 208452 3046 208610 3052
rect 208400 2994 208452 3000
rect 204996 2916 205048 2922
rect 204996 2858 205048 2864
rect 206192 2916 206244 2922
rect 206192 2858 206244 2864
rect 205088 2848 205140 2854
rect 205088 2790 205140 2796
rect 204168 1352 204220 1358
rect 204168 1294 204220 1300
rect 205100 480 205128 2790
rect 206204 480 206232 2858
rect 207388 1352 207440 1358
rect 207388 1294 207440 1300
rect 207400 480 207428 1294
rect 197882 326 198320 354
rect 197882 -960 197994 326
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 354 208666 480
rect 208964 354 208992 3062
rect 209424 3046 209714 3074
rect 210528 3046 210818 3074
rect 211632 3046 211922 3074
rect 213880 3068 214130 3074
rect 213828 3062 214130 3068
rect 209424 2990 209452 3046
rect 209412 2984 209464 2990
rect 209412 2926 209464 2932
rect 209780 2984 209832 2990
rect 209780 2926 209832 2932
rect 209792 480 209820 2926
rect 210528 2854 210556 3046
rect 211632 2922 211660 3046
rect 212172 2984 212224 2990
rect 212172 2926 212224 2932
rect 211620 2916 211672 2922
rect 211620 2858 211672 2864
rect 210516 2848 210568 2854
rect 210516 2790 210568 2796
rect 210976 2848 211028 2854
rect 210976 2790 211028 2796
rect 210988 480 211016 2790
rect 212184 480 212212 2926
rect 213012 1358 213040 3060
rect 213840 3046 214130 3062
rect 213368 2916 213420 2922
rect 213368 2858 213420 2864
rect 213000 1352 213052 1358
rect 213000 1294 213052 1300
rect 213380 480 213408 2858
rect 214484 480 214512 3130
rect 215668 3120 215720 3126
rect 214944 3058 215234 3074
rect 219360 3074 219388 3130
rect 215668 3062 215720 3068
rect 214932 3052 215234 3058
rect 214984 3046 215234 3052
rect 214932 2994 214984 3000
rect 215680 480 215708 3062
rect 216048 3046 216338 3074
rect 217152 3046 217442 3074
rect 218060 3052 218112 3058
rect 216048 2854 216076 3046
rect 217152 2990 217180 3046
rect 218060 2994 218112 3000
rect 218256 3046 218546 3074
rect 219360 3046 219650 3074
rect 217140 2984 217192 2990
rect 217140 2926 217192 2932
rect 216036 2848 216088 2854
rect 216036 2790 216088 2796
rect 216864 2848 216916 2854
rect 216864 2790 216916 2796
rect 216876 480 216904 2790
rect 218072 480 218100 2994
rect 218256 2922 218284 3046
rect 218244 2916 218296 2922
rect 218244 2858 218296 2864
rect 219256 2916 219308 2922
rect 219256 2858 219308 2864
rect 219268 480 219296 2858
rect 208554 326 208992 354
rect 208554 -960 208666 326
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220280 218 220308 3130
rect 220452 3120 220504 3126
rect 221556 3120 221608 3126
rect 220504 3068 220754 3074
rect 220452 3062 220754 3068
rect 225972 3120 226024 3126
rect 221556 3062 221608 3068
rect 220464 3046 220754 3062
rect 221568 480 221596 3062
rect 221844 2854 221872 3060
rect 222672 3058 222962 3074
rect 222660 3052 222962 3058
rect 222712 3046 222962 3052
rect 223500 3046 224066 3074
rect 226024 3068 226274 3074
rect 225972 3062 226274 3068
rect 225512 3052 225564 3058
rect 222660 2994 222712 3000
rect 222752 2984 222804 2990
rect 222752 2926 222804 2932
rect 221832 2848 221884 2854
rect 221832 2790 221884 2796
rect 222764 480 222792 2926
rect 223500 2922 223528 3046
rect 225984 3046 226274 3062
rect 225512 2994 225564 3000
rect 223488 2916 223540 2922
rect 223488 2858 223540 2864
rect 223948 2848 224000 2854
rect 223948 2790 224000 2796
rect 223960 480 223988 2790
rect 220422 218 220534 480
rect 220280 190 220534 218
rect 220422 -960 220534 190
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 354 225226 480
rect 225524 354 225552 2994
rect 227364 2990 227392 3060
rect 227352 2984 227404 2990
rect 227352 2926 227404 2932
rect 227536 2984 227588 2990
rect 227536 2926 227588 2932
rect 226340 2916 226392 2922
rect 226340 2858 226392 2864
rect 226352 480 226380 2858
rect 227548 480 227576 2926
rect 228468 2854 228496 3060
rect 229296 3058 229586 3074
rect 229284 3052 229586 3058
rect 229336 3046 229586 3052
rect 229284 2994 229336 3000
rect 228456 2848 228508 2854
rect 228456 2790 228508 2796
rect 228732 2848 228784 2854
rect 228732 2790 228784 2796
rect 228744 480 228772 2790
rect 229848 480 229876 3130
rect 231032 3120 231084 3126
rect 231032 3062 231084 3068
rect 234804 3120 234856 3126
rect 530032 3120 530084 3126
rect 234856 3068 235106 3074
rect 234804 3062 235106 3068
rect 230676 2922 230704 3060
rect 230664 2916 230716 2922
rect 230664 2858 230716 2864
rect 231044 480 231072 3062
rect 231780 2990 231808 3060
rect 231768 2984 231820 2990
rect 231768 2926 231820 2932
rect 232228 2916 232280 2922
rect 232228 2858 232280 2864
rect 232240 480 232268 2858
rect 232884 2854 232912 3060
rect 233424 3052 233476 3058
rect 234816 3046 235106 3062
rect 233424 2994 233476 3000
rect 232872 2848 232924 2854
rect 232872 2790 232924 2796
rect 233436 480 233464 2994
rect 234620 2984 234672 2990
rect 234620 2926 234672 2932
rect 234632 480 234660 2926
rect 236196 2922 236224 3060
rect 237024 3058 237314 3074
rect 237012 3052 237314 3058
rect 237064 3046 237314 3052
rect 238116 3052 238168 3058
rect 237012 2994 237064 3000
rect 238116 2994 238168 3000
rect 236184 2916 236236 2922
rect 236184 2858 236236 2864
rect 237012 2916 237064 2922
rect 237012 2858 237064 2864
rect 235816 2848 235868 2854
rect 235816 2790 235868 2796
rect 235828 480 235856 2790
rect 237024 480 237052 2858
rect 238128 480 238156 2994
rect 238404 2990 238432 3060
rect 238392 2984 238444 2990
rect 238392 2926 238444 2932
rect 239312 2984 239364 2990
rect 239312 2926 239364 2932
rect 239324 480 239352 2926
rect 239508 2854 239536 3060
rect 240612 2922 240640 3060
rect 241532 3058 241730 3074
rect 241520 3052 241730 3058
rect 241572 3046 241730 3052
rect 241520 2994 241572 3000
rect 242820 2990 242848 3060
rect 242808 2984 242860 2990
rect 242808 2926 242860 2932
rect 242900 2984 242952 2990
rect 242900 2926 242952 2932
rect 240600 2916 240652 2922
rect 240600 2858 240652 2864
rect 242072 2916 242124 2922
rect 242072 2858 242124 2864
rect 239496 2848 239548 2854
rect 239496 2790 239548 2796
rect 240508 2848 240560 2854
rect 240508 2790 240560 2796
rect 240520 480 240548 2790
rect 225114 326 225552 354
rect 225114 -960 225226 326
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 354 241786 480
rect 242084 354 242112 2858
rect 242912 480 242940 2926
rect 243924 2854 243952 3060
rect 245028 2922 245056 3060
rect 246132 2990 246160 3060
rect 246120 2984 246172 2990
rect 246120 2926 246172 2932
rect 246396 2984 246448 2990
rect 246396 2926 246448 2932
rect 245016 2916 245068 2922
rect 245016 2858 245068 2864
rect 245200 2916 245252 2922
rect 245200 2858 245252 2864
rect 243912 2848 243964 2854
rect 243912 2790 243964 2796
rect 244096 2848 244148 2854
rect 244096 2790 244148 2796
rect 244108 480 244136 2790
rect 245212 480 245240 2858
rect 246408 480 246436 2926
rect 247236 2854 247264 3060
rect 248340 2922 248368 3060
rect 248788 3052 248840 3058
rect 248788 2994 248840 3000
rect 248328 2916 248380 2922
rect 248328 2858 248380 2864
rect 247224 2848 247276 2854
rect 247224 2790 247276 2796
rect 247592 2848 247644 2854
rect 247592 2790 247644 2796
rect 247604 480 247632 2790
rect 248800 480 248828 2994
rect 249444 2990 249472 3060
rect 249432 2984 249484 2990
rect 249432 2926 249484 2932
rect 249984 2916 250036 2922
rect 249984 2858 250036 2864
rect 249996 480 250024 2858
rect 250548 2854 250576 3060
rect 251376 3058 251666 3074
rect 251364 3052 251666 3058
rect 251416 3046 251666 3052
rect 251364 2994 251416 3000
rect 252756 2922 252784 3060
rect 253480 2984 253532 2990
rect 253480 2926 253532 2932
rect 252744 2916 252796 2922
rect 252744 2858 252796 2864
rect 250536 2848 250588 2854
rect 250536 2790 250588 2796
rect 252376 2848 252428 2854
rect 252376 2790 252428 2796
rect 251180 808 251232 814
rect 251180 750 251232 756
rect 251192 480 251220 750
rect 252388 480 252416 2790
rect 253492 480 253520 2926
rect 253860 814 253888 3060
rect 254676 2916 254728 2922
rect 254676 2858 254728 2864
rect 253848 808 253900 814
rect 253848 750 253900 756
rect 254688 480 254716 2858
rect 254964 2854 254992 3060
rect 256068 2990 256096 3060
rect 256056 2984 256108 2990
rect 256056 2926 256108 2932
rect 257172 2922 257200 3060
rect 257160 2916 257212 2922
rect 257160 2858 257212 2864
rect 258276 2854 258304 3060
rect 254952 2848 255004 2854
rect 254952 2790 255004 2796
rect 255872 2848 255924 2854
rect 255872 2790 255924 2796
rect 258264 2848 258316 2854
rect 258264 2790 258316 2796
rect 255884 480 255912 2790
rect 259380 1358 259408 3060
rect 257068 1352 257120 1358
rect 257068 1294 257120 1300
rect 259368 1352 259420 1358
rect 259368 1294 259420 1300
rect 259460 1352 259512 1358
rect 259460 1294 259512 1300
rect 257080 480 257108 1294
rect 258264 1284 258316 1290
rect 258264 1226 258316 1232
rect 258276 480 258304 1226
rect 259472 480 259500 1294
rect 260484 1290 260512 3060
rect 260656 2848 260708 2854
rect 260656 2790 260708 2796
rect 260472 1284 260524 1290
rect 260472 1226 260524 1232
rect 260668 480 260696 2790
rect 261588 1358 261616 3060
rect 261760 2916 261812 2922
rect 261760 2858 261812 2864
rect 261576 1352 261628 1358
rect 261576 1294 261628 1300
rect 261772 480 261800 2858
rect 262692 2854 262720 3060
rect 263796 2922 263824 3060
rect 263784 2916 263836 2922
rect 263784 2858 263836 2864
rect 262680 2848 262732 2854
rect 262680 2790 262732 2796
rect 264900 1358 264928 3060
rect 262956 1352 263008 1358
rect 262956 1294 263008 1300
rect 264888 1352 264940 1358
rect 264888 1294 264940 1300
rect 265348 1352 265400 1358
rect 265348 1294 265400 1300
rect 262968 480 262996 1294
rect 264152 1284 264204 1290
rect 264152 1226 264204 1232
rect 264164 480 264192 1226
rect 265360 480 265388 1294
rect 266004 1290 266032 3060
rect 267108 1358 267136 3060
rect 267096 1352 267148 1358
rect 267096 1294 267148 1300
rect 267740 1352 267792 1358
rect 267740 1294 267792 1300
rect 265992 1284 266044 1290
rect 265992 1226 266044 1232
rect 266544 1284 266596 1290
rect 266544 1226 266596 1232
rect 266556 480 266584 1226
rect 267752 480 267780 1294
rect 268212 1290 268240 3060
rect 269316 1358 269344 3060
rect 269304 1352 269356 1358
rect 269304 1294 269356 1300
rect 268200 1284 268252 1290
rect 268200 1226 268252 1232
rect 270040 1284 270092 1290
rect 270040 1226 270092 1232
rect 268844 1216 268896 1222
rect 268844 1158 268896 1164
rect 268856 480 268884 1158
rect 270052 480 270080 1226
rect 270420 1222 270448 3060
rect 271236 1352 271288 1358
rect 271236 1294 271288 1300
rect 270408 1216 270460 1222
rect 270408 1158 270460 1164
rect 271248 480 271276 1294
rect 271524 1290 271552 3060
rect 272628 1358 272656 3060
rect 272616 1352 272668 1358
rect 272616 1294 272668 1300
rect 273628 1352 273680 1358
rect 273628 1294 273680 1300
rect 271512 1284 271564 1290
rect 271512 1226 271564 1232
rect 272432 1284 272484 1290
rect 272432 1226 272484 1232
rect 272444 480 272472 1226
rect 273640 480 273668 1294
rect 273732 1290 273760 3060
rect 274836 1358 274864 3060
rect 275296 3046 275954 3074
rect 276124 3046 277058 3074
rect 274824 1352 274876 1358
rect 274824 1294 274876 1300
rect 273720 1284 273772 1290
rect 273720 1226 273772 1232
rect 241674 326 242112 354
rect 241674 -960 241786 326
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 354 274906 480
rect 275296 354 275324 3046
rect 276124 1578 276152 3046
rect 276032 1550 276152 1578
rect 276032 480 276060 1550
rect 278148 1358 278176 3060
rect 278792 3046 279266 3074
rect 277124 1352 277176 1358
rect 277124 1294 277176 1300
rect 278136 1352 278188 1358
rect 278136 1294 278188 1300
rect 277136 480 277164 1294
rect 274794 326 275324 354
rect 274794 -960 274906 326
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 354 278402 480
rect 278792 354 278820 3046
rect 280356 1358 280384 3060
rect 281184 3046 281474 3074
rect 281920 3046 282578 3074
rect 283392 3046 283682 3074
rect 284312 3046 284786 3074
rect 285416 3046 285890 3074
rect 279516 1352 279568 1358
rect 279516 1294 279568 1300
rect 280344 1352 280396 1358
rect 280344 1294 280396 1300
rect 279528 480 279556 1294
rect 278290 326 278820 354
rect 278290 -960 278402 326
rect 279486 -960 279598 480
rect 280682 354 280794 480
rect 281184 354 281212 3046
rect 281920 480 281948 3046
rect 280682 326 281212 354
rect 280682 -960 280794 326
rect 281878 -960 281990 480
rect 283074 354 283186 480
rect 283392 354 283420 3046
rect 284312 480 284340 3046
rect 285416 480 285444 3046
rect 283074 326 283420 354
rect 283074 -960 283186 326
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 354 286682 480
rect 286980 354 287008 3060
rect 287808 3046 288098 3074
rect 289004 3046 289202 3074
rect 290200 3046 290306 3074
rect 287808 480 287836 3046
rect 289004 480 289032 3046
rect 290200 480 290228 3046
rect 291396 480 291424 3060
rect 292592 480 292620 3060
rect 293696 480 293724 3060
rect 294814 3046 294920 3074
rect 295918 3046 296116 3074
rect 297022 3046 297312 3074
rect 294892 480 294920 3046
rect 296088 480 296116 3046
rect 297284 480 297312 3046
rect 286570 326 287008 354
rect 286570 -960 286682 326
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 3060
rect 299230 3046 299704 3074
rect 300334 3046 300808 3074
rect 301438 3046 301728 3074
rect 302542 3046 303200 3074
rect 303646 3046 303936 3074
rect 299676 480 299704 3046
rect 300780 480 300808 3046
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301700 354 301728 3046
rect 303172 480 303200 3046
rect 301934 354 302046 480
rect 301700 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 3046
rect 304736 2854 304764 3060
rect 305854 3046 306328 3074
rect 304724 2848 304776 2854
rect 304724 2790 304776 2796
rect 305552 2848 305604 2854
rect 305552 2790 305604 2796
rect 305564 480 305592 2790
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306300 354 306328 3046
rect 306944 2854 306972 3060
rect 308062 3046 308996 3074
rect 306932 2848 306984 2854
rect 306932 2790 306984 2796
rect 307944 2848 307996 2854
rect 307944 2790 307996 2796
rect 307956 480 307984 2790
rect 308968 1578 308996 3046
rect 309152 2854 309180 3060
rect 310256 2990 310284 3060
rect 310244 2984 310296 2990
rect 310244 2926 310296 2932
rect 311360 2854 311388 3060
rect 311440 2984 311492 2990
rect 311440 2926 311492 2932
rect 309140 2848 309192 2854
rect 309140 2790 309192 2796
rect 310244 2848 310296 2854
rect 310244 2790 310296 2796
rect 311348 2848 311400 2854
rect 311348 2790 311400 2796
rect 308968 1550 309088 1578
rect 309060 480 309088 1550
rect 310256 480 310284 2790
rect 311452 480 311480 2926
rect 312464 2922 312492 3060
rect 312452 2916 312504 2922
rect 312452 2858 312504 2864
rect 313568 2854 313596 3060
rect 314580 2922 314608 3060
rect 313832 2916 313884 2922
rect 313832 2858 313884 2864
rect 314568 2916 314620 2922
rect 314568 2858 314620 2864
rect 312636 2848 312688 2854
rect 312636 2790 312688 2796
rect 313556 2848 313608 2854
rect 313556 2790 313608 2796
rect 312648 480 312676 2790
rect 313844 480 313872 2858
rect 315776 2854 315804 3060
rect 316880 2922 316908 3060
rect 316224 2916 316276 2922
rect 316224 2858 316276 2864
rect 316868 2916 316920 2922
rect 316868 2858 316920 2864
rect 315028 2848 315080 2854
rect 315028 2790 315080 2796
rect 315764 2848 315816 2854
rect 315764 2790 315816 2796
rect 315040 480 315068 2790
rect 316236 480 316264 2858
rect 317984 2854 318012 3060
rect 319088 2922 319116 3060
rect 318524 2916 318576 2922
rect 318524 2858 318576 2864
rect 319076 2916 319128 2922
rect 319076 2858 319128 2864
rect 317328 2848 317380 2854
rect 317328 2790 317380 2796
rect 317972 2848 318024 2854
rect 317972 2790 318024 2796
rect 317340 480 317368 2790
rect 318536 480 318564 2858
rect 320100 2854 320128 3060
rect 321296 2922 321324 3060
rect 320916 2916 320968 2922
rect 320916 2858 320968 2864
rect 321284 2916 321336 2922
rect 321284 2858 321336 2864
rect 319720 2848 319772 2854
rect 319720 2790 319772 2796
rect 320088 2848 320140 2854
rect 320088 2790 320140 2796
rect 319732 480 319760 2790
rect 320928 480 320956 2858
rect 322400 2854 322428 3060
rect 323504 2922 323532 3060
rect 323308 2916 323360 2922
rect 323308 2858 323360 2864
rect 323492 2916 323544 2922
rect 323492 2858 323544 2864
rect 322112 2848 322164 2854
rect 322112 2790 322164 2796
rect 322388 2848 322440 2854
rect 322388 2790 322440 2796
rect 322124 480 322152 2790
rect 323320 480 323348 2858
rect 324608 2854 324636 3060
rect 325712 2990 325740 3060
rect 326830 3046 327028 3074
rect 325700 2984 325752 2990
rect 325700 2926 325752 2932
rect 325608 2916 325660 2922
rect 325608 2858 325660 2864
rect 324412 2848 324464 2854
rect 324412 2790 324464 2796
rect 324596 2848 324648 2854
rect 324596 2790 324648 2796
rect 324424 480 324452 2790
rect 325620 480 325648 2858
rect 327000 2854 327028 3046
rect 327920 2922 327948 3060
rect 329024 2990 329052 3060
rect 328000 2984 328052 2990
rect 328000 2926 328052 2932
rect 329012 2984 329064 2990
rect 329012 2926 329064 2932
rect 327908 2916 327960 2922
rect 327908 2858 327960 2864
rect 326804 2848 326856 2854
rect 326804 2790 326856 2796
rect 326988 2848 327040 2854
rect 326988 2790 327040 2796
rect 326816 480 326844 2790
rect 328012 480 328040 2926
rect 330128 2854 330156 3060
rect 331246 3058 331352 3074
rect 331246 3052 331364 3058
rect 331246 3046 331312 3052
rect 331312 2994 331364 3000
rect 332336 2990 332364 3060
rect 331588 2984 331640 2990
rect 331588 2926 331640 2932
rect 332324 2984 332376 2990
rect 332324 2926 332376 2932
rect 330392 2916 330444 2922
rect 330392 2858 330444 2864
rect 329196 2848 329248 2854
rect 329196 2790 329248 2796
rect 330116 2848 330168 2854
rect 330116 2790 330168 2796
rect 329208 480 329236 2790
rect 330404 480 330432 2858
rect 331600 480 331628 2926
rect 333440 2922 333468 3060
rect 334558 3058 334848 3074
rect 333888 3052 333940 3058
rect 334558 3052 334860 3058
rect 334558 3046 334808 3052
rect 333888 2994 333940 3000
rect 334808 2994 334860 3000
rect 333428 2916 333480 2922
rect 333428 2858 333480 2864
rect 332692 2848 332744 2854
rect 332692 2790 332744 2796
rect 332704 480 332732 2790
rect 333900 480 333928 2994
rect 335084 2984 335136 2990
rect 335084 2926 335136 2932
rect 335096 480 335124 2926
rect 335648 2854 335676 3060
rect 336280 2916 336332 2922
rect 336280 2858 336332 2864
rect 335636 2848 335688 2854
rect 335636 2790 335688 2796
rect 336292 480 336320 2858
rect 336660 1358 336688 3060
rect 337476 3052 337528 3058
rect 337476 2994 337528 3000
rect 336648 1352 336700 1358
rect 336648 1294 336700 1300
rect 337488 480 337516 2994
rect 337856 882 337884 3060
rect 338960 2854 338988 3060
rect 340064 2922 340092 3060
rect 341168 2990 341196 3060
rect 341156 2984 341208 2990
rect 341156 2926 341208 2932
rect 340052 2916 340104 2922
rect 340052 2858 340104 2864
rect 338672 2848 338724 2854
rect 338672 2790 338724 2796
rect 338948 2848 339000 2854
rect 338948 2790 339000 2796
rect 342076 2848 342128 2854
rect 342076 2790 342128 2796
rect 337844 876 337896 882
rect 337844 818 337896 824
rect 338684 480 338712 2790
rect 339868 1352 339920 1358
rect 339868 1294 339920 1300
rect 339880 480 339908 1294
rect 342088 1170 342116 2790
rect 342180 1358 342208 3060
rect 342996 2916 343048 2922
rect 342996 2858 343048 2864
rect 342168 1352 342220 1358
rect 342168 1294 342220 1300
rect 342088 1142 342208 1170
rect 340972 876 341024 882
rect 340972 818 341024 824
rect 340984 480 341012 818
rect 342180 480 342208 1142
rect 306718 354 306830 480
rect 306300 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343008 354 343036 2858
rect 343376 1290 343404 3060
rect 344494 3046 344784 3074
rect 344560 2984 344612 2990
rect 344560 2926 344612 2932
rect 343364 1284 343416 1290
rect 343364 1226 343416 1232
rect 344572 480 344600 2926
rect 343334 354 343446 480
rect 343008 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 344756 134 344784 3046
rect 345584 1018 345612 3060
rect 346688 2854 346716 3060
rect 346676 2848 346728 2854
rect 346676 2790 346728 2796
rect 345756 1352 345808 1358
rect 345756 1294 345808 1300
rect 345572 1012 345624 1018
rect 345572 954 345624 960
rect 345768 480 345796 1294
rect 346952 1284 347004 1290
rect 346952 1226 347004 1232
rect 346964 480 346992 1226
rect 347700 882 347728 3060
rect 348896 1358 348924 3060
rect 348884 1352 348936 1358
rect 348884 1294 348936 1300
rect 350000 1290 350028 3060
rect 350448 2848 350500 2854
rect 350448 2790 350500 2796
rect 349988 1284 350040 1290
rect 349988 1226 350040 1232
rect 349252 1012 349304 1018
rect 349252 954 349304 960
rect 347688 876 347740 882
rect 347688 818 347740 824
rect 349264 480 349292 954
rect 350460 480 350488 2790
rect 351104 1018 351132 3060
rect 352208 1154 352236 3060
rect 353220 2854 353248 3060
rect 353208 2848 353260 2854
rect 353208 2790 353260 2796
rect 352840 1352 352892 1358
rect 352840 1294 352892 1300
rect 352196 1148 352248 1154
rect 352196 1090 352248 1096
rect 351092 1012 351144 1018
rect 351092 954 351144 960
rect 351644 876 351696 882
rect 351644 818 351696 824
rect 351656 480 351684 818
rect 352852 480 352880 1294
rect 354036 1284 354088 1290
rect 354036 1226 354088 1232
rect 354048 480 354076 1226
rect 344744 128 344796 134
rect 344744 70 344796 76
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 82 348138 480
rect 348240 128 348292 134
rect 348026 76 348240 82
rect 348026 70 348292 76
rect 348026 54 348280 70
rect 348026 -960 348138 54
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 354416 134 354444 3060
rect 355520 1086 355548 3060
rect 356624 1358 356652 3060
rect 357532 2848 357584 2854
rect 357532 2790 357584 2796
rect 356612 1352 356664 1358
rect 356612 1294 356664 1300
rect 356336 1148 356388 1154
rect 356336 1090 356388 1096
rect 355508 1080 355560 1086
rect 355508 1022 355560 1028
rect 355232 1012 355284 1018
rect 355232 954 355284 960
rect 355244 480 355272 954
rect 356348 480 356376 1090
rect 357544 480 357572 2790
rect 357728 1290 357756 3060
rect 357716 1284 357768 1290
rect 357716 1226 357768 1232
rect 358740 950 358768 3060
rect 359936 1222 359964 3060
rect 359924 1216 359976 1222
rect 359924 1158 359976 1164
rect 361040 1154 361068 3060
rect 361120 1352 361172 1358
rect 361120 1294 361172 1300
rect 361028 1148 361080 1154
rect 361028 1090 361080 1096
rect 359924 1080 359976 1086
rect 359924 1022 359976 1028
rect 358728 944 358780 950
rect 358728 886 358780 892
rect 359936 480 359964 1022
rect 361132 480 361160 1294
rect 362144 1018 362172 3060
rect 362316 1284 362368 1290
rect 362316 1226 362368 1232
rect 362132 1012 362184 1018
rect 362132 954 362184 960
rect 362328 480 362356 1226
rect 354404 128 354456 134
rect 354404 70 354456 76
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 82 358810 480
rect 358912 128 358964 134
rect 358698 76 358912 82
rect 358698 70 358964 76
rect 358698 54 358952 70
rect 358698 -960 358810 54
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363248 66 363276 3060
rect 364260 1358 364288 3060
rect 364248 1352 364300 1358
rect 364248 1294 364300 1300
rect 365456 1290 365484 3060
rect 365444 1284 365496 1290
rect 365444 1226 365496 1232
rect 364616 1216 364668 1222
rect 364616 1158 364668 1164
rect 363512 944 363564 950
rect 363512 886 363564 892
rect 363524 480 363552 886
rect 364628 480 364656 1158
rect 366560 1154 366588 3060
rect 365444 1148 365496 1154
rect 365444 1090 365496 1096
rect 366548 1148 366600 1154
rect 366548 1090 366600 1096
rect 363236 60 363288 66
rect 363236 2 363288 8
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365456 354 365484 1090
rect 367664 1086 367692 3060
rect 368768 1222 368796 3060
rect 369780 1358 369808 3060
rect 369400 1352 369452 1358
rect 369400 1294 369452 1300
rect 369768 1352 369820 1358
rect 369768 1294 369820 1300
rect 368756 1216 368808 1222
rect 368756 1158 368808 1164
rect 367652 1080 367704 1086
rect 367652 1022 367704 1028
rect 367008 1012 367060 1018
rect 367008 954 367060 960
rect 367020 480 367048 954
rect 369412 480 369440 1294
rect 370976 1290 371004 3060
rect 372094 3046 372384 3074
rect 372356 2854 372384 3046
rect 372344 2848 372396 2854
rect 372344 2790 372396 2796
rect 370228 1284 370280 1290
rect 370228 1226 370280 1232
rect 370964 1284 371016 1290
rect 370964 1226 371016 1232
rect 365782 354 365894 480
rect 365456 326 365894 354
rect 365782 -960 365894 326
rect 366978 -960 367090 480
rect 368174 82 368286 480
rect 367848 66 368286 82
rect 367836 60 368286 66
rect 367888 54 368286 60
rect 367836 2 367888 8
rect 368174 -960 368286 54
rect 369370 -960 369482 480
rect 370240 354 370268 1226
rect 371332 1148 371384 1154
rect 371332 1090 371384 1096
rect 370566 354 370678 480
rect 370240 326 370678 354
rect 371344 354 371372 1090
rect 372896 1080 372948 1086
rect 372896 1022 372948 1028
rect 372908 480 372936 1022
rect 373184 1018 373212 3060
rect 374288 1222 374316 3060
rect 375208 3046 375314 3074
rect 373908 1216 373960 1222
rect 373908 1158 373960 1164
rect 374276 1216 374328 1222
rect 374276 1158 374328 1164
rect 373172 1012 373224 1018
rect 373172 954 373224 960
rect 371670 354 371782 480
rect 371344 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 373920 354 373948 1158
rect 375208 1154 375236 3046
rect 376496 1358 376524 3060
rect 375288 1352 375340 1358
rect 375288 1294 375340 1300
rect 376484 1352 376536 1358
rect 376484 1294 376536 1300
rect 375196 1148 375248 1154
rect 375196 1090 375248 1096
rect 375300 480 375328 1294
rect 376116 1284 376168 1290
rect 376116 1226 376168 1232
rect 374062 354 374174 480
rect 373920 326 374174 354
rect 374062 -960 374174 326
rect 375258 -960 375370 480
rect 376128 354 376156 1226
rect 377600 1086 377628 3060
rect 377680 2848 377732 2854
rect 377680 2790 377732 2796
rect 377588 1080 377640 1086
rect 377588 1022 377640 1028
rect 377692 480 377720 2790
rect 378704 1290 378732 3060
rect 378692 1284 378744 1290
rect 378692 1226 378744 1232
rect 379808 1222 379836 3060
rect 379612 1216 379664 1222
rect 379612 1158 379664 1164
rect 379796 1216 379848 1222
rect 379796 1158 379848 1164
rect 378508 1012 378560 1018
rect 378508 954 378560 960
rect 376454 354 376566 480
rect 376128 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378520 354 378548 954
rect 378846 354 378958 480
rect 378520 326 378958 354
rect 379624 354 379652 1158
rect 379950 354 380062 480
rect 379624 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 380820 202 380848 3060
rect 381176 1148 381228 1154
rect 381176 1090 381228 1096
rect 381188 480 381216 1090
rect 380808 196 380860 202
rect 380808 138 380860 144
rect 381146 -960 381258 480
rect 382016 338 382044 3060
rect 382372 1352 382424 1358
rect 382372 1294 382424 1300
rect 382384 480 382412 1294
rect 382004 332 382056 338
rect 382004 274 382056 280
rect 382342 -960 382454 480
rect 383120 134 383148 3060
rect 384224 1358 384252 3060
rect 384212 1352 384264 1358
rect 384212 1294 384264 1300
rect 384396 1284 384448 1290
rect 384396 1226 384448 1232
rect 383568 1080 383620 1086
rect 383568 1022 383620 1028
rect 383580 480 383608 1022
rect 383108 128 383160 134
rect 383108 70 383160 76
rect 383538 -960 383650 480
rect 384408 354 384436 1226
rect 385328 1154 385356 3060
rect 385960 1216 386012 1222
rect 385960 1158 386012 1164
rect 385316 1148 385368 1154
rect 385316 1090 385368 1096
rect 385972 480 386000 1158
rect 386340 746 386368 3060
rect 387536 1290 387564 3060
rect 387524 1284 387576 1290
rect 387524 1226 387576 1232
rect 386328 740 386380 746
rect 386328 682 386380 688
rect 388640 610 388668 3060
rect 388628 604 388680 610
rect 388628 546 388680 552
rect 384734 354 384846 480
rect 384408 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 387126 218 387238 480
rect 388230 354 388342 480
rect 387904 338 388342 354
rect 387892 332 388342 338
rect 387944 326 388342 332
rect 387892 274 387944 280
rect 386800 202 387238 218
rect 386788 196 387238 202
rect 386840 190 387238 196
rect 386788 138 386840 144
rect 387126 -960 387238 190
rect 388230 -960 388342 326
rect 389426 82 389538 480
rect 389744 338 389772 3060
rect 390652 1352 390704 1358
rect 390652 1294 390704 1300
rect 390664 480 390692 1294
rect 389732 332 389784 338
rect 389732 274 389784 280
rect 389640 128 389692 134
rect 389426 76 389640 82
rect 389426 70 389692 76
rect 389426 54 389680 70
rect 389426 -960 389538 54
rect 390622 -960 390734 480
rect 390848 270 390876 3060
rect 391676 3046 391874 3074
rect 390836 264 390888 270
rect 390836 206 390888 212
rect 391676 202 391704 3046
rect 391848 1148 391900 1154
rect 391848 1090 391900 1096
rect 391860 480 391888 1090
rect 392676 740 392728 746
rect 392676 682 392728 688
rect 391664 196 391716 202
rect 391664 138 391716 144
rect 391818 -960 391930 480
rect 392688 354 392716 682
rect 393056 678 393084 3060
rect 394160 1358 394188 3060
rect 394148 1352 394200 1358
rect 394148 1294 394200 1300
rect 394240 1284 394292 1290
rect 394240 1226 394292 1232
rect 393044 672 393096 678
rect 393044 614 393096 620
rect 394252 480 394280 1226
rect 395264 1222 395292 3060
rect 396368 1290 396396 3060
rect 396356 1284 396408 1290
rect 396356 1226 396408 1232
rect 395252 1216 395304 1222
rect 395252 1158 395304 1164
rect 397380 1154 397408 3060
rect 397368 1148 397420 1154
rect 397368 1090 397420 1096
rect 395344 604 395396 610
rect 395344 546 395396 552
rect 395356 480 395384 546
rect 393014 354 393126 480
rect 392688 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 354 396622 480
rect 396184 338 396622 354
rect 396172 332 396622 338
rect 396224 326 396622 332
rect 396172 274 396224 280
rect 396510 -960 396622 326
rect 397706 218 397818 480
rect 397920 264 397972 270
rect 397706 212 397920 218
rect 397706 206 397972 212
rect 397706 190 397960 206
rect 397706 -960 397818 190
rect 398576 134 398604 3060
rect 398902 218 399014 480
rect 398760 202 399014 218
rect 398748 196 399014 202
rect 398800 190 399014 196
rect 398748 138 398800 144
rect 398564 128 398616 134
rect 398564 70 398616 76
rect 398902 -960 399014 190
rect 399680 66 399708 3060
rect 400784 678 400812 3060
rect 401324 1352 401376 1358
rect 401324 1294 401376 1300
rect 400128 672 400180 678
rect 400128 614 400180 620
rect 400772 672 400824 678
rect 400772 614 400824 620
rect 400140 480 400168 614
rect 401336 480 401364 1294
rect 399668 60 399720 66
rect 399668 2 399720 8
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 401888 474 401916 3060
rect 402520 1216 402572 1222
rect 402520 1158 402572 1164
rect 402532 480 402560 1158
rect 401876 468 401928 474
rect 401876 410 401928 416
rect 402490 -960 402602 480
rect 402900 270 402928 3060
rect 404096 1290 404124 3060
rect 403624 1284 403676 1290
rect 403624 1226 403676 1232
rect 404084 1284 404136 1290
rect 404084 1226 404136 1232
rect 403636 480 403664 1226
rect 404820 1148 404872 1154
rect 404820 1090 404872 1096
rect 404832 480 404860 1090
rect 402888 264 402940 270
rect 402888 206 402940 212
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405200 202 405228 3060
rect 406304 1358 406332 3060
rect 406292 1352 406344 1358
rect 406292 1294 406344 1300
rect 405188 196 405240 202
rect 405188 138 405240 144
rect 405986 82 406098 480
rect 406200 128 406252 134
rect 405986 76 406200 82
rect 407182 82 407294 480
rect 407408 406 407436 3060
rect 408420 746 408448 3060
rect 408408 740 408460 746
rect 408408 682 408460 688
rect 409616 678 409644 3060
rect 409604 672 409656 678
rect 409604 614 409656 620
rect 408408 604 408460 610
rect 408408 546 408460 552
rect 408420 480 408448 546
rect 407396 400 407448 406
rect 407396 342 407448 348
rect 405986 70 406252 76
rect 405986 54 406240 70
rect 407040 66 407294 82
rect 407028 60 407294 66
rect 405986 -960 406098 54
rect 407080 54 407294 60
rect 407028 2 407080 8
rect 407182 -960 407294 54
rect 408378 -960 408490 480
rect 409236 468 409288 474
rect 409236 410 409288 416
rect 409248 354 409276 410
rect 409574 354 409686 480
rect 409248 326 409686 354
rect 409574 -960 409686 326
rect 410628 66 410656 3060
rect 411838 3046 412128 3074
rect 411904 1284 411956 1290
rect 411904 1226 411956 1232
rect 411916 480 411944 1226
rect 410770 218 410882 480
rect 410984 264 411036 270
rect 410770 212 410984 218
rect 410770 206 411036 212
rect 410770 190 411024 206
rect 410616 60 410668 66
rect 410616 2 410668 8
rect 410770 -960 410882 190
rect 411874 -960 411986 480
rect 412100 134 412128 3046
rect 412928 1154 412956 3060
rect 412916 1148 412968 1154
rect 412916 1090 412968 1096
rect 413070 218 413182 480
rect 413940 338 413968 3060
rect 414296 1352 414348 1358
rect 414296 1294 414348 1300
rect 414308 480 414336 1294
rect 413928 332 413980 338
rect 413928 274 413980 280
rect 412836 202 413182 218
rect 412824 196 413182 202
rect 412876 190 413182 196
rect 412824 138 412876 144
rect 412088 128 412140 134
rect 412088 70 412140 76
rect 413070 -960 413182 190
rect 414266 -960 414378 480
rect 415136 270 415164 3060
rect 416240 1018 416268 3060
rect 416228 1012 416280 1018
rect 416228 954 416280 960
rect 416688 740 416740 746
rect 416688 682 416740 688
rect 416700 480 416728 682
rect 415308 400 415360 406
rect 415462 354 415574 480
rect 415360 348 415574 354
rect 415308 342 415574 348
rect 415320 326 415574 342
rect 415124 264 415176 270
rect 415124 206 415176 212
rect 415462 -960 415574 326
rect 416658 -960 416770 480
rect 417344 406 417372 3060
rect 418448 678 418476 3060
rect 417884 672 417936 678
rect 417884 614 417936 620
rect 418436 672 418488 678
rect 418436 614 418488 620
rect 417896 480 417924 614
rect 417332 400 417384 406
rect 417332 342 417384 348
rect 417854 -960 417966 480
rect 418958 82 419070 480
rect 419460 202 419488 3060
rect 420656 542 420684 3060
rect 421380 1148 421432 1154
rect 421380 1090 421432 1096
rect 420644 536 420696 542
rect 419448 196 419500 202
rect 419448 138 419500 144
rect 418632 66 419070 82
rect 418620 60 419070 66
rect 418672 54 419070 60
rect 418620 2 418672 8
rect 418958 -960 419070 54
rect 420154 82 420266 480
rect 420644 478 420696 484
rect 421392 480 421420 1090
rect 420368 128 420420 134
rect 420154 76 420368 82
rect 420154 70 420420 76
rect 420154 54 420408 70
rect 420154 -960 420266 54
rect 421350 -960 421462 480
rect 421760 66 421788 3060
rect 422546 354 422658 480
rect 422546 338 422800 354
rect 422546 332 422812 338
rect 422546 326 422760 332
rect 421748 60 421800 66
rect 421748 2 421800 8
rect 422546 -960 422658 326
rect 422760 274 422812 280
rect 422864 134 422892 3060
rect 423968 746 423996 3060
rect 424796 3046 424994 3074
rect 423956 740 424008 746
rect 423956 682 424008 688
rect 423588 264 423640 270
rect 423742 218 423854 480
rect 424796 474 424824 3046
rect 424968 1012 425020 1018
rect 424968 954 425020 960
rect 424980 480 425008 954
rect 426176 610 426204 3060
rect 427294 3046 427584 3074
rect 428398 3046 428688 3074
rect 427268 672 427320 678
rect 427268 614 427320 620
rect 426164 604 426216 610
rect 426164 546 426216 552
rect 427280 480 427308 614
rect 424784 468 424836 474
rect 424784 410 424836 416
rect 423640 212 423854 218
rect 423588 206 423854 212
rect 423600 190 423854 206
rect 422852 128 422904 134
rect 422852 70 422904 76
rect 423742 -960 423854 190
rect 424938 -960 425050 480
rect 425796 400 425848 406
rect 426134 354 426246 480
rect 425848 348 426246 354
rect 425796 342 426246 348
rect 425808 326 426246 342
rect 426134 -960 426246 326
rect 427238 -960 427350 480
rect 427556 338 427584 3046
rect 427544 332 427596 338
rect 427544 274 427596 280
rect 428434 218 428546 480
rect 428660 406 428688 3046
rect 429488 542 429516 3060
rect 430500 1290 430528 3060
rect 430488 1284 430540 1290
rect 430488 1226 430540 1232
rect 429292 536 429344 542
rect 429292 478 429344 484
rect 429476 536 429528 542
rect 429476 478 429528 484
rect 428648 400 428700 406
rect 428648 342 428700 348
rect 429304 354 429332 478
rect 429630 354 429742 480
rect 429304 326 429742 354
rect 428434 202 428688 218
rect 428434 196 428700 202
rect 428434 190 428648 196
rect 428434 -960 428546 190
rect 428648 138 428700 144
rect 429630 -960 429742 326
rect 430826 82 430938 480
rect 431696 202 431724 3060
rect 431684 196 431736 202
rect 431684 138 431736 144
rect 431868 128 431920 134
rect 430826 66 431080 82
rect 432022 82 432134 480
rect 432800 270 432828 3060
rect 433248 740 433300 746
rect 433248 682 433300 688
rect 433260 480 433288 682
rect 432788 264 432840 270
rect 432788 206 432840 212
rect 431920 76 432134 82
rect 431868 70 432134 76
rect 430826 60 431092 66
rect 430826 54 431040 60
rect 430826 -960 430938 54
rect 431880 54 432134 70
rect 431040 2 431092 8
rect 432022 -960 432134 54
rect 433218 -960 433330 480
rect 433904 134 433932 3060
rect 434076 468 434128 474
rect 434076 410 434128 416
rect 434088 354 434116 410
rect 434414 354 434526 480
rect 435008 474 435036 3060
rect 436020 1358 436048 3060
rect 436008 1352 436060 1358
rect 436008 1294 436060 1300
rect 437216 1154 437244 3060
rect 437204 1148 437256 1154
rect 437204 1090 437256 1096
rect 438320 814 438348 3060
rect 438308 808 438360 814
rect 438308 750 438360 756
rect 435548 604 435600 610
rect 435548 546 435600 552
rect 439136 604 439188 610
rect 439136 546 439188 552
rect 435560 480 435588 546
rect 439148 480 439176 546
rect 434996 468 435048 474
rect 434996 410 435048 416
rect 434088 326 434526 354
rect 433892 128 433944 134
rect 433892 70 433944 76
rect 434414 -960 434526 326
rect 435518 -960 435630 480
rect 436714 354 436826 480
rect 437572 400 437624 406
rect 436714 338 436968 354
rect 437910 354 438022 480
rect 437624 348 438022 354
rect 437572 342 438022 348
rect 436714 332 436980 338
rect 436714 326 436928 332
rect 436714 -960 436826 326
rect 437584 326 438022 342
rect 436928 274 436980 280
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 439424 66 439452 3060
rect 439964 1284 440016 1290
rect 439964 1226 440016 1232
rect 439976 354 440004 1226
rect 440302 354 440414 480
rect 439976 326 440414 354
rect 440528 338 440556 3060
rect 441540 882 441568 3060
rect 441528 876 441580 882
rect 441528 818 441580 824
rect 442736 678 442764 3060
rect 443840 1222 443868 3060
rect 443828 1216 443880 1222
rect 443828 1158 443880 1164
rect 444944 950 444972 3060
rect 445852 1352 445904 1358
rect 445852 1294 445904 1300
rect 444932 944 444984 950
rect 444932 886 444984 892
rect 442724 672 442776 678
rect 441356 598 441568 626
rect 442724 614 442776 620
rect 441356 354 441384 598
rect 441540 480 441568 598
rect 439412 60 439464 66
rect 439412 2 439464 8
rect 440302 -960 440414 326
rect 440516 332 440568 338
rect 440516 274 440568 280
rect 441264 326 441384 354
rect 441264 202 441292 326
rect 441252 196 441304 202
rect 441252 138 441304 144
rect 441498 -960 441610 480
rect 442602 218 442714 480
rect 442816 264 442868 270
rect 442602 212 442816 218
rect 442602 206 442868 212
rect 442602 190 442856 206
rect 442602 -960 442714 190
rect 443460 128 443512 134
rect 443798 82 443910 480
rect 443512 76 443910 82
rect 443460 70 443910 76
rect 443472 54 443910 70
rect 443798 -960 443910 54
rect 444994 354 445106 480
rect 445208 468 445260 474
rect 445208 410 445260 416
rect 445220 354 445248 410
rect 444994 326 445248 354
rect 445864 354 445892 1294
rect 446048 746 446076 3060
rect 447060 1290 447088 3060
rect 447048 1284 447100 1290
rect 447048 1226 447100 1232
rect 447416 1148 447468 1154
rect 447416 1090 447468 1096
rect 446036 740 446088 746
rect 446036 682 446088 688
rect 447428 480 447456 1090
rect 448256 1018 448284 3060
rect 448244 1012 448296 1018
rect 448244 954 448296 960
rect 449360 814 449388 3060
rect 450464 1358 450492 3060
rect 450452 1352 450504 1358
rect 450452 1294 450504 1300
rect 451568 1086 451596 3060
rect 451556 1080 451608 1086
rect 451556 1022 451608 1028
rect 451740 876 451792 882
rect 451740 818 451792 824
rect 448244 808 448296 814
rect 448244 750 448296 756
rect 449348 808 449400 814
rect 449348 750 449400 756
rect 446190 354 446302 480
rect 445864 326 446302 354
rect 444994 -960 445106 326
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448256 354 448284 750
rect 448582 354 448694 480
rect 448256 326 448694 354
rect 448582 -960 448694 326
rect 449778 82 449890 480
rect 450882 354 450994 480
rect 451752 354 451780 818
rect 452078 354 452190 480
rect 450882 338 451136 354
rect 450882 332 451148 338
rect 450882 326 451096 332
rect 449778 66 450032 82
rect 449778 60 450044 66
rect 449778 54 449992 60
rect 449778 -960 449890 54
rect 449992 2 450044 8
rect 450882 -960 450994 326
rect 451752 326 452190 354
rect 451096 274 451148 280
rect 452078 -960 452190 326
rect 452580 66 452608 3060
rect 453304 672 453356 678
rect 453304 614 453356 620
rect 453316 480 453344 614
rect 452568 60 452620 66
rect 452568 2 452620 8
rect 453274 -960 453386 480
rect 453776 202 453804 3060
rect 454132 1216 454184 1222
rect 454132 1158 454184 1164
rect 454144 354 454172 1158
rect 454880 882 454908 3060
rect 455984 950 456012 3060
rect 456432 1284 456484 1290
rect 456432 1226 456484 1232
rect 455696 944 455748 950
rect 455696 886 455748 892
rect 455972 944 456024 950
rect 455972 886 456024 892
rect 454868 876 454920 882
rect 454868 818 454920 824
rect 455708 480 455736 886
rect 454470 354 454582 480
rect 454144 326 454582 354
rect 453764 196 453816 202
rect 453764 138 453816 144
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456444 270 456472 1226
rect 457088 1222 457116 3060
rect 457916 3046 458114 3074
rect 459310 3046 459508 3074
rect 460414 3046 460612 3074
rect 461518 3046 461808 3074
rect 457076 1216 457128 1222
rect 457076 1158 457128 1164
rect 456524 740 456576 746
rect 456524 682 456576 688
rect 456536 354 456564 682
rect 456862 354 456974 480
rect 457916 474 457944 3046
rect 459192 1012 459244 1018
rect 459192 954 459244 960
rect 459204 480 459232 954
rect 457904 468 457956 474
rect 457904 410 457956 416
rect 456536 326 456974 354
rect 456432 264 456484 270
rect 456432 206 456484 212
rect 456862 -960 456974 326
rect 458058 218 458170 480
rect 458272 264 458324 270
rect 458058 212 458272 218
rect 458058 206 458324 212
rect 458058 190 458312 206
rect 458058 -960 458170 190
rect 459162 -960 459274 480
rect 459480 406 459508 3046
rect 460020 808 460072 814
rect 460020 750 460072 756
rect 459468 400 459520 406
rect 459468 342 459520 348
rect 460032 354 460060 750
rect 460358 354 460470 480
rect 460032 326 460470 354
rect 460358 -960 460470 326
rect 460584 270 460612 3046
rect 461584 1352 461636 1358
rect 461584 1294 461636 1300
rect 461596 480 461624 1294
rect 461780 542 461808 3046
rect 462608 1358 462636 3060
rect 462596 1352 462648 1358
rect 462596 1294 462648 1300
rect 462412 1080 462464 1086
rect 462412 1022 462464 1028
rect 461768 536 461820 542
rect 460572 264 460624 270
rect 460572 206 460624 212
rect 461554 -960 461666 480
rect 461768 478 461820 484
rect 462424 354 462452 1022
rect 462750 354 462862 480
rect 462424 326 462862 354
rect 462750 -960 462862 326
rect 463620 134 463648 3060
rect 464816 610 464844 3060
rect 464804 604 464856 610
rect 464804 546 464856 552
rect 463608 128 463660 134
rect 463608 70 463660 76
rect 463946 82 464058 480
rect 465142 218 465254 480
rect 465000 202 465254 218
rect 464988 196 465254 202
rect 465040 190 465254 196
rect 464988 138 465040 144
rect 463946 66 464200 82
rect 463946 60 464212 66
rect 463946 54 464160 60
rect 463946 -960 464058 54
rect 464160 2 464212 8
rect 465142 -960 465254 190
rect 465828 66 465856 3060
rect 465908 876 465960 882
rect 465908 818 465960 824
rect 465920 354 465948 818
rect 466246 354 466358 480
rect 465920 326 466358 354
rect 467024 338 467052 3060
rect 467472 944 467524 950
rect 467472 886 467524 892
rect 467484 480 467512 886
rect 468128 678 468156 3060
rect 469140 1222 469168 3060
rect 468300 1216 468352 1222
rect 468300 1158 468352 1164
rect 469128 1216 469180 1222
rect 469128 1158 469180 1164
rect 468116 672 468168 678
rect 468116 614 468168 620
rect 465816 60 465868 66
rect 465816 2 465868 8
rect 466246 -960 466358 326
rect 467012 332 467064 338
rect 467012 274 467064 280
rect 467442 -960 467554 480
rect 468312 354 468340 1158
rect 468638 354 468750 480
rect 468312 326 468750 354
rect 468638 -960 468750 326
rect 469834 354 469946 480
rect 470336 474 470364 3060
rect 470048 468 470100 474
rect 470048 410 470100 416
rect 470324 468 470376 474
rect 470324 410 470376 416
rect 470060 354 470088 410
rect 469834 326 470088 354
rect 470784 400 470836 406
rect 471030 354 471142 480
rect 470836 348 471142 354
rect 470784 342 471142 348
rect 470796 326 471142 342
rect 469834 -960 469946 326
rect 471030 -960 471142 326
rect 471440 202 471468 3060
rect 472226 218 472338 480
rect 472544 406 472572 3060
rect 473452 604 473504 610
rect 473452 546 473504 552
rect 473464 480 473492 546
rect 473648 542 473676 3060
rect 474188 1352 474240 1358
rect 474188 1294 474240 1300
rect 473636 536 473688 542
rect 472532 400 472584 406
rect 472532 342 472584 348
rect 472440 264 472492 270
rect 472226 212 472440 218
rect 472226 206 472492 212
rect 471428 196 471480 202
rect 471428 138 471480 144
rect 472226 190 472480 206
rect 472226 -960 472338 190
rect 473422 -960 473534 480
rect 473636 478 473688 484
rect 474200 354 474228 1294
rect 474660 1290 474688 3060
rect 475856 1358 475884 3060
rect 476974 3046 477264 3074
rect 478078 3046 478368 3074
rect 479182 3046 479564 3074
rect 475844 1352 475896 1358
rect 475844 1294 475896 1300
rect 474648 1284 474700 1290
rect 474648 1226 474700 1232
rect 476948 672 477000 678
rect 476948 614 477000 620
rect 476960 480 476988 614
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 82 475834 480
rect 475936 128 475988 134
rect 475722 76 475936 82
rect 475722 70 475988 76
rect 475722 54 475976 70
rect 475722 -960 475834 54
rect 476918 -960 477030 480
rect 477236 134 477264 3046
rect 477224 128 477276 134
rect 477224 70 477276 76
rect 478114 82 478226 480
rect 478340 270 478368 3046
rect 479310 354 479422 480
rect 478984 338 479422 354
rect 479536 338 479564 3046
rect 480180 950 480208 3060
rect 481390 3046 481588 3074
rect 529966 3068 530032 3074
rect 546684 3120 546736 3126
rect 529966 3062 530084 3068
rect 481364 1216 481416 1222
rect 481364 1158 481416 1164
rect 480168 944 480220 950
rect 480168 886 480220 892
rect 480536 740 480588 746
rect 480536 682 480588 688
rect 480548 480 480576 682
rect 478972 332 479422 338
rect 479024 326 479422 332
rect 478972 274 479024 280
rect 478328 264 478380 270
rect 478328 206 478380 212
rect 478114 66 478368 82
rect 478114 60 478380 66
rect 478114 54 478328 60
rect 478114 -960 478226 54
rect 478328 2 478380 8
rect 479310 -960 479422 326
rect 479524 332 479576 338
rect 479524 274 479576 280
rect 480506 -960 480618 480
rect 481376 354 481404 1158
rect 481560 678 481588 3046
rect 482480 1018 482508 3060
rect 482468 1012 482520 1018
rect 482468 954 482520 960
rect 483584 814 483612 3060
rect 483572 808 483624 814
rect 483572 750 483624 756
rect 481548 672 481600 678
rect 481548 614 481600 620
rect 481702 354 481814 480
rect 482468 468 482520 474
rect 482468 410 482520 416
rect 481376 326 481814 354
rect 482480 354 482508 410
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 481702 -960 481814 326
rect 482806 -960 482918 326
rect 484002 218 484114 480
rect 484002 202 484256 218
rect 484002 196 484268 202
rect 484002 190 484216 196
rect 484002 -960 484114 190
rect 484216 138 484268 144
rect 484688 66 484716 3060
rect 485700 1154 485728 3060
rect 485688 1148 485740 1154
rect 485688 1090 485740 1096
rect 486424 604 486476 610
rect 486424 546 486476 552
rect 486436 480 486464 546
rect 486896 542 486924 3060
rect 487252 1284 487304 1290
rect 487252 1226 487304 1232
rect 486884 536 486936 542
rect 484860 400 484912 406
rect 485198 354 485310 480
rect 484912 348 485310 354
rect 484860 342 485310 348
rect 484872 326 485310 342
rect 484676 60 484728 66
rect 484676 2 484728 8
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 486884 478 486936 484
rect 487264 354 487292 1226
rect 488000 746 488028 3060
rect 488816 1352 488868 1358
rect 488816 1294 488868 1300
rect 487988 740 488040 746
rect 487988 682 488040 688
rect 488828 480 488856 1294
rect 489104 1086 489132 3060
rect 490208 1222 490236 3060
rect 490196 1216 490248 1222
rect 490196 1158 490248 1164
rect 489092 1080 489144 1086
rect 489092 1022 489144 1028
rect 491220 610 491248 3060
rect 492416 882 492444 3060
rect 493520 1358 493548 3060
rect 493508 1352 493560 1358
rect 493508 1294 493560 1300
rect 494624 950 494652 3060
rect 495728 1018 495756 3060
rect 495532 1012 495584 1018
rect 495532 954 495584 960
rect 495716 1012 495768 1018
rect 495716 954 495768 960
rect 493140 944 493192 950
rect 493140 886 493192 892
rect 494612 944 494664 950
rect 494612 886 494664 892
rect 492404 876 492456 882
rect 492404 818 492456 824
rect 491208 604 491260 610
rect 491208 546 491260 552
rect 487590 354 487702 480
rect 487264 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 82 490002 480
rect 490748 264 490800 270
rect 491086 218 491198 480
rect 490800 212 491198 218
rect 490748 206 491198 212
rect 490760 190 491198 206
rect 490104 128 490156 134
rect 489890 76 490104 82
rect 489890 70 490156 76
rect 489890 54 490144 70
rect 489890 -960 490002 54
rect 491086 -960 491198 190
rect 492282 354 492394 480
rect 493152 354 493180 886
rect 494704 672 494756 678
rect 494704 614 494756 620
rect 494716 480 494744 614
rect 493478 354 493590 480
rect 492282 338 492536 354
rect 492282 332 492548 338
rect 492282 326 492496 332
rect 492282 -960 492394 326
rect 493152 326 493590 354
rect 492496 274 492548 280
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495544 354 495572 954
rect 495870 354 495982 480
rect 496740 406 496768 3060
rect 497096 808 497148 814
rect 497096 750 497148 756
rect 497108 480 497136 750
rect 497936 678 497964 3060
rect 499040 1290 499068 3060
rect 500144 1358 500172 3060
rect 500040 1352 500092 1358
rect 500040 1294 500092 1300
rect 500132 1352 500184 1358
rect 500132 1294 500184 1300
rect 499028 1284 499080 1290
rect 499028 1226 499080 1232
rect 499028 1148 499080 1154
rect 499028 1090 499080 1096
rect 497924 672 497976 678
rect 497924 614 497976 620
rect 495544 326 495982 354
rect 496728 400 496780 406
rect 496728 342 496780 348
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 82 498282 480
rect 499040 354 499068 1090
rect 499366 354 499478 480
rect 500052 474 500080 1294
rect 500408 1148 500460 1154
rect 500408 1090 500460 1096
rect 500420 678 500448 1090
rect 500408 672 500460 678
rect 500408 614 500460 620
rect 500592 604 500644 610
rect 500592 546 500644 552
rect 500604 480 500632 546
rect 501248 542 501276 3060
rect 502260 814 502288 3060
rect 503456 1086 503484 3060
rect 503812 1216 503864 1222
rect 503812 1158 503864 1164
rect 502984 1080 503036 1086
rect 502984 1022 503036 1028
rect 503444 1080 503496 1086
rect 503444 1022 503496 1028
rect 502248 808 502300 814
rect 502248 750 502300 756
rect 501420 740 501472 746
rect 501420 682 501472 688
rect 501236 536 501288 542
rect 500040 468 500092 474
rect 500040 410 500092 416
rect 499040 326 499478 354
rect 498170 66 498424 82
rect 498170 60 498436 66
rect 498170 54 498384 60
rect 498170 -960 498282 54
rect 498384 2 498436 8
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501236 478 501288 484
rect 501432 354 501460 682
rect 502996 480 503024 1022
rect 501758 354 501870 480
rect 501432 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503824 354 503852 1158
rect 504560 746 504588 3060
rect 504548 740 504600 746
rect 504548 682 504600 688
rect 505376 672 505428 678
rect 505376 614 505428 620
rect 505388 480 505416 614
rect 504150 354 504262 480
rect 503824 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 505664 338 505692 3060
rect 506480 876 506532 882
rect 506480 818 506532 824
rect 506492 480 506520 818
rect 505652 332 505704 338
rect 505652 274 505704 280
rect 506450 -960 506562 480
rect 506768 66 506796 3060
rect 507032 1352 507084 1358
rect 507032 1294 507084 1300
rect 507044 814 507072 1294
rect 507032 808 507084 814
rect 507032 750 507084 756
rect 507780 626 507808 3060
rect 508872 944 508924 950
rect 508872 886 508924 892
rect 507780 598 507900 626
rect 507308 468 507360 474
rect 507308 410 507360 416
rect 507320 354 507348 410
rect 507646 354 507758 480
rect 507872 474 507900 598
rect 508884 480 508912 886
rect 508976 882 509004 3060
rect 509700 1012 509752 1018
rect 509700 954 509752 960
rect 508964 876 509016 882
rect 508964 818 509016 824
rect 507860 468 507912 474
rect 507860 410 507912 416
rect 507320 326 507758 354
rect 506756 60 506808 66
rect 506756 2 506808 8
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509712 354 509740 954
rect 510080 950 510108 3060
rect 511184 1154 511212 3060
rect 512288 1290 512316 3060
rect 512276 1284 512328 1290
rect 512276 1226 512328 1232
rect 511172 1148 511224 1154
rect 511172 1090 511224 1096
rect 512092 1080 512144 1086
rect 512092 1022 512144 1028
rect 510068 944 510120 950
rect 510068 886 510120 892
rect 510038 354 510150 480
rect 509712 326 510150 354
rect 510038 -960 510150 326
rect 511234 354 511346 480
rect 511448 400 511500 406
rect 511234 348 511448 354
rect 511234 342 511500 348
rect 512104 354 512132 1022
rect 512430 354 512542 480
rect 511234 326 511488 342
rect 512104 326 512542 354
rect 511234 -960 511346 326
rect 512430 -960 512542 326
rect 513300 134 513328 3060
rect 513380 1216 513432 1222
rect 513380 1158 513432 1164
rect 513392 354 513420 1158
rect 513534 354 513646 480
rect 514496 406 514524 3060
rect 514760 808 514812 814
rect 514760 750 514812 756
rect 514772 480 514800 750
rect 513392 326 513646 354
rect 514484 400 514536 406
rect 514484 342 514536 348
rect 513288 128 513340 134
rect 513288 70 513340 76
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515508 270 515536 3060
rect 516704 1358 516732 3060
rect 516692 1352 516744 1358
rect 516692 1294 516744 1300
rect 517808 1222 517836 3060
rect 517796 1216 517848 1222
rect 517796 1158 517848 1164
rect 517980 1012 518032 1018
rect 517980 954 518032 960
rect 517152 740 517204 746
rect 517152 682 517204 688
rect 515588 536 515640 542
rect 515588 478 515640 484
rect 517164 480 517192 682
rect 515600 354 515628 478
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515496 264 515548 270
rect 515496 206 515548 212
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517992 354 518020 954
rect 518820 542 518848 3060
rect 519544 604 519596 610
rect 519544 546 519596 552
rect 518808 536 518860 542
rect 518318 354 518430 480
rect 518808 478 518860 484
rect 519556 480 519584 546
rect 517992 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520016 202 520044 3060
rect 520710 354 520822 480
rect 520384 338 520822 354
rect 521120 338 521148 3060
rect 522224 610 522252 3060
rect 522212 604 522264 610
rect 522212 546 522264 552
rect 520372 332 520822 338
rect 520424 326 520822 332
rect 520372 274 520424 280
rect 520004 196 520056 202
rect 520004 138 520056 144
rect 520710 -960 520822 326
rect 521108 332 521160 338
rect 521108 274 521160 280
rect 521814 82 521926 480
rect 521672 66 521926 82
rect 521660 60 521926 66
rect 521712 54 521926 60
rect 521660 2 521712 8
rect 521814 -960 521926 54
rect 523010 354 523122 480
rect 523224 468 523276 474
rect 523224 410 523276 416
rect 523236 354 523264 410
rect 523010 326 523264 354
rect 523010 -960 523122 326
rect 523328 66 523356 3060
rect 523868 876 523920 882
rect 523868 818 523920 824
rect 523880 354 523908 818
rect 524340 746 524368 3060
rect 525432 944 525484 950
rect 525432 886 525484 892
rect 524328 740 524380 746
rect 524328 682 524380 688
rect 525444 480 525472 886
rect 525536 678 525564 3060
rect 526640 2922 526668 3060
rect 526628 2916 526680 2922
rect 526628 2858 526680 2864
rect 526260 1148 526312 1154
rect 526260 1090 526312 1096
rect 525524 672 525576 678
rect 525524 614 525576 620
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 523316 60 523368 66
rect 523316 2 523368 8
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526272 354 526300 1090
rect 527744 814 527772 3060
rect 527824 1284 527876 1290
rect 527824 1226 527876 1232
rect 527732 808 527784 814
rect 527732 750 527784 756
rect 527836 480 527864 1226
rect 526598 354 526710 480
rect 526272 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528848 474 528876 3060
rect 529966 3046 530072 3062
rect 528836 468 528888 474
rect 528836 410 528888 416
rect 528744 128 528796 134
rect 528990 82 529102 480
rect 529940 400 529992 406
rect 530094 354 530206 480
rect 529992 348 530206 354
rect 529940 342 530206 348
rect 529952 326 530206 342
rect 528796 76 529102 82
rect 528744 70 529102 76
rect 528756 54 529102 70
rect 528990 -960 529102 54
rect 530094 -960 530206 326
rect 531056 134 531084 3060
rect 532056 1352 532108 1358
rect 532056 1294 532108 1300
rect 531290 218 531402 480
rect 532068 354 532096 1294
rect 532160 950 532188 3060
rect 532148 944 532200 950
rect 532148 886 532200 892
rect 532486 354 532598 480
rect 533264 406 533292 3060
rect 533712 1216 533764 1222
rect 533712 1158 533764 1164
rect 533724 480 533752 1158
rect 534368 1018 534396 3060
rect 534356 1012 534408 1018
rect 534356 954 534408 960
rect 534540 536 534592 542
rect 532068 326 532598 354
rect 533252 400 533304 406
rect 533252 342 533304 348
rect 531504 264 531556 270
rect 531290 212 531504 218
rect 531290 206 531556 212
rect 531290 190 531544 206
rect 531044 128 531096 134
rect 531044 70 531096 76
rect 531290 -960 531402 190
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534540 478 534592 484
rect 534552 354 534580 478
rect 534878 354 534990 480
rect 534552 326 534990 354
rect 534878 -960 534990 326
rect 535380 270 535408 3060
rect 536576 2990 536604 3060
rect 536564 2984 536616 2990
rect 536564 2926 536616 2932
rect 535368 264 535420 270
rect 535368 206 535420 212
rect 536074 218 536186 480
rect 537178 354 537290 480
rect 537178 338 537432 354
rect 537178 332 537444 338
rect 537178 326 537392 332
rect 536074 202 536328 218
rect 536074 196 536340 202
rect 536074 190 536288 196
rect 536074 -960 536186 190
rect 536288 138 536340 144
rect 537178 -960 537290 326
rect 537392 274 537444 280
rect 537680 202 537708 3060
rect 538404 604 538456 610
rect 538404 546 538456 552
rect 538416 480 538444 546
rect 537668 196 537720 202
rect 537668 138 537720 144
rect 538374 -960 538486 480
rect 538784 338 538812 3060
rect 539888 1358 539916 3060
rect 539876 1352 539928 1358
rect 539876 1294 539928 1300
rect 540900 746 540928 3060
rect 540796 740 540848 746
rect 540796 682 540848 688
rect 540888 740 540940 746
rect 540888 682 540940 688
rect 540808 480 540836 682
rect 541992 672 542044 678
rect 541992 614 542044 620
rect 542004 480 542032 614
rect 542096 610 542124 3060
rect 543214 3058 543504 3074
rect 543214 3052 543516 3058
rect 543214 3046 543464 3052
rect 544318 3046 544608 3074
rect 564348 3120 564400 3126
rect 546684 3062 546736 3068
rect 543464 2994 543516 3000
rect 542820 2916 542872 2922
rect 542820 2858 542872 2864
rect 542084 604 542136 610
rect 542084 546 542136 552
rect 538772 332 538824 338
rect 538772 274 538824 280
rect 539570 82 539682 480
rect 539570 66 539824 82
rect 539570 60 539836 66
rect 539570 54 539784 60
rect 539570 -960 539682 54
rect 539784 2 539836 8
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542832 354 542860 2858
rect 544384 808 544436 814
rect 544384 750 544436 756
rect 544396 480 544424 750
rect 544580 542 544608 3046
rect 545408 678 545436 3060
rect 545396 672 545448 678
rect 545396 614 545448 620
rect 544568 536 544620 542
rect 543158 354 543270 480
rect 542832 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 544568 478 544620 484
rect 545458 354 545570 480
rect 545672 468 545724 474
rect 545672 410 545724 416
rect 545684 354 545712 410
rect 545458 326 545712 354
rect 545458 -960 545570 326
rect 546420 66 546448 3060
rect 546500 2848 546552 2854
rect 546500 2790 546552 2796
rect 546512 1358 546540 2790
rect 546500 1352 546552 1358
rect 546500 1294 546552 1300
rect 546696 480 546724 3062
rect 547616 814 547644 3060
rect 547604 808 547656 814
rect 547604 750 547656 756
rect 546408 60 546460 66
rect 546408 2 546460 8
rect 546654 -960 546766 480
rect 547850 82 547962 480
rect 548720 474 548748 3060
rect 549824 2922 549852 3060
rect 549812 2916 549864 2922
rect 549812 2858 549864 2864
rect 549076 944 549128 950
rect 549076 886 549128 892
rect 549088 480 549116 886
rect 550928 882 550956 3060
rect 551468 1012 551520 1018
rect 551468 954 551520 960
rect 550916 876 550968 882
rect 550916 818 550968 824
rect 551480 480 551508 954
rect 548708 468 548760 474
rect 548708 410 548760 416
rect 548064 128 548116 134
rect 547850 76 548064 82
rect 547850 70 548116 76
rect 547850 54 548104 70
rect 547850 -960 547962 54
rect 549046 -960 549158 480
rect 550242 354 550354 480
rect 550456 400 550508 406
rect 550242 348 550456 354
rect 550242 342 550508 348
rect 550242 326 550496 342
rect 550242 -960 550354 326
rect 551438 -960 551550 480
rect 551940 134 551968 3060
rect 553768 2984 553820 2990
rect 553768 2926 553820 2932
rect 553780 480 553808 2926
rect 552634 218 552746 480
rect 552848 264 552900 270
rect 552634 212 552848 218
rect 552634 206 552900 212
rect 552634 190 552888 206
rect 551928 128 551980 134
rect 551928 70 551980 76
rect 552634 -960 552746 190
rect 553738 -960 553850 480
rect 554240 270 554268 3060
rect 554228 264 554280 270
rect 554934 218 555046 480
rect 555344 406 555372 3060
rect 557184 3046 557474 3074
rect 558670 3046 558868 3074
rect 555332 400 555384 406
rect 555332 342 555384 348
rect 556130 354 556242 480
rect 554228 206 554280 212
rect 554792 202 555046 218
rect 554780 196 555046 202
rect 554832 190 555046 196
rect 554780 138 554832 144
rect 554934 -960 555046 190
rect 556130 338 556384 354
rect 557184 338 557212 3046
rect 557356 2848 557408 2854
rect 557356 2790 557408 2796
rect 557368 480 557396 2790
rect 558552 740 558604 746
rect 558552 682 558604 688
rect 558564 480 558592 682
rect 556130 332 556396 338
rect 556130 326 556344 332
rect 556130 -960 556242 326
rect 556344 274 556396 280
rect 557172 332 557224 338
rect 557172 274 557224 280
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 558840 202 558868 3046
rect 560484 3052 560536 3058
rect 560484 2994 560536 3000
rect 559748 604 559800 610
rect 559748 546 559800 552
rect 559760 480 559788 546
rect 558828 196 558880 202
rect 558828 138 558880 144
rect 559718 -960 559830 480
rect 560496 354 560524 2994
rect 560864 2990 560892 3060
rect 561982 3058 562272 3074
rect 564190 3068 564348 3074
rect 564190 3062 564400 3068
rect 561982 3052 562284 3058
rect 561982 3046 562232 3052
rect 562232 2994 562284 3000
rect 560852 2984 560904 2990
rect 560852 2926 560904 2932
rect 562980 2854 563008 3060
rect 564190 3046 564388 3062
rect 568028 2916 568080 2922
rect 568028 2858 568080 2864
rect 562968 2848 563020 2854
rect 562968 2790 563020 2796
rect 565636 808 565688 814
rect 565636 750 565688 756
rect 563244 672 563296 678
rect 563244 614 563296 620
rect 562048 604 562100 610
rect 562048 546 562100 552
rect 562060 480 562088 546
rect 563256 480 563284 614
rect 565648 480 565676 750
rect 568040 480 568068 2858
rect 569132 876 569184 882
rect 569132 818 569184 824
rect 569144 480 569172 818
rect 571536 480 571564 3198
rect 575112 3188 575164 3194
rect 575112 3130 575164 3136
rect 575124 480 575152 3130
rect 578620 480 578648 3266
rect 583392 3120 583444 3126
rect 583392 3062 583444 3068
rect 581000 3052 581052 3058
rect 581000 2994 581052 3000
rect 579804 2984 579856 2990
rect 579804 2926 579856 2932
rect 579816 480 579844 2926
rect 581012 480 581040 2994
rect 582196 2848 582248 2854
rect 582196 2790 582248 2796
rect 582208 480 582236 2790
rect 583404 480 583432 3062
rect 560822 354 560934 480
rect 560496 326 560934 354
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 82 564522 480
rect 564410 66 564664 82
rect 564410 60 564676 66
rect 564410 54 564624 60
rect 564410 -960 564522 54
rect 564624 2 564676 8
rect 565606 -960 565718 480
rect 566802 354 566914 480
rect 567016 468 567068 474
rect 567016 410 567068 416
rect 567028 354 567056 410
rect 566802 326 567056 354
rect 566802 -960 566914 326
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 82 570410 480
rect 570512 128 570564 134
rect 570298 76 570512 82
rect 570298 70 570564 76
rect 570298 54 570552 70
rect 570298 -960 570410 54
rect 571494 -960 571606 480
rect 572690 218 572802 480
rect 573548 400 573600 406
rect 573886 354 573998 480
rect 573600 348 573998 354
rect 573548 342 573998 348
rect 573560 326 573998 342
rect 572904 264 572956 270
rect 572690 212 572904 218
rect 572690 206 572956 212
rect 572690 190 572944 206
rect 572690 -960 572802 190
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 354 576390 480
rect 575952 338 576390 354
rect 575940 332 576390 338
rect 575992 326 576390 332
rect 575940 274 575992 280
rect 576278 -960 576390 326
rect 577382 218 577494 480
rect 577148 202 577494 218
rect 577136 196 577494 202
rect 577188 190 577494 196
rect 577136 138 577188 144
rect 577382 -960 577494 190
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2042 697312 2098 697368
rect 581642 697176 581698 697232
rect 581642 691464 581698 691520
rect 2042 690784 2098 690840
rect 1030 684256 1086 684312
rect 582378 683848 582434 683904
rect 582378 678408 582434 678464
rect 1030 678000 1086 678056
rect 1030 671200 1086 671256
rect 582378 670656 582434 670712
rect 582378 665352 582434 665408
rect 1030 665216 1086 665272
rect 18 657600 74 657656
rect 582378 657328 582434 657384
rect 18 652432 74 652488
rect 582378 652296 582434 652352
rect 1306 645088 1362 645144
rect 581642 644000 581698 644056
rect 1306 639648 1362 639704
rect 581642 639240 581698 639296
rect 1306 632032 1362 632088
rect 582378 630808 582434 630864
rect 1306 626864 1362 626920
rect 582378 626184 582434 626240
rect 18 618568 74 618624
rect 581642 617480 581698 617536
rect 18 613944 74 614000
rect 581642 613128 581698 613184
rect 846 606056 902 606112
rect 581642 604152 581698 604208
rect 846 601296 902 601352
rect 581642 600072 581698 600128
rect 2778 593000 2834 593056
rect 581642 590960 581698 591016
rect 2778 588512 2834 588568
rect 581642 587016 581698 587072
rect 2778 579944 2834 580000
rect 581642 577632 581698 577688
rect 2778 575728 2834 575784
rect 581642 573960 581698 574016
rect 2778 566888 2834 566944
rect 582378 564304 582434 564360
rect 2778 562944 2834 563000
rect 582378 560904 582434 560960
rect 2778 553832 2834 553888
rect 581642 551112 581698 551168
rect 2778 550160 2834 550216
rect 581642 547712 581698 547768
rect 1398 540776 1454 540832
rect 582378 537784 582434 537840
rect 1398 537376 1454 537432
rect 582378 534792 582434 534848
rect 1490 527856 1546 527912
rect 1490 524592 1546 524648
rect 582378 524456 582434 524512
rect 582378 521736 582434 521792
rect 2778 514800 2834 514856
rect 2778 511808 2834 511864
rect 582378 511264 582434 511320
rect 582378 508680 582434 508736
rect 1582 501744 1638 501800
rect 1582 499024 1638 499080
rect 581642 497936 581698 497992
rect 581642 495624 581698 495680
rect 1582 488688 1638 488744
rect 1582 486240 1638 486296
rect 582378 484608 582434 484664
rect 582378 482568 582434 482624
rect 2778 475632 2834 475688
rect 2778 473456 2834 473512
rect 581642 471416 581698 471472
rect 581642 469512 581698 469568
rect 1582 462576 1638 462632
rect 1582 460672 1638 460728
rect 581642 458088 581698 458144
rect 581642 456456 581698 456512
rect 2778 449520 2834 449576
rect 2778 447888 2834 447944
rect 2778 436600 2834 436656
rect 2778 435104 2834 435160
rect 2778 423544 2834 423600
rect 2778 422320 2834 422376
rect 1306 294344 1362 294400
rect 1306 293120 1362 293176
rect 2778 281560 2834 281616
rect 2778 280064 2834 280120
rect 1306 268776 1362 268832
rect 1306 267144 1362 267200
rect 582378 260480 582434 260536
rect 582378 258848 582434 258904
rect 1306 255992 1362 256048
rect 1306 254088 1362 254144
rect 580906 247016 580962 247072
rect 580906 245520 580962 245576
rect 2778 243208 2834 243264
rect 2778 241032 2834 241088
rect 582378 234368 582434 234424
rect 582378 232328 582434 232384
rect 2778 230560 2834 230616
rect 2778 227976 2834 228032
rect 580906 220904 580962 220960
rect 580906 219000 580962 219056
rect 2778 217640 2834 217696
rect 2778 214920 2834 214976
rect 582378 208256 582434 208312
rect 582378 205672 582434 205728
rect 2778 204856 2834 204912
rect 2778 201864 2834 201920
rect 580906 194656 580962 194712
rect 580906 192480 580962 192536
rect 1306 192072 1362 192128
rect 1306 188808 1362 188864
rect 580906 182416 580962 182472
rect 2778 179288 2834 179344
rect 580906 179152 580962 179208
rect 2778 175888 2834 175944
rect 580906 168544 580962 168600
rect 2778 166504 2834 166560
rect 580906 165824 580962 165880
rect 2778 162832 2834 162888
rect 580906 156304 580962 156360
rect 1306 153720 1362 153776
rect 580906 152632 580962 152688
rect 1306 149776 1362 149832
rect 580906 142568 580962 142624
rect 570 140936 626 140992
rect 580906 139304 580962 139360
rect 570 136720 626 136776
rect 580906 130192 580962 130248
rect 754 128152 810 128208
rect 580906 125976 580962 126032
rect 754 123664 810 123720
rect 579894 116320 579950 116376
rect 1306 115368 1362 115424
rect 579894 112784 579950 112840
rect 1306 110608 1362 110664
rect 580906 103536 580962 103592
rect 1582 102584 1638 102640
rect 580906 99456 580962 99512
rect 1582 97552 1638 97608
rect 580906 90208 580962 90264
rect 1582 89800 1638 89856
rect 580906 86128 580962 86184
rect 1582 84632 1638 84688
rect 579894 77288 579950 77344
rect 1582 77016 1638 77072
rect 579894 72936 579950 72992
rect 1582 71576 1638 71632
rect 1490 64232 1546 64288
rect 580906 64096 580962 64152
rect 580906 59608 580962 59664
rect 1490 58520 1546 58576
rect 2778 51448 2834 51504
rect 580906 51040 580962 51096
rect 580906 46280 580962 46336
rect 2778 45464 2834 45520
rect 2778 38664 2834 38720
rect 580906 37984 580962 38040
rect 580906 33088 580962 33144
rect 2778 32408 2834 32464
rect 1490 25880 1546 25936
rect 580906 24928 580962 24984
rect 580906 19760 580962 19816
rect 1490 19352 1546 19408
rect 2778 13096 2834 13152
rect 579894 12688 579950 12744
rect 579894 6568 579950 6624
rect 2778 6432 2834 6488
rect 5446 176 5502 232
rect 6274 40 6330 96
rect 12162 448 12218 504
rect 13726 312 13782 368
rect 23938 176 23994 232
rect 25042 40 25098 96
rect 25686 176 25742 232
rect 28906 584 28962 640
rect 30838 448 30894 504
rect 31942 312 31998 368
rect 37002 40 37058 96
rect 42706 176 42762 232
rect 46294 584 46350 640
rect 46846 176 46902 232
rect 54022 40 54078 96
rect 62854 176 62910 232
<< metal3 >>
rect -960 697370 480 697460
rect 2037 697370 2103 697373
rect -960 697368 2103 697370
rect -960 697312 2042 697368
rect 2098 697312 2103 697368
rect -960 697310 2103 697312
rect -960 697220 480 697310
rect 2037 697307 2103 697310
rect 581637 697234 581703 697237
rect 583520 697234 584960 697324
rect 581637 697232 584960 697234
rect 581637 697176 581642 697232
rect 581698 697176 584960 697232
rect 581637 697174 584960 697176
rect 581637 697171 581703 697174
rect 583520 697084 584960 697174
rect 581637 691522 581703 691525
rect 580796 691520 581703 691522
rect 580796 691464 581642 691520
rect 581698 691464 581703 691520
rect 580796 691462 581703 691464
rect 581637 691459 581703 691462
rect 2037 690842 2103 690845
rect 2037 690840 3220 690842
rect 2037 690784 2042 690840
rect 2098 690784 3220 690840
rect 2037 690782 3220 690784
rect 2037 690779 2103 690782
rect -960 684314 480 684404
rect 1025 684314 1091 684317
rect -960 684312 1091 684314
rect -960 684256 1030 684312
rect 1086 684256 1091 684312
rect -960 684254 1091 684256
rect -960 684164 480 684254
rect 1025 684251 1091 684254
rect 582373 683906 582439 683909
rect 583520 683906 584960 683996
rect 582373 683904 584960 683906
rect 582373 683848 582378 683904
rect 582434 683848 584960 683904
rect 582373 683846 584960 683848
rect 582373 683843 582439 683846
rect 583520 683756 584960 683846
rect 582373 678466 582439 678469
rect 580796 678464 582439 678466
rect 580796 678408 582378 678464
rect 582434 678408 582439 678464
rect 580796 678406 582439 678408
rect 582373 678403 582439 678406
rect 1025 678058 1091 678061
rect 1025 678056 3220 678058
rect 1025 678000 1030 678056
rect 1086 678000 3220 678056
rect 1025 677998 3220 678000
rect 1025 677995 1091 677998
rect -960 671258 480 671348
rect 1025 671258 1091 671261
rect -960 671256 1091 671258
rect -960 671200 1030 671256
rect 1086 671200 1091 671256
rect -960 671198 1091 671200
rect -960 671108 480 671198
rect 1025 671195 1091 671198
rect 582373 670714 582439 670717
rect 583520 670714 584960 670804
rect 582373 670712 584960 670714
rect 582373 670656 582378 670712
rect 582434 670656 584960 670712
rect 582373 670654 584960 670656
rect 582373 670651 582439 670654
rect 583520 670564 584960 670654
rect 582373 665410 582439 665413
rect 580796 665408 582439 665410
rect 580796 665352 582378 665408
rect 582434 665352 582439 665408
rect 580796 665350 582439 665352
rect 582373 665347 582439 665350
rect 1025 665274 1091 665277
rect 1025 665272 3220 665274
rect 1025 665216 1030 665272
rect 1086 665216 3220 665272
rect 1025 665214 3220 665216
rect 1025 665211 1091 665214
rect -960 658202 480 658292
rect -960 658142 674 658202
rect -960 658066 480 658142
rect 614 658066 674 658142
rect -960 658052 674 658066
rect 62 658006 674 658052
rect 62 657661 122 658006
rect 13 657656 122 657661
rect 13 657600 18 657656
rect 74 657600 122 657656
rect 13 657598 122 657600
rect 13 657595 79 657598
rect 582373 657386 582439 657389
rect 583520 657386 584960 657476
rect 582373 657384 584960 657386
rect 582373 657328 582378 657384
rect 582434 657328 584960 657384
rect 582373 657326 584960 657328
rect 582373 657323 582439 657326
rect 583520 657236 584960 657326
rect 13 652490 79 652493
rect 13 652488 3220 652490
rect 13 652432 18 652488
rect 74 652432 3220 652488
rect 13 652430 3220 652432
rect 13 652427 79 652430
rect 582373 652354 582439 652357
rect 580796 652352 582439 652354
rect 580796 652296 582378 652352
rect 582434 652296 582439 652352
rect 580796 652294 582439 652296
rect 582373 652291 582439 652294
rect -960 645146 480 645236
rect 1301 645146 1367 645149
rect -960 645144 1367 645146
rect -960 645088 1306 645144
rect 1362 645088 1367 645144
rect -960 645086 1367 645088
rect -960 644996 480 645086
rect 1301 645083 1367 645086
rect 581637 644058 581703 644061
rect 583520 644058 584960 644148
rect 581637 644056 584960 644058
rect 581637 644000 581642 644056
rect 581698 644000 584960 644056
rect 581637 643998 584960 644000
rect 581637 643995 581703 643998
rect 583520 643908 584960 643998
rect 1301 639706 1367 639709
rect 1301 639704 3220 639706
rect 1301 639648 1306 639704
rect 1362 639648 3220 639704
rect 1301 639646 3220 639648
rect 1301 639643 1367 639646
rect 581637 639298 581703 639301
rect 580796 639296 581703 639298
rect 580796 639240 581642 639296
rect 581698 639240 581703 639296
rect 580796 639238 581703 639240
rect 581637 639235 581703 639238
rect -960 632090 480 632180
rect 1301 632090 1367 632093
rect -960 632088 1367 632090
rect -960 632032 1306 632088
rect 1362 632032 1367 632088
rect -960 632030 1367 632032
rect -960 631940 480 632030
rect 1301 632027 1367 632030
rect 582373 630866 582439 630869
rect 583520 630866 584960 630956
rect 582373 630864 584960 630866
rect 582373 630808 582378 630864
rect 582434 630808 584960 630864
rect 582373 630806 584960 630808
rect 582373 630803 582439 630806
rect 583520 630716 584960 630806
rect 1301 626922 1367 626925
rect 1301 626920 3220 626922
rect 1301 626864 1306 626920
rect 1362 626864 3220 626920
rect 1301 626862 3220 626864
rect 1301 626859 1367 626862
rect 582373 626242 582439 626245
rect 580796 626240 582439 626242
rect 580796 626184 582378 626240
rect 582434 626184 582439 626240
rect 580796 626182 582439 626184
rect 582373 626179 582439 626182
rect -960 619170 480 619260
rect -960 619110 674 619170
rect -960 619034 480 619110
rect 614 619034 674 619110
rect -960 619020 674 619034
rect 62 618974 674 619020
rect 62 618629 122 618974
rect 13 618624 122 618629
rect 13 618568 18 618624
rect 74 618568 122 618624
rect 13 618566 122 618568
rect 13 618563 79 618566
rect 581637 617538 581703 617541
rect 583520 617538 584960 617628
rect 581637 617536 584960 617538
rect 581637 617480 581642 617536
rect 581698 617480 584960 617536
rect 581637 617478 584960 617480
rect 581637 617475 581703 617478
rect 583520 617388 584960 617478
rect 13 614002 79 614005
rect 13 614000 3220 614002
rect 13 613944 18 614000
rect 74 613944 3220 614000
rect 13 613942 3220 613944
rect 13 613939 79 613942
rect 581637 613186 581703 613189
rect 580796 613184 581703 613186
rect 580796 613128 581642 613184
rect 581698 613128 581703 613184
rect 580796 613126 581703 613128
rect 581637 613123 581703 613126
rect -960 606114 480 606204
rect 841 606114 907 606117
rect -960 606112 907 606114
rect -960 606056 846 606112
rect 902 606056 907 606112
rect -960 606054 907 606056
rect -960 605964 480 606054
rect 841 606051 907 606054
rect 581637 604210 581703 604213
rect 583520 604210 584960 604300
rect 581637 604208 584960 604210
rect 581637 604152 581642 604208
rect 581698 604152 584960 604208
rect 581637 604150 584960 604152
rect 581637 604147 581703 604150
rect 583520 604060 584960 604150
rect 841 601354 907 601357
rect 841 601352 3220 601354
rect 841 601296 846 601352
rect 902 601296 3220 601352
rect 841 601294 3220 601296
rect 841 601291 907 601294
rect 581637 600130 581703 600133
rect 580796 600128 581703 600130
rect 580796 600072 581642 600128
rect 581698 600072 581703 600128
rect 580796 600070 581703 600072
rect 581637 600067 581703 600070
rect -960 593058 480 593148
rect 2773 593058 2839 593061
rect -960 593056 2839 593058
rect -960 593000 2778 593056
rect 2834 593000 2839 593056
rect -960 592998 2839 593000
rect -960 592908 480 592998
rect 2773 592995 2839 592998
rect 581637 591018 581703 591021
rect 583520 591018 584960 591108
rect 581637 591016 584960 591018
rect 581637 590960 581642 591016
rect 581698 590960 584960 591016
rect 581637 590958 584960 590960
rect 581637 590955 581703 590958
rect 583520 590868 584960 590958
rect 2773 588570 2839 588573
rect 2773 588568 3220 588570
rect 2773 588512 2778 588568
rect 2834 588512 3220 588568
rect 2773 588510 3220 588512
rect 2773 588507 2839 588510
rect 581637 587074 581703 587077
rect 580796 587072 581703 587074
rect 580796 587016 581642 587072
rect 581698 587016 581703 587072
rect 580796 587014 581703 587016
rect 581637 587011 581703 587014
rect -960 580002 480 580092
rect 2773 580002 2839 580005
rect -960 580000 2839 580002
rect -960 579944 2778 580000
rect 2834 579944 2839 580000
rect -960 579942 2839 579944
rect -960 579852 480 579942
rect 2773 579939 2839 579942
rect 581637 577690 581703 577693
rect 583520 577690 584960 577780
rect 581637 577688 584960 577690
rect 581637 577632 581642 577688
rect 581698 577632 584960 577688
rect 581637 577630 584960 577632
rect 581637 577627 581703 577630
rect 583520 577540 584960 577630
rect 2773 575786 2839 575789
rect 2773 575784 3220 575786
rect 2773 575728 2778 575784
rect 2834 575728 3220 575784
rect 2773 575726 3220 575728
rect 2773 575723 2839 575726
rect 581637 574018 581703 574021
rect 580796 574016 581703 574018
rect 580796 573960 581642 574016
rect 581698 573960 581703 574016
rect 580796 573958 581703 573960
rect 581637 573955 581703 573958
rect -960 566946 480 567036
rect 2773 566946 2839 566949
rect -960 566944 2839 566946
rect -960 566888 2778 566944
rect 2834 566888 2839 566944
rect -960 566886 2839 566888
rect -960 566796 480 566886
rect 2773 566883 2839 566886
rect 582373 564362 582439 564365
rect 583520 564362 584960 564452
rect 582373 564360 584960 564362
rect 582373 564304 582378 564360
rect 582434 564304 584960 564360
rect 582373 564302 584960 564304
rect 582373 564299 582439 564302
rect 583520 564212 584960 564302
rect 2773 563002 2839 563005
rect 2773 563000 3220 563002
rect 2773 562944 2778 563000
rect 2834 562944 3220 563000
rect 2773 562942 3220 562944
rect 2773 562939 2839 562942
rect 582373 560962 582439 560965
rect 580796 560960 582439 560962
rect 580796 560904 582378 560960
rect 582434 560904 582439 560960
rect 580796 560902 582439 560904
rect 582373 560899 582439 560902
rect -960 553890 480 553980
rect 2773 553890 2839 553893
rect -960 553888 2839 553890
rect -960 553832 2778 553888
rect 2834 553832 2839 553888
rect -960 553830 2839 553832
rect -960 553740 480 553830
rect 2773 553827 2839 553830
rect 581637 551170 581703 551173
rect 583520 551170 584960 551260
rect 581637 551168 584960 551170
rect 581637 551112 581642 551168
rect 581698 551112 584960 551168
rect 581637 551110 584960 551112
rect 581637 551107 581703 551110
rect 583520 551020 584960 551110
rect 2773 550218 2839 550221
rect 2773 550216 3220 550218
rect 2773 550160 2778 550216
rect 2834 550160 3220 550216
rect 2773 550158 3220 550160
rect 2773 550155 2839 550158
rect 581637 547770 581703 547773
rect 580796 547768 581703 547770
rect 580796 547712 581642 547768
rect 581698 547712 581703 547768
rect 580796 547710 581703 547712
rect 581637 547707 581703 547710
rect -960 540834 480 540924
rect 1393 540834 1459 540837
rect -960 540832 1459 540834
rect -960 540776 1398 540832
rect 1454 540776 1459 540832
rect -960 540774 1459 540776
rect -960 540684 480 540774
rect 1393 540771 1459 540774
rect 582373 537842 582439 537845
rect 583520 537842 584960 537932
rect 582373 537840 584960 537842
rect 582373 537784 582378 537840
rect 582434 537784 584960 537840
rect 582373 537782 584960 537784
rect 582373 537779 582439 537782
rect 583520 537692 584960 537782
rect 1393 537434 1459 537437
rect 1393 537432 3220 537434
rect 1393 537376 1398 537432
rect 1454 537376 3220 537432
rect 1393 537374 3220 537376
rect 1393 537371 1459 537374
rect 582373 534850 582439 534853
rect 580796 534848 582439 534850
rect 580796 534792 582378 534848
rect 582434 534792 582439 534848
rect 580796 534790 582439 534792
rect 582373 534787 582439 534790
rect -960 527914 480 528004
rect 1485 527914 1551 527917
rect -960 527912 1551 527914
rect -960 527856 1490 527912
rect 1546 527856 1551 527912
rect -960 527854 1551 527856
rect -960 527764 480 527854
rect 1485 527851 1551 527854
rect 1485 524650 1551 524653
rect 1485 524648 3220 524650
rect 1485 524592 1490 524648
rect 1546 524592 3220 524648
rect 1485 524590 3220 524592
rect 1485 524587 1551 524590
rect 582373 524514 582439 524517
rect 583520 524514 584960 524604
rect 582373 524512 584960 524514
rect 582373 524456 582378 524512
rect 582434 524456 584960 524512
rect 582373 524454 584960 524456
rect 582373 524451 582439 524454
rect 583520 524364 584960 524454
rect 582373 521794 582439 521797
rect 580796 521792 582439 521794
rect 580796 521736 582378 521792
rect 582434 521736 582439 521792
rect 580796 521734 582439 521736
rect 582373 521731 582439 521734
rect -960 514858 480 514948
rect 2773 514858 2839 514861
rect -960 514856 2839 514858
rect -960 514800 2778 514856
rect 2834 514800 2839 514856
rect -960 514798 2839 514800
rect -960 514708 480 514798
rect 2773 514795 2839 514798
rect 2773 511866 2839 511869
rect 2773 511864 3220 511866
rect 2773 511808 2778 511864
rect 2834 511808 3220 511864
rect 2773 511806 3220 511808
rect 2773 511803 2839 511806
rect 582373 511322 582439 511325
rect 583520 511322 584960 511412
rect 582373 511320 584960 511322
rect 582373 511264 582378 511320
rect 582434 511264 584960 511320
rect 582373 511262 584960 511264
rect 582373 511259 582439 511262
rect 583520 511172 584960 511262
rect 582373 508738 582439 508741
rect 580796 508736 582439 508738
rect 580796 508680 582378 508736
rect 582434 508680 582439 508736
rect 580796 508678 582439 508680
rect 582373 508675 582439 508678
rect -960 501802 480 501892
rect 1577 501802 1643 501805
rect -960 501800 1643 501802
rect -960 501744 1582 501800
rect 1638 501744 1643 501800
rect -960 501742 1643 501744
rect -960 501652 480 501742
rect 1577 501739 1643 501742
rect 1577 499082 1643 499085
rect 1577 499080 3220 499082
rect 1577 499024 1582 499080
rect 1638 499024 3220 499080
rect 1577 499022 3220 499024
rect 1577 499019 1643 499022
rect 581637 497994 581703 497997
rect 583520 497994 584960 498084
rect 581637 497992 584960 497994
rect 581637 497936 581642 497992
rect 581698 497936 584960 497992
rect 581637 497934 584960 497936
rect 581637 497931 581703 497934
rect 583520 497844 584960 497934
rect 581637 495682 581703 495685
rect 580796 495680 581703 495682
rect 580796 495624 581642 495680
rect 581698 495624 581703 495680
rect 580796 495622 581703 495624
rect 581637 495619 581703 495622
rect -960 488746 480 488836
rect 1577 488746 1643 488749
rect -960 488744 1643 488746
rect -960 488688 1582 488744
rect 1638 488688 1643 488744
rect -960 488686 1643 488688
rect -960 488596 480 488686
rect 1577 488683 1643 488686
rect 1577 486298 1643 486301
rect 1577 486296 3220 486298
rect 1577 486240 1582 486296
rect 1638 486240 3220 486296
rect 1577 486238 3220 486240
rect 1577 486235 1643 486238
rect 582373 484666 582439 484669
rect 583520 484666 584960 484756
rect 582373 484664 584960 484666
rect 582373 484608 582378 484664
rect 582434 484608 584960 484664
rect 582373 484606 584960 484608
rect 582373 484603 582439 484606
rect 583520 484516 584960 484606
rect 582373 482626 582439 482629
rect 580796 482624 582439 482626
rect 580796 482568 582378 482624
rect 582434 482568 582439 482624
rect 580796 482566 582439 482568
rect 582373 482563 582439 482566
rect -960 475690 480 475780
rect 2773 475690 2839 475693
rect -960 475688 2839 475690
rect -960 475632 2778 475688
rect 2834 475632 2839 475688
rect -960 475630 2839 475632
rect -960 475540 480 475630
rect 2773 475627 2839 475630
rect 2773 473514 2839 473517
rect 2773 473512 3220 473514
rect 2773 473456 2778 473512
rect 2834 473456 3220 473512
rect 2773 473454 3220 473456
rect 2773 473451 2839 473454
rect 581637 471474 581703 471477
rect 583520 471474 584960 471564
rect 581637 471472 584960 471474
rect 581637 471416 581642 471472
rect 581698 471416 584960 471472
rect 581637 471414 584960 471416
rect 581637 471411 581703 471414
rect 583520 471324 584960 471414
rect 581637 469570 581703 469573
rect 580796 469568 581703 469570
rect 580796 469512 581642 469568
rect 581698 469512 581703 469568
rect 580796 469510 581703 469512
rect 581637 469507 581703 469510
rect -960 462634 480 462724
rect 1577 462634 1643 462637
rect -960 462632 1643 462634
rect -960 462576 1582 462632
rect 1638 462576 1643 462632
rect -960 462574 1643 462576
rect -960 462484 480 462574
rect 1577 462571 1643 462574
rect 1577 460730 1643 460733
rect 1577 460728 3220 460730
rect 1577 460672 1582 460728
rect 1638 460672 3220 460728
rect 1577 460670 3220 460672
rect 1577 460667 1643 460670
rect 581637 458146 581703 458149
rect 583520 458146 584960 458236
rect 581637 458144 584960 458146
rect 581637 458088 581642 458144
rect 581698 458088 584960 458144
rect 581637 458086 584960 458088
rect 581637 458083 581703 458086
rect 583520 457996 584960 458086
rect 581637 456514 581703 456517
rect 580796 456512 581703 456514
rect 580796 456456 581642 456512
rect 581698 456456 581703 456512
rect 580796 456454 581703 456456
rect 581637 456451 581703 456454
rect -960 449578 480 449668
rect 2773 449578 2839 449581
rect -960 449576 2839 449578
rect -960 449520 2778 449576
rect 2834 449520 2839 449576
rect -960 449518 2839 449520
rect -960 449428 480 449518
rect 2773 449515 2839 449518
rect 2773 447946 2839 447949
rect 2773 447944 3220 447946
rect 2773 447888 2778 447944
rect 2834 447888 3220 447944
rect 2773 447886 3220 447888
rect 2773 447883 2839 447886
rect 583520 444818 584960 444908
rect 583342 444758 584960 444818
rect 583342 444682 583402 444758
rect 583520 444682 584960 444758
rect 583342 444668 584960 444682
rect 583342 444622 583586 444668
rect 583526 444138 583586 444622
rect 580766 444078 583586 444138
rect 580766 443428 580826 444078
rect -960 436658 480 436748
rect 2773 436658 2839 436661
rect -960 436656 2839 436658
rect -960 436600 2778 436656
rect 2834 436600 2839 436656
rect -960 436598 2839 436600
rect -960 436508 480 436598
rect 2773 436595 2839 436598
rect 2773 435162 2839 435165
rect 2773 435160 3220 435162
rect 2773 435104 2778 435160
rect 2834 435104 3220 435160
rect 2773 435102 3220 435104
rect 2773 435099 2839 435102
rect 583520 431626 584960 431716
rect 583342 431566 584960 431626
rect 583342 431490 583402 431566
rect 583520 431490 584960 431566
rect 583342 431476 584960 431490
rect 583342 431430 583586 431476
rect 583526 431082 583586 431430
rect 580766 431022 583586 431082
rect 580766 430372 580826 431022
rect -960 423602 480 423692
rect 2773 423602 2839 423605
rect -960 423600 2839 423602
rect -960 423544 2778 423600
rect 2834 423544 2839 423600
rect -960 423542 2839 423544
rect -960 423452 480 423542
rect 2773 423539 2839 423542
rect 2773 422378 2839 422381
rect 2773 422376 3220 422378
rect 2773 422320 2778 422376
rect 2834 422320 3220 422376
rect 2773 422318 3220 422320
rect 2773 422315 2839 422318
rect 583520 418298 584960 418388
rect 583342 418238 584960 418298
rect 583342 418162 583402 418238
rect 583520 418162 584960 418238
rect 583342 418148 584960 418162
rect 583342 418102 583586 418148
rect 583526 417754 583586 418102
rect 580766 417694 583586 417754
rect 580766 417316 580826 417694
rect -960 410546 480 410636
rect -960 410486 3250 410546
rect -960 410396 480 410486
rect 3190 409564 3250 410486
rect 583520 404970 584960 405060
rect 580766 404910 584960 404970
rect 580766 404260 580826 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect -960 397430 3250 397490
rect -960 397340 480 397430
rect 3190 396780 3250 397430
rect 583520 391778 584960 391868
rect 580766 391718 584960 391778
rect 580766 391204 580826 391718
rect 583520 391628 584960 391718
rect -960 384434 480 384524
rect -960 384374 3250 384434
rect -960 384284 480 384374
rect 3190 383996 3250 384374
rect 583520 378450 584960 378540
rect 580766 378390 584960 378450
rect 580766 378148 580826 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect -960 371318 3250 371378
rect -960 371228 480 371318
rect 3190 371212 3250 371318
rect 583520 365122 584960 365212
rect 580796 365062 584960 365122
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect -960 358398 3220 358458
rect -960 358308 480 358398
rect 583520 351930 584960 352020
rect 580796 351870 584960 351930
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 1534 345478 3220 345538
rect 1534 345402 1594 345478
rect -960 345342 1594 345402
rect -960 345252 480 345342
rect 580766 338602 580826 338844
rect 583520 338602 584960 338692
rect 580766 338542 584960 338602
rect 583520 338452 584960 338542
rect -960 332346 480 332436
rect 3190 332346 3250 332724
rect -960 332286 3250 332346
rect -960 332196 480 332286
rect 580766 325274 580826 325788
rect 583520 325274 584960 325364
rect 580766 325214 584960 325274
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3190 319290 3250 319940
rect -960 319230 3250 319290
rect -960 319140 480 319230
rect 580766 312082 580826 312732
rect 583520 312082 584960 312172
rect 580766 312022 584960 312082
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3190 306234 3250 307156
rect -960 306174 3250 306234
rect -960 306084 480 306174
rect 580766 299298 580826 299676
rect 580766 299238 583586 299298
rect 583526 298890 583586 299238
rect 583342 298844 583586 298890
rect 583342 298830 584960 298844
rect 583342 298754 583402 298830
rect 583520 298754 584960 298830
rect 583342 298694 584960 298754
rect 583520 298604 584960 298694
rect 1301 294402 1367 294405
rect 1301 294400 3220 294402
rect 1301 294344 1306 294400
rect 1362 294344 3220 294400
rect 1301 294342 3220 294344
rect 1301 294339 1367 294342
rect -960 293178 480 293268
rect 1301 293178 1367 293181
rect -960 293176 1367 293178
rect -960 293120 1306 293176
rect 1362 293120 1367 293176
rect -960 293118 1367 293120
rect -960 293028 480 293118
rect 1301 293115 1367 293118
rect 580766 285970 580826 286620
rect 580766 285910 583586 285970
rect 583526 285562 583586 285910
rect 583342 285516 583586 285562
rect 583342 285502 584960 285516
rect 583342 285426 583402 285502
rect 583520 285426 584960 285502
rect 583342 285366 584960 285426
rect 583520 285276 584960 285366
rect 2773 281618 2839 281621
rect 2773 281616 3220 281618
rect 2773 281560 2778 281616
rect 2834 281560 3220 281616
rect 2773 281558 3220 281560
rect 2773 281555 2839 281558
rect -960 280122 480 280212
rect 2773 280122 2839 280125
rect -960 280120 2839 280122
rect -960 280064 2778 280120
rect 2834 280064 2839 280120
rect -960 280062 2839 280064
rect -960 279972 480 280062
rect 2773 280059 2839 280062
rect 580766 272914 580826 273564
rect 580766 272854 583586 272914
rect 583526 272370 583586 272854
rect 583342 272324 583586 272370
rect 583342 272310 584960 272324
rect 583342 272234 583402 272310
rect 583520 272234 584960 272310
rect 583342 272174 584960 272234
rect 583520 272084 584960 272174
rect 1301 268834 1367 268837
rect 1301 268832 3220 268834
rect 1301 268776 1306 268832
rect 1362 268776 3220 268832
rect 1301 268774 3220 268776
rect 1301 268771 1367 268774
rect -960 267202 480 267292
rect 1301 267202 1367 267205
rect -960 267200 1367 267202
rect -960 267144 1306 267200
rect 1362 267144 1367 267200
rect -960 267142 1367 267144
rect -960 267052 480 267142
rect 1301 267139 1367 267142
rect 582373 260538 582439 260541
rect 580796 260536 582439 260538
rect 580796 260480 582378 260536
rect 582434 260480 582439 260536
rect 580796 260478 582439 260480
rect 582373 260475 582439 260478
rect 582373 258906 582439 258909
rect 583520 258906 584960 258996
rect 582373 258904 584960 258906
rect 582373 258848 582378 258904
rect 582434 258848 584960 258904
rect 582373 258846 584960 258848
rect 582373 258843 582439 258846
rect 583520 258756 584960 258846
rect 1301 256050 1367 256053
rect 1301 256048 3220 256050
rect 1301 255992 1306 256048
rect 1362 255992 3220 256048
rect 1301 255990 3220 255992
rect 1301 255987 1367 255990
rect -960 254146 480 254236
rect 1301 254146 1367 254149
rect -960 254144 1367 254146
rect -960 254088 1306 254144
rect 1362 254088 1367 254144
rect -960 254086 1367 254088
rect -960 253996 480 254086
rect 1301 254083 1367 254086
rect 580766 247074 580826 247452
rect 580901 247074 580967 247077
rect 580766 247072 580967 247074
rect 580766 247016 580906 247072
rect 580962 247016 580967 247072
rect 580766 247014 580967 247016
rect 580901 247011 580967 247014
rect 580901 245578 580967 245581
rect 583520 245578 584960 245668
rect 580901 245576 584960 245578
rect 580901 245520 580906 245576
rect 580962 245520 584960 245576
rect 580901 245518 584960 245520
rect 580901 245515 580967 245518
rect 583520 245428 584960 245518
rect 2773 243266 2839 243269
rect 2773 243264 3220 243266
rect 2773 243208 2778 243264
rect 2834 243208 3220 243264
rect 2773 243206 3220 243208
rect 2773 243203 2839 243206
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 582373 234426 582439 234429
rect 580796 234424 582439 234426
rect 580796 234368 582378 234424
rect 582434 234368 582439 234424
rect 580796 234366 582439 234368
rect 582373 234363 582439 234366
rect 582373 232386 582439 232389
rect 583520 232386 584960 232476
rect 582373 232384 584960 232386
rect 582373 232328 582378 232384
rect 582434 232328 584960 232384
rect 582373 232326 584960 232328
rect 582373 232323 582439 232326
rect 583520 232236 584960 232326
rect 2773 230618 2839 230621
rect 2773 230616 3220 230618
rect 2773 230560 2778 230616
rect 2834 230560 3220 230616
rect 2773 230558 3220 230560
rect 2773 230555 2839 230558
rect -960 228034 480 228124
rect 2773 228034 2839 228037
rect -960 228032 2839 228034
rect -960 227976 2778 228032
rect 2834 227976 2839 228032
rect -960 227974 2839 227976
rect -960 227884 480 227974
rect 2773 227971 2839 227974
rect 580766 220962 580826 221340
rect 580901 220962 580967 220965
rect 580766 220960 580967 220962
rect 580766 220904 580906 220960
rect 580962 220904 580967 220960
rect 580766 220902 580967 220904
rect 580901 220899 580967 220902
rect 580901 219058 580967 219061
rect 583520 219058 584960 219148
rect 580901 219056 584960 219058
rect 580901 219000 580906 219056
rect 580962 219000 584960 219056
rect 580901 218998 584960 219000
rect 580901 218995 580967 218998
rect 583520 218908 584960 218998
rect 2773 217698 2839 217701
rect 2773 217696 3220 217698
rect 2773 217640 2778 217696
rect 2834 217640 3220 217696
rect 2773 217638 3220 217640
rect 2773 217635 2839 217638
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 582373 208314 582439 208317
rect 580796 208312 582439 208314
rect 580796 208256 582378 208312
rect 582434 208256 582439 208312
rect 580796 208254 582439 208256
rect 582373 208251 582439 208254
rect 582373 205730 582439 205733
rect 583520 205730 584960 205820
rect 582373 205728 584960 205730
rect 582373 205672 582378 205728
rect 582434 205672 584960 205728
rect 582373 205670 584960 205672
rect 582373 205667 582439 205670
rect 583520 205580 584960 205670
rect 2773 204914 2839 204917
rect 2773 204912 3220 204914
rect 2773 204856 2778 204912
rect 2834 204856 3220 204912
rect 2773 204854 3220 204856
rect 2773 204851 2839 204854
rect -960 201922 480 202012
rect 2773 201922 2839 201925
rect -960 201920 2839 201922
rect -960 201864 2778 201920
rect 2834 201864 2839 201920
rect -960 201862 2839 201864
rect -960 201772 480 201862
rect 2773 201859 2839 201862
rect 580766 194714 580826 195228
rect 580901 194714 580967 194717
rect 580766 194712 580967 194714
rect 580766 194656 580906 194712
rect 580962 194656 580967 194712
rect 580766 194654 580967 194656
rect 580901 194651 580967 194654
rect 580901 192538 580967 192541
rect 583520 192538 584960 192628
rect 580901 192536 584960 192538
rect 580901 192480 580906 192536
rect 580962 192480 584960 192536
rect 580901 192478 584960 192480
rect 580901 192475 580967 192478
rect 583520 192388 584960 192478
rect 1301 192130 1367 192133
rect 1301 192128 3220 192130
rect 1301 192072 1306 192128
rect 1362 192072 3220 192128
rect 1301 192070 3220 192072
rect 1301 192067 1367 192070
rect -960 188866 480 188956
rect 1301 188866 1367 188869
rect -960 188864 1367 188866
rect -960 188808 1306 188864
rect 1362 188808 1367 188864
rect -960 188806 1367 188808
rect -960 188716 480 188806
rect 1301 188803 1367 188806
rect 580901 182474 580967 182477
rect 580766 182472 580967 182474
rect 580766 182416 580906 182472
rect 580962 182416 580967 182472
rect 580766 182414 580967 182416
rect 580766 182308 580826 182414
rect 580901 182411 580967 182414
rect 2773 179346 2839 179349
rect 2773 179344 3220 179346
rect 2773 179288 2778 179344
rect 2834 179288 3220 179344
rect 2773 179286 3220 179288
rect 2773 179283 2839 179286
rect 580901 179210 580967 179213
rect 583520 179210 584960 179300
rect 580901 179208 584960 179210
rect 580901 179152 580906 179208
rect 580962 179152 584960 179208
rect 580901 179150 584960 179152
rect 580901 179147 580967 179150
rect 583520 179060 584960 179150
rect -960 175946 480 176036
rect 2773 175946 2839 175949
rect -960 175944 2839 175946
rect -960 175888 2778 175944
rect 2834 175888 2839 175944
rect -960 175886 2839 175888
rect -960 175796 480 175886
rect 2773 175883 2839 175886
rect 580766 168602 580826 169116
rect 580901 168602 580967 168605
rect 580766 168600 580967 168602
rect 580766 168544 580906 168600
rect 580962 168544 580967 168600
rect 580766 168542 580967 168544
rect 580901 168539 580967 168542
rect 2773 166562 2839 166565
rect 2773 166560 3220 166562
rect 2773 166504 2778 166560
rect 2834 166504 3220 166560
rect 2773 166502 3220 166504
rect 2773 166499 2839 166502
rect 580901 165882 580967 165885
rect 583520 165882 584960 165972
rect 580901 165880 584960 165882
rect 580901 165824 580906 165880
rect 580962 165824 584960 165880
rect 580901 165822 584960 165824
rect 580901 165819 580967 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 2773 162890 2839 162893
rect -960 162888 2839 162890
rect -960 162832 2778 162888
rect 2834 162832 2839 162888
rect -960 162830 2839 162832
rect -960 162740 480 162830
rect 2773 162827 2839 162830
rect 580901 156362 580967 156365
rect 580766 156360 580967 156362
rect 580766 156304 580906 156360
rect 580962 156304 580967 156360
rect 580766 156302 580967 156304
rect 580766 156196 580826 156302
rect 580901 156299 580967 156302
rect 1301 153778 1367 153781
rect 1301 153776 3220 153778
rect 1301 153720 1306 153776
rect 1362 153720 3220 153776
rect 1301 153718 3220 153720
rect 1301 153715 1367 153718
rect 580901 152690 580967 152693
rect 583520 152690 584960 152780
rect 580901 152688 584960 152690
rect 580901 152632 580906 152688
rect 580962 152632 584960 152688
rect 580901 152630 584960 152632
rect 580901 152627 580967 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 1301 149834 1367 149837
rect -960 149832 1367 149834
rect -960 149776 1306 149832
rect 1362 149776 1367 149832
rect -960 149774 1367 149776
rect -960 149684 480 149774
rect 1301 149771 1367 149774
rect 580766 142626 580826 143004
rect 580901 142626 580967 142629
rect 580766 142624 580967 142626
rect 580766 142568 580906 142624
rect 580962 142568 580967 142624
rect 580766 142566 580967 142568
rect 580901 142563 580967 142566
rect 565 140994 631 140997
rect 565 140992 3220 140994
rect 565 140936 570 140992
rect 626 140936 3220 140992
rect 565 140934 3220 140936
rect 565 140931 631 140934
rect 580901 139362 580967 139365
rect 583520 139362 584960 139452
rect 580901 139360 584960 139362
rect 580901 139304 580906 139360
rect 580962 139304 584960 139360
rect 580901 139302 584960 139304
rect 580901 139299 580967 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 565 136778 631 136781
rect -960 136776 631 136778
rect -960 136720 570 136776
rect 626 136720 631 136776
rect -960 136718 631 136720
rect -960 136628 480 136718
rect 565 136715 631 136718
rect 580901 130250 580967 130253
rect 580766 130248 580967 130250
rect 580766 130192 580906 130248
rect 580962 130192 580967 130248
rect 580766 130190 580967 130192
rect 580766 130084 580826 130190
rect 580901 130187 580967 130190
rect 749 128210 815 128213
rect 749 128208 3220 128210
rect 749 128152 754 128208
rect 810 128152 3220 128208
rect 749 128150 3220 128152
rect 749 128147 815 128150
rect 580901 126034 580967 126037
rect 583520 126034 584960 126124
rect 580901 126032 584960 126034
rect 580901 125976 580906 126032
rect 580962 125976 584960 126032
rect 580901 125974 584960 125976
rect 580901 125971 580967 125974
rect 583520 125884 584960 125974
rect -960 123722 480 123812
rect 749 123722 815 123725
rect -960 123720 815 123722
rect -960 123664 754 123720
rect 810 123664 815 123720
rect -960 123662 815 123664
rect -960 123572 480 123662
rect 749 123659 815 123662
rect 579889 116378 579955 116381
rect 580030 116378 580090 116892
rect 579889 116376 580090 116378
rect 579889 116320 579894 116376
rect 579950 116320 580090 116376
rect 579889 116318 580090 116320
rect 579889 116315 579955 116318
rect 1301 115426 1367 115429
rect 1301 115424 3220 115426
rect 1301 115368 1306 115424
rect 1362 115368 3220 115424
rect 1301 115366 3220 115368
rect 1301 115363 1367 115366
rect 579889 112842 579955 112845
rect 583520 112842 584960 112932
rect 579889 112840 584960 112842
rect 579889 112784 579894 112840
rect 579950 112784 584960 112840
rect 579889 112782 584960 112784
rect 579889 112779 579955 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 1301 110666 1367 110669
rect -960 110664 1367 110666
rect -960 110608 1306 110664
rect 1362 110608 1367 110664
rect -960 110606 1367 110608
rect -960 110516 480 110606
rect 1301 110603 1367 110606
rect 580766 103594 580826 103836
rect 580901 103594 580967 103597
rect 580766 103592 580967 103594
rect 580766 103536 580906 103592
rect 580962 103536 580967 103592
rect 580766 103534 580967 103536
rect 580901 103531 580967 103534
rect 1577 102642 1643 102645
rect 1577 102640 3220 102642
rect 1577 102584 1582 102640
rect 1638 102584 3220 102640
rect 1577 102582 3220 102584
rect 1577 102579 1643 102582
rect 580901 99514 580967 99517
rect 583520 99514 584960 99604
rect 580901 99512 584960 99514
rect 580901 99456 580906 99512
rect 580962 99456 584960 99512
rect 580901 99454 584960 99456
rect 580901 99451 580967 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 1577 97610 1643 97613
rect -960 97608 1643 97610
rect -960 97552 1582 97608
rect 1638 97552 1643 97608
rect -960 97550 1643 97552
rect -960 97460 480 97550
rect 1577 97547 1643 97550
rect 580766 90266 580826 90780
rect 580901 90266 580967 90269
rect 580766 90264 580967 90266
rect 580766 90208 580906 90264
rect 580962 90208 580967 90264
rect 580766 90206 580967 90208
rect 580901 90203 580967 90206
rect 1577 89858 1643 89861
rect 1577 89856 3220 89858
rect 1577 89800 1582 89856
rect 1638 89800 3220 89856
rect 1577 89798 3220 89800
rect 1577 89795 1643 89798
rect 580901 86186 580967 86189
rect 583520 86186 584960 86276
rect 580901 86184 584960 86186
rect 580901 86128 580906 86184
rect 580962 86128 584960 86184
rect 580901 86126 584960 86128
rect 580901 86123 580967 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 1577 84690 1643 84693
rect -960 84688 1643 84690
rect -960 84632 1582 84688
rect 1638 84632 1643 84688
rect -960 84630 1643 84632
rect -960 84540 480 84630
rect 1577 84627 1643 84630
rect 579889 77346 579955 77349
rect 580030 77346 580090 77724
rect 579889 77344 580090 77346
rect 579889 77288 579894 77344
rect 579950 77288 580090 77344
rect 579889 77286 580090 77288
rect 579889 77283 579955 77286
rect 1577 77074 1643 77077
rect 1577 77072 3220 77074
rect 1577 77016 1582 77072
rect 1638 77016 3220 77072
rect 1577 77014 3220 77016
rect 1577 77011 1643 77014
rect 579889 72994 579955 72997
rect 583520 72994 584960 73084
rect 579889 72992 584960 72994
rect 579889 72936 579894 72992
rect 579950 72936 584960 72992
rect 579889 72934 584960 72936
rect 579889 72931 579955 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 1577 71634 1643 71637
rect -960 71632 1643 71634
rect -960 71576 1582 71632
rect 1638 71576 1643 71632
rect -960 71574 1643 71576
rect -960 71484 480 71574
rect 1577 71571 1643 71574
rect 1485 64290 1551 64293
rect 1485 64288 3220 64290
rect 1485 64232 1490 64288
rect 1546 64232 3220 64288
rect 1485 64230 3220 64232
rect 1485 64227 1551 64230
rect 580766 64154 580826 64668
rect 580901 64154 580967 64157
rect 580766 64152 580967 64154
rect 580766 64096 580906 64152
rect 580962 64096 580967 64152
rect 580766 64094 580967 64096
rect 580901 64091 580967 64094
rect 580901 59666 580967 59669
rect 583520 59666 584960 59756
rect 580901 59664 584960 59666
rect 580901 59608 580906 59664
rect 580962 59608 584960 59664
rect 580901 59606 584960 59608
rect 580901 59603 580967 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 1485 58578 1551 58581
rect -960 58576 1551 58578
rect -960 58520 1490 58576
rect 1546 58520 1551 58576
rect -960 58518 1551 58520
rect -960 58428 480 58518
rect 1485 58515 1551 58518
rect 2773 51506 2839 51509
rect 2773 51504 3220 51506
rect 2773 51448 2778 51504
rect 2834 51448 3220 51504
rect 2773 51446 3220 51448
rect 2773 51443 2839 51446
rect 580766 51098 580826 51612
rect 580901 51098 580967 51101
rect 580766 51096 580967 51098
rect 580766 51040 580906 51096
rect 580962 51040 580967 51096
rect 580766 51038 580967 51040
rect 580901 51035 580967 51038
rect 580901 46338 580967 46341
rect 583520 46338 584960 46428
rect 580901 46336 584960 46338
rect 580901 46280 580906 46336
rect 580962 46280 584960 46336
rect 580901 46278 584960 46280
rect 580901 46275 580967 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 2773 45522 2839 45525
rect -960 45520 2839 45522
rect -960 45464 2778 45520
rect 2834 45464 2839 45520
rect -960 45462 2839 45464
rect -960 45372 480 45462
rect 2773 45459 2839 45462
rect 2773 38722 2839 38725
rect 2773 38720 3220 38722
rect 2773 38664 2778 38720
rect 2834 38664 3220 38720
rect 2773 38662 3220 38664
rect 2773 38659 2839 38662
rect 580766 38042 580826 38556
rect 580901 38042 580967 38045
rect 580766 38040 580967 38042
rect 580766 37984 580906 38040
rect 580962 37984 580967 38040
rect 580766 37982 580967 37984
rect 580901 37979 580967 37982
rect 580901 33146 580967 33149
rect 583520 33146 584960 33236
rect 580901 33144 584960 33146
rect 580901 33088 580906 33144
rect 580962 33088 584960 33144
rect 580901 33086 584960 33088
rect 580901 33083 580967 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2773 32466 2839 32469
rect -960 32464 2839 32466
rect -960 32408 2778 32464
rect 2834 32408 2839 32464
rect -960 32406 2839 32408
rect -960 32316 480 32406
rect 2773 32403 2839 32406
rect 1485 25938 1551 25941
rect 1485 25936 3220 25938
rect 1485 25880 1490 25936
rect 1546 25880 3220 25936
rect 1485 25878 3220 25880
rect 1485 25875 1551 25878
rect 580766 24986 580826 25500
rect 580901 24986 580967 24989
rect 580766 24984 580967 24986
rect 580766 24928 580906 24984
rect 580962 24928 580967 24984
rect 580766 24926 580967 24928
rect 580901 24923 580967 24926
rect 580901 19818 580967 19821
rect 583520 19818 584960 19908
rect 580901 19816 584960 19818
rect 580901 19760 580906 19816
rect 580962 19760 584960 19816
rect 580901 19758 584960 19760
rect 580901 19755 580967 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 1485 19410 1551 19413
rect -960 19408 1551 19410
rect -960 19352 1490 19408
rect 1546 19352 1551 19408
rect -960 19350 1551 19352
rect -960 19260 480 19350
rect 1485 19347 1551 19350
rect 2773 13154 2839 13157
rect 2773 13152 3220 13154
rect 2773 13096 2778 13152
rect 2834 13096 3220 13152
rect 2773 13094 3220 13096
rect 2773 13091 2839 13094
rect 579889 12746 579955 12749
rect 579889 12744 580090 12746
rect 579889 12688 579894 12744
rect 579950 12688 580090 12744
rect 579889 12686 580090 12688
rect 579889 12683 579955 12686
rect 580030 12580 580090 12686
rect 579889 6626 579955 6629
rect 583520 6626 584960 6716
rect 579889 6624 584960 6626
rect -960 6490 480 6580
rect 579889 6568 579894 6624
rect 579950 6568 584960 6624
rect 579889 6566 584960 6568
rect 579889 6563 579955 6566
rect 2773 6490 2839 6493
rect -960 6488 2839 6490
rect -960 6432 2778 6488
rect 2834 6432 2839 6488
rect 583520 6476 584960 6566
rect -960 6430 2839 6432
rect -960 6340 480 6430
rect 2773 6427 2839 6430
rect 28901 642 28967 645
rect 46289 642 46355 645
rect 28901 640 46355 642
rect 28901 584 28906 640
rect 28962 584 46294 640
rect 46350 584 46355 640
rect 28901 582 46355 584
rect 28901 579 28967 582
rect 46289 579 46355 582
rect 12157 506 12223 509
rect 30833 506 30899 509
rect 12157 504 30899 506
rect 12157 448 12162 504
rect 12218 448 30838 504
rect 30894 448 30899 504
rect 12157 446 30899 448
rect 12157 443 12223 446
rect 30833 443 30899 446
rect 13721 370 13787 373
rect 31937 370 32003 373
rect 13721 368 32003 370
rect 13721 312 13726 368
rect 13782 312 31942 368
rect 31998 312 32003 368
rect 13721 310 32003 312
rect 13721 307 13787 310
rect 31937 307 32003 310
rect 5441 234 5507 237
rect 23933 234 23999 237
rect 5441 232 23999 234
rect 5441 176 5446 232
rect 5502 176 23938 232
rect 23994 176 23999 232
rect 5441 174 23999 176
rect 5441 171 5507 174
rect 23933 171 23999 174
rect 25681 234 25747 237
rect 42701 234 42767 237
rect 25681 232 42767 234
rect 25681 176 25686 232
rect 25742 176 42706 232
rect 42762 176 42767 232
rect 25681 174 42767 176
rect 25681 171 25747 174
rect 42701 171 42767 174
rect 46841 234 46907 237
rect 62849 234 62915 237
rect 46841 232 62915 234
rect 46841 176 46846 232
rect 46902 176 62854 232
rect 62910 176 62915 232
rect 46841 174 62915 176
rect 46841 171 46907 174
rect 62849 171 62915 174
rect 6269 98 6335 101
rect 25037 98 25103 101
rect 6269 96 25103 98
rect 6269 40 6274 96
rect 6330 40 25042 96
rect 25098 40 25103 96
rect 6269 38 25103 40
rect 6269 35 6335 38
rect 25037 35 25103 38
rect 36997 98 37063 101
rect 54017 98 54083 101
rect 36997 96 54083 98
rect 36997 40 37002 96
rect 37058 40 54022 96
rect 54078 40 54083 96
rect 36997 38 54083 40
rect 36997 35 37063 38
rect 54017 35 54083 38
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 -7066 -8106 711002
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 -6106 -7146 710042
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 -5146 -6186 709082
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 -4186 -5226 708122
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 -3226 -4266 707162
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 -2266 -3306 706202
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 700174 -2346 705242
rect -2966 699938 -2934 700174
rect -2698 699938 -2614 700174
rect -2378 699938 -2346 700174
rect -2966 699854 -2346 699938
rect -2966 699618 -2934 699854
rect -2698 699618 -2614 699854
rect -2378 699618 -2346 699854
rect -2966 664174 -2346 699618
rect -2966 663938 -2934 664174
rect -2698 663938 -2614 664174
rect -2378 663938 -2346 664174
rect -2966 663854 -2346 663938
rect -2966 663618 -2934 663854
rect -2698 663618 -2614 663854
rect -2378 663618 -2346 663854
rect -2966 628174 -2346 663618
rect -2966 627938 -2934 628174
rect -2698 627938 -2614 628174
rect -2378 627938 -2346 628174
rect -2966 627854 -2346 627938
rect -2966 627618 -2934 627854
rect -2698 627618 -2614 627854
rect -2378 627618 -2346 627854
rect -2966 592174 -2346 627618
rect -2966 591938 -2934 592174
rect -2698 591938 -2614 592174
rect -2378 591938 -2346 592174
rect -2966 591854 -2346 591938
rect -2966 591618 -2934 591854
rect -2698 591618 -2614 591854
rect -2378 591618 -2346 591854
rect -2966 556174 -2346 591618
rect -2966 555938 -2934 556174
rect -2698 555938 -2614 556174
rect -2378 555938 -2346 556174
rect -2966 555854 -2346 555938
rect -2966 555618 -2934 555854
rect -2698 555618 -2614 555854
rect -2378 555618 -2346 555854
rect -2966 520174 -2346 555618
rect -2966 519938 -2934 520174
rect -2698 519938 -2614 520174
rect -2378 519938 -2346 520174
rect -2966 519854 -2346 519938
rect -2966 519618 -2934 519854
rect -2698 519618 -2614 519854
rect -2378 519618 -2346 519854
rect -2966 484174 -2346 519618
rect -2966 483938 -2934 484174
rect -2698 483938 -2614 484174
rect -2378 483938 -2346 484174
rect -2966 483854 -2346 483938
rect -2966 483618 -2934 483854
rect -2698 483618 -2614 483854
rect -2378 483618 -2346 483854
rect -2966 448174 -2346 483618
rect -2966 447938 -2934 448174
rect -2698 447938 -2614 448174
rect -2378 447938 -2346 448174
rect -2966 447854 -2346 447938
rect -2966 447618 -2934 447854
rect -2698 447618 -2614 447854
rect -2378 447618 -2346 447854
rect -2966 412174 -2346 447618
rect -2966 411938 -2934 412174
rect -2698 411938 -2614 412174
rect -2378 411938 -2346 412174
rect -2966 411854 -2346 411938
rect -2966 411618 -2934 411854
rect -2698 411618 -2614 411854
rect -2378 411618 -2346 411854
rect -2966 376174 -2346 411618
rect -2966 375938 -2934 376174
rect -2698 375938 -2614 376174
rect -2378 375938 -2346 376174
rect -2966 375854 -2346 375938
rect -2966 375618 -2934 375854
rect -2698 375618 -2614 375854
rect -2378 375618 -2346 375854
rect -2966 340174 -2346 375618
rect -2966 339938 -2934 340174
rect -2698 339938 -2614 340174
rect -2378 339938 -2346 340174
rect -2966 339854 -2346 339938
rect -2966 339618 -2934 339854
rect -2698 339618 -2614 339854
rect -2378 339618 -2346 339854
rect -2966 304174 -2346 339618
rect -2966 303938 -2934 304174
rect -2698 303938 -2614 304174
rect -2378 303938 -2346 304174
rect -2966 303854 -2346 303938
rect -2966 303618 -2934 303854
rect -2698 303618 -2614 303854
rect -2378 303618 -2346 303854
rect -2966 268174 -2346 303618
rect -2966 267938 -2934 268174
rect -2698 267938 -2614 268174
rect -2378 267938 -2346 268174
rect -2966 267854 -2346 267938
rect -2966 267618 -2934 267854
rect -2698 267618 -2614 267854
rect -2378 267618 -2346 267854
rect -2966 232174 -2346 267618
rect -2966 231938 -2934 232174
rect -2698 231938 -2614 232174
rect -2378 231938 -2346 232174
rect -2966 231854 -2346 231938
rect -2966 231618 -2934 231854
rect -2698 231618 -2614 231854
rect -2378 231618 -2346 231854
rect -2966 196174 -2346 231618
rect -2966 195938 -2934 196174
rect -2698 195938 -2614 196174
rect -2378 195938 -2346 196174
rect -2966 195854 -2346 195938
rect -2966 195618 -2934 195854
rect -2698 195618 -2614 195854
rect -2378 195618 -2346 195854
rect -2966 160174 -2346 195618
rect -2966 159938 -2934 160174
rect -2698 159938 -2614 160174
rect -2378 159938 -2346 160174
rect -2966 159854 -2346 159938
rect -2966 159618 -2934 159854
rect -2698 159618 -2614 159854
rect -2378 159618 -2346 159854
rect -2966 124174 -2346 159618
rect -2966 123938 -2934 124174
rect -2698 123938 -2614 124174
rect -2378 123938 -2346 124174
rect -2966 123854 -2346 123938
rect -2966 123618 -2934 123854
rect -2698 123618 -2614 123854
rect -2378 123618 -2346 123854
rect -2966 88174 -2346 123618
rect -2966 87938 -2934 88174
rect -2698 87938 -2614 88174
rect -2378 87938 -2346 88174
rect -2966 87854 -2346 87938
rect -2966 87618 -2934 87854
rect -2698 87618 -2614 87854
rect -2378 87618 -2346 87854
rect -2966 52174 -2346 87618
rect -2966 51938 -2934 52174
rect -2698 51938 -2614 52174
rect -2378 51938 -2346 52174
rect -2966 51854 -2346 51938
rect -2966 51618 -2934 51854
rect -2698 51618 -2614 51854
rect -2378 51618 -2346 51854
rect -2966 16174 -2346 51618
rect -2966 15938 -2934 16174
rect -2698 15938 -2614 16174
rect -2378 15938 -2346 16174
rect -2966 15854 -2346 15938
rect -2966 15618 -2934 15854
rect -2698 15618 -2614 15854
rect -2378 15618 -2346 15854
rect -2966 -1306 -2346 15618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 696454 -1386 704282
rect -2006 696218 -1974 696454
rect -1738 696218 -1654 696454
rect -1418 696218 -1386 696454
rect -2006 696134 -1386 696218
rect -2006 695898 -1974 696134
rect -1738 695898 -1654 696134
rect -1418 695898 -1386 696134
rect -2006 660454 -1386 695898
rect -2006 660218 -1974 660454
rect -1738 660218 -1654 660454
rect -1418 660218 -1386 660454
rect -2006 660134 -1386 660218
rect -2006 659898 -1974 660134
rect -1738 659898 -1654 660134
rect -1418 659898 -1386 660134
rect -2006 624454 -1386 659898
rect -2006 624218 -1974 624454
rect -1738 624218 -1654 624454
rect -1418 624218 -1386 624454
rect -2006 624134 -1386 624218
rect -2006 623898 -1974 624134
rect -1738 623898 -1654 624134
rect -1418 623898 -1386 624134
rect -2006 588454 -1386 623898
rect -2006 588218 -1974 588454
rect -1738 588218 -1654 588454
rect -1418 588218 -1386 588454
rect -2006 588134 -1386 588218
rect -2006 587898 -1974 588134
rect -1738 587898 -1654 588134
rect -1418 587898 -1386 588134
rect -2006 552454 -1386 587898
rect -2006 552218 -1974 552454
rect -1738 552218 -1654 552454
rect -1418 552218 -1386 552454
rect -2006 552134 -1386 552218
rect -2006 551898 -1974 552134
rect -1738 551898 -1654 552134
rect -1418 551898 -1386 552134
rect -2006 516454 -1386 551898
rect -2006 516218 -1974 516454
rect -1738 516218 -1654 516454
rect -1418 516218 -1386 516454
rect -2006 516134 -1386 516218
rect -2006 515898 -1974 516134
rect -1738 515898 -1654 516134
rect -1418 515898 -1386 516134
rect -2006 480454 -1386 515898
rect -2006 480218 -1974 480454
rect -1738 480218 -1654 480454
rect -1418 480218 -1386 480454
rect -2006 480134 -1386 480218
rect -2006 479898 -1974 480134
rect -1738 479898 -1654 480134
rect -1418 479898 -1386 480134
rect -2006 444454 -1386 479898
rect -2006 444218 -1974 444454
rect -1738 444218 -1654 444454
rect -1418 444218 -1386 444454
rect -2006 444134 -1386 444218
rect -2006 443898 -1974 444134
rect -1738 443898 -1654 444134
rect -1418 443898 -1386 444134
rect -2006 408454 -1386 443898
rect -2006 408218 -1974 408454
rect -1738 408218 -1654 408454
rect -1418 408218 -1386 408454
rect -2006 408134 -1386 408218
rect -2006 407898 -1974 408134
rect -1738 407898 -1654 408134
rect -1418 407898 -1386 408134
rect -2006 372454 -1386 407898
rect -2006 372218 -1974 372454
rect -1738 372218 -1654 372454
rect -1418 372218 -1386 372454
rect -2006 372134 -1386 372218
rect -2006 371898 -1974 372134
rect -1738 371898 -1654 372134
rect -1418 371898 -1386 372134
rect -2006 336454 -1386 371898
rect -2006 336218 -1974 336454
rect -1738 336218 -1654 336454
rect -1418 336218 -1386 336454
rect -2006 336134 -1386 336218
rect -2006 335898 -1974 336134
rect -1738 335898 -1654 336134
rect -1418 335898 -1386 336134
rect -2006 300454 -1386 335898
rect -2006 300218 -1974 300454
rect -1738 300218 -1654 300454
rect -1418 300218 -1386 300454
rect -2006 300134 -1386 300218
rect -2006 299898 -1974 300134
rect -1738 299898 -1654 300134
rect -1418 299898 -1386 300134
rect -2006 264454 -1386 299898
rect -2006 264218 -1974 264454
rect -1738 264218 -1654 264454
rect -1418 264218 -1386 264454
rect -2006 264134 -1386 264218
rect -2006 263898 -1974 264134
rect -1738 263898 -1654 264134
rect -1418 263898 -1386 264134
rect -2006 228454 -1386 263898
rect -2006 228218 -1974 228454
rect -1738 228218 -1654 228454
rect -1418 228218 -1386 228454
rect -2006 228134 -1386 228218
rect -2006 227898 -1974 228134
rect -1738 227898 -1654 228134
rect -1418 227898 -1386 228134
rect -2006 192454 -1386 227898
rect -2006 192218 -1974 192454
rect -1738 192218 -1654 192454
rect -1418 192218 -1386 192454
rect -2006 192134 -1386 192218
rect -2006 191898 -1974 192134
rect -1738 191898 -1654 192134
rect -1418 191898 -1386 192134
rect -2006 156454 -1386 191898
rect -2006 156218 -1974 156454
rect -1738 156218 -1654 156454
rect -1418 156218 -1386 156454
rect -2006 156134 -1386 156218
rect -2006 155898 -1974 156134
rect -1738 155898 -1654 156134
rect -1418 155898 -1386 156134
rect -2006 120454 -1386 155898
rect -2006 120218 -1974 120454
rect -1738 120218 -1654 120454
rect -1418 120218 -1386 120454
rect -2006 120134 -1386 120218
rect -2006 119898 -1974 120134
rect -1738 119898 -1654 120134
rect -1418 119898 -1386 120134
rect -2006 84454 -1386 119898
rect -2006 84218 -1974 84454
rect -1738 84218 -1654 84454
rect -1418 84218 -1386 84454
rect -2006 84134 -1386 84218
rect -2006 83898 -1974 84134
rect -1738 83898 -1654 84134
rect -1418 83898 -1386 84134
rect -2006 48454 -1386 83898
rect -2006 48218 -1974 48454
rect -1738 48218 -1654 48454
rect -1418 48218 -1386 48454
rect -2006 48134 -1386 48218
rect -2006 47898 -1974 48134
rect -1738 47898 -1654 48134
rect -1418 47898 -1386 48134
rect -2006 12454 -1386 47898
rect -2006 12218 -1974 12454
rect -1738 12218 -1654 12454
rect -1418 12218 -1386 12454
rect -2006 12134 -1386 12218
rect -2006 11898 -1974 12134
rect -1738 11898 -1654 12134
rect -1418 11898 -1386 12134
rect -2006 -346 -1386 11898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 696454 2414 704282
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 700085 6134 705242
rect 5514 699849 5546 700085
rect 5782 699849 5866 700085
rect 6102 699849 6134 700085
rect 5514 699728 6134 699849
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 700085 42134 705242
rect 41514 699849 41546 700085
rect 41782 699849 41866 700085
rect 42102 699849 42134 700085
rect 41514 699728 42134 699849
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 700085 78134 705242
rect 77514 699849 77546 700085
rect 77782 699849 77866 700085
rect 78102 699849 78134 700085
rect 77514 699728 78134 699849
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 700085 114134 705242
rect 113514 699849 113546 700085
rect 113782 699849 113866 700085
rect 114102 699849 114134 700085
rect 113514 699728 114134 699849
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 700085 150134 705242
rect 149514 699849 149546 700085
rect 149782 699849 149866 700085
rect 150102 699849 150134 700085
rect 149514 699728 150134 699849
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 700085 186134 705242
rect 185514 699849 185546 700085
rect 185782 699849 185866 700085
rect 186102 699849 186134 700085
rect 185514 699728 186134 699849
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 700085 222134 705242
rect 221514 699849 221546 700085
rect 221782 699849 221866 700085
rect 222102 699849 222134 700085
rect 221514 699728 222134 699849
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 700085 258134 705242
rect 257514 699849 257546 700085
rect 257782 699849 257866 700085
rect 258102 699849 258134 700085
rect 257514 699728 258134 699849
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 700085 294134 705242
rect 293514 699849 293546 700085
rect 293782 699849 293866 700085
rect 294102 699849 294134 700085
rect 293514 699728 294134 699849
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 700085 330134 705242
rect 329514 699849 329546 700085
rect 329782 699849 329866 700085
rect 330102 699849 330134 700085
rect 329514 699728 330134 699849
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 700085 366134 705242
rect 365514 699849 365546 700085
rect 365782 699849 365866 700085
rect 366102 699849 366134 700085
rect 365514 699728 366134 699849
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 700085 402134 705242
rect 401514 699849 401546 700085
rect 401782 699849 401866 700085
rect 402102 699849 402134 700085
rect 401514 699728 402134 699849
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 700085 438134 705242
rect 437514 699849 437546 700085
rect 437782 699849 437866 700085
rect 438102 699849 438134 700085
rect 437514 699728 438134 699849
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 700085 474134 705242
rect 473514 699849 473546 700085
rect 473782 699849 473866 700085
rect 474102 699849 474134 700085
rect 473514 699728 474134 699849
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 700085 510134 705242
rect 509514 699849 509546 700085
rect 509782 699849 509866 700085
rect 510102 699849 510134 700085
rect 509514 699728 510134 699849
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 700085 546134 705242
rect 545514 699849 545546 700085
rect 545782 699849 545866 700085
rect 546102 699849 546134 700085
rect 545514 699728 546134 699849
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 696454 578414 704282
rect 1794 696218 1826 696454
rect 2062 696218 2146 696454
rect 2382 696218 2414 696454
rect 1794 696134 2414 696218
rect 1794 695898 1826 696134
rect 2062 695898 2146 696134
rect 2382 695898 2414 696134
rect 5794 696218 5826 696454
rect 6062 696218 6146 696454
rect 6382 696218 6414 696454
rect 5794 696134 6414 696218
rect 5794 695898 5826 696134
rect 6062 695898 6146 696134
rect 6382 695898 6414 696134
rect 41794 696218 41826 696454
rect 42062 696218 42146 696454
rect 42382 696218 42414 696454
rect 41794 696134 42414 696218
rect 41794 695898 41826 696134
rect 42062 695898 42146 696134
rect 42382 695898 42414 696134
rect 77794 696218 77826 696454
rect 78062 696218 78146 696454
rect 78382 696218 78414 696454
rect 77794 696134 78414 696218
rect 77794 695898 77826 696134
rect 78062 695898 78146 696134
rect 78382 695898 78414 696134
rect 113794 696218 113826 696454
rect 114062 696218 114146 696454
rect 114382 696218 114414 696454
rect 113794 696134 114414 696218
rect 113794 695898 113826 696134
rect 114062 695898 114146 696134
rect 114382 695898 114414 696134
rect 149794 696218 149826 696454
rect 150062 696218 150146 696454
rect 150382 696218 150414 696454
rect 149794 696134 150414 696218
rect 149794 695898 149826 696134
rect 150062 695898 150146 696134
rect 150382 695898 150414 696134
rect 185794 696218 185826 696454
rect 186062 696218 186146 696454
rect 186382 696218 186414 696454
rect 185794 696134 186414 696218
rect 185794 695898 185826 696134
rect 186062 695898 186146 696134
rect 186382 695898 186414 696134
rect 221794 696218 221826 696454
rect 222062 696218 222146 696454
rect 222382 696218 222414 696454
rect 221794 696134 222414 696218
rect 221794 695898 221826 696134
rect 222062 695898 222146 696134
rect 222382 695898 222414 696134
rect 257794 696218 257826 696454
rect 258062 696218 258146 696454
rect 258382 696218 258414 696454
rect 257794 696134 258414 696218
rect 257794 695898 257826 696134
rect 258062 695898 258146 696134
rect 258382 695898 258414 696134
rect 293794 696218 293826 696454
rect 294062 696218 294146 696454
rect 294382 696218 294414 696454
rect 293794 696134 294414 696218
rect 293794 695898 293826 696134
rect 294062 695898 294146 696134
rect 294382 695898 294414 696134
rect 329794 696218 329826 696454
rect 330062 696218 330146 696454
rect 330382 696218 330414 696454
rect 329794 696134 330414 696218
rect 329794 695898 329826 696134
rect 330062 695898 330146 696134
rect 330382 695898 330414 696134
rect 365794 696218 365826 696454
rect 366062 696218 366146 696454
rect 366382 696218 366414 696454
rect 365794 696134 366414 696218
rect 365794 695898 365826 696134
rect 366062 695898 366146 696134
rect 366382 695898 366414 696134
rect 401794 696218 401826 696454
rect 402062 696218 402146 696454
rect 402382 696218 402414 696454
rect 401794 696134 402414 696218
rect 401794 695898 401826 696134
rect 402062 695898 402146 696134
rect 402382 695898 402414 696134
rect 437794 696218 437826 696454
rect 438062 696218 438146 696454
rect 438382 696218 438414 696454
rect 437794 696134 438414 696218
rect 437794 695898 437826 696134
rect 438062 695898 438146 696134
rect 438382 695898 438414 696134
rect 473794 696218 473826 696454
rect 474062 696218 474146 696454
rect 474382 696218 474414 696454
rect 473794 696134 474414 696218
rect 473794 695898 473826 696134
rect 474062 695898 474146 696134
rect 474382 695898 474414 696134
rect 509794 696218 509826 696454
rect 510062 696218 510146 696454
rect 510382 696218 510414 696454
rect 509794 696134 510414 696218
rect 509794 695898 509826 696134
rect 510062 695898 510146 696134
rect 510382 695898 510414 696134
rect 545794 696218 545826 696454
rect 546062 696218 546146 696454
rect 546382 696218 546414 696454
rect 545794 696134 546414 696218
rect 545794 695898 545826 696134
rect 546062 695898 546146 696134
rect 546382 695898 546414 696134
rect 577794 696218 577826 696454
rect 578062 696218 578146 696454
rect 578382 696218 578414 696454
rect 577794 696134 578414 696218
rect 577794 695898 577826 696134
rect 578062 695898 578146 696134
rect 578382 695898 578414 696134
rect 1794 660454 2414 695898
rect 9514 663938 9546 664174
rect 9782 663938 9866 664174
rect 10102 663938 10134 664174
rect 9514 663854 10134 663938
rect 9514 663618 9546 663854
rect 9782 663618 9866 663854
rect 10102 663618 10134 663854
rect 189514 663938 189546 664174
rect 189782 663938 189866 664174
rect 190102 663938 190134 664174
rect 189514 663854 190134 663938
rect 189514 663618 189546 663854
rect 189782 663618 189866 663854
rect 190102 663618 190134 663854
rect 369514 663938 369546 664174
rect 369782 663938 369866 664174
rect 370102 663938 370134 664174
rect 369514 663854 370134 663938
rect 369514 663618 369546 663854
rect 369782 663618 369866 663854
rect 370102 663618 370134 663854
rect 405514 663938 405546 664174
rect 405782 663938 405866 664174
rect 406102 663938 406134 664174
rect 405514 663854 406134 663938
rect 405514 663618 405546 663854
rect 405782 663618 405866 663854
rect 406102 663618 406134 663854
rect 572342 663938 572374 664174
rect 572610 663938 572694 664174
rect 572930 663938 572962 664174
rect 572342 663854 572962 663938
rect 572342 663618 572374 663854
rect 572610 663618 572694 663854
rect 572930 663618 572962 663854
rect 577794 660454 578414 695898
rect 1794 660218 1826 660454
rect 2062 660218 2146 660454
rect 2382 660218 2414 660454
rect 1794 660134 2414 660218
rect 1794 659898 1826 660134
rect 2062 659898 2146 660134
rect 2382 659898 2414 660134
rect 5794 660218 5826 660454
rect 6062 660218 6146 660454
rect 6382 660218 6414 660454
rect 5794 660134 6414 660218
rect 5794 659898 5826 660134
rect 6062 659898 6146 660134
rect 6382 659898 6414 660134
rect 185794 660218 185826 660454
rect 186062 660218 186146 660454
rect 186382 660218 186414 660454
rect 185794 660134 186414 660218
rect 185794 659898 185826 660134
rect 186062 659898 186146 660134
rect 186382 659898 186414 660134
rect 365794 660218 365826 660454
rect 366062 660218 366146 660454
rect 366382 660218 366414 660454
rect 365794 660134 366414 660218
rect 365794 659898 365826 660134
rect 366062 659898 366146 660134
rect 366382 659898 366414 660134
rect 401794 660218 401826 660454
rect 402062 660218 402146 660454
rect 402382 660218 402414 660454
rect 401794 660134 402414 660218
rect 401794 659898 401826 660134
rect 402062 659898 402146 660134
rect 402382 659898 402414 660134
rect 568478 660218 568510 660454
rect 568746 660218 568830 660454
rect 569066 660218 569098 660454
rect 568478 660134 569098 660218
rect 568478 659898 568510 660134
rect 568746 659898 568830 660134
rect 569066 659898 569098 660134
rect 577794 660218 577826 660454
rect 578062 660218 578146 660454
rect 578382 660218 578414 660454
rect 577794 660134 578414 660218
rect 577794 659898 577826 660134
rect 578062 659898 578146 660134
rect 578382 659898 578414 660134
rect 1794 624454 2414 659898
rect 9514 627938 9546 628174
rect 9782 627938 9866 628174
rect 10102 627938 10134 628174
rect 9514 627854 10134 627938
rect 9514 627618 9546 627854
rect 9782 627618 9866 627854
rect 10102 627618 10134 627854
rect 189514 627938 189546 628174
rect 189782 627938 189866 628174
rect 190102 627938 190134 628174
rect 189514 627854 190134 627938
rect 189514 627618 189546 627854
rect 189782 627618 189866 627854
rect 190102 627618 190134 627854
rect 369514 627938 369546 628174
rect 369782 627938 369866 628174
rect 370102 627938 370134 628174
rect 369514 627854 370134 627938
rect 369514 627618 369546 627854
rect 369782 627618 369866 627854
rect 370102 627618 370134 627854
rect 405514 627938 405546 628174
rect 405782 627938 405866 628174
rect 406102 627938 406134 628174
rect 405514 627854 406134 627938
rect 405514 627618 405546 627854
rect 405782 627618 405866 627854
rect 406102 627618 406134 627854
rect 572342 627938 572374 628174
rect 572610 627938 572694 628174
rect 572930 627938 572962 628174
rect 572342 627854 572962 627938
rect 572342 627618 572374 627854
rect 572610 627618 572694 627854
rect 572930 627618 572962 627854
rect 577794 624454 578414 659898
rect 1794 624218 1826 624454
rect 2062 624218 2146 624454
rect 2382 624218 2414 624454
rect 1794 624134 2414 624218
rect 1794 623898 1826 624134
rect 2062 623898 2146 624134
rect 2382 623898 2414 624134
rect 5794 624218 5826 624454
rect 6062 624218 6146 624454
rect 6382 624218 6414 624454
rect 5794 624134 6414 624218
rect 5794 623898 5826 624134
rect 6062 623898 6146 624134
rect 6382 623898 6414 624134
rect 185794 624218 185826 624454
rect 186062 624218 186146 624454
rect 186382 624218 186414 624454
rect 185794 624134 186414 624218
rect 185794 623898 185826 624134
rect 186062 623898 186146 624134
rect 186382 623898 186414 624134
rect 365794 624218 365826 624454
rect 366062 624218 366146 624454
rect 366382 624218 366414 624454
rect 365794 624134 366414 624218
rect 365794 623898 365826 624134
rect 366062 623898 366146 624134
rect 366382 623898 366414 624134
rect 401794 624218 401826 624454
rect 402062 624218 402146 624454
rect 402382 624218 402414 624454
rect 401794 624134 402414 624218
rect 401794 623898 401826 624134
rect 402062 623898 402146 624134
rect 402382 623898 402414 624134
rect 568478 624218 568510 624454
rect 568746 624218 568830 624454
rect 569066 624218 569098 624454
rect 568478 624134 569098 624218
rect 568478 623898 568510 624134
rect 568746 623898 568830 624134
rect 569066 623898 569098 624134
rect 577794 624218 577826 624454
rect 578062 624218 578146 624454
rect 578382 624218 578414 624454
rect 577794 624134 578414 624218
rect 577794 623898 577826 624134
rect 578062 623898 578146 624134
rect 578382 623898 578414 624134
rect 1794 588454 2414 623898
rect 9514 591938 9546 592174
rect 9782 591938 9866 592174
rect 10102 591938 10134 592174
rect 9514 591854 10134 591938
rect 9514 591618 9546 591854
rect 9782 591618 9866 591854
rect 10102 591618 10134 591854
rect 45514 591938 45546 592174
rect 45782 591938 45866 592174
rect 46102 591938 46134 592174
rect 45514 591854 46134 591938
rect 45514 591618 45546 591854
rect 45782 591618 45866 591854
rect 46102 591618 46134 591854
rect 81514 591938 81546 592174
rect 81782 591938 81866 592174
rect 82102 591938 82134 592174
rect 81514 591854 82134 591938
rect 81514 591618 81546 591854
rect 81782 591618 81866 591854
rect 82102 591618 82134 591854
rect 117514 591938 117546 592174
rect 117782 591938 117866 592174
rect 118102 591938 118134 592174
rect 117514 591854 118134 591938
rect 117514 591618 117546 591854
rect 117782 591618 117866 591854
rect 118102 591618 118134 591854
rect 153514 591938 153546 592174
rect 153782 591938 153866 592174
rect 154102 591938 154134 592174
rect 153514 591854 154134 591938
rect 153514 591618 153546 591854
rect 153782 591618 153866 591854
rect 154102 591618 154134 591854
rect 189514 591938 189546 592174
rect 189782 591938 189866 592174
rect 190102 591938 190134 592174
rect 189514 591854 190134 591938
rect 189514 591618 189546 591854
rect 189782 591618 189866 591854
rect 190102 591618 190134 591854
rect 225514 591938 225546 592174
rect 225782 591938 225866 592174
rect 226102 591938 226134 592174
rect 225514 591854 226134 591938
rect 225514 591618 225546 591854
rect 225782 591618 225866 591854
rect 226102 591618 226134 591854
rect 261514 591938 261546 592174
rect 261782 591938 261866 592174
rect 262102 591938 262134 592174
rect 261514 591854 262134 591938
rect 261514 591618 261546 591854
rect 261782 591618 261866 591854
rect 262102 591618 262134 591854
rect 297514 591938 297546 592174
rect 297782 591938 297866 592174
rect 298102 591938 298134 592174
rect 297514 591854 298134 591938
rect 297514 591618 297546 591854
rect 297782 591618 297866 591854
rect 298102 591618 298134 591854
rect 333514 591938 333546 592174
rect 333782 591938 333866 592174
rect 334102 591938 334134 592174
rect 333514 591854 334134 591938
rect 333514 591618 333546 591854
rect 333782 591618 333866 591854
rect 334102 591618 334134 591854
rect 369514 591938 369546 592174
rect 369782 591938 369866 592174
rect 370102 591938 370134 592174
rect 369514 591854 370134 591938
rect 369514 591618 369546 591854
rect 369782 591618 369866 591854
rect 370102 591618 370134 591854
rect 405514 591938 405546 592174
rect 405782 591938 405866 592174
rect 406102 591938 406134 592174
rect 405514 591854 406134 591938
rect 405514 591618 405546 591854
rect 405782 591618 405866 591854
rect 406102 591618 406134 591854
rect 441514 591938 441546 592174
rect 441782 591938 441866 592174
rect 442102 591938 442134 592174
rect 441514 591854 442134 591938
rect 441514 591618 441546 591854
rect 441782 591618 441866 591854
rect 442102 591618 442134 591854
rect 477514 591938 477546 592174
rect 477782 591938 477866 592174
rect 478102 591938 478134 592174
rect 477514 591854 478134 591938
rect 477514 591618 477546 591854
rect 477782 591618 477866 591854
rect 478102 591618 478134 591854
rect 513514 591938 513546 592174
rect 513782 591938 513866 592174
rect 514102 591938 514134 592174
rect 513514 591854 514134 591938
rect 513514 591618 513546 591854
rect 513782 591618 513866 591854
rect 514102 591618 514134 591854
rect 549514 591938 549546 592174
rect 549782 591938 549866 592174
rect 550102 591938 550134 592174
rect 549514 591854 550134 591938
rect 549514 591618 549546 591854
rect 549782 591618 549866 591854
rect 550102 591618 550134 591854
rect 577794 588454 578414 623898
rect 1794 588218 1826 588454
rect 2062 588218 2146 588454
rect 2382 588218 2414 588454
rect 1794 588134 2414 588218
rect 1794 587898 1826 588134
rect 2062 587898 2146 588134
rect 2382 587898 2414 588134
rect 5794 588218 5826 588454
rect 6062 588218 6146 588454
rect 6382 588218 6414 588454
rect 5794 588134 6414 588218
rect 5794 587898 5826 588134
rect 6062 587898 6146 588134
rect 6382 587898 6414 588134
rect 41794 588218 41826 588454
rect 42062 588218 42146 588454
rect 42382 588218 42414 588454
rect 41794 588134 42414 588218
rect 41794 587898 41826 588134
rect 42062 587898 42146 588134
rect 42382 587898 42414 588134
rect 77794 588218 77826 588454
rect 78062 588218 78146 588454
rect 78382 588218 78414 588454
rect 77794 588134 78414 588218
rect 77794 587898 77826 588134
rect 78062 587898 78146 588134
rect 78382 587898 78414 588134
rect 113794 588218 113826 588454
rect 114062 588218 114146 588454
rect 114382 588218 114414 588454
rect 113794 588134 114414 588218
rect 113794 587898 113826 588134
rect 114062 587898 114146 588134
rect 114382 587898 114414 588134
rect 149794 588218 149826 588454
rect 150062 588218 150146 588454
rect 150382 588218 150414 588454
rect 149794 588134 150414 588218
rect 149794 587898 149826 588134
rect 150062 587898 150146 588134
rect 150382 587898 150414 588134
rect 185794 588218 185826 588454
rect 186062 588218 186146 588454
rect 186382 588218 186414 588454
rect 185794 588134 186414 588218
rect 185794 587898 185826 588134
rect 186062 587898 186146 588134
rect 186382 587898 186414 588134
rect 221794 588218 221826 588454
rect 222062 588218 222146 588454
rect 222382 588218 222414 588454
rect 221794 588134 222414 588218
rect 221794 587898 221826 588134
rect 222062 587898 222146 588134
rect 222382 587898 222414 588134
rect 257794 588218 257826 588454
rect 258062 588218 258146 588454
rect 258382 588218 258414 588454
rect 257794 588134 258414 588218
rect 257794 587898 257826 588134
rect 258062 587898 258146 588134
rect 258382 587898 258414 588134
rect 293794 588218 293826 588454
rect 294062 588218 294146 588454
rect 294382 588218 294414 588454
rect 293794 588134 294414 588218
rect 293794 587898 293826 588134
rect 294062 587898 294146 588134
rect 294382 587898 294414 588134
rect 329794 588218 329826 588454
rect 330062 588218 330146 588454
rect 330382 588218 330414 588454
rect 329794 588134 330414 588218
rect 329794 587898 329826 588134
rect 330062 587898 330146 588134
rect 330382 587898 330414 588134
rect 365794 588218 365826 588454
rect 366062 588218 366146 588454
rect 366382 588218 366414 588454
rect 365794 588134 366414 588218
rect 365794 587898 365826 588134
rect 366062 587898 366146 588134
rect 366382 587898 366414 588134
rect 401794 588218 401826 588454
rect 402062 588218 402146 588454
rect 402382 588218 402414 588454
rect 401794 588134 402414 588218
rect 401794 587898 401826 588134
rect 402062 587898 402146 588134
rect 402382 587898 402414 588134
rect 437794 588218 437826 588454
rect 438062 588218 438146 588454
rect 438382 588218 438414 588454
rect 437794 588134 438414 588218
rect 437794 587898 437826 588134
rect 438062 587898 438146 588134
rect 438382 587898 438414 588134
rect 473794 588218 473826 588454
rect 474062 588218 474146 588454
rect 474382 588218 474414 588454
rect 473794 588134 474414 588218
rect 473794 587898 473826 588134
rect 474062 587898 474146 588134
rect 474382 587898 474414 588134
rect 509794 588218 509826 588454
rect 510062 588218 510146 588454
rect 510382 588218 510414 588454
rect 509794 588134 510414 588218
rect 509794 587898 509826 588134
rect 510062 587898 510146 588134
rect 510382 587898 510414 588134
rect 545794 588218 545826 588454
rect 546062 588218 546146 588454
rect 546382 588218 546414 588454
rect 545794 588134 546414 588218
rect 545794 587898 545826 588134
rect 546062 587898 546146 588134
rect 546382 587898 546414 588134
rect 577794 588218 577826 588454
rect 578062 588218 578146 588454
rect 578382 588218 578414 588454
rect 577794 588134 578414 588218
rect 577794 587898 577826 588134
rect 578062 587898 578146 588134
rect 578382 587898 578414 588134
rect 1794 552454 2414 587898
rect 9514 555938 9546 556174
rect 9782 555938 9866 556174
rect 10102 555938 10134 556174
rect 9514 555854 10134 555938
rect 9514 555618 9546 555854
rect 9782 555618 9866 555854
rect 10102 555618 10134 555854
rect 189514 555938 189546 556174
rect 189782 555938 189866 556174
rect 190102 555938 190134 556174
rect 189514 555854 190134 555938
rect 189514 555618 189546 555854
rect 189782 555618 189866 555854
rect 190102 555618 190134 555854
rect 225514 555938 225546 556174
rect 225782 555938 225866 556174
rect 226102 555938 226134 556174
rect 225514 555854 226134 555938
rect 225514 555618 225546 555854
rect 225782 555618 225866 555854
rect 226102 555618 226134 555854
rect 261514 555938 261546 556174
rect 261782 555938 261866 556174
rect 262102 555938 262134 556174
rect 261514 555854 262134 555938
rect 261514 555618 261546 555854
rect 261782 555618 261866 555854
rect 262102 555618 262134 555854
rect 297514 555938 297546 556174
rect 297782 555938 297866 556174
rect 298102 555938 298134 556174
rect 297514 555854 298134 555938
rect 297514 555618 297546 555854
rect 297782 555618 297866 555854
rect 298102 555618 298134 555854
rect 333514 555938 333546 556174
rect 333782 555938 333866 556174
rect 334102 555938 334134 556174
rect 333514 555854 334134 555938
rect 333514 555618 333546 555854
rect 333782 555618 333866 555854
rect 334102 555618 334134 555854
rect 369514 555938 369546 556174
rect 369782 555938 369866 556174
rect 370102 555938 370134 556174
rect 369514 555854 370134 555938
rect 369514 555618 369546 555854
rect 369782 555618 369866 555854
rect 370102 555618 370134 555854
rect 405514 555938 405546 556174
rect 405782 555938 405866 556174
rect 406102 555938 406134 556174
rect 405514 555854 406134 555938
rect 405514 555618 405546 555854
rect 405782 555618 405866 555854
rect 406102 555618 406134 555854
rect 572342 555938 572374 556174
rect 572610 555938 572694 556174
rect 572930 555938 572962 556174
rect 572342 555854 572962 555938
rect 572342 555618 572374 555854
rect 572610 555618 572694 555854
rect 572930 555618 572962 555854
rect 577794 552454 578414 587898
rect 1794 552218 1826 552454
rect 2062 552218 2146 552454
rect 2382 552218 2414 552454
rect 1794 552134 2414 552218
rect 1794 551898 1826 552134
rect 2062 551898 2146 552134
rect 2382 551898 2414 552134
rect 5794 552218 5826 552454
rect 6062 552218 6146 552454
rect 6382 552218 6414 552454
rect 5794 552134 6414 552218
rect 5794 551898 5826 552134
rect 6062 551898 6146 552134
rect 6382 551898 6414 552134
rect 185794 552218 185826 552454
rect 186062 552218 186146 552454
rect 186382 552218 186414 552454
rect 185794 552134 186414 552218
rect 185794 551898 185826 552134
rect 186062 551898 186146 552134
rect 186382 551898 186414 552134
rect 221794 552218 221826 552454
rect 222062 552218 222146 552454
rect 222382 552218 222414 552454
rect 221794 552134 222414 552218
rect 221794 551898 221826 552134
rect 222062 551898 222146 552134
rect 222382 551898 222414 552134
rect 257794 552218 257826 552454
rect 258062 552218 258146 552454
rect 258382 552218 258414 552454
rect 257794 552134 258414 552218
rect 257794 551898 257826 552134
rect 258062 551898 258146 552134
rect 258382 551898 258414 552134
rect 293794 552218 293826 552454
rect 294062 552218 294146 552454
rect 294382 552218 294414 552454
rect 293794 552134 294414 552218
rect 293794 551898 293826 552134
rect 294062 551898 294146 552134
rect 294382 551898 294414 552134
rect 329794 552218 329826 552454
rect 330062 552218 330146 552454
rect 330382 552218 330414 552454
rect 329794 552134 330414 552218
rect 329794 551898 329826 552134
rect 330062 551898 330146 552134
rect 330382 551898 330414 552134
rect 365794 552218 365826 552454
rect 366062 552218 366146 552454
rect 366382 552218 366414 552454
rect 365794 552134 366414 552218
rect 365794 551898 365826 552134
rect 366062 551898 366146 552134
rect 366382 551898 366414 552134
rect 401794 552218 401826 552454
rect 402062 552218 402146 552454
rect 402382 552218 402414 552454
rect 401794 552134 402414 552218
rect 401794 551898 401826 552134
rect 402062 551898 402146 552134
rect 402382 551898 402414 552134
rect 568478 552218 568510 552454
rect 568746 552218 568830 552454
rect 569066 552218 569098 552454
rect 568478 552134 569098 552218
rect 568478 551898 568510 552134
rect 568746 551898 568830 552134
rect 569066 551898 569098 552134
rect 577794 552218 577826 552454
rect 578062 552218 578146 552454
rect 578382 552218 578414 552454
rect 577794 552134 578414 552218
rect 577794 551898 577826 552134
rect 578062 551898 578146 552134
rect 578382 551898 578414 552134
rect 1794 516454 2414 551898
rect 9514 519938 9546 520174
rect 9782 519938 9866 520174
rect 10102 519938 10134 520174
rect 9514 519854 10134 519938
rect 9514 519618 9546 519854
rect 9782 519618 9866 519854
rect 10102 519618 10134 519854
rect 189514 519938 189546 520174
rect 189782 519938 189866 520174
rect 190102 519938 190134 520174
rect 189514 519854 190134 519938
rect 189514 519618 189546 519854
rect 189782 519618 189866 519854
rect 190102 519618 190134 519854
rect 225514 519938 225546 520174
rect 225782 519938 225866 520174
rect 226102 519938 226134 520174
rect 225514 519854 226134 519938
rect 225514 519618 225546 519854
rect 225782 519618 225866 519854
rect 226102 519618 226134 519854
rect 261514 519938 261546 520174
rect 261782 519938 261866 520174
rect 262102 519938 262134 520174
rect 261514 519854 262134 519938
rect 261514 519618 261546 519854
rect 261782 519618 261866 519854
rect 262102 519618 262134 519854
rect 297514 519938 297546 520174
rect 297782 519938 297866 520174
rect 298102 519938 298134 520174
rect 297514 519854 298134 519938
rect 297514 519618 297546 519854
rect 297782 519618 297866 519854
rect 298102 519618 298134 519854
rect 333514 519938 333546 520174
rect 333782 519938 333866 520174
rect 334102 519938 334134 520174
rect 333514 519854 334134 519938
rect 333514 519618 333546 519854
rect 333782 519618 333866 519854
rect 334102 519618 334134 519854
rect 369514 519938 369546 520174
rect 369782 519938 369866 520174
rect 370102 519938 370134 520174
rect 369514 519854 370134 519938
rect 369514 519618 369546 519854
rect 369782 519618 369866 519854
rect 370102 519618 370134 519854
rect 405514 519938 405546 520174
rect 405782 519938 405866 520174
rect 406102 519938 406134 520174
rect 405514 519854 406134 519938
rect 405514 519618 405546 519854
rect 405782 519618 405866 519854
rect 406102 519618 406134 519854
rect 572342 519938 572374 520174
rect 572610 519938 572694 520174
rect 572930 519938 572962 520174
rect 572342 519854 572962 519938
rect 572342 519618 572374 519854
rect 572610 519618 572694 519854
rect 572930 519618 572962 519854
rect 577794 516454 578414 551898
rect 1794 516218 1826 516454
rect 2062 516218 2146 516454
rect 2382 516218 2414 516454
rect 1794 516134 2414 516218
rect 1794 515898 1826 516134
rect 2062 515898 2146 516134
rect 2382 515898 2414 516134
rect 5794 516218 5826 516454
rect 6062 516218 6146 516454
rect 6382 516218 6414 516454
rect 5794 516134 6414 516218
rect 5794 515898 5826 516134
rect 6062 515898 6146 516134
rect 6382 515898 6414 516134
rect 185794 516218 185826 516454
rect 186062 516218 186146 516454
rect 186382 516218 186414 516454
rect 185794 516134 186414 516218
rect 185794 515898 185826 516134
rect 186062 515898 186146 516134
rect 186382 515898 186414 516134
rect 221794 516218 221826 516454
rect 222062 516218 222146 516454
rect 222382 516218 222414 516454
rect 221794 516134 222414 516218
rect 221794 515898 221826 516134
rect 222062 515898 222146 516134
rect 222382 515898 222414 516134
rect 257794 516218 257826 516454
rect 258062 516218 258146 516454
rect 258382 516218 258414 516454
rect 257794 516134 258414 516218
rect 257794 515898 257826 516134
rect 258062 515898 258146 516134
rect 258382 515898 258414 516134
rect 293794 516218 293826 516454
rect 294062 516218 294146 516454
rect 294382 516218 294414 516454
rect 293794 516134 294414 516218
rect 293794 515898 293826 516134
rect 294062 515898 294146 516134
rect 294382 515898 294414 516134
rect 329794 516218 329826 516454
rect 330062 516218 330146 516454
rect 330382 516218 330414 516454
rect 329794 516134 330414 516218
rect 329794 515898 329826 516134
rect 330062 515898 330146 516134
rect 330382 515898 330414 516134
rect 365794 516218 365826 516454
rect 366062 516218 366146 516454
rect 366382 516218 366414 516454
rect 365794 516134 366414 516218
rect 365794 515898 365826 516134
rect 366062 515898 366146 516134
rect 366382 515898 366414 516134
rect 401794 516218 401826 516454
rect 402062 516218 402146 516454
rect 402382 516218 402414 516454
rect 401794 516134 402414 516218
rect 401794 515898 401826 516134
rect 402062 515898 402146 516134
rect 402382 515898 402414 516134
rect 568478 516218 568510 516454
rect 568746 516218 568830 516454
rect 569066 516218 569098 516454
rect 568478 516134 569098 516218
rect 568478 515898 568510 516134
rect 568746 515898 568830 516134
rect 569066 515898 569098 516134
rect 577794 516218 577826 516454
rect 578062 516218 578146 516454
rect 578382 516218 578414 516454
rect 577794 516134 578414 516218
rect 577794 515898 577826 516134
rect 578062 515898 578146 516134
rect 578382 515898 578414 516134
rect 1794 480454 2414 515898
rect 9514 483938 9546 484174
rect 9782 483938 9866 484174
rect 10102 483938 10134 484174
rect 9514 483854 10134 483938
rect 9514 483618 9546 483854
rect 9782 483618 9866 483854
rect 10102 483618 10134 483854
rect 45514 483938 45546 484174
rect 45782 483938 45866 484174
rect 46102 483938 46134 484174
rect 45514 483854 46134 483938
rect 45514 483618 45546 483854
rect 45782 483618 45866 483854
rect 46102 483618 46134 483854
rect 81514 483938 81546 484174
rect 81782 483938 81866 484174
rect 82102 483938 82134 484174
rect 81514 483854 82134 483938
rect 81514 483618 81546 483854
rect 81782 483618 81866 483854
rect 82102 483618 82134 483854
rect 117514 483938 117546 484174
rect 117782 483938 117866 484174
rect 118102 483938 118134 484174
rect 117514 483854 118134 483938
rect 117514 483618 117546 483854
rect 117782 483618 117866 483854
rect 118102 483618 118134 483854
rect 153514 483938 153546 484174
rect 153782 483938 153866 484174
rect 154102 483938 154134 484174
rect 153514 483854 154134 483938
rect 153514 483618 153546 483854
rect 153782 483618 153866 483854
rect 154102 483618 154134 483854
rect 189514 483938 189546 484174
rect 189782 483938 189866 484174
rect 190102 483938 190134 484174
rect 189514 483854 190134 483938
rect 189514 483618 189546 483854
rect 189782 483618 189866 483854
rect 190102 483618 190134 483854
rect 225514 483938 225546 484174
rect 225782 483938 225866 484174
rect 226102 483938 226134 484174
rect 225514 483854 226134 483938
rect 225514 483618 225546 483854
rect 225782 483618 225866 483854
rect 226102 483618 226134 483854
rect 261514 483938 261546 484174
rect 261782 483938 261866 484174
rect 262102 483938 262134 484174
rect 261514 483854 262134 483938
rect 261514 483618 261546 483854
rect 261782 483618 261866 483854
rect 262102 483618 262134 483854
rect 297514 483938 297546 484174
rect 297782 483938 297866 484174
rect 298102 483938 298134 484174
rect 297514 483854 298134 483938
rect 297514 483618 297546 483854
rect 297782 483618 297866 483854
rect 298102 483618 298134 483854
rect 333514 483938 333546 484174
rect 333782 483938 333866 484174
rect 334102 483938 334134 484174
rect 333514 483854 334134 483938
rect 333514 483618 333546 483854
rect 333782 483618 333866 483854
rect 334102 483618 334134 483854
rect 369514 483938 369546 484174
rect 369782 483938 369866 484174
rect 370102 483938 370134 484174
rect 369514 483854 370134 483938
rect 369514 483618 369546 483854
rect 369782 483618 369866 483854
rect 370102 483618 370134 483854
rect 405514 483938 405546 484174
rect 405782 483938 405866 484174
rect 406102 483938 406134 484174
rect 405514 483854 406134 483938
rect 405514 483618 405546 483854
rect 405782 483618 405866 483854
rect 406102 483618 406134 483854
rect 441514 483938 441546 484174
rect 441782 483938 441866 484174
rect 442102 483938 442134 484174
rect 441514 483854 442134 483938
rect 441514 483618 441546 483854
rect 441782 483618 441866 483854
rect 442102 483618 442134 483854
rect 477514 483938 477546 484174
rect 477782 483938 477866 484174
rect 478102 483938 478134 484174
rect 477514 483854 478134 483938
rect 477514 483618 477546 483854
rect 477782 483618 477866 483854
rect 478102 483618 478134 483854
rect 513514 483938 513546 484174
rect 513782 483938 513866 484174
rect 514102 483938 514134 484174
rect 513514 483854 514134 483938
rect 513514 483618 513546 483854
rect 513782 483618 513866 483854
rect 514102 483618 514134 483854
rect 549514 483938 549546 484174
rect 549782 483938 549866 484174
rect 550102 483938 550134 484174
rect 549514 483854 550134 483938
rect 549514 483618 549546 483854
rect 549782 483618 549866 483854
rect 550102 483618 550134 483854
rect 577794 480454 578414 515898
rect 1794 480218 1826 480454
rect 2062 480218 2146 480454
rect 2382 480218 2414 480454
rect 1794 480134 2414 480218
rect 1794 479898 1826 480134
rect 2062 479898 2146 480134
rect 2382 479898 2414 480134
rect 5794 480218 5826 480454
rect 6062 480218 6146 480454
rect 6382 480218 6414 480454
rect 5794 480134 6414 480218
rect 5794 479898 5826 480134
rect 6062 479898 6146 480134
rect 6382 479898 6414 480134
rect 41794 480218 41826 480454
rect 42062 480218 42146 480454
rect 42382 480218 42414 480454
rect 41794 480134 42414 480218
rect 41794 479898 41826 480134
rect 42062 479898 42146 480134
rect 42382 479898 42414 480134
rect 77794 480218 77826 480454
rect 78062 480218 78146 480454
rect 78382 480218 78414 480454
rect 77794 480134 78414 480218
rect 77794 479898 77826 480134
rect 78062 479898 78146 480134
rect 78382 479898 78414 480134
rect 113794 480218 113826 480454
rect 114062 480218 114146 480454
rect 114382 480218 114414 480454
rect 113794 480134 114414 480218
rect 113794 479898 113826 480134
rect 114062 479898 114146 480134
rect 114382 479898 114414 480134
rect 149794 480218 149826 480454
rect 150062 480218 150146 480454
rect 150382 480218 150414 480454
rect 149794 480134 150414 480218
rect 149794 479898 149826 480134
rect 150062 479898 150146 480134
rect 150382 479898 150414 480134
rect 185794 480218 185826 480454
rect 186062 480218 186146 480454
rect 186382 480218 186414 480454
rect 185794 480134 186414 480218
rect 185794 479898 185826 480134
rect 186062 479898 186146 480134
rect 186382 479898 186414 480134
rect 221794 480218 221826 480454
rect 222062 480218 222146 480454
rect 222382 480218 222414 480454
rect 221794 480134 222414 480218
rect 221794 479898 221826 480134
rect 222062 479898 222146 480134
rect 222382 479898 222414 480134
rect 257794 480218 257826 480454
rect 258062 480218 258146 480454
rect 258382 480218 258414 480454
rect 257794 480134 258414 480218
rect 257794 479898 257826 480134
rect 258062 479898 258146 480134
rect 258382 479898 258414 480134
rect 293794 480218 293826 480454
rect 294062 480218 294146 480454
rect 294382 480218 294414 480454
rect 293794 480134 294414 480218
rect 293794 479898 293826 480134
rect 294062 479898 294146 480134
rect 294382 479898 294414 480134
rect 329794 480218 329826 480454
rect 330062 480218 330146 480454
rect 330382 480218 330414 480454
rect 329794 480134 330414 480218
rect 329794 479898 329826 480134
rect 330062 479898 330146 480134
rect 330382 479898 330414 480134
rect 365794 480218 365826 480454
rect 366062 480218 366146 480454
rect 366382 480218 366414 480454
rect 365794 480134 366414 480218
rect 365794 479898 365826 480134
rect 366062 479898 366146 480134
rect 366382 479898 366414 480134
rect 401794 480218 401826 480454
rect 402062 480218 402146 480454
rect 402382 480218 402414 480454
rect 401794 480134 402414 480218
rect 401794 479898 401826 480134
rect 402062 479898 402146 480134
rect 402382 479898 402414 480134
rect 437794 480218 437826 480454
rect 438062 480218 438146 480454
rect 438382 480218 438414 480454
rect 437794 480134 438414 480218
rect 437794 479898 437826 480134
rect 438062 479898 438146 480134
rect 438382 479898 438414 480134
rect 473794 480218 473826 480454
rect 474062 480218 474146 480454
rect 474382 480218 474414 480454
rect 473794 480134 474414 480218
rect 473794 479898 473826 480134
rect 474062 479898 474146 480134
rect 474382 479898 474414 480134
rect 509794 480218 509826 480454
rect 510062 480218 510146 480454
rect 510382 480218 510414 480454
rect 509794 480134 510414 480218
rect 509794 479898 509826 480134
rect 510062 479898 510146 480134
rect 510382 479898 510414 480134
rect 545794 480218 545826 480454
rect 546062 480218 546146 480454
rect 546382 480218 546414 480454
rect 545794 480134 546414 480218
rect 545794 479898 545826 480134
rect 546062 479898 546146 480134
rect 546382 479898 546414 480134
rect 577794 480218 577826 480454
rect 578062 480218 578146 480454
rect 578382 480218 578414 480454
rect 577794 480134 578414 480218
rect 577794 479898 577826 480134
rect 578062 479898 578146 480134
rect 578382 479898 578414 480134
rect 1794 444454 2414 479898
rect 9514 447938 9546 448174
rect 9782 447938 9866 448174
rect 10102 447938 10134 448174
rect 9514 447854 10134 447938
rect 9514 447618 9546 447854
rect 9782 447618 9866 447854
rect 10102 447618 10134 447854
rect 189514 447938 189546 448174
rect 189782 447938 189866 448174
rect 190102 447938 190134 448174
rect 189514 447854 190134 447938
rect 189514 447618 189546 447854
rect 189782 447618 189866 447854
rect 190102 447618 190134 447854
rect 225514 447938 225546 448174
rect 225782 447938 225866 448174
rect 226102 447938 226134 448174
rect 225514 447854 226134 447938
rect 225514 447618 225546 447854
rect 225782 447618 225866 447854
rect 226102 447618 226134 447854
rect 261514 447938 261546 448174
rect 261782 447938 261866 448174
rect 262102 447938 262134 448174
rect 261514 447854 262134 447938
rect 261514 447618 261546 447854
rect 261782 447618 261866 447854
rect 262102 447618 262134 447854
rect 297514 447938 297546 448174
rect 297782 447938 297866 448174
rect 298102 447938 298134 448174
rect 297514 447854 298134 447938
rect 297514 447618 297546 447854
rect 297782 447618 297866 447854
rect 298102 447618 298134 447854
rect 333514 447938 333546 448174
rect 333782 447938 333866 448174
rect 334102 447938 334134 448174
rect 333514 447854 334134 447938
rect 333514 447618 333546 447854
rect 333782 447618 333866 447854
rect 334102 447618 334134 447854
rect 369514 447938 369546 448174
rect 369782 447938 369866 448174
rect 370102 447938 370134 448174
rect 369514 447854 370134 447938
rect 369514 447618 369546 447854
rect 369782 447618 369866 447854
rect 370102 447618 370134 447854
rect 405514 447938 405546 448174
rect 405782 447938 405866 448174
rect 406102 447938 406134 448174
rect 405514 447854 406134 447938
rect 405514 447618 405546 447854
rect 405782 447618 405866 447854
rect 406102 447618 406134 447854
rect 572342 447938 572374 448174
rect 572610 447938 572694 448174
rect 572930 447938 572962 448174
rect 572342 447854 572962 447938
rect 572342 447618 572374 447854
rect 572610 447618 572694 447854
rect 572930 447618 572962 447854
rect 577794 444454 578414 479898
rect 1794 444218 1826 444454
rect 2062 444218 2146 444454
rect 2382 444218 2414 444454
rect 1794 444134 2414 444218
rect 1794 443898 1826 444134
rect 2062 443898 2146 444134
rect 2382 443898 2414 444134
rect 5794 444218 5826 444454
rect 6062 444218 6146 444454
rect 6382 444218 6414 444454
rect 5794 444134 6414 444218
rect 5794 443898 5826 444134
rect 6062 443898 6146 444134
rect 6382 443898 6414 444134
rect 185794 444218 185826 444454
rect 186062 444218 186146 444454
rect 186382 444218 186414 444454
rect 185794 444134 186414 444218
rect 185794 443898 185826 444134
rect 186062 443898 186146 444134
rect 186382 443898 186414 444134
rect 221794 444218 221826 444454
rect 222062 444218 222146 444454
rect 222382 444218 222414 444454
rect 221794 444134 222414 444218
rect 221794 443898 221826 444134
rect 222062 443898 222146 444134
rect 222382 443898 222414 444134
rect 257794 444218 257826 444454
rect 258062 444218 258146 444454
rect 258382 444218 258414 444454
rect 257794 444134 258414 444218
rect 257794 443898 257826 444134
rect 258062 443898 258146 444134
rect 258382 443898 258414 444134
rect 293794 444218 293826 444454
rect 294062 444218 294146 444454
rect 294382 444218 294414 444454
rect 293794 444134 294414 444218
rect 293794 443898 293826 444134
rect 294062 443898 294146 444134
rect 294382 443898 294414 444134
rect 329794 444218 329826 444454
rect 330062 444218 330146 444454
rect 330382 444218 330414 444454
rect 329794 444134 330414 444218
rect 329794 443898 329826 444134
rect 330062 443898 330146 444134
rect 330382 443898 330414 444134
rect 365794 444218 365826 444454
rect 366062 444218 366146 444454
rect 366382 444218 366414 444454
rect 365794 444134 366414 444218
rect 365794 443898 365826 444134
rect 366062 443898 366146 444134
rect 366382 443898 366414 444134
rect 401794 444218 401826 444454
rect 402062 444218 402146 444454
rect 402382 444218 402414 444454
rect 401794 444134 402414 444218
rect 401794 443898 401826 444134
rect 402062 443898 402146 444134
rect 402382 443898 402414 444134
rect 568478 444218 568510 444454
rect 568746 444218 568830 444454
rect 569066 444218 569098 444454
rect 568478 444134 569098 444218
rect 568478 443898 568510 444134
rect 568746 443898 568830 444134
rect 569066 443898 569098 444134
rect 577794 444218 577826 444454
rect 578062 444218 578146 444454
rect 578382 444218 578414 444454
rect 577794 444134 578414 444218
rect 577794 443898 577826 444134
rect 578062 443898 578146 444134
rect 578382 443898 578414 444134
rect 1794 408454 2414 443898
rect 9514 411938 9546 412174
rect 9782 411938 9866 412174
rect 10102 411938 10134 412174
rect 9514 411854 10134 411938
rect 9514 411618 9546 411854
rect 9782 411618 9866 411854
rect 10102 411618 10134 411854
rect 189514 411938 189546 412174
rect 189782 411938 189866 412174
rect 190102 411938 190134 412174
rect 189514 411854 190134 411938
rect 189514 411618 189546 411854
rect 189782 411618 189866 411854
rect 190102 411618 190134 411854
rect 225514 411938 225546 412174
rect 225782 411938 225866 412174
rect 226102 411938 226134 412174
rect 225514 411854 226134 411938
rect 225514 411618 225546 411854
rect 225782 411618 225866 411854
rect 226102 411618 226134 411854
rect 261514 411938 261546 412174
rect 261782 411938 261866 412174
rect 262102 411938 262134 412174
rect 261514 411854 262134 411938
rect 261514 411618 261546 411854
rect 261782 411618 261866 411854
rect 262102 411618 262134 411854
rect 297514 411938 297546 412174
rect 297782 411938 297866 412174
rect 298102 411938 298134 412174
rect 297514 411854 298134 411938
rect 297514 411618 297546 411854
rect 297782 411618 297866 411854
rect 298102 411618 298134 411854
rect 333514 411938 333546 412174
rect 333782 411938 333866 412174
rect 334102 411938 334134 412174
rect 333514 411854 334134 411938
rect 333514 411618 333546 411854
rect 333782 411618 333866 411854
rect 334102 411618 334134 411854
rect 369514 411938 369546 412174
rect 369782 411938 369866 412174
rect 370102 411938 370134 412174
rect 369514 411854 370134 411938
rect 369514 411618 369546 411854
rect 369782 411618 369866 411854
rect 370102 411618 370134 411854
rect 405514 411938 405546 412174
rect 405782 411938 405866 412174
rect 406102 411938 406134 412174
rect 405514 411854 406134 411938
rect 405514 411618 405546 411854
rect 405782 411618 405866 411854
rect 406102 411618 406134 411854
rect 572342 411938 572374 412174
rect 572610 411938 572694 412174
rect 572930 411938 572962 412174
rect 572342 411854 572962 411938
rect 572342 411618 572374 411854
rect 572610 411618 572694 411854
rect 572930 411618 572962 411854
rect 577794 408454 578414 443898
rect 1794 408218 1826 408454
rect 2062 408218 2146 408454
rect 2382 408218 2414 408454
rect 1794 408134 2414 408218
rect 1794 407898 1826 408134
rect 2062 407898 2146 408134
rect 2382 407898 2414 408134
rect 5794 408218 5826 408454
rect 6062 408218 6146 408454
rect 6382 408218 6414 408454
rect 5794 408134 6414 408218
rect 5794 407898 5826 408134
rect 6062 407898 6146 408134
rect 6382 407898 6414 408134
rect 185794 408218 185826 408454
rect 186062 408218 186146 408454
rect 186382 408218 186414 408454
rect 185794 408134 186414 408218
rect 185794 407898 185826 408134
rect 186062 407898 186146 408134
rect 186382 407898 186414 408134
rect 221794 408218 221826 408454
rect 222062 408218 222146 408454
rect 222382 408218 222414 408454
rect 221794 408134 222414 408218
rect 221794 407898 221826 408134
rect 222062 407898 222146 408134
rect 222382 407898 222414 408134
rect 257794 408218 257826 408454
rect 258062 408218 258146 408454
rect 258382 408218 258414 408454
rect 257794 408134 258414 408218
rect 257794 407898 257826 408134
rect 258062 407898 258146 408134
rect 258382 407898 258414 408134
rect 293794 408218 293826 408454
rect 294062 408218 294146 408454
rect 294382 408218 294414 408454
rect 293794 408134 294414 408218
rect 293794 407898 293826 408134
rect 294062 407898 294146 408134
rect 294382 407898 294414 408134
rect 329794 408218 329826 408454
rect 330062 408218 330146 408454
rect 330382 408218 330414 408454
rect 329794 408134 330414 408218
rect 329794 407898 329826 408134
rect 330062 407898 330146 408134
rect 330382 407898 330414 408134
rect 365794 408218 365826 408454
rect 366062 408218 366146 408454
rect 366382 408218 366414 408454
rect 365794 408134 366414 408218
rect 365794 407898 365826 408134
rect 366062 407898 366146 408134
rect 366382 407898 366414 408134
rect 401794 408218 401826 408454
rect 402062 408218 402146 408454
rect 402382 408218 402414 408454
rect 401794 408134 402414 408218
rect 401794 407898 401826 408134
rect 402062 407898 402146 408134
rect 402382 407898 402414 408134
rect 568478 408218 568510 408454
rect 568746 408218 568830 408454
rect 569066 408218 569098 408454
rect 568478 408134 569098 408218
rect 568478 407898 568510 408134
rect 568746 407898 568830 408134
rect 569066 407898 569098 408134
rect 577794 408218 577826 408454
rect 578062 408218 578146 408454
rect 578382 408218 578414 408454
rect 577794 408134 578414 408218
rect 577794 407898 577826 408134
rect 578062 407898 578146 408134
rect 578382 407898 578414 408134
rect 1794 372454 2414 407898
rect 9514 375938 9546 376174
rect 9782 375938 9866 376174
rect 10102 375938 10134 376174
rect 9514 375854 10134 375938
rect 9514 375618 9546 375854
rect 9782 375618 9866 375854
rect 10102 375618 10134 375854
rect 189514 375938 189546 376174
rect 189782 375938 189866 376174
rect 190102 375938 190134 376174
rect 189514 375854 190134 375938
rect 189514 375618 189546 375854
rect 189782 375618 189866 375854
rect 190102 375618 190134 375854
rect 225514 375938 225546 376174
rect 225782 375938 225866 376174
rect 226102 375938 226134 376174
rect 225514 375854 226134 375938
rect 225514 375618 225546 375854
rect 225782 375618 225866 375854
rect 226102 375618 226134 375854
rect 261514 375938 261546 376174
rect 261782 375938 261866 376174
rect 262102 375938 262134 376174
rect 261514 375854 262134 375938
rect 261514 375618 261546 375854
rect 261782 375618 261866 375854
rect 262102 375618 262134 375854
rect 297514 375938 297546 376174
rect 297782 375938 297866 376174
rect 298102 375938 298134 376174
rect 297514 375854 298134 375938
rect 297514 375618 297546 375854
rect 297782 375618 297866 375854
rect 298102 375618 298134 375854
rect 333514 375938 333546 376174
rect 333782 375938 333866 376174
rect 334102 375938 334134 376174
rect 333514 375854 334134 375938
rect 333514 375618 333546 375854
rect 333782 375618 333866 375854
rect 334102 375618 334134 375854
rect 369514 375938 369546 376174
rect 369782 375938 369866 376174
rect 370102 375938 370134 376174
rect 369514 375854 370134 375938
rect 369514 375618 369546 375854
rect 369782 375618 369866 375854
rect 370102 375618 370134 375854
rect 405514 375938 405546 376174
rect 405782 375938 405866 376174
rect 406102 375938 406134 376174
rect 405514 375854 406134 375938
rect 405514 375618 405546 375854
rect 405782 375618 405866 375854
rect 406102 375618 406134 375854
rect 572342 375938 572374 376174
rect 572610 375938 572694 376174
rect 572930 375938 572962 376174
rect 572342 375854 572962 375938
rect 572342 375618 572374 375854
rect 572610 375618 572694 375854
rect 572930 375618 572962 375854
rect 577794 372454 578414 407898
rect 1794 372218 1826 372454
rect 2062 372218 2146 372454
rect 2382 372218 2414 372454
rect 1794 372134 2414 372218
rect 1794 371898 1826 372134
rect 2062 371898 2146 372134
rect 2382 371898 2414 372134
rect 5794 372218 5826 372454
rect 6062 372218 6146 372454
rect 6382 372218 6414 372454
rect 5794 372134 6414 372218
rect 5794 371898 5826 372134
rect 6062 371898 6146 372134
rect 6382 371898 6414 372134
rect 185794 372218 185826 372454
rect 186062 372218 186146 372454
rect 186382 372218 186414 372454
rect 185794 372134 186414 372218
rect 185794 371898 185826 372134
rect 186062 371898 186146 372134
rect 186382 371898 186414 372134
rect 221794 372218 221826 372454
rect 222062 372218 222146 372454
rect 222382 372218 222414 372454
rect 221794 372134 222414 372218
rect 221794 371898 221826 372134
rect 222062 371898 222146 372134
rect 222382 371898 222414 372134
rect 257794 372218 257826 372454
rect 258062 372218 258146 372454
rect 258382 372218 258414 372454
rect 257794 372134 258414 372218
rect 257794 371898 257826 372134
rect 258062 371898 258146 372134
rect 258382 371898 258414 372134
rect 293794 372218 293826 372454
rect 294062 372218 294146 372454
rect 294382 372218 294414 372454
rect 293794 372134 294414 372218
rect 293794 371898 293826 372134
rect 294062 371898 294146 372134
rect 294382 371898 294414 372134
rect 329794 372218 329826 372454
rect 330062 372218 330146 372454
rect 330382 372218 330414 372454
rect 329794 372134 330414 372218
rect 329794 371898 329826 372134
rect 330062 371898 330146 372134
rect 330382 371898 330414 372134
rect 365794 372218 365826 372454
rect 366062 372218 366146 372454
rect 366382 372218 366414 372454
rect 365794 372134 366414 372218
rect 365794 371898 365826 372134
rect 366062 371898 366146 372134
rect 366382 371898 366414 372134
rect 401794 372218 401826 372454
rect 402062 372218 402146 372454
rect 402382 372218 402414 372454
rect 401794 372134 402414 372218
rect 401794 371898 401826 372134
rect 402062 371898 402146 372134
rect 402382 371898 402414 372134
rect 568478 372218 568510 372454
rect 568746 372218 568830 372454
rect 569066 372218 569098 372454
rect 568478 372134 569098 372218
rect 568478 371898 568510 372134
rect 568746 371898 568830 372134
rect 569066 371898 569098 372134
rect 577794 372218 577826 372454
rect 578062 372218 578146 372454
rect 578382 372218 578414 372454
rect 577794 372134 578414 372218
rect 577794 371898 577826 372134
rect 578062 371898 578146 372134
rect 578382 371898 578414 372134
rect 1794 336454 2414 371898
rect 9514 339938 9546 340174
rect 9782 339938 9866 340174
rect 10102 339938 10134 340174
rect 9514 339854 10134 339938
rect 9514 339618 9546 339854
rect 9782 339618 9866 339854
rect 10102 339618 10134 339854
rect 189514 339938 189546 340174
rect 189782 339938 189866 340174
rect 190102 339938 190134 340174
rect 189514 339854 190134 339938
rect 189514 339618 189546 339854
rect 189782 339618 189866 339854
rect 190102 339618 190134 339854
rect 225514 339938 225546 340174
rect 225782 339938 225866 340174
rect 226102 339938 226134 340174
rect 225514 339854 226134 339938
rect 225514 339618 225546 339854
rect 225782 339618 225866 339854
rect 226102 339618 226134 339854
rect 261514 339938 261546 340174
rect 261782 339938 261866 340174
rect 262102 339938 262134 340174
rect 261514 339854 262134 339938
rect 261514 339618 261546 339854
rect 261782 339618 261866 339854
rect 262102 339618 262134 339854
rect 297514 339938 297546 340174
rect 297782 339938 297866 340174
rect 298102 339938 298134 340174
rect 297514 339854 298134 339938
rect 297514 339618 297546 339854
rect 297782 339618 297866 339854
rect 298102 339618 298134 339854
rect 333514 339938 333546 340174
rect 333782 339938 333866 340174
rect 334102 339938 334134 340174
rect 333514 339854 334134 339938
rect 333514 339618 333546 339854
rect 333782 339618 333866 339854
rect 334102 339618 334134 339854
rect 369514 339938 369546 340174
rect 369782 339938 369866 340174
rect 370102 339938 370134 340174
rect 369514 339854 370134 339938
rect 369514 339618 369546 339854
rect 369782 339618 369866 339854
rect 370102 339618 370134 339854
rect 405514 339938 405546 340174
rect 405782 339938 405866 340174
rect 406102 339938 406134 340174
rect 405514 339854 406134 339938
rect 405514 339618 405546 339854
rect 405782 339618 405866 339854
rect 406102 339618 406134 339854
rect 572342 339938 572374 340174
rect 572610 339938 572694 340174
rect 572930 339938 572962 340174
rect 572342 339854 572962 339938
rect 572342 339618 572374 339854
rect 572610 339618 572694 339854
rect 572930 339618 572962 339854
rect 577794 336454 578414 371898
rect 1794 336218 1826 336454
rect 2062 336218 2146 336454
rect 2382 336218 2414 336454
rect 1794 336134 2414 336218
rect 1794 335898 1826 336134
rect 2062 335898 2146 336134
rect 2382 335898 2414 336134
rect 5794 336218 5826 336454
rect 6062 336218 6146 336454
rect 6382 336218 6414 336454
rect 5794 336134 6414 336218
rect 5794 335898 5826 336134
rect 6062 335898 6146 336134
rect 6382 335898 6414 336134
rect 185794 336218 185826 336454
rect 186062 336218 186146 336454
rect 186382 336218 186414 336454
rect 185794 336134 186414 336218
rect 185794 335898 185826 336134
rect 186062 335898 186146 336134
rect 186382 335898 186414 336134
rect 221794 336218 221826 336454
rect 222062 336218 222146 336454
rect 222382 336218 222414 336454
rect 221794 336134 222414 336218
rect 221794 335898 221826 336134
rect 222062 335898 222146 336134
rect 222382 335898 222414 336134
rect 257794 336218 257826 336454
rect 258062 336218 258146 336454
rect 258382 336218 258414 336454
rect 257794 336134 258414 336218
rect 257794 335898 257826 336134
rect 258062 335898 258146 336134
rect 258382 335898 258414 336134
rect 293794 336218 293826 336454
rect 294062 336218 294146 336454
rect 294382 336218 294414 336454
rect 293794 336134 294414 336218
rect 293794 335898 293826 336134
rect 294062 335898 294146 336134
rect 294382 335898 294414 336134
rect 329794 336218 329826 336454
rect 330062 336218 330146 336454
rect 330382 336218 330414 336454
rect 329794 336134 330414 336218
rect 329794 335898 329826 336134
rect 330062 335898 330146 336134
rect 330382 335898 330414 336134
rect 365794 336218 365826 336454
rect 366062 336218 366146 336454
rect 366382 336218 366414 336454
rect 365794 336134 366414 336218
rect 365794 335898 365826 336134
rect 366062 335898 366146 336134
rect 366382 335898 366414 336134
rect 401794 336218 401826 336454
rect 402062 336218 402146 336454
rect 402382 336218 402414 336454
rect 401794 336134 402414 336218
rect 401794 335898 401826 336134
rect 402062 335898 402146 336134
rect 402382 335898 402414 336134
rect 568478 336218 568510 336454
rect 568746 336218 568830 336454
rect 569066 336218 569098 336454
rect 568478 336134 569098 336218
rect 568478 335898 568510 336134
rect 568746 335898 568830 336134
rect 569066 335898 569098 336134
rect 577794 336218 577826 336454
rect 578062 336218 578146 336454
rect 578382 336218 578414 336454
rect 577794 336134 578414 336218
rect 577794 335898 577826 336134
rect 578062 335898 578146 336134
rect 578382 335898 578414 336134
rect 1794 300454 2414 335898
rect 9514 303938 9546 304174
rect 9782 303938 9866 304174
rect 10102 303938 10134 304174
rect 9514 303854 10134 303938
rect 9514 303618 9546 303854
rect 9782 303618 9866 303854
rect 10102 303618 10134 303854
rect 189514 303938 189546 304174
rect 189782 303938 189866 304174
rect 190102 303938 190134 304174
rect 189514 303854 190134 303938
rect 189514 303618 189546 303854
rect 189782 303618 189866 303854
rect 190102 303618 190134 303854
rect 225514 303938 225546 304174
rect 225782 303938 225866 304174
rect 226102 303938 226134 304174
rect 225514 303854 226134 303938
rect 225514 303618 225546 303854
rect 225782 303618 225866 303854
rect 226102 303618 226134 303854
rect 261514 303938 261546 304174
rect 261782 303938 261866 304174
rect 262102 303938 262134 304174
rect 261514 303854 262134 303938
rect 261514 303618 261546 303854
rect 261782 303618 261866 303854
rect 262102 303618 262134 303854
rect 297514 303938 297546 304174
rect 297782 303938 297866 304174
rect 298102 303938 298134 304174
rect 297514 303854 298134 303938
rect 297514 303618 297546 303854
rect 297782 303618 297866 303854
rect 298102 303618 298134 303854
rect 333514 303938 333546 304174
rect 333782 303938 333866 304174
rect 334102 303938 334134 304174
rect 333514 303854 334134 303938
rect 333514 303618 333546 303854
rect 333782 303618 333866 303854
rect 334102 303618 334134 303854
rect 369514 303938 369546 304174
rect 369782 303938 369866 304174
rect 370102 303938 370134 304174
rect 369514 303854 370134 303938
rect 369514 303618 369546 303854
rect 369782 303618 369866 303854
rect 370102 303618 370134 303854
rect 405514 303938 405546 304174
rect 405782 303938 405866 304174
rect 406102 303938 406134 304174
rect 405514 303854 406134 303938
rect 405514 303618 405546 303854
rect 405782 303618 405866 303854
rect 406102 303618 406134 303854
rect 572342 303938 572374 304174
rect 572610 303938 572694 304174
rect 572930 303938 572962 304174
rect 572342 303854 572962 303938
rect 572342 303618 572374 303854
rect 572610 303618 572694 303854
rect 572930 303618 572962 303854
rect 577794 300454 578414 335898
rect 1794 300218 1826 300454
rect 2062 300218 2146 300454
rect 2382 300218 2414 300454
rect 1794 300134 2414 300218
rect 1794 299898 1826 300134
rect 2062 299898 2146 300134
rect 2382 299898 2414 300134
rect 5794 300218 5826 300454
rect 6062 300218 6146 300454
rect 6382 300218 6414 300454
rect 5794 300134 6414 300218
rect 5794 299898 5826 300134
rect 6062 299898 6146 300134
rect 6382 299898 6414 300134
rect 185794 300218 185826 300454
rect 186062 300218 186146 300454
rect 186382 300218 186414 300454
rect 185794 300134 186414 300218
rect 185794 299898 185826 300134
rect 186062 299898 186146 300134
rect 186382 299898 186414 300134
rect 221794 300218 221826 300454
rect 222062 300218 222146 300454
rect 222382 300218 222414 300454
rect 221794 300134 222414 300218
rect 221794 299898 221826 300134
rect 222062 299898 222146 300134
rect 222382 299898 222414 300134
rect 257794 300218 257826 300454
rect 258062 300218 258146 300454
rect 258382 300218 258414 300454
rect 257794 300134 258414 300218
rect 257794 299898 257826 300134
rect 258062 299898 258146 300134
rect 258382 299898 258414 300134
rect 293794 300218 293826 300454
rect 294062 300218 294146 300454
rect 294382 300218 294414 300454
rect 293794 300134 294414 300218
rect 293794 299898 293826 300134
rect 294062 299898 294146 300134
rect 294382 299898 294414 300134
rect 329794 300218 329826 300454
rect 330062 300218 330146 300454
rect 330382 300218 330414 300454
rect 329794 300134 330414 300218
rect 329794 299898 329826 300134
rect 330062 299898 330146 300134
rect 330382 299898 330414 300134
rect 365794 300218 365826 300454
rect 366062 300218 366146 300454
rect 366382 300218 366414 300454
rect 365794 300134 366414 300218
rect 365794 299898 365826 300134
rect 366062 299898 366146 300134
rect 366382 299898 366414 300134
rect 401794 300218 401826 300454
rect 402062 300218 402146 300454
rect 402382 300218 402414 300454
rect 401794 300134 402414 300218
rect 401794 299898 401826 300134
rect 402062 299898 402146 300134
rect 402382 299898 402414 300134
rect 568478 300218 568510 300454
rect 568746 300218 568830 300454
rect 569066 300218 569098 300454
rect 568478 300134 569098 300218
rect 568478 299898 568510 300134
rect 568746 299898 568830 300134
rect 569066 299898 569098 300134
rect 577794 300218 577826 300454
rect 578062 300218 578146 300454
rect 578382 300218 578414 300454
rect 577794 300134 578414 300218
rect 577794 299898 577826 300134
rect 578062 299898 578146 300134
rect 578382 299898 578414 300134
rect 1794 264454 2414 299898
rect 9514 267938 9546 268174
rect 9782 267938 9866 268174
rect 10102 267938 10134 268174
rect 9514 267854 10134 267938
rect 9514 267618 9546 267854
rect 9782 267618 9866 267854
rect 10102 267618 10134 267854
rect 189514 267938 189546 268174
rect 189782 267938 189866 268174
rect 190102 267938 190134 268174
rect 189514 267854 190134 267938
rect 189514 267618 189546 267854
rect 189782 267618 189866 267854
rect 190102 267618 190134 267854
rect 225514 267938 225546 268174
rect 225782 267938 225866 268174
rect 226102 267938 226134 268174
rect 225514 267854 226134 267938
rect 225514 267618 225546 267854
rect 225782 267618 225866 267854
rect 226102 267618 226134 267854
rect 261514 267938 261546 268174
rect 261782 267938 261866 268174
rect 262102 267938 262134 268174
rect 261514 267854 262134 267938
rect 261514 267618 261546 267854
rect 261782 267618 261866 267854
rect 262102 267618 262134 267854
rect 297514 267938 297546 268174
rect 297782 267938 297866 268174
rect 298102 267938 298134 268174
rect 297514 267854 298134 267938
rect 297514 267618 297546 267854
rect 297782 267618 297866 267854
rect 298102 267618 298134 267854
rect 333514 267938 333546 268174
rect 333782 267938 333866 268174
rect 334102 267938 334134 268174
rect 333514 267854 334134 267938
rect 333514 267618 333546 267854
rect 333782 267618 333866 267854
rect 334102 267618 334134 267854
rect 369514 267938 369546 268174
rect 369782 267938 369866 268174
rect 370102 267938 370134 268174
rect 369514 267854 370134 267938
rect 369514 267618 369546 267854
rect 369782 267618 369866 267854
rect 370102 267618 370134 267854
rect 405514 267938 405546 268174
rect 405782 267938 405866 268174
rect 406102 267938 406134 268174
rect 405514 267854 406134 267938
rect 405514 267618 405546 267854
rect 405782 267618 405866 267854
rect 406102 267618 406134 267854
rect 572342 267938 572374 268174
rect 572610 267938 572694 268174
rect 572930 267938 572962 268174
rect 572342 267854 572962 267938
rect 572342 267618 572374 267854
rect 572610 267618 572694 267854
rect 572930 267618 572962 267854
rect 577794 264454 578414 299898
rect 1794 264218 1826 264454
rect 2062 264218 2146 264454
rect 2382 264218 2414 264454
rect 1794 264134 2414 264218
rect 1794 263898 1826 264134
rect 2062 263898 2146 264134
rect 2382 263898 2414 264134
rect 5794 264218 5826 264454
rect 6062 264218 6146 264454
rect 6382 264218 6414 264454
rect 5794 264134 6414 264218
rect 5794 263898 5826 264134
rect 6062 263898 6146 264134
rect 6382 263898 6414 264134
rect 185794 264218 185826 264454
rect 186062 264218 186146 264454
rect 186382 264218 186414 264454
rect 185794 264134 186414 264218
rect 185794 263898 185826 264134
rect 186062 263898 186146 264134
rect 186382 263898 186414 264134
rect 221794 264218 221826 264454
rect 222062 264218 222146 264454
rect 222382 264218 222414 264454
rect 221794 264134 222414 264218
rect 221794 263898 221826 264134
rect 222062 263898 222146 264134
rect 222382 263898 222414 264134
rect 257794 264218 257826 264454
rect 258062 264218 258146 264454
rect 258382 264218 258414 264454
rect 257794 264134 258414 264218
rect 257794 263898 257826 264134
rect 258062 263898 258146 264134
rect 258382 263898 258414 264134
rect 293794 264218 293826 264454
rect 294062 264218 294146 264454
rect 294382 264218 294414 264454
rect 293794 264134 294414 264218
rect 293794 263898 293826 264134
rect 294062 263898 294146 264134
rect 294382 263898 294414 264134
rect 329794 264218 329826 264454
rect 330062 264218 330146 264454
rect 330382 264218 330414 264454
rect 329794 264134 330414 264218
rect 329794 263898 329826 264134
rect 330062 263898 330146 264134
rect 330382 263898 330414 264134
rect 365794 264218 365826 264454
rect 366062 264218 366146 264454
rect 366382 264218 366414 264454
rect 365794 264134 366414 264218
rect 365794 263898 365826 264134
rect 366062 263898 366146 264134
rect 366382 263898 366414 264134
rect 401794 264218 401826 264454
rect 402062 264218 402146 264454
rect 402382 264218 402414 264454
rect 401794 264134 402414 264218
rect 401794 263898 401826 264134
rect 402062 263898 402146 264134
rect 402382 263898 402414 264134
rect 568478 264218 568510 264454
rect 568746 264218 568830 264454
rect 569066 264218 569098 264454
rect 568478 264134 569098 264218
rect 568478 263898 568510 264134
rect 568746 263898 568830 264134
rect 569066 263898 569098 264134
rect 577794 264218 577826 264454
rect 578062 264218 578146 264454
rect 578382 264218 578414 264454
rect 577794 264134 578414 264218
rect 577794 263898 577826 264134
rect 578062 263898 578146 264134
rect 578382 263898 578414 264134
rect 1794 228454 2414 263898
rect 9514 231938 9546 232174
rect 9782 231938 9866 232174
rect 10102 231938 10134 232174
rect 9514 231854 10134 231938
rect 9514 231618 9546 231854
rect 9782 231618 9866 231854
rect 10102 231618 10134 231854
rect 45514 231938 45546 232174
rect 45782 231938 45866 232174
rect 46102 231938 46134 232174
rect 45514 231854 46134 231938
rect 45514 231618 45546 231854
rect 45782 231618 45866 231854
rect 46102 231618 46134 231854
rect 81514 231938 81546 232174
rect 81782 231938 81866 232174
rect 82102 231938 82134 232174
rect 81514 231854 82134 231938
rect 81514 231618 81546 231854
rect 81782 231618 81866 231854
rect 82102 231618 82134 231854
rect 117514 231938 117546 232174
rect 117782 231938 117866 232174
rect 118102 231938 118134 232174
rect 117514 231854 118134 231938
rect 117514 231618 117546 231854
rect 117782 231618 117866 231854
rect 118102 231618 118134 231854
rect 153514 231938 153546 232174
rect 153782 231938 153866 232174
rect 154102 231938 154134 232174
rect 153514 231854 154134 231938
rect 153514 231618 153546 231854
rect 153782 231618 153866 231854
rect 154102 231618 154134 231854
rect 189514 231938 189546 232174
rect 189782 231938 189866 232174
rect 190102 231938 190134 232174
rect 189514 231854 190134 231938
rect 189514 231618 189546 231854
rect 189782 231618 189866 231854
rect 190102 231618 190134 231854
rect 225514 231938 225546 232174
rect 225782 231938 225866 232174
rect 226102 231938 226134 232174
rect 225514 231854 226134 231938
rect 225514 231618 225546 231854
rect 225782 231618 225866 231854
rect 226102 231618 226134 231854
rect 261514 231938 261546 232174
rect 261782 231938 261866 232174
rect 262102 231938 262134 232174
rect 261514 231854 262134 231938
rect 261514 231618 261546 231854
rect 261782 231618 261866 231854
rect 262102 231618 262134 231854
rect 297514 231938 297546 232174
rect 297782 231938 297866 232174
rect 298102 231938 298134 232174
rect 297514 231854 298134 231938
rect 297514 231618 297546 231854
rect 297782 231618 297866 231854
rect 298102 231618 298134 231854
rect 333514 231938 333546 232174
rect 333782 231938 333866 232174
rect 334102 231938 334134 232174
rect 333514 231854 334134 231938
rect 333514 231618 333546 231854
rect 333782 231618 333866 231854
rect 334102 231618 334134 231854
rect 369514 231938 369546 232174
rect 369782 231938 369866 232174
rect 370102 231938 370134 232174
rect 369514 231854 370134 231938
rect 369514 231618 369546 231854
rect 369782 231618 369866 231854
rect 370102 231618 370134 231854
rect 405514 231938 405546 232174
rect 405782 231938 405866 232174
rect 406102 231938 406134 232174
rect 405514 231854 406134 231938
rect 405514 231618 405546 231854
rect 405782 231618 405866 231854
rect 406102 231618 406134 231854
rect 441514 231938 441546 232174
rect 441782 231938 441866 232174
rect 442102 231938 442134 232174
rect 441514 231854 442134 231938
rect 441514 231618 441546 231854
rect 441782 231618 441866 231854
rect 442102 231618 442134 231854
rect 477514 231938 477546 232174
rect 477782 231938 477866 232174
rect 478102 231938 478134 232174
rect 477514 231854 478134 231938
rect 477514 231618 477546 231854
rect 477782 231618 477866 231854
rect 478102 231618 478134 231854
rect 513514 231938 513546 232174
rect 513782 231938 513866 232174
rect 514102 231938 514134 232174
rect 513514 231854 514134 231938
rect 513514 231618 513546 231854
rect 513782 231618 513866 231854
rect 514102 231618 514134 231854
rect 549514 231938 549546 232174
rect 549782 231938 549866 232174
rect 550102 231938 550134 232174
rect 549514 231854 550134 231938
rect 549514 231618 549546 231854
rect 549782 231618 549866 231854
rect 550102 231618 550134 231854
rect 577794 228454 578414 263898
rect 1794 228218 1826 228454
rect 2062 228218 2146 228454
rect 2382 228218 2414 228454
rect 1794 228134 2414 228218
rect 1794 227898 1826 228134
rect 2062 227898 2146 228134
rect 2382 227898 2414 228134
rect 5794 228218 5826 228454
rect 6062 228218 6146 228454
rect 6382 228218 6414 228454
rect 5794 228134 6414 228218
rect 5794 227898 5826 228134
rect 6062 227898 6146 228134
rect 6382 227898 6414 228134
rect 41794 228218 41826 228454
rect 42062 228218 42146 228454
rect 42382 228218 42414 228454
rect 41794 228134 42414 228218
rect 41794 227898 41826 228134
rect 42062 227898 42146 228134
rect 42382 227898 42414 228134
rect 77794 228218 77826 228454
rect 78062 228218 78146 228454
rect 78382 228218 78414 228454
rect 77794 228134 78414 228218
rect 77794 227898 77826 228134
rect 78062 227898 78146 228134
rect 78382 227898 78414 228134
rect 113794 228218 113826 228454
rect 114062 228218 114146 228454
rect 114382 228218 114414 228454
rect 113794 228134 114414 228218
rect 113794 227898 113826 228134
rect 114062 227898 114146 228134
rect 114382 227898 114414 228134
rect 149794 228218 149826 228454
rect 150062 228218 150146 228454
rect 150382 228218 150414 228454
rect 149794 228134 150414 228218
rect 149794 227898 149826 228134
rect 150062 227898 150146 228134
rect 150382 227898 150414 228134
rect 185794 228218 185826 228454
rect 186062 228218 186146 228454
rect 186382 228218 186414 228454
rect 185794 228134 186414 228218
rect 185794 227898 185826 228134
rect 186062 227898 186146 228134
rect 186382 227898 186414 228134
rect 221794 228218 221826 228454
rect 222062 228218 222146 228454
rect 222382 228218 222414 228454
rect 221794 228134 222414 228218
rect 221794 227898 221826 228134
rect 222062 227898 222146 228134
rect 222382 227898 222414 228134
rect 257794 228218 257826 228454
rect 258062 228218 258146 228454
rect 258382 228218 258414 228454
rect 257794 228134 258414 228218
rect 257794 227898 257826 228134
rect 258062 227898 258146 228134
rect 258382 227898 258414 228134
rect 293794 228218 293826 228454
rect 294062 228218 294146 228454
rect 294382 228218 294414 228454
rect 293794 228134 294414 228218
rect 293794 227898 293826 228134
rect 294062 227898 294146 228134
rect 294382 227898 294414 228134
rect 329794 228218 329826 228454
rect 330062 228218 330146 228454
rect 330382 228218 330414 228454
rect 329794 228134 330414 228218
rect 329794 227898 329826 228134
rect 330062 227898 330146 228134
rect 330382 227898 330414 228134
rect 365794 228218 365826 228454
rect 366062 228218 366146 228454
rect 366382 228218 366414 228454
rect 365794 228134 366414 228218
rect 365794 227898 365826 228134
rect 366062 227898 366146 228134
rect 366382 227898 366414 228134
rect 401794 228218 401826 228454
rect 402062 228218 402146 228454
rect 402382 228218 402414 228454
rect 401794 228134 402414 228218
rect 401794 227898 401826 228134
rect 402062 227898 402146 228134
rect 402382 227898 402414 228134
rect 437794 228218 437826 228454
rect 438062 228218 438146 228454
rect 438382 228218 438414 228454
rect 437794 228134 438414 228218
rect 437794 227898 437826 228134
rect 438062 227898 438146 228134
rect 438382 227898 438414 228134
rect 473794 228218 473826 228454
rect 474062 228218 474146 228454
rect 474382 228218 474414 228454
rect 473794 228134 474414 228218
rect 473794 227898 473826 228134
rect 474062 227898 474146 228134
rect 474382 227898 474414 228134
rect 509794 228218 509826 228454
rect 510062 228218 510146 228454
rect 510382 228218 510414 228454
rect 509794 228134 510414 228218
rect 509794 227898 509826 228134
rect 510062 227898 510146 228134
rect 510382 227898 510414 228134
rect 545794 228218 545826 228454
rect 546062 228218 546146 228454
rect 546382 228218 546414 228454
rect 545794 228134 546414 228218
rect 577794 228218 577826 228454
rect 578062 228218 578146 228454
rect 578382 228218 578414 228454
rect 545794 227898 545826 228134
rect 546062 227898 546146 228134
rect 546382 227898 546414 228134
rect 568478 228139 569098 228176
rect 568478 227903 568510 228139
rect 568746 227903 568830 228139
rect 569066 227903 569098 228139
rect 1794 192454 2414 227898
rect 568478 227866 569098 227903
rect 577794 228134 578414 228218
rect 577794 227898 577826 228134
rect 578062 227898 578146 228134
rect 578382 227898 578414 228134
rect 9514 195938 9546 196174
rect 9782 195938 9866 196174
rect 10102 195938 10134 196174
rect 9514 195854 10134 195938
rect 9514 195618 9546 195854
rect 9782 195618 9866 195854
rect 10102 195618 10134 195854
rect 189514 195938 189546 196174
rect 189782 195938 189866 196174
rect 190102 195938 190134 196174
rect 189514 195854 190134 195938
rect 189514 195618 189546 195854
rect 189782 195618 189866 195854
rect 190102 195618 190134 195854
rect 225514 195938 225546 196174
rect 225782 195938 225866 196174
rect 226102 195938 226134 196174
rect 225514 195854 226134 195938
rect 225514 195618 225546 195854
rect 225782 195618 225866 195854
rect 226102 195618 226134 195854
rect 261514 195938 261546 196174
rect 261782 195938 261866 196174
rect 262102 195938 262134 196174
rect 261514 195854 262134 195938
rect 261514 195618 261546 195854
rect 261782 195618 261866 195854
rect 262102 195618 262134 195854
rect 297514 195938 297546 196174
rect 297782 195938 297866 196174
rect 298102 195938 298134 196174
rect 297514 195854 298134 195938
rect 297514 195618 297546 195854
rect 297782 195618 297866 195854
rect 298102 195618 298134 195854
rect 333514 195938 333546 196174
rect 333782 195938 333866 196174
rect 334102 195938 334134 196174
rect 333514 195854 334134 195938
rect 333514 195618 333546 195854
rect 333782 195618 333866 195854
rect 334102 195618 334134 195854
rect 369514 195938 369546 196174
rect 369782 195938 369866 196174
rect 370102 195938 370134 196174
rect 369514 195854 370134 195938
rect 369514 195618 369546 195854
rect 369782 195618 369866 195854
rect 370102 195618 370134 195854
rect 405514 195938 405546 196174
rect 405782 195938 405866 196174
rect 406102 195938 406134 196174
rect 405514 195854 406134 195938
rect 405514 195618 405546 195854
rect 405782 195618 405866 195854
rect 406102 195618 406134 195854
rect 572342 195938 572374 196174
rect 572610 195938 572694 196174
rect 572930 195938 572962 196174
rect 572342 195854 572962 195938
rect 572342 195618 572374 195854
rect 572610 195618 572694 195854
rect 572930 195618 572962 195854
rect 577794 192454 578414 227898
rect 1794 192218 1826 192454
rect 2062 192218 2146 192454
rect 2382 192218 2414 192454
rect 1794 192134 2414 192218
rect 1794 191898 1826 192134
rect 2062 191898 2146 192134
rect 2382 191898 2414 192134
rect 5794 192218 5826 192454
rect 6062 192218 6146 192454
rect 6382 192218 6414 192454
rect 5794 192134 6414 192218
rect 5794 191898 5826 192134
rect 6062 191898 6146 192134
rect 6382 191898 6414 192134
rect 185794 192218 185826 192454
rect 186062 192218 186146 192454
rect 186382 192218 186414 192454
rect 185794 192134 186414 192218
rect 185794 191898 185826 192134
rect 186062 191898 186146 192134
rect 186382 191898 186414 192134
rect 221794 192218 221826 192454
rect 222062 192218 222146 192454
rect 222382 192218 222414 192454
rect 221794 192134 222414 192218
rect 221794 191898 221826 192134
rect 222062 191898 222146 192134
rect 222382 191898 222414 192134
rect 257794 192218 257826 192454
rect 258062 192218 258146 192454
rect 258382 192218 258414 192454
rect 257794 192134 258414 192218
rect 257794 191898 257826 192134
rect 258062 191898 258146 192134
rect 258382 191898 258414 192134
rect 293794 192218 293826 192454
rect 294062 192218 294146 192454
rect 294382 192218 294414 192454
rect 293794 192134 294414 192218
rect 293794 191898 293826 192134
rect 294062 191898 294146 192134
rect 294382 191898 294414 192134
rect 329794 192218 329826 192454
rect 330062 192218 330146 192454
rect 330382 192218 330414 192454
rect 329794 192134 330414 192218
rect 329794 191898 329826 192134
rect 330062 191898 330146 192134
rect 330382 191898 330414 192134
rect 365794 192218 365826 192454
rect 366062 192218 366146 192454
rect 366382 192218 366414 192454
rect 365794 192134 366414 192218
rect 365794 191898 365826 192134
rect 366062 191898 366146 192134
rect 366382 191898 366414 192134
rect 401794 192218 401826 192454
rect 402062 192218 402146 192454
rect 402382 192218 402414 192454
rect 401794 192134 402414 192218
rect 401794 191898 401826 192134
rect 402062 191898 402146 192134
rect 402382 191898 402414 192134
rect 568478 192218 568510 192454
rect 568746 192218 568830 192454
rect 569066 192218 569098 192454
rect 568478 192134 569098 192218
rect 568478 191898 568510 192134
rect 568746 191898 568830 192134
rect 569066 191898 569098 192134
rect 577794 192218 577826 192454
rect 578062 192218 578146 192454
rect 578382 192218 578414 192454
rect 577794 192134 578414 192218
rect 577794 191898 577826 192134
rect 578062 191898 578146 192134
rect 578382 191898 578414 192134
rect 1794 156454 2414 191898
rect 9514 159938 9546 160174
rect 9782 159938 9866 160174
rect 10102 159938 10134 160174
rect 9514 159854 10134 159938
rect 9514 159618 9546 159854
rect 9782 159618 9866 159854
rect 10102 159618 10134 159854
rect 189514 159938 189546 160174
rect 189782 159938 189866 160174
rect 190102 159938 190134 160174
rect 189514 159854 190134 159938
rect 189514 159618 189546 159854
rect 189782 159618 189866 159854
rect 190102 159618 190134 159854
rect 225514 159938 225546 160174
rect 225782 159938 225866 160174
rect 226102 159938 226134 160174
rect 225514 159854 226134 159938
rect 225514 159618 225546 159854
rect 225782 159618 225866 159854
rect 226102 159618 226134 159854
rect 261514 159938 261546 160174
rect 261782 159938 261866 160174
rect 262102 159938 262134 160174
rect 261514 159854 262134 159938
rect 261514 159618 261546 159854
rect 261782 159618 261866 159854
rect 262102 159618 262134 159854
rect 297514 159938 297546 160174
rect 297782 159938 297866 160174
rect 298102 159938 298134 160174
rect 297514 159854 298134 159938
rect 297514 159618 297546 159854
rect 297782 159618 297866 159854
rect 298102 159618 298134 159854
rect 333514 159938 333546 160174
rect 333782 159938 333866 160174
rect 334102 159938 334134 160174
rect 333514 159854 334134 159938
rect 333514 159618 333546 159854
rect 333782 159618 333866 159854
rect 334102 159618 334134 159854
rect 369514 159938 369546 160174
rect 369782 159938 369866 160174
rect 370102 159938 370134 160174
rect 369514 159854 370134 159938
rect 369514 159618 369546 159854
rect 369782 159618 369866 159854
rect 370102 159618 370134 159854
rect 405514 159938 405546 160174
rect 405782 159938 405866 160174
rect 406102 159938 406134 160174
rect 405514 159854 406134 159938
rect 405514 159618 405546 159854
rect 405782 159618 405866 159854
rect 406102 159618 406134 159854
rect 572342 159938 572374 160174
rect 572610 159938 572694 160174
rect 572930 159938 572962 160174
rect 572342 159854 572962 159938
rect 572342 159618 572374 159854
rect 572610 159618 572694 159854
rect 572930 159618 572962 159854
rect 577794 156454 578414 191898
rect 1794 156218 1826 156454
rect 2062 156218 2146 156454
rect 2382 156218 2414 156454
rect 1794 156134 2414 156218
rect 1794 155898 1826 156134
rect 2062 155898 2146 156134
rect 2382 155898 2414 156134
rect 5794 156218 5826 156454
rect 6062 156218 6146 156454
rect 6382 156218 6414 156454
rect 5794 156134 6414 156218
rect 5794 155898 5826 156134
rect 6062 155898 6146 156134
rect 6382 155898 6414 156134
rect 185794 156218 185826 156454
rect 186062 156218 186146 156454
rect 186382 156218 186414 156454
rect 185794 156134 186414 156218
rect 185794 155898 185826 156134
rect 186062 155898 186146 156134
rect 186382 155898 186414 156134
rect 221794 156218 221826 156454
rect 222062 156218 222146 156454
rect 222382 156218 222414 156454
rect 221794 156134 222414 156218
rect 221794 155898 221826 156134
rect 222062 155898 222146 156134
rect 222382 155898 222414 156134
rect 257794 156218 257826 156454
rect 258062 156218 258146 156454
rect 258382 156218 258414 156454
rect 257794 156134 258414 156218
rect 257794 155898 257826 156134
rect 258062 155898 258146 156134
rect 258382 155898 258414 156134
rect 293794 156218 293826 156454
rect 294062 156218 294146 156454
rect 294382 156218 294414 156454
rect 293794 156134 294414 156218
rect 293794 155898 293826 156134
rect 294062 155898 294146 156134
rect 294382 155898 294414 156134
rect 329794 156218 329826 156454
rect 330062 156218 330146 156454
rect 330382 156218 330414 156454
rect 329794 156134 330414 156218
rect 329794 155898 329826 156134
rect 330062 155898 330146 156134
rect 330382 155898 330414 156134
rect 365794 156218 365826 156454
rect 366062 156218 366146 156454
rect 366382 156218 366414 156454
rect 365794 156134 366414 156218
rect 365794 155898 365826 156134
rect 366062 155898 366146 156134
rect 366382 155898 366414 156134
rect 401794 156218 401826 156454
rect 402062 156218 402146 156454
rect 402382 156218 402414 156454
rect 401794 156134 402414 156218
rect 401794 155898 401826 156134
rect 402062 155898 402146 156134
rect 402382 155898 402414 156134
rect 568478 156218 568510 156454
rect 568746 156218 568830 156454
rect 569066 156218 569098 156454
rect 568478 156134 569098 156218
rect 568478 155898 568510 156134
rect 568746 155898 568830 156134
rect 569066 155898 569098 156134
rect 577794 156218 577826 156454
rect 578062 156218 578146 156454
rect 578382 156218 578414 156454
rect 577794 156134 578414 156218
rect 577794 155898 577826 156134
rect 578062 155898 578146 156134
rect 578382 155898 578414 156134
rect 1794 120454 2414 155898
rect 9514 123938 9546 124174
rect 9782 123938 9866 124174
rect 10102 123938 10134 124174
rect 9514 123854 10134 123938
rect 9514 123618 9546 123854
rect 9782 123618 9866 123854
rect 10102 123618 10134 123854
rect 45514 123938 45546 124174
rect 45782 123938 45866 124174
rect 46102 123938 46134 124174
rect 45514 123854 46134 123938
rect 45514 123618 45546 123854
rect 45782 123618 45866 123854
rect 46102 123618 46134 123854
rect 81514 123938 81546 124174
rect 81782 123938 81866 124174
rect 82102 123938 82134 124174
rect 81514 123854 82134 123938
rect 81514 123618 81546 123854
rect 81782 123618 81866 123854
rect 82102 123618 82134 123854
rect 117514 123938 117546 124174
rect 117782 123938 117866 124174
rect 118102 123938 118134 124174
rect 117514 123854 118134 123938
rect 117514 123618 117546 123854
rect 117782 123618 117866 123854
rect 118102 123618 118134 123854
rect 153514 123938 153546 124174
rect 153782 123938 153866 124174
rect 154102 123938 154134 124174
rect 153514 123854 154134 123938
rect 153514 123618 153546 123854
rect 153782 123618 153866 123854
rect 154102 123618 154134 123854
rect 189514 123938 189546 124174
rect 189782 123938 189866 124174
rect 190102 123938 190134 124174
rect 189514 123854 190134 123938
rect 189514 123618 189546 123854
rect 189782 123618 189866 123854
rect 190102 123618 190134 123854
rect 225514 123938 225546 124174
rect 225782 123938 225866 124174
rect 226102 123938 226134 124174
rect 225514 123854 226134 123938
rect 225514 123618 225546 123854
rect 225782 123618 225866 123854
rect 226102 123618 226134 123854
rect 261514 123938 261546 124174
rect 261782 123938 261866 124174
rect 262102 123938 262134 124174
rect 261514 123854 262134 123938
rect 261514 123618 261546 123854
rect 261782 123618 261866 123854
rect 262102 123618 262134 123854
rect 297514 123938 297546 124174
rect 297782 123938 297866 124174
rect 298102 123938 298134 124174
rect 297514 123854 298134 123938
rect 297514 123618 297546 123854
rect 297782 123618 297866 123854
rect 298102 123618 298134 123854
rect 333514 123938 333546 124174
rect 333782 123938 333866 124174
rect 334102 123938 334134 124174
rect 333514 123854 334134 123938
rect 333514 123618 333546 123854
rect 333782 123618 333866 123854
rect 334102 123618 334134 123854
rect 369514 123938 369546 124174
rect 369782 123938 369866 124174
rect 370102 123938 370134 124174
rect 369514 123854 370134 123938
rect 369514 123618 369546 123854
rect 369782 123618 369866 123854
rect 370102 123618 370134 123854
rect 405514 123938 405546 124174
rect 405782 123938 405866 124174
rect 406102 123938 406134 124174
rect 405514 123854 406134 123938
rect 405514 123618 405546 123854
rect 405782 123618 405866 123854
rect 406102 123618 406134 123854
rect 441514 123938 441546 124174
rect 441782 123938 441866 124174
rect 442102 123938 442134 124174
rect 441514 123854 442134 123938
rect 441514 123618 441546 123854
rect 441782 123618 441866 123854
rect 442102 123618 442134 123854
rect 477514 123938 477546 124174
rect 477782 123938 477866 124174
rect 478102 123938 478134 124174
rect 477514 123854 478134 123938
rect 477514 123618 477546 123854
rect 477782 123618 477866 123854
rect 478102 123618 478134 123854
rect 513514 123938 513546 124174
rect 513782 123938 513866 124174
rect 514102 123938 514134 124174
rect 513514 123854 514134 123938
rect 513514 123618 513546 123854
rect 513782 123618 513866 123854
rect 514102 123618 514134 123854
rect 549514 123938 549546 124174
rect 549782 123938 549866 124174
rect 550102 123938 550134 124174
rect 549514 123854 550134 123938
rect 549514 123618 549546 123854
rect 549782 123618 549866 123854
rect 550102 123618 550134 123854
rect 577794 120454 578414 155898
rect 1794 120218 1826 120454
rect 2062 120218 2146 120454
rect 2382 120218 2414 120454
rect 1794 120134 2414 120218
rect 1794 119898 1826 120134
rect 2062 119898 2146 120134
rect 2382 119898 2414 120134
rect 5794 120218 5826 120454
rect 6062 120218 6146 120454
rect 6382 120218 6414 120454
rect 5794 120134 6414 120218
rect 5794 119898 5826 120134
rect 6062 119898 6146 120134
rect 6382 119898 6414 120134
rect 41794 120218 41826 120454
rect 42062 120218 42146 120454
rect 42382 120218 42414 120454
rect 41794 120134 42414 120218
rect 41794 119898 41826 120134
rect 42062 119898 42146 120134
rect 42382 119898 42414 120134
rect 77794 120218 77826 120454
rect 78062 120218 78146 120454
rect 78382 120218 78414 120454
rect 77794 120134 78414 120218
rect 77794 119898 77826 120134
rect 78062 119898 78146 120134
rect 78382 119898 78414 120134
rect 113794 120218 113826 120454
rect 114062 120218 114146 120454
rect 114382 120218 114414 120454
rect 113794 120134 114414 120218
rect 113794 119898 113826 120134
rect 114062 119898 114146 120134
rect 114382 119898 114414 120134
rect 149794 120218 149826 120454
rect 150062 120218 150146 120454
rect 150382 120218 150414 120454
rect 149794 120134 150414 120218
rect 149794 119898 149826 120134
rect 150062 119898 150146 120134
rect 150382 119898 150414 120134
rect 185794 120218 185826 120454
rect 186062 120218 186146 120454
rect 186382 120218 186414 120454
rect 185794 120134 186414 120218
rect 185794 119898 185826 120134
rect 186062 119898 186146 120134
rect 186382 119898 186414 120134
rect 221794 120218 221826 120454
rect 222062 120218 222146 120454
rect 222382 120218 222414 120454
rect 221794 120134 222414 120218
rect 221794 119898 221826 120134
rect 222062 119898 222146 120134
rect 222382 119898 222414 120134
rect 257794 120218 257826 120454
rect 258062 120218 258146 120454
rect 258382 120218 258414 120454
rect 257794 120134 258414 120218
rect 257794 119898 257826 120134
rect 258062 119898 258146 120134
rect 258382 119898 258414 120134
rect 293794 120218 293826 120454
rect 294062 120218 294146 120454
rect 294382 120218 294414 120454
rect 293794 120134 294414 120218
rect 293794 119898 293826 120134
rect 294062 119898 294146 120134
rect 294382 119898 294414 120134
rect 329794 120218 329826 120454
rect 330062 120218 330146 120454
rect 330382 120218 330414 120454
rect 329794 120134 330414 120218
rect 329794 119898 329826 120134
rect 330062 119898 330146 120134
rect 330382 119898 330414 120134
rect 365794 120218 365826 120454
rect 366062 120218 366146 120454
rect 366382 120218 366414 120454
rect 365794 120134 366414 120218
rect 365794 119898 365826 120134
rect 366062 119898 366146 120134
rect 366382 119898 366414 120134
rect 401794 120218 401826 120454
rect 402062 120218 402146 120454
rect 402382 120218 402414 120454
rect 401794 120134 402414 120218
rect 401794 119898 401826 120134
rect 402062 119898 402146 120134
rect 402382 119898 402414 120134
rect 437794 120218 437826 120454
rect 438062 120218 438146 120454
rect 438382 120218 438414 120454
rect 437794 120134 438414 120218
rect 437794 119898 437826 120134
rect 438062 119898 438146 120134
rect 438382 119898 438414 120134
rect 473794 120218 473826 120454
rect 474062 120218 474146 120454
rect 474382 120218 474414 120454
rect 473794 120134 474414 120218
rect 473794 119898 473826 120134
rect 474062 119898 474146 120134
rect 474382 119898 474414 120134
rect 509794 120218 509826 120454
rect 510062 120218 510146 120454
rect 510382 120218 510414 120454
rect 509794 120134 510414 120218
rect 509794 119898 509826 120134
rect 510062 119898 510146 120134
rect 510382 119898 510414 120134
rect 545794 120218 545826 120454
rect 546062 120218 546146 120454
rect 546382 120218 546414 120454
rect 545794 120134 546414 120218
rect 545794 119898 545826 120134
rect 546062 119898 546146 120134
rect 546382 119898 546414 120134
rect 577794 120218 577826 120454
rect 578062 120218 578146 120454
rect 578382 120218 578414 120454
rect 577794 120134 578414 120218
rect 577794 119898 577826 120134
rect 578062 119898 578146 120134
rect 578382 119898 578414 120134
rect 1794 84454 2414 119898
rect 9514 87938 9546 88174
rect 9782 87938 9866 88174
rect 10102 87938 10134 88174
rect 9514 87854 10134 87938
rect 9514 87618 9546 87854
rect 9782 87618 9866 87854
rect 10102 87618 10134 87854
rect 189514 87938 189546 88174
rect 189782 87938 189866 88174
rect 190102 87938 190134 88174
rect 189514 87854 190134 87938
rect 189514 87618 189546 87854
rect 189782 87618 189866 87854
rect 190102 87618 190134 87854
rect 369514 87938 369546 88174
rect 369782 87938 369866 88174
rect 370102 87938 370134 88174
rect 369514 87854 370134 87938
rect 369514 87618 369546 87854
rect 369782 87618 369866 87854
rect 370102 87618 370134 87854
rect 405514 87938 405546 88174
rect 405782 87938 405866 88174
rect 406102 87938 406134 88174
rect 405514 87854 406134 87938
rect 405514 87618 405546 87854
rect 405782 87618 405866 87854
rect 406102 87618 406134 87854
rect 572342 87938 572374 88174
rect 572610 87938 572694 88174
rect 572930 87938 572962 88174
rect 572342 87854 572962 87938
rect 572342 87618 572374 87854
rect 572610 87618 572694 87854
rect 572930 87618 572962 87854
rect 577794 84454 578414 119898
rect 1794 84218 1826 84454
rect 2062 84218 2146 84454
rect 2382 84218 2414 84454
rect 1794 84134 2414 84218
rect 1794 83898 1826 84134
rect 2062 83898 2146 84134
rect 2382 83898 2414 84134
rect 5794 84218 5826 84454
rect 6062 84218 6146 84454
rect 6382 84218 6414 84454
rect 5794 84134 6414 84218
rect 5794 83898 5826 84134
rect 6062 83898 6146 84134
rect 6382 83898 6414 84134
rect 185794 84218 185826 84454
rect 186062 84218 186146 84454
rect 186382 84218 186414 84454
rect 185794 84134 186414 84218
rect 185794 83898 185826 84134
rect 186062 83898 186146 84134
rect 186382 83898 186414 84134
rect 365794 84218 365826 84454
rect 366062 84218 366146 84454
rect 366382 84218 366414 84454
rect 365794 84134 366414 84218
rect 365794 83898 365826 84134
rect 366062 83898 366146 84134
rect 366382 83898 366414 84134
rect 401794 84218 401826 84454
rect 402062 84218 402146 84454
rect 402382 84218 402414 84454
rect 401794 84134 402414 84218
rect 401794 83898 401826 84134
rect 402062 83898 402146 84134
rect 402382 83898 402414 84134
rect 568478 84218 568510 84454
rect 568746 84218 568830 84454
rect 569066 84218 569098 84454
rect 568478 84134 569098 84218
rect 568478 83898 568510 84134
rect 568746 83898 568830 84134
rect 569066 83898 569098 84134
rect 577794 84218 577826 84454
rect 578062 84218 578146 84454
rect 578382 84218 578414 84454
rect 577794 84134 578414 84218
rect 577794 83898 577826 84134
rect 578062 83898 578146 84134
rect 578382 83898 578414 84134
rect 1794 48454 2414 83898
rect 9514 51938 9546 52174
rect 9782 51938 9866 52174
rect 10102 51938 10134 52174
rect 9514 51854 10134 51938
rect 9514 51618 9546 51854
rect 9782 51618 9866 51854
rect 10102 51618 10134 51854
rect 189514 51938 189546 52174
rect 189782 51938 189866 52174
rect 190102 51938 190134 52174
rect 189514 51854 190134 51938
rect 189514 51618 189546 51854
rect 189782 51618 189866 51854
rect 190102 51618 190134 51854
rect 369514 51938 369546 52174
rect 369782 51938 369866 52174
rect 370102 51938 370134 52174
rect 369514 51854 370134 51938
rect 369514 51618 369546 51854
rect 369782 51618 369866 51854
rect 370102 51618 370134 51854
rect 405514 51938 405546 52174
rect 405782 51938 405866 52174
rect 406102 51938 406134 52174
rect 405514 51854 406134 51938
rect 405514 51618 405546 51854
rect 405782 51618 405866 51854
rect 406102 51618 406134 51854
rect 572342 51938 572374 52174
rect 572610 51938 572694 52174
rect 572930 51938 572962 52174
rect 572342 51854 572962 51938
rect 572342 51618 572374 51854
rect 572610 51618 572694 51854
rect 572930 51618 572962 51854
rect 577794 48454 578414 83898
rect 1794 48218 1826 48454
rect 2062 48218 2146 48454
rect 2382 48218 2414 48454
rect 1794 48134 2414 48218
rect 1794 47898 1826 48134
rect 2062 47898 2146 48134
rect 2382 47898 2414 48134
rect 5794 48218 5826 48454
rect 6062 48218 6146 48454
rect 6382 48218 6414 48454
rect 5794 48134 6414 48218
rect 5794 47898 5826 48134
rect 6062 47898 6146 48134
rect 6382 47898 6414 48134
rect 185794 48218 185826 48454
rect 186062 48218 186146 48454
rect 186382 48218 186414 48454
rect 185794 48134 186414 48218
rect 185794 47898 185826 48134
rect 186062 47898 186146 48134
rect 186382 47898 186414 48134
rect 365794 48218 365826 48454
rect 366062 48218 366146 48454
rect 366382 48218 366414 48454
rect 365794 48134 366414 48218
rect 365794 47898 365826 48134
rect 366062 47898 366146 48134
rect 366382 47898 366414 48134
rect 401794 48218 401826 48454
rect 402062 48218 402146 48454
rect 402382 48218 402414 48454
rect 401794 48134 402414 48218
rect 401794 47898 401826 48134
rect 402062 47898 402146 48134
rect 402382 47898 402414 48134
rect 568478 48218 568510 48454
rect 568746 48218 568830 48454
rect 569066 48218 569098 48454
rect 568478 48134 569098 48218
rect 568478 47898 568510 48134
rect 568746 47898 568830 48134
rect 569066 47898 569098 48134
rect 577794 48218 577826 48454
rect 578062 48218 578146 48454
rect 578382 48218 578414 48454
rect 577794 48134 578414 48218
rect 577794 47898 577826 48134
rect 578062 47898 578146 48134
rect 578382 47898 578414 48134
rect 1794 12454 2414 47898
rect 9514 15938 9546 16174
rect 9782 15938 9866 16174
rect 10102 15938 10134 16174
rect 9514 15854 10134 15938
rect 9514 15618 9546 15854
rect 9782 15618 9866 15854
rect 10102 15618 10134 15854
rect 45514 15938 45546 16174
rect 45782 15938 45866 16174
rect 46102 15938 46134 16174
rect 45514 15854 46134 15938
rect 45514 15618 45546 15854
rect 45782 15618 45866 15854
rect 46102 15618 46134 15854
rect 81514 15938 81546 16174
rect 81782 15938 81866 16174
rect 82102 15938 82134 16174
rect 81514 15854 82134 15938
rect 81514 15618 81546 15854
rect 81782 15618 81866 15854
rect 82102 15618 82134 15854
rect 117514 15938 117546 16174
rect 117782 15938 117866 16174
rect 118102 15938 118134 16174
rect 117514 15854 118134 15938
rect 117514 15618 117546 15854
rect 117782 15618 117866 15854
rect 118102 15618 118134 15854
rect 153514 15938 153546 16174
rect 153782 15938 153866 16174
rect 154102 15938 154134 16174
rect 153514 15854 154134 15938
rect 153514 15618 153546 15854
rect 153782 15618 153866 15854
rect 154102 15618 154134 15854
rect 189514 15938 189546 16174
rect 189782 15938 189866 16174
rect 190102 15938 190134 16174
rect 189514 15854 190134 15938
rect 189514 15618 189546 15854
rect 189782 15618 189866 15854
rect 190102 15618 190134 15854
rect 225514 15938 225546 16174
rect 225782 15938 225866 16174
rect 226102 15938 226134 16174
rect 225514 15854 226134 15938
rect 225514 15618 225546 15854
rect 225782 15618 225866 15854
rect 226102 15618 226134 15854
rect 261514 15938 261546 16174
rect 261782 15938 261866 16174
rect 262102 15938 262134 16174
rect 261514 15854 262134 15938
rect 261514 15618 261546 15854
rect 261782 15618 261866 15854
rect 262102 15618 262134 15854
rect 297514 15938 297546 16174
rect 297782 15938 297866 16174
rect 298102 15938 298134 16174
rect 297514 15854 298134 15938
rect 297514 15618 297546 15854
rect 297782 15618 297866 15854
rect 298102 15618 298134 15854
rect 333514 15938 333546 16174
rect 333782 15938 333866 16174
rect 334102 15938 334134 16174
rect 333514 15854 334134 15938
rect 333514 15618 333546 15854
rect 333782 15618 333866 15854
rect 334102 15618 334134 15854
rect 369514 15938 369546 16174
rect 369782 15938 369866 16174
rect 370102 15938 370134 16174
rect 369514 15854 370134 15938
rect 369514 15618 369546 15854
rect 369782 15618 369866 15854
rect 370102 15618 370134 15854
rect 405514 15938 405546 16174
rect 405782 15938 405866 16174
rect 406102 15938 406134 16174
rect 405514 15854 406134 15938
rect 405514 15618 405546 15854
rect 405782 15618 405866 15854
rect 406102 15618 406134 15854
rect 441514 15938 441546 16174
rect 441782 15938 441866 16174
rect 442102 15938 442134 16174
rect 441514 15854 442134 15938
rect 441514 15618 441546 15854
rect 441782 15618 441866 15854
rect 442102 15618 442134 15854
rect 477514 15938 477546 16174
rect 477782 15938 477866 16174
rect 478102 15938 478134 16174
rect 477514 15854 478134 15938
rect 477514 15618 477546 15854
rect 477782 15618 477866 15854
rect 478102 15618 478134 15854
rect 513514 15938 513546 16174
rect 513782 15938 513866 16174
rect 514102 15938 514134 16174
rect 513514 15854 514134 15938
rect 513514 15618 513546 15854
rect 513782 15618 513866 15854
rect 514102 15618 514134 15854
rect 549514 15938 549546 16174
rect 549782 15938 549866 16174
rect 550102 15938 550134 16174
rect 549514 15854 550134 15938
rect 549514 15618 549546 15854
rect 549782 15618 549866 15854
rect 550102 15618 550134 15854
rect 577794 12454 578414 47898
rect 1794 12218 1826 12454
rect 2062 12218 2146 12454
rect 2382 12218 2414 12454
rect 1794 12134 2414 12218
rect 1794 11898 1826 12134
rect 2062 11898 2146 12134
rect 2382 11898 2414 12134
rect 5794 12218 5826 12454
rect 6062 12218 6146 12454
rect 6382 12218 6414 12454
rect 5794 12134 6414 12218
rect 5794 11898 5826 12134
rect 6062 11898 6146 12134
rect 6382 11898 6414 12134
rect 41794 12218 41826 12454
rect 42062 12218 42146 12454
rect 42382 12218 42414 12454
rect 41794 12134 42414 12218
rect 41794 11898 41826 12134
rect 42062 11898 42146 12134
rect 42382 11898 42414 12134
rect 77794 12218 77826 12454
rect 78062 12218 78146 12454
rect 78382 12218 78414 12454
rect 77794 12134 78414 12218
rect 77794 11898 77826 12134
rect 78062 11898 78146 12134
rect 78382 11898 78414 12134
rect 113794 12218 113826 12454
rect 114062 12218 114146 12454
rect 114382 12218 114414 12454
rect 113794 12134 114414 12218
rect 113794 11898 113826 12134
rect 114062 11898 114146 12134
rect 114382 11898 114414 12134
rect 149794 12218 149826 12454
rect 150062 12218 150146 12454
rect 150382 12218 150414 12454
rect 149794 12134 150414 12218
rect 149794 11898 149826 12134
rect 150062 11898 150146 12134
rect 150382 11898 150414 12134
rect 185794 12218 185826 12454
rect 186062 12218 186146 12454
rect 186382 12218 186414 12454
rect 185794 12134 186414 12218
rect 185794 11898 185826 12134
rect 186062 11898 186146 12134
rect 186382 11898 186414 12134
rect 221794 12218 221826 12454
rect 222062 12218 222146 12454
rect 222382 12218 222414 12454
rect 221794 12134 222414 12218
rect 221794 11898 221826 12134
rect 222062 11898 222146 12134
rect 222382 11898 222414 12134
rect 257794 12218 257826 12454
rect 258062 12218 258146 12454
rect 258382 12218 258414 12454
rect 257794 12134 258414 12218
rect 257794 11898 257826 12134
rect 258062 11898 258146 12134
rect 258382 11898 258414 12134
rect 293794 12218 293826 12454
rect 294062 12218 294146 12454
rect 294382 12218 294414 12454
rect 293794 12134 294414 12218
rect 293794 11898 293826 12134
rect 294062 11898 294146 12134
rect 294382 11898 294414 12134
rect 329794 12218 329826 12454
rect 330062 12218 330146 12454
rect 330382 12218 330414 12454
rect 329794 12134 330414 12218
rect 329794 11898 329826 12134
rect 330062 11898 330146 12134
rect 330382 11898 330414 12134
rect 365794 12218 365826 12454
rect 366062 12218 366146 12454
rect 366382 12218 366414 12454
rect 365794 12134 366414 12218
rect 365794 11898 365826 12134
rect 366062 11898 366146 12134
rect 366382 11898 366414 12134
rect 401794 12218 401826 12454
rect 402062 12218 402146 12454
rect 402382 12218 402414 12454
rect 401794 12134 402414 12218
rect 401794 11898 401826 12134
rect 402062 11898 402146 12134
rect 402382 11898 402414 12134
rect 437794 12218 437826 12454
rect 438062 12218 438146 12454
rect 438382 12218 438414 12454
rect 437794 12134 438414 12218
rect 437794 11898 437826 12134
rect 438062 11898 438146 12134
rect 438382 11898 438414 12134
rect 473794 12218 473826 12454
rect 474062 12218 474146 12454
rect 474382 12218 474414 12454
rect 473794 12134 474414 12218
rect 473794 11898 473826 12134
rect 474062 11898 474146 12134
rect 474382 11898 474414 12134
rect 509794 12218 509826 12454
rect 510062 12218 510146 12454
rect 510382 12218 510414 12454
rect 509794 12134 510414 12218
rect 509794 11898 509826 12134
rect 510062 11898 510146 12134
rect 510382 11898 510414 12134
rect 545794 12218 545826 12454
rect 546062 12218 546146 12454
rect 546382 12218 546414 12454
rect 545794 12134 546414 12218
rect 545794 11898 545826 12134
rect 546062 11898 546146 12134
rect 546382 11898 546414 12134
rect 577794 12218 577826 12454
rect 578062 12218 578146 12454
rect 578382 12218 578414 12454
rect 577794 12134 578414 12218
rect 577794 11898 577826 12134
rect 578062 11898 578146 12134
rect 578382 11898 578414 12134
rect 1794 -346 2414 11898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 577794 -346 578414 11898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 700174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 699938 581546 700174
rect 581782 699938 581866 700174
rect 582102 699938 582134 700174
rect 581514 699854 582134 699938
rect 581514 699618 581546 699854
rect 581782 699618 581866 699854
rect 582102 699618 582134 699854
rect 581514 664174 582134 699618
rect 581514 663938 581546 664174
rect 581782 663938 581866 664174
rect 582102 663938 582134 664174
rect 581514 663854 582134 663938
rect 581514 663618 581546 663854
rect 581782 663618 581866 663854
rect 582102 663618 582134 663854
rect 581514 628174 582134 663618
rect 581514 627938 581546 628174
rect 581782 627938 581866 628174
rect 582102 627938 582134 628174
rect 581514 627854 582134 627938
rect 581514 627618 581546 627854
rect 581782 627618 581866 627854
rect 582102 627618 582134 627854
rect 581514 592174 582134 627618
rect 581514 591938 581546 592174
rect 581782 591938 581866 592174
rect 582102 591938 582134 592174
rect 581514 591854 582134 591938
rect 581514 591618 581546 591854
rect 581782 591618 581866 591854
rect 582102 591618 582134 591854
rect 581514 556174 582134 591618
rect 581514 555938 581546 556174
rect 581782 555938 581866 556174
rect 582102 555938 582134 556174
rect 581514 555854 582134 555938
rect 581514 555618 581546 555854
rect 581782 555618 581866 555854
rect 582102 555618 582134 555854
rect 581514 520174 582134 555618
rect 581514 519938 581546 520174
rect 581782 519938 581866 520174
rect 582102 519938 582134 520174
rect 581514 519854 582134 519938
rect 581514 519618 581546 519854
rect 581782 519618 581866 519854
rect 582102 519618 582134 519854
rect 581514 484174 582134 519618
rect 581514 483938 581546 484174
rect 581782 483938 581866 484174
rect 582102 483938 582134 484174
rect 581514 483854 582134 483938
rect 581514 483618 581546 483854
rect 581782 483618 581866 483854
rect 582102 483618 582134 483854
rect 581514 448174 582134 483618
rect 581514 447938 581546 448174
rect 581782 447938 581866 448174
rect 582102 447938 582134 448174
rect 581514 447854 582134 447938
rect 581514 447618 581546 447854
rect 581782 447618 581866 447854
rect 582102 447618 582134 447854
rect 581514 412174 582134 447618
rect 581514 411938 581546 412174
rect 581782 411938 581866 412174
rect 582102 411938 582134 412174
rect 581514 411854 582134 411938
rect 581514 411618 581546 411854
rect 581782 411618 581866 411854
rect 582102 411618 582134 411854
rect 581514 376174 582134 411618
rect 581514 375938 581546 376174
rect 581782 375938 581866 376174
rect 582102 375938 582134 376174
rect 581514 375854 582134 375938
rect 581514 375618 581546 375854
rect 581782 375618 581866 375854
rect 582102 375618 582134 375854
rect 581514 340174 582134 375618
rect 581514 339938 581546 340174
rect 581782 339938 581866 340174
rect 582102 339938 582134 340174
rect 581514 339854 582134 339938
rect 581514 339618 581546 339854
rect 581782 339618 581866 339854
rect 582102 339618 582134 339854
rect 581514 304174 582134 339618
rect 581514 303938 581546 304174
rect 581782 303938 581866 304174
rect 582102 303938 582134 304174
rect 581514 303854 582134 303938
rect 581514 303618 581546 303854
rect 581782 303618 581866 303854
rect 582102 303618 582134 303854
rect 581514 268174 582134 303618
rect 581514 267938 581546 268174
rect 581782 267938 581866 268174
rect 582102 267938 582134 268174
rect 581514 267854 582134 267938
rect 581514 267618 581546 267854
rect 581782 267618 581866 267854
rect 582102 267618 582134 267854
rect 581514 232174 582134 267618
rect 581514 231938 581546 232174
rect 581782 231938 581866 232174
rect 582102 231938 582134 232174
rect 581514 231854 582134 231938
rect 581514 231618 581546 231854
rect 581782 231618 581866 231854
rect 582102 231618 582134 231854
rect 581514 196174 582134 231618
rect 581514 195938 581546 196174
rect 581782 195938 581866 196174
rect 582102 195938 582134 196174
rect 581514 195854 582134 195938
rect 581514 195618 581546 195854
rect 581782 195618 581866 195854
rect 582102 195618 582134 195854
rect 581514 160174 582134 195618
rect 581514 159938 581546 160174
rect 581782 159938 581866 160174
rect 582102 159938 582134 160174
rect 581514 159854 582134 159938
rect 581514 159618 581546 159854
rect 581782 159618 581866 159854
rect 582102 159618 582134 159854
rect 581514 124174 582134 159618
rect 581514 123938 581546 124174
rect 581782 123938 581866 124174
rect 582102 123938 582134 124174
rect 581514 123854 582134 123938
rect 581514 123618 581546 123854
rect 581782 123618 581866 123854
rect 582102 123618 582134 123854
rect 581514 88174 582134 123618
rect 581514 87938 581546 88174
rect 581782 87938 581866 88174
rect 582102 87938 582134 88174
rect 581514 87854 582134 87938
rect 581514 87618 581546 87854
rect 581782 87618 581866 87854
rect 582102 87618 582134 87854
rect 581514 52174 582134 87618
rect 581514 51938 581546 52174
rect 581782 51938 581866 52174
rect 582102 51938 582134 52174
rect 581514 51854 582134 51938
rect 581514 51618 581546 51854
rect 581782 51618 581866 51854
rect 582102 51618 582134 51854
rect 581514 16174 582134 51618
rect 581514 15938 581546 16174
rect 581782 15938 581866 16174
rect 582102 15938 582134 16174
rect 581514 15854 582134 15938
rect 581514 15618 581546 15854
rect 581782 15618 581866 15854
rect 582102 15618 582134 15854
rect 581514 -1306 582134 15618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 696454 585930 704282
rect 585310 696218 585342 696454
rect 585578 696218 585662 696454
rect 585898 696218 585930 696454
rect 585310 696134 585930 696218
rect 585310 695898 585342 696134
rect 585578 695898 585662 696134
rect 585898 695898 585930 696134
rect 585310 660454 585930 695898
rect 585310 660218 585342 660454
rect 585578 660218 585662 660454
rect 585898 660218 585930 660454
rect 585310 660134 585930 660218
rect 585310 659898 585342 660134
rect 585578 659898 585662 660134
rect 585898 659898 585930 660134
rect 585310 624454 585930 659898
rect 585310 624218 585342 624454
rect 585578 624218 585662 624454
rect 585898 624218 585930 624454
rect 585310 624134 585930 624218
rect 585310 623898 585342 624134
rect 585578 623898 585662 624134
rect 585898 623898 585930 624134
rect 585310 588454 585930 623898
rect 585310 588218 585342 588454
rect 585578 588218 585662 588454
rect 585898 588218 585930 588454
rect 585310 588134 585930 588218
rect 585310 587898 585342 588134
rect 585578 587898 585662 588134
rect 585898 587898 585930 588134
rect 585310 552454 585930 587898
rect 585310 552218 585342 552454
rect 585578 552218 585662 552454
rect 585898 552218 585930 552454
rect 585310 552134 585930 552218
rect 585310 551898 585342 552134
rect 585578 551898 585662 552134
rect 585898 551898 585930 552134
rect 585310 516454 585930 551898
rect 585310 516218 585342 516454
rect 585578 516218 585662 516454
rect 585898 516218 585930 516454
rect 585310 516134 585930 516218
rect 585310 515898 585342 516134
rect 585578 515898 585662 516134
rect 585898 515898 585930 516134
rect 585310 480454 585930 515898
rect 585310 480218 585342 480454
rect 585578 480218 585662 480454
rect 585898 480218 585930 480454
rect 585310 480134 585930 480218
rect 585310 479898 585342 480134
rect 585578 479898 585662 480134
rect 585898 479898 585930 480134
rect 585310 444454 585930 479898
rect 585310 444218 585342 444454
rect 585578 444218 585662 444454
rect 585898 444218 585930 444454
rect 585310 444134 585930 444218
rect 585310 443898 585342 444134
rect 585578 443898 585662 444134
rect 585898 443898 585930 444134
rect 585310 408454 585930 443898
rect 585310 408218 585342 408454
rect 585578 408218 585662 408454
rect 585898 408218 585930 408454
rect 585310 408134 585930 408218
rect 585310 407898 585342 408134
rect 585578 407898 585662 408134
rect 585898 407898 585930 408134
rect 585310 372454 585930 407898
rect 585310 372218 585342 372454
rect 585578 372218 585662 372454
rect 585898 372218 585930 372454
rect 585310 372134 585930 372218
rect 585310 371898 585342 372134
rect 585578 371898 585662 372134
rect 585898 371898 585930 372134
rect 585310 336454 585930 371898
rect 585310 336218 585342 336454
rect 585578 336218 585662 336454
rect 585898 336218 585930 336454
rect 585310 336134 585930 336218
rect 585310 335898 585342 336134
rect 585578 335898 585662 336134
rect 585898 335898 585930 336134
rect 585310 300454 585930 335898
rect 585310 300218 585342 300454
rect 585578 300218 585662 300454
rect 585898 300218 585930 300454
rect 585310 300134 585930 300218
rect 585310 299898 585342 300134
rect 585578 299898 585662 300134
rect 585898 299898 585930 300134
rect 585310 264454 585930 299898
rect 585310 264218 585342 264454
rect 585578 264218 585662 264454
rect 585898 264218 585930 264454
rect 585310 264134 585930 264218
rect 585310 263898 585342 264134
rect 585578 263898 585662 264134
rect 585898 263898 585930 264134
rect 585310 228454 585930 263898
rect 585310 228218 585342 228454
rect 585578 228218 585662 228454
rect 585898 228218 585930 228454
rect 585310 228134 585930 228218
rect 585310 227898 585342 228134
rect 585578 227898 585662 228134
rect 585898 227898 585930 228134
rect 585310 192454 585930 227898
rect 585310 192218 585342 192454
rect 585578 192218 585662 192454
rect 585898 192218 585930 192454
rect 585310 192134 585930 192218
rect 585310 191898 585342 192134
rect 585578 191898 585662 192134
rect 585898 191898 585930 192134
rect 585310 156454 585930 191898
rect 585310 156218 585342 156454
rect 585578 156218 585662 156454
rect 585898 156218 585930 156454
rect 585310 156134 585930 156218
rect 585310 155898 585342 156134
rect 585578 155898 585662 156134
rect 585898 155898 585930 156134
rect 585310 120454 585930 155898
rect 585310 120218 585342 120454
rect 585578 120218 585662 120454
rect 585898 120218 585930 120454
rect 585310 120134 585930 120218
rect 585310 119898 585342 120134
rect 585578 119898 585662 120134
rect 585898 119898 585930 120134
rect 585310 84454 585930 119898
rect 585310 84218 585342 84454
rect 585578 84218 585662 84454
rect 585898 84218 585930 84454
rect 585310 84134 585930 84218
rect 585310 83898 585342 84134
rect 585578 83898 585662 84134
rect 585898 83898 585930 84134
rect 585310 48454 585930 83898
rect 585310 48218 585342 48454
rect 585578 48218 585662 48454
rect 585898 48218 585930 48454
rect 585310 48134 585930 48218
rect 585310 47898 585342 48134
rect 585578 47898 585662 48134
rect 585898 47898 585930 48134
rect 585310 12454 585930 47898
rect 585310 12218 585342 12454
rect 585578 12218 585662 12454
rect 585898 12218 585930 12454
rect 585310 12134 585930 12218
rect 585310 11898 585342 12134
rect 585578 11898 585662 12134
rect 585898 11898 585930 12134
rect 585310 -346 585930 11898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 700174 586890 705242
rect 586270 699938 586302 700174
rect 586538 699938 586622 700174
rect 586858 699938 586890 700174
rect 586270 699854 586890 699938
rect 586270 699618 586302 699854
rect 586538 699618 586622 699854
rect 586858 699618 586890 699854
rect 586270 664174 586890 699618
rect 586270 663938 586302 664174
rect 586538 663938 586622 664174
rect 586858 663938 586890 664174
rect 586270 663854 586890 663938
rect 586270 663618 586302 663854
rect 586538 663618 586622 663854
rect 586858 663618 586890 663854
rect 586270 628174 586890 663618
rect 586270 627938 586302 628174
rect 586538 627938 586622 628174
rect 586858 627938 586890 628174
rect 586270 627854 586890 627938
rect 586270 627618 586302 627854
rect 586538 627618 586622 627854
rect 586858 627618 586890 627854
rect 586270 592174 586890 627618
rect 586270 591938 586302 592174
rect 586538 591938 586622 592174
rect 586858 591938 586890 592174
rect 586270 591854 586890 591938
rect 586270 591618 586302 591854
rect 586538 591618 586622 591854
rect 586858 591618 586890 591854
rect 586270 556174 586890 591618
rect 586270 555938 586302 556174
rect 586538 555938 586622 556174
rect 586858 555938 586890 556174
rect 586270 555854 586890 555938
rect 586270 555618 586302 555854
rect 586538 555618 586622 555854
rect 586858 555618 586890 555854
rect 586270 520174 586890 555618
rect 586270 519938 586302 520174
rect 586538 519938 586622 520174
rect 586858 519938 586890 520174
rect 586270 519854 586890 519938
rect 586270 519618 586302 519854
rect 586538 519618 586622 519854
rect 586858 519618 586890 519854
rect 586270 484174 586890 519618
rect 586270 483938 586302 484174
rect 586538 483938 586622 484174
rect 586858 483938 586890 484174
rect 586270 483854 586890 483938
rect 586270 483618 586302 483854
rect 586538 483618 586622 483854
rect 586858 483618 586890 483854
rect 586270 448174 586890 483618
rect 586270 447938 586302 448174
rect 586538 447938 586622 448174
rect 586858 447938 586890 448174
rect 586270 447854 586890 447938
rect 586270 447618 586302 447854
rect 586538 447618 586622 447854
rect 586858 447618 586890 447854
rect 586270 412174 586890 447618
rect 586270 411938 586302 412174
rect 586538 411938 586622 412174
rect 586858 411938 586890 412174
rect 586270 411854 586890 411938
rect 586270 411618 586302 411854
rect 586538 411618 586622 411854
rect 586858 411618 586890 411854
rect 586270 376174 586890 411618
rect 586270 375938 586302 376174
rect 586538 375938 586622 376174
rect 586858 375938 586890 376174
rect 586270 375854 586890 375938
rect 586270 375618 586302 375854
rect 586538 375618 586622 375854
rect 586858 375618 586890 375854
rect 586270 340174 586890 375618
rect 586270 339938 586302 340174
rect 586538 339938 586622 340174
rect 586858 339938 586890 340174
rect 586270 339854 586890 339938
rect 586270 339618 586302 339854
rect 586538 339618 586622 339854
rect 586858 339618 586890 339854
rect 586270 304174 586890 339618
rect 586270 303938 586302 304174
rect 586538 303938 586622 304174
rect 586858 303938 586890 304174
rect 586270 303854 586890 303938
rect 586270 303618 586302 303854
rect 586538 303618 586622 303854
rect 586858 303618 586890 303854
rect 586270 268174 586890 303618
rect 586270 267938 586302 268174
rect 586538 267938 586622 268174
rect 586858 267938 586890 268174
rect 586270 267854 586890 267938
rect 586270 267618 586302 267854
rect 586538 267618 586622 267854
rect 586858 267618 586890 267854
rect 586270 232174 586890 267618
rect 586270 231938 586302 232174
rect 586538 231938 586622 232174
rect 586858 231938 586890 232174
rect 586270 231854 586890 231938
rect 586270 231618 586302 231854
rect 586538 231618 586622 231854
rect 586858 231618 586890 231854
rect 586270 196174 586890 231618
rect 586270 195938 586302 196174
rect 586538 195938 586622 196174
rect 586858 195938 586890 196174
rect 586270 195854 586890 195938
rect 586270 195618 586302 195854
rect 586538 195618 586622 195854
rect 586858 195618 586890 195854
rect 586270 160174 586890 195618
rect 586270 159938 586302 160174
rect 586538 159938 586622 160174
rect 586858 159938 586890 160174
rect 586270 159854 586890 159938
rect 586270 159618 586302 159854
rect 586538 159618 586622 159854
rect 586858 159618 586890 159854
rect 586270 124174 586890 159618
rect 586270 123938 586302 124174
rect 586538 123938 586622 124174
rect 586858 123938 586890 124174
rect 586270 123854 586890 123938
rect 586270 123618 586302 123854
rect 586538 123618 586622 123854
rect 586858 123618 586890 123854
rect 586270 88174 586890 123618
rect 586270 87938 586302 88174
rect 586538 87938 586622 88174
rect 586858 87938 586890 88174
rect 586270 87854 586890 87938
rect 586270 87618 586302 87854
rect 586538 87618 586622 87854
rect 586858 87618 586890 87854
rect 586270 52174 586890 87618
rect 586270 51938 586302 52174
rect 586538 51938 586622 52174
rect 586858 51938 586890 52174
rect 586270 51854 586890 51938
rect 586270 51618 586302 51854
rect 586538 51618 586622 51854
rect 586858 51618 586890 51854
rect 586270 16174 586890 51618
rect 586270 15938 586302 16174
rect 586538 15938 586622 16174
rect 586858 15938 586890 16174
rect 586270 15854 586890 15938
rect 586270 15618 586302 15854
rect 586538 15618 586622 15854
rect 586858 15618 586890 15854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 15618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 -2266 587850 706202
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 -3226 588810 707162
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 -4186 589770 708122
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 -5146 590730 709082
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 -6106 591690 710042
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 -7066 592650 711002
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 699938 -2698 700174
rect -2614 699938 -2378 700174
rect -2934 699618 -2698 699854
rect -2614 699618 -2378 699854
rect -2934 663938 -2698 664174
rect -2614 663938 -2378 664174
rect -2934 663618 -2698 663854
rect -2614 663618 -2378 663854
rect -2934 627938 -2698 628174
rect -2614 627938 -2378 628174
rect -2934 627618 -2698 627854
rect -2614 627618 -2378 627854
rect -2934 591938 -2698 592174
rect -2614 591938 -2378 592174
rect -2934 591618 -2698 591854
rect -2614 591618 -2378 591854
rect -2934 555938 -2698 556174
rect -2614 555938 -2378 556174
rect -2934 555618 -2698 555854
rect -2614 555618 -2378 555854
rect -2934 519938 -2698 520174
rect -2614 519938 -2378 520174
rect -2934 519618 -2698 519854
rect -2614 519618 -2378 519854
rect -2934 483938 -2698 484174
rect -2614 483938 -2378 484174
rect -2934 483618 -2698 483854
rect -2614 483618 -2378 483854
rect -2934 447938 -2698 448174
rect -2614 447938 -2378 448174
rect -2934 447618 -2698 447854
rect -2614 447618 -2378 447854
rect -2934 411938 -2698 412174
rect -2614 411938 -2378 412174
rect -2934 411618 -2698 411854
rect -2614 411618 -2378 411854
rect -2934 375938 -2698 376174
rect -2614 375938 -2378 376174
rect -2934 375618 -2698 375854
rect -2614 375618 -2378 375854
rect -2934 339938 -2698 340174
rect -2614 339938 -2378 340174
rect -2934 339618 -2698 339854
rect -2614 339618 -2378 339854
rect -2934 303938 -2698 304174
rect -2614 303938 -2378 304174
rect -2934 303618 -2698 303854
rect -2614 303618 -2378 303854
rect -2934 267938 -2698 268174
rect -2614 267938 -2378 268174
rect -2934 267618 -2698 267854
rect -2614 267618 -2378 267854
rect -2934 231938 -2698 232174
rect -2614 231938 -2378 232174
rect -2934 231618 -2698 231854
rect -2614 231618 -2378 231854
rect -2934 195938 -2698 196174
rect -2614 195938 -2378 196174
rect -2934 195618 -2698 195854
rect -2614 195618 -2378 195854
rect -2934 159938 -2698 160174
rect -2614 159938 -2378 160174
rect -2934 159618 -2698 159854
rect -2614 159618 -2378 159854
rect -2934 123938 -2698 124174
rect -2614 123938 -2378 124174
rect -2934 123618 -2698 123854
rect -2614 123618 -2378 123854
rect -2934 87938 -2698 88174
rect -2614 87938 -2378 88174
rect -2934 87618 -2698 87854
rect -2614 87618 -2378 87854
rect -2934 51938 -2698 52174
rect -2614 51938 -2378 52174
rect -2934 51618 -2698 51854
rect -2614 51618 -2378 51854
rect -2934 15938 -2698 16174
rect -2614 15938 -2378 16174
rect -2934 15618 -2698 15854
rect -2614 15618 -2378 15854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 696218 -1738 696454
rect -1654 696218 -1418 696454
rect -1974 695898 -1738 696134
rect -1654 695898 -1418 696134
rect -1974 660218 -1738 660454
rect -1654 660218 -1418 660454
rect -1974 659898 -1738 660134
rect -1654 659898 -1418 660134
rect -1974 624218 -1738 624454
rect -1654 624218 -1418 624454
rect -1974 623898 -1738 624134
rect -1654 623898 -1418 624134
rect -1974 588218 -1738 588454
rect -1654 588218 -1418 588454
rect -1974 587898 -1738 588134
rect -1654 587898 -1418 588134
rect -1974 552218 -1738 552454
rect -1654 552218 -1418 552454
rect -1974 551898 -1738 552134
rect -1654 551898 -1418 552134
rect -1974 516218 -1738 516454
rect -1654 516218 -1418 516454
rect -1974 515898 -1738 516134
rect -1654 515898 -1418 516134
rect -1974 480218 -1738 480454
rect -1654 480218 -1418 480454
rect -1974 479898 -1738 480134
rect -1654 479898 -1418 480134
rect -1974 444218 -1738 444454
rect -1654 444218 -1418 444454
rect -1974 443898 -1738 444134
rect -1654 443898 -1418 444134
rect -1974 408218 -1738 408454
rect -1654 408218 -1418 408454
rect -1974 407898 -1738 408134
rect -1654 407898 -1418 408134
rect -1974 372218 -1738 372454
rect -1654 372218 -1418 372454
rect -1974 371898 -1738 372134
rect -1654 371898 -1418 372134
rect -1974 336218 -1738 336454
rect -1654 336218 -1418 336454
rect -1974 335898 -1738 336134
rect -1654 335898 -1418 336134
rect -1974 300218 -1738 300454
rect -1654 300218 -1418 300454
rect -1974 299898 -1738 300134
rect -1654 299898 -1418 300134
rect -1974 264218 -1738 264454
rect -1654 264218 -1418 264454
rect -1974 263898 -1738 264134
rect -1654 263898 -1418 264134
rect -1974 228218 -1738 228454
rect -1654 228218 -1418 228454
rect -1974 227898 -1738 228134
rect -1654 227898 -1418 228134
rect -1974 192218 -1738 192454
rect -1654 192218 -1418 192454
rect -1974 191898 -1738 192134
rect -1654 191898 -1418 192134
rect -1974 156218 -1738 156454
rect -1654 156218 -1418 156454
rect -1974 155898 -1738 156134
rect -1654 155898 -1418 156134
rect -1974 120218 -1738 120454
rect -1654 120218 -1418 120454
rect -1974 119898 -1738 120134
rect -1654 119898 -1418 120134
rect -1974 84218 -1738 84454
rect -1654 84218 -1418 84454
rect -1974 83898 -1738 84134
rect -1654 83898 -1418 84134
rect -1974 48218 -1738 48454
rect -1654 48218 -1418 48454
rect -1974 47898 -1738 48134
rect -1654 47898 -1418 48134
rect -1974 12218 -1738 12454
rect -1654 12218 -1418 12454
rect -1974 11898 -1738 12134
rect -1654 11898 -1418 12134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 699849 5782 700085
rect 5866 699849 6102 700085
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 699849 41782 700085
rect 41866 699849 42102 700085
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 699849 77782 700085
rect 77866 699849 78102 700085
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 699849 113782 700085
rect 113866 699849 114102 700085
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 699849 149782 700085
rect 149866 699849 150102 700085
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 699849 185782 700085
rect 185866 699849 186102 700085
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 699849 221782 700085
rect 221866 699849 222102 700085
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 699849 257782 700085
rect 257866 699849 258102 700085
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 699849 293782 700085
rect 293866 699849 294102 700085
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 699849 329782 700085
rect 329866 699849 330102 700085
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 699849 365782 700085
rect 365866 699849 366102 700085
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 699849 401782 700085
rect 401866 699849 402102 700085
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 699849 437782 700085
rect 437866 699849 438102 700085
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 699849 473782 700085
rect 473866 699849 474102 700085
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 699849 509782 700085
rect 509866 699849 510102 700085
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 699849 545782 700085
rect 545866 699849 546102 700085
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 1826 696218 2062 696454
rect 2146 696218 2382 696454
rect 1826 695898 2062 696134
rect 2146 695898 2382 696134
rect 5826 696218 6062 696454
rect 6146 696218 6382 696454
rect 5826 695898 6062 696134
rect 6146 695898 6382 696134
rect 41826 696218 42062 696454
rect 42146 696218 42382 696454
rect 41826 695898 42062 696134
rect 42146 695898 42382 696134
rect 77826 696218 78062 696454
rect 78146 696218 78382 696454
rect 77826 695898 78062 696134
rect 78146 695898 78382 696134
rect 113826 696218 114062 696454
rect 114146 696218 114382 696454
rect 113826 695898 114062 696134
rect 114146 695898 114382 696134
rect 149826 696218 150062 696454
rect 150146 696218 150382 696454
rect 149826 695898 150062 696134
rect 150146 695898 150382 696134
rect 185826 696218 186062 696454
rect 186146 696218 186382 696454
rect 185826 695898 186062 696134
rect 186146 695898 186382 696134
rect 221826 696218 222062 696454
rect 222146 696218 222382 696454
rect 221826 695898 222062 696134
rect 222146 695898 222382 696134
rect 257826 696218 258062 696454
rect 258146 696218 258382 696454
rect 257826 695898 258062 696134
rect 258146 695898 258382 696134
rect 293826 696218 294062 696454
rect 294146 696218 294382 696454
rect 293826 695898 294062 696134
rect 294146 695898 294382 696134
rect 329826 696218 330062 696454
rect 330146 696218 330382 696454
rect 329826 695898 330062 696134
rect 330146 695898 330382 696134
rect 365826 696218 366062 696454
rect 366146 696218 366382 696454
rect 365826 695898 366062 696134
rect 366146 695898 366382 696134
rect 401826 696218 402062 696454
rect 402146 696218 402382 696454
rect 401826 695898 402062 696134
rect 402146 695898 402382 696134
rect 437826 696218 438062 696454
rect 438146 696218 438382 696454
rect 437826 695898 438062 696134
rect 438146 695898 438382 696134
rect 473826 696218 474062 696454
rect 474146 696218 474382 696454
rect 473826 695898 474062 696134
rect 474146 695898 474382 696134
rect 509826 696218 510062 696454
rect 510146 696218 510382 696454
rect 509826 695898 510062 696134
rect 510146 695898 510382 696134
rect 545826 696218 546062 696454
rect 546146 696218 546382 696454
rect 545826 695898 546062 696134
rect 546146 695898 546382 696134
rect 577826 696218 578062 696454
rect 578146 696218 578382 696454
rect 577826 695898 578062 696134
rect 578146 695898 578382 696134
rect 9546 663938 9782 664174
rect 9866 663938 10102 664174
rect 9546 663618 9782 663854
rect 9866 663618 10102 663854
rect 189546 663938 189782 664174
rect 189866 663938 190102 664174
rect 189546 663618 189782 663854
rect 189866 663618 190102 663854
rect 369546 663938 369782 664174
rect 369866 663938 370102 664174
rect 369546 663618 369782 663854
rect 369866 663618 370102 663854
rect 405546 663938 405782 664174
rect 405866 663938 406102 664174
rect 405546 663618 405782 663854
rect 405866 663618 406102 663854
rect 572374 663938 572610 664174
rect 572694 663938 572930 664174
rect 572374 663618 572610 663854
rect 572694 663618 572930 663854
rect 1826 660218 2062 660454
rect 2146 660218 2382 660454
rect 1826 659898 2062 660134
rect 2146 659898 2382 660134
rect 5826 660218 6062 660454
rect 6146 660218 6382 660454
rect 5826 659898 6062 660134
rect 6146 659898 6382 660134
rect 185826 660218 186062 660454
rect 186146 660218 186382 660454
rect 185826 659898 186062 660134
rect 186146 659898 186382 660134
rect 365826 660218 366062 660454
rect 366146 660218 366382 660454
rect 365826 659898 366062 660134
rect 366146 659898 366382 660134
rect 401826 660218 402062 660454
rect 402146 660218 402382 660454
rect 401826 659898 402062 660134
rect 402146 659898 402382 660134
rect 568510 660218 568746 660454
rect 568830 660218 569066 660454
rect 568510 659898 568746 660134
rect 568830 659898 569066 660134
rect 577826 660218 578062 660454
rect 578146 660218 578382 660454
rect 577826 659898 578062 660134
rect 578146 659898 578382 660134
rect 9546 627938 9782 628174
rect 9866 627938 10102 628174
rect 9546 627618 9782 627854
rect 9866 627618 10102 627854
rect 189546 627938 189782 628174
rect 189866 627938 190102 628174
rect 189546 627618 189782 627854
rect 189866 627618 190102 627854
rect 369546 627938 369782 628174
rect 369866 627938 370102 628174
rect 369546 627618 369782 627854
rect 369866 627618 370102 627854
rect 405546 627938 405782 628174
rect 405866 627938 406102 628174
rect 405546 627618 405782 627854
rect 405866 627618 406102 627854
rect 572374 627938 572610 628174
rect 572694 627938 572930 628174
rect 572374 627618 572610 627854
rect 572694 627618 572930 627854
rect 1826 624218 2062 624454
rect 2146 624218 2382 624454
rect 1826 623898 2062 624134
rect 2146 623898 2382 624134
rect 5826 624218 6062 624454
rect 6146 624218 6382 624454
rect 5826 623898 6062 624134
rect 6146 623898 6382 624134
rect 185826 624218 186062 624454
rect 186146 624218 186382 624454
rect 185826 623898 186062 624134
rect 186146 623898 186382 624134
rect 365826 624218 366062 624454
rect 366146 624218 366382 624454
rect 365826 623898 366062 624134
rect 366146 623898 366382 624134
rect 401826 624218 402062 624454
rect 402146 624218 402382 624454
rect 401826 623898 402062 624134
rect 402146 623898 402382 624134
rect 568510 624218 568746 624454
rect 568830 624218 569066 624454
rect 568510 623898 568746 624134
rect 568830 623898 569066 624134
rect 577826 624218 578062 624454
rect 578146 624218 578382 624454
rect 577826 623898 578062 624134
rect 578146 623898 578382 624134
rect 9546 591938 9782 592174
rect 9866 591938 10102 592174
rect 9546 591618 9782 591854
rect 9866 591618 10102 591854
rect 45546 591938 45782 592174
rect 45866 591938 46102 592174
rect 45546 591618 45782 591854
rect 45866 591618 46102 591854
rect 81546 591938 81782 592174
rect 81866 591938 82102 592174
rect 81546 591618 81782 591854
rect 81866 591618 82102 591854
rect 117546 591938 117782 592174
rect 117866 591938 118102 592174
rect 117546 591618 117782 591854
rect 117866 591618 118102 591854
rect 153546 591938 153782 592174
rect 153866 591938 154102 592174
rect 153546 591618 153782 591854
rect 153866 591618 154102 591854
rect 189546 591938 189782 592174
rect 189866 591938 190102 592174
rect 189546 591618 189782 591854
rect 189866 591618 190102 591854
rect 225546 591938 225782 592174
rect 225866 591938 226102 592174
rect 225546 591618 225782 591854
rect 225866 591618 226102 591854
rect 261546 591938 261782 592174
rect 261866 591938 262102 592174
rect 261546 591618 261782 591854
rect 261866 591618 262102 591854
rect 297546 591938 297782 592174
rect 297866 591938 298102 592174
rect 297546 591618 297782 591854
rect 297866 591618 298102 591854
rect 333546 591938 333782 592174
rect 333866 591938 334102 592174
rect 333546 591618 333782 591854
rect 333866 591618 334102 591854
rect 369546 591938 369782 592174
rect 369866 591938 370102 592174
rect 369546 591618 369782 591854
rect 369866 591618 370102 591854
rect 405546 591938 405782 592174
rect 405866 591938 406102 592174
rect 405546 591618 405782 591854
rect 405866 591618 406102 591854
rect 441546 591938 441782 592174
rect 441866 591938 442102 592174
rect 441546 591618 441782 591854
rect 441866 591618 442102 591854
rect 477546 591938 477782 592174
rect 477866 591938 478102 592174
rect 477546 591618 477782 591854
rect 477866 591618 478102 591854
rect 513546 591938 513782 592174
rect 513866 591938 514102 592174
rect 513546 591618 513782 591854
rect 513866 591618 514102 591854
rect 549546 591938 549782 592174
rect 549866 591938 550102 592174
rect 549546 591618 549782 591854
rect 549866 591618 550102 591854
rect 1826 588218 2062 588454
rect 2146 588218 2382 588454
rect 1826 587898 2062 588134
rect 2146 587898 2382 588134
rect 5826 588218 6062 588454
rect 6146 588218 6382 588454
rect 5826 587898 6062 588134
rect 6146 587898 6382 588134
rect 41826 588218 42062 588454
rect 42146 588218 42382 588454
rect 41826 587898 42062 588134
rect 42146 587898 42382 588134
rect 77826 588218 78062 588454
rect 78146 588218 78382 588454
rect 77826 587898 78062 588134
rect 78146 587898 78382 588134
rect 113826 588218 114062 588454
rect 114146 588218 114382 588454
rect 113826 587898 114062 588134
rect 114146 587898 114382 588134
rect 149826 588218 150062 588454
rect 150146 588218 150382 588454
rect 149826 587898 150062 588134
rect 150146 587898 150382 588134
rect 185826 588218 186062 588454
rect 186146 588218 186382 588454
rect 185826 587898 186062 588134
rect 186146 587898 186382 588134
rect 221826 588218 222062 588454
rect 222146 588218 222382 588454
rect 221826 587898 222062 588134
rect 222146 587898 222382 588134
rect 257826 588218 258062 588454
rect 258146 588218 258382 588454
rect 257826 587898 258062 588134
rect 258146 587898 258382 588134
rect 293826 588218 294062 588454
rect 294146 588218 294382 588454
rect 293826 587898 294062 588134
rect 294146 587898 294382 588134
rect 329826 588218 330062 588454
rect 330146 588218 330382 588454
rect 329826 587898 330062 588134
rect 330146 587898 330382 588134
rect 365826 588218 366062 588454
rect 366146 588218 366382 588454
rect 365826 587898 366062 588134
rect 366146 587898 366382 588134
rect 401826 588218 402062 588454
rect 402146 588218 402382 588454
rect 401826 587898 402062 588134
rect 402146 587898 402382 588134
rect 437826 588218 438062 588454
rect 438146 588218 438382 588454
rect 437826 587898 438062 588134
rect 438146 587898 438382 588134
rect 473826 588218 474062 588454
rect 474146 588218 474382 588454
rect 473826 587898 474062 588134
rect 474146 587898 474382 588134
rect 509826 588218 510062 588454
rect 510146 588218 510382 588454
rect 509826 587898 510062 588134
rect 510146 587898 510382 588134
rect 545826 588218 546062 588454
rect 546146 588218 546382 588454
rect 545826 587898 546062 588134
rect 546146 587898 546382 588134
rect 577826 588218 578062 588454
rect 578146 588218 578382 588454
rect 577826 587898 578062 588134
rect 578146 587898 578382 588134
rect 9546 555938 9782 556174
rect 9866 555938 10102 556174
rect 9546 555618 9782 555854
rect 9866 555618 10102 555854
rect 189546 555938 189782 556174
rect 189866 555938 190102 556174
rect 189546 555618 189782 555854
rect 189866 555618 190102 555854
rect 225546 555938 225782 556174
rect 225866 555938 226102 556174
rect 225546 555618 225782 555854
rect 225866 555618 226102 555854
rect 261546 555938 261782 556174
rect 261866 555938 262102 556174
rect 261546 555618 261782 555854
rect 261866 555618 262102 555854
rect 297546 555938 297782 556174
rect 297866 555938 298102 556174
rect 297546 555618 297782 555854
rect 297866 555618 298102 555854
rect 333546 555938 333782 556174
rect 333866 555938 334102 556174
rect 333546 555618 333782 555854
rect 333866 555618 334102 555854
rect 369546 555938 369782 556174
rect 369866 555938 370102 556174
rect 369546 555618 369782 555854
rect 369866 555618 370102 555854
rect 405546 555938 405782 556174
rect 405866 555938 406102 556174
rect 405546 555618 405782 555854
rect 405866 555618 406102 555854
rect 572374 555938 572610 556174
rect 572694 555938 572930 556174
rect 572374 555618 572610 555854
rect 572694 555618 572930 555854
rect 1826 552218 2062 552454
rect 2146 552218 2382 552454
rect 1826 551898 2062 552134
rect 2146 551898 2382 552134
rect 5826 552218 6062 552454
rect 6146 552218 6382 552454
rect 5826 551898 6062 552134
rect 6146 551898 6382 552134
rect 185826 552218 186062 552454
rect 186146 552218 186382 552454
rect 185826 551898 186062 552134
rect 186146 551898 186382 552134
rect 221826 552218 222062 552454
rect 222146 552218 222382 552454
rect 221826 551898 222062 552134
rect 222146 551898 222382 552134
rect 257826 552218 258062 552454
rect 258146 552218 258382 552454
rect 257826 551898 258062 552134
rect 258146 551898 258382 552134
rect 293826 552218 294062 552454
rect 294146 552218 294382 552454
rect 293826 551898 294062 552134
rect 294146 551898 294382 552134
rect 329826 552218 330062 552454
rect 330146 552218 330382 552454
rect 329826 551898 330062 552134
rect 330146 551898 330382 552134
rect 365826 552218 366062 552454
rect 366146 552218 366382 552454
rect 365826 551898 366062 552134
rect 366146 551898 366382 552134
rect 401826 552218 402062 552454
rect 402146 552218 402382 552454
rect 401826 551898 402062 552134
rect 402146 551898 402382 552134
rect 568510 552218 568746 552454
rect 568830 552218 569066 552454
rect 568510 551898 568746 552134
rect 568830 551898 569066 552134
rect 577826 552218 578062 552454
rect 578146 552218 578382 552454
rect 577826 551898 578062 552134
rect 578146 551898 578382 552134
rect 9546 519938 9782 520174
rect 9866 519938 10102 520174
rect 9546 519618 9782 519854
rect 9866 519618 10102 519854
rect 189546 519938 189782 520174
rect 189866 519938 190102 520174
rect 189546 519618 189782 519854
rect 189866 519618 190102 519854
rect 225546 519938 225782 520174
rect 225866 519938 226102 520174
rect 225546 519618 225782 519854
rect 225866 519618 226102 519854
rect 261546 519938 261782 520174
rect 261866 519938 262102 520174
rect 261546 519618 261782 519854
rect 261866 519618 262102 519854
rect 297546 519938 297782 520174
rect 297866 519938 298102 520174
rect 297546 519618 297782 519854
rect 297866 519618 298102 519854
rect 333546 519938 333782 520174
rect 333866 519938 334102 520174
rect 333546 519618 333782 519854
rect 333866 519618 334102 519854
rect 369546 519938 369782 520174
rect 369866 519938 370102 520174
rect 369546 519618 369782 519854
rect 369866 519618 370102 519854
rect 405546 519938 405782 520174
rect 405866 519938 406102 520174
rect 405546 519618 405782 519854
rect 405866 519618 406102 519854
rect 572374 519938 572610 520174
rect 572694 519938 572930 520174
rect 572374 519618 572610 519854
rect 572694 519618 572930 519854
rect 1826 516218 2062 516454
rect 2146 516218 2382 516454
rect 1826 515898 2062 516134
rect 2146 515898 2382 516134
rect 5826 516218 6062 516454
rect 6146 516218 6382 516454
rect 5826 515898 6062 516134
rect 6146 515898 6382 516134
rect 185826 516218 186062 516454
rect 186146 516218 186382 516454
rect 185826 515898 186062 516134
rect 186146 515898 186382 516134
rect 221826 516218 222062 516454
rect 222146 516218 222382 516454
rect 221826 515898 222062 516134
rect 222146 515898 222382 516134
rect 257826 516218 258062 516454
rect 258146 516218 258382 516454
rect 257826 515898 258062 516134
rect 258146 515898 258382 516134
rect 293826 516218 294062 516454
rect 294146 516218 294382 516454
rect 293826 515898 294062 516134
rect 294146 515898 294382 516134
rect 329826 516218 330062 516454
rect 330146 516218 330382 516454
rect 329826 515898 330062 516134
rect 330146 515898 330382 516134
rect 365826 516218 366062 516454
rect 366146 516218 366382 516454
rect 365826 515898 366062 516134
rect 366146 515898 366382 516134
rect 401826 516218 402062 516454
rect 402146 516218 402382 516454
rect 401826 515898 402062 516134
rect 402146 515898 402382 516134
rect 568510 516218 568746 516454
rect 568830 516218 569066 516454
rect 568510 515898 568746 516134
rect 568830 515898 569066 516134
rect 577826 516218 578062 516454
rect 578146 516218 578382 516454
rect 577826 515898 578062 516134
rect 578146 515898 578382 516134
rect 9546 483938 9782 484174
rect 9866 483938 10102 484174
rect 9546 483618 9782 483854
rect 9866 483618 10102 483854
rect 45546 483938 45782 484174
rect 45866 483938 46102 484174
rect 45546 483618 45782 483854
rect 45866 483618 46102 483854
rect 81546 483938 81782 484174
rect 81866 483938 82102 484174
rect 81546 483618 81782 483854
rect 81866 483618 82102 483854
rect 117546 483938 117782 484174
rect 117866 483938 118102 484174
rect 117546 483618 117782 483854
rect 117866 483618 118102 483854
rect 153546 483938 153782 484174
rect 153866 483938 154102 484174
rect 153546 483618 153782 483854
rect 153866 483618 154102 483854
rect 189546 483938 189782 484174
rect 189866 483938 190102 484174
rect 189546 483618 189782 483854
rect 189866 483618 190102 483854
rect 225546 483938 225782 484174
rect 225866 483938 226102 484174
rect 225546 483618 225782 483854
rect 225866 483618 226102 483854
rect 261546 483938 261782 484174
rect 261866 483938 262102 484174
rect 261546 483618 261782 483854
rect 261866 483618 262102 483854
rect 297546 483938 297782 484174
rect 297866 483938 298102 484174
rect 297546 483618 297782 483854
rect 297866 483618 298102 483854
rect 333546 483938 333782 484174
rect 333866 483938 334102 484174
rect 333546 483618 333782 483854
rect 333866 483618 334102 483854
rect 369546 483938 369782 484174
rect 369866 483938 370102 484174
rect 369546 483618 369782 483854
rect 369866 483618 370102 483854
rect 405546 483938 405782 484174
rect 405866 483938 406102 484174
rect 405546 483618 405782 483854
rect 405866 483618 406102 483854
rect 441546 483938 441782 484174
rect 441866 483938 442102 484174
rect 441546 483618 441782 483854
rect 441866 483618 442102 483854
rect 477546 483938 477782 484174
rect 477866 483938 478102 484174
rect 477546 483618 477782 483854
rect 477866 483618 478102 483854
rect 513546 483938 513782 484174
rect 513866 483938 514102 484174
rect 513546 483618 513782 483854
rect 513866 483618 514102 483854
rect 549546 483938 549782 484174
rect 549866 483938 550102 484174
rect 549546 483618 549782 483854
rect 549866 483618 550102 483854
rect 1826 480218 2062 480454
rect 2146 480218 2382 480454
rect 1826 479898 2062 480134
rect 2146 479898 2382 480134
rect 5826 480218 6062 480454
rect 6146 480218 6382 480454
rect 5826 479898 6062 480134
rect 6146 479898 6382 480134
rect 41826 480218 42062 480454
rect 42146 480218 42382 480454
rect 41826 479898 42062 480134
rect 42146 479898 42382 480134
rect 77826 480218 78062 480454
rect 78146 480218 78382 480454
rect 77826 479898 78062 480134
rect 78146 479898 78382 480134
rect 113826 480218 114062 480454
rect 114146 480218 114382 480454
rect 113826 479898 114062 480134
rect 114146 479898 114382 480134
rect 149826 480218 150062 480454
rect 150146 480218 150382 480454
rect 149826 479898 150062 480134
rect 150146 479898 150382 480134
rect 185826 480218 186062 480454
rect 186146 480218 186382 480454
rect 185826 479898 186062 480134
rect 186146 479898 186382 480134
rect 221826 480218 222062 480454
rect 222146 480218 222382 480454
rect 221826 479898 222062 480134
rect 222146 479898 222382 480134
rect 257826 480218 258062 480454
rect 258146 480218 258382 480454
rect 257826 479898 258062 480134
rect 258146 479898 258382 480134
rect 293826 480218 294062 480454
rect 294146 480218 294382 480454
rect 293826 479898 294062 480134
rect 294146 479898 294382 480134
rect 329826 480218 330062 480454
rect 330146 480218 330382 480454
rect 329826 479898 330062 480134
rect 330146 479898 330382 480134
rect 365826 480218 366062 480454
rect 366146 480218 366382 480454
rect 365826 479898 366062 480134
rect 366146 479898 366382 480134
rect 401826 480218 402062 480454
rect 402146 480218 402382 480454
rect 401826 479898 402062 480134
rect 402146 479898 402382 480134
rect 437826 480218 438062 480454
rect 438146 480218 438382 480454
rect 437826 479898 438062 480134
rect 438146 479898 438382 480134
rect 473826 480218 474062 480454
rect 474146 480218 474382 480454
rect 473826 479898 474062 480134
rect 474146 479898 474382 480134
rect 509826 480218 510062 480454
rect 510146 480218 510382 480454
rect 509826 479898 510062 480134
rect 510146 479898 510382 480134
rect 545826 480218 546062 480454
rect 546146 480218 546382 480454
rect 545826 479898 546062 480134
rect 546146 479898 546382 480134
rect 577826 480218 578062 480454
rect 578146 480218 578382 480454
rect 577826 479898 578062 480134
rect 578146 479898 578382 480134
rect 9546 447938 9782 448174
rect 9866 447938 10102 448174
rect 9546 447618 9782 447854
rect 9866 447618 10102 447854
rect 189546 447938 189782 448174
rect 189866 447938 190102 448174
rect 189546 447618 189782 447854
rect 189866 447618 190102 447854
rect 225546 447938 225782 448174
rect 225866 447938 226102 448174
rect 225546 447618 225782 447854
rect 225866 447618 226102 447854
rect 261546 447938 261782 448174
rect 261866 447938 262102 448174
rect 261546 447618 261782 447854
rect 261866 447618 262102 447854
rect 297546 447938 297782 448174
rect 297866 447938 298102 448174
rect 297546 447618 297782 447854
rect 297866 447618 298102 447854
rect 333546 447938 333782 448174
rect 333866 447938 334102 448174
rect 333546 447618 333782 447854
rect 333866 447618 334102 447854
rect 369546 447938 369782 448174
rect 369866 447938 370102 448174
rect 369546 447618 369782 447854
rect 369866 447618 370102 447854
rect 405546 447938 405782 448174
rect 405866 447938 406102 448174
rect 405546 447618 405782 447854
rect 405866 447618 406102 447854
rect 572374 447938 572610 448174
rect 572694 447938 572930 448174
rect 572374 447618 572610 447854
rect 572694 447618 572930 447854
rect 1826 444218 2062 444454
rect 2146 444218 2382 444454
rect 1826 443898 2062 444134
rect 2146 443898 2382 444134
rect 5826 444218 6062 444454
rect 6146 444218 6382 444454
rect 5826 443898 6062 444134
rect 6146 443898 6382 444134
rect 185826 444218 186062 444454
rect 186146 444218 186382 444454
rect 185826 443898 186062 444134
rect 186146 443898 186382 444134
rect 221826 444218 222062 444454
rect 222146 444218 222382 444454
rect 221826 443898 222062 444134
rect 222146 443898 222382 444134
rect 257826 444218 258062 444454
rect 258146 444218 258382 444454
rect 257826 443898 258062 444134
rect 258146 443898 258382 444134
rect 293826 444218 294062 444454
rect 294146 444218 294382 444454
rect 293826 443898 294062 444134
rect 294146 443898 294382 444134
rect 329826 444218 330062 444454
rect 330146 444218 330382 444454
rect 329826 443898 330062 444134
rect 330146 443898 330382 444134
rect 365826 444218 366062 444454
rect 366146 444218 366382 444454
rect 365826 443898 366062 444134
rect 366146 443898 366382 444134
rect 401826 444218 402062 444454
rect 402146 444218 402382 444454
rect 401826 443898 402062 444134
rect 402146 443898 402382 444134
rect 568510 444218 568746 444454
rect 568830 444218 569066 444454
rect 568510 443898 568746 444134
rect 568830 443898 569066 444134
rect 577826 444218 578062 444454
rect 578146 444218 578382 444454
rect 577826 443898 578062 444134
rect 578146 443898 578382 444134
rect 9546 411938 9782 412174
rect 9866 411938 10102 412174
rect 9546 411618 9782 411854
rect 9866 411618 10102 411854
rect 189546 411938 189782 412174
rect 189866 411938 190102 412174
rect 189546 411618 189782 411854
rect 189866 411618 190102 411854
rect 225546 411938 225782 412174
rect 225866 411938 226102 412174
rect 225546 411618 225782 411854
rect 225866 411618 226102 411854
rect 261546 411938 261782 412174
rect 261866 411938 262102 412174
rect 261546 411618 261782 411854
rect 261866 411618 262102 411854
rect 297546 411938 297782 412174
rect 297866 411938 298102 412174
rect 297546 411618 297782 411854
rect 297866 411618 298102 411854
rect 333546 411938 333782 412174
rect 333866 411938 334102 412174
rect 333546 411618 333782 411854
rect 333866 411618 334102 411854
rect 369546 411938 369782 412174
rect 369866 411938 370102 412174
rect 369546 411618 369782 411854
rect 369866 411618 370102 411854
rect 405546 411938 405782 412174
rect 405866 411938 406102 412174
rect 405546 411618 405782 411854
rect 405866 411618 406102 411854
rect 572374 411938 572610 412174
rect 572694 411938 572930 412174
rect 572374 411618 572610 411854
rect 572694 411618 572930 411854
rect 1826 408218 2062 408454
rect 2146 408218 2382 408454
rect 1826 407898 2062 408134
rect 2146 407898 2382 408134
rect 5826 408218 6062 408454
rect 6146 408218 6382 408454
rect 5826 407898 6062 408134
rect 6146 407898 6382 408134
rect 185826 408218 186062 408454
rect 186146 408218 186382 408454
rect 185826 407898 186062 408134
rect 186146 407898 186382 408134
rect 221826 408218 222062 408454
rect 222146 408218 222382 408454
rect 221826 407898 222062 408134
rect 222146 407898 222382 408134
rect 257826 408218 258062 408454
rect 258146 408218 258382 408454
rect 257826 407898 258062 408134
rect 258146 407898 258382 408134
rect 293826 408218 294062 408454
rect 294146 408218 294382 408454
rect 293826 407898 294062 408134
rect 294146 407898 294382 408134
rect 329826 408218 330062 408454
rect 330146 408218 330382 408454
rect 329826 407898 330062 408134
rect 330146 407898 330382 408134
rect 365826 408218 366062 408454
rect 366146 408218 366382 408454
rect 365826 407898 366062 408134
rect 366146 407898 366382 408134
rect 401826 408218 402062 408454
rect 402146 408218 402382 408454
rect 401826 407898 402062 408134
rect 402146 407898 402382 408134
rect 568510 408218 568746 408454
rect 568830 408218 569066 408454
rect 568510 407898 568746 408134
rect 568830 407898 569066 408134
rect 577826 408218 578062 408454
rect 578146 408218 578382 408454
rect 577826 407898 578062 408134
rect 578146 407898 578382 408134
rect 9546 375938 9782 376174
rect 9866 375938 10102 376174
rect 9546 375618 9782 375854
rect 9866 375618 10102 375854
rect 189546 375938 189782 376174
rect 189866 375938 190102 376174
rect 189546 375618 189782 375854
rect 189866 375618 190102 375854
rect 225546 375938 225782 376174
rect 225866 375938 226102 376174
rect 225546 375618 225782 375854
rect 225866 375618 226102 375854
rect 261546 375938 261782 376174
rect 261866 375938 262102 376174
rect 261546 375618 261782 375854
rect 261866 375618 262102 375854
rect 297546 375938 297782 376174
rect 297866 375938 298102 376174
rect 297546 375618 297782 375854
rect 297866 375618 298102 375854
rect 333546 375938 333782 376174
rect 333866 375938 334102 376174
rect 333546 375618 333782 375854
rect 333866 375618 334102 375854
rect 369546 375938 369782 376174
rect 369866 375938 370102 376174
rect 369546 375618 369782 375854
rect 369866 375618 370102 375854
rect 405546 375938 405782 376174
rect 405866 375938 406102 376174
rect 405546 375618 405782 375854
rect 405866 375618 406102 375854
rect 572374 375938 572610 376174
rect 572694 375938 572930 376174
rect 572374 375618 572610 375854
rect 572694 375618 572930 375854
rect 1826 372218 2062 372454
rect 2146 372218 2382 372454
rect 1826 371898 2062 372134
rect 2146 371898 2382 372134
rect 5826 372218 6062 372454
rect 6146 372218 6382 372454
rect 5826 371898 6062 372134
rect 6146 371898 6382 372134
rect 185826 372218 186062 372454
rect 186146 372218 186382 372454
rect 185826 371898 186062 372134
rect 186146 371898 186382 372134
rect 221826 372218 222062 372454
rect 222146 372218 222382 372454
rect 221826 371898 222062 372134
rect 222146 371898 222382 372134
rect 257826 372218 258062 372454
rect 258146 372218 258382 372454
rect 257826 371898 258062 372134
rect 258146 371898 258382 372134
rect 293826 372218 294062 372454
rect 294146 372218 294382 372454
rect 293826 371898 294062 372134
rect 294146 371898 294382 372134
rect 329826 372218 330062 372454
rect 330146 372218 330382 372454
rect 329826 371898 330062 372134
rect 330146 371898 330382 372134
rect 365826 372218 366062 372454
rect 366146 372218 366382 372454
rect 365826 371898 366062 372134
rect 366146 371898 366382 372134
rect 401826 372218 402062 372454
rect 402146 372218 402382 372454
rect 401826 371898 402062 372134
rect 402146 371898 402382 372134
rect 568510 372218 568746 372454
rect 568830 372218 569066 372454
rect 568510 371898 568746 372134
rect 568830 371898 569066 372134
rect 577826 372218 578062 372454
rect 578146 372218 578382 372454
rect 577826 371898 578062 372134
rect 578146 371898 578382 372134
rect 9546 339938 9782 340174
rect 9866 339938 10102 340174
rect 9546 339618 9782 339854
rect 9866 339618 10102 339854
rect 189546 339938 189782 340174
rect 189866 339938 190102 340174
rect 189546 339618 189782 339854
rect 189866 339618 190102 339854
rect 225546 339938 225782 340174
rect 225866 339938 226102 340174
rect 225546 339618 225782 339854
rect 225866 339618 226102 339854
rect 261546 339938 261782 340174
rect 261866 339938 262102 340174
rect 261546 339618 261782 339854
rect 261866 339618 262102 339854
rect 297546 339938 297782 340174
rect 297866 339938 298102 340174
rect 297546 339618 297782 339854
rect 297866 339618 298102 339854
rect 333546 339938 333782 340174
rect 333866 339938 334102 340174
rect 333546 339618 333782 339854
rect 333866 339618 334102 339854
rect 369546 339938 369782 340174
rect 369866 339938 370102 340174
rect 369546 339618 369782 339854
rect 369866 339618 370102 339854
rect 405546 339938 405782 340174
rect 405866 339938 406102 340174
rect 405546 339618 405782 339854
rect 405866 339618 406102 339854
rect 572374 339938 572610 340174
rect 572694 339938 572930 340174
rect 572374 339618 572610 339854
rect 572694 339618 572930 339854
rect 1826 336218 2062 336454
rect 2146 336218 2382 336454
rect 1826 335898 2062 336134
rect 2146 335898 2382 336134
rect 5826 336218 6062 336454
rect 6146 336218 6382 336454
rect 5826 335898 6062 336134
rect 6146 335898 6382 336134
rect 185826 336218 186062 336454
rect 186146 336218 186382 336454
rect 185826 335898 186062 336134
rect 186146 335898 186382 336134
rect 221826 336218 222062 336454
rect 222146 336218 222382 336454
rect 221826 335898 222062 336134
rect 222146 335898 222382 336134
rect 257826 336218 258062 336454
rect 258146 336218 258382 336454
rect 257826 335898 258062 336134
rect 258146 335898 258382 336134
rect 293826 336218 294062 336454
rect 294146 336218 294382 336454
rect 293826 335898 294062 336134
rect 294146 335898 294382 336134
rect 329826 336218 330062 336454
rect 330146 336218 330382 336454
rect 329826 335898 330062 336134
rect 330146 335898 330382 336134
rect 365826 336218 366062 336454
rect 366146 336218 366382 336454
rect 365826 335898 366062 336134
rect 366146 335898 366382 336134
rect 401826 336218 402062 336454
rect 402146 336218 402382 336454
rect 401826 335898 402062 336134
rect 402146 335898 402382 336134
rect 568510 336218 568746 336454
rect 568830 336218 569066 336454
rect 568510 335898 568746 336134
rect 568830 335898 569066 336134
rect 577826 336218 578062 336454
rect 578146 336218 578382 336454
rect 577826 335898 578062 336134
rect 578146 335898 578382 336134
rect 9546 303938 9782 304174
rect 9866 303938 10102 304174
rect 9546 303618 9782 303854
rect 9866 303618 10102 303854
rect 189546 303938 189782 304174
rect 189866 303938 190102 304174
rect 189546 303618 189782 303854
rect 189866 303618 190102 303854
rect 225546 303938 225782 304174
rect 225866 303938 226102 304174
rect 225546 303618 225782 303854
rect 225866 303618 226102 303854
rect 261546 303938 261782 304174
rect 261866 303938 262102 304174
rect 261546 303618 261782 303854
rect 261866 303618 262102 303854
rect 297546 303938 297782 304174
rect 297866 303938 298102 304174
rect 297546 303618 297782 303854
rect 297866 303618 298102 303854
rect 333546 303938 333782 304174
rect 333866 303938 334102 304174
rect 333546 303618 333782 303854
rect 333866 303618 334102 303854
rect 369546 303938 369782 304174
rect 369866 303938 370102 304174
rect 369546 303618 369782 303854
rect 369866 303618 370102 303854
rect 405546 303938 405782 304174
rect 405866 303938 406102 304174
rect 405546 303618 405782 303854
rect 405866 303618 406102 303854
rect 572374 303938 572610 304174
rect 572694 303938 572930 304174
rect 572374 303618 572610 303854
rect 572694 303618 572930 303854
rect 1826 300218 2062 300454
rect 2146 300218 2382 300454
rect 1826 299898 2062 300134
rect 2146 299898 2382 300134
rect 5826 300218 6062 300454
rect 6146 300218 6382 300454
rect 5826 299898 6062 300134
rect 6146 299898 6382 300134
rect 185826 300218 186062 300454
rect 186146 300218 186382 300454
rect 185826 299898 186062 300134
rect 186146 299898 186382 300134
rect 221826 300218 222062 300454
rect 222146 300218 222382 300454
rect 221826 299898 222062 300134
rect 222146 299898 222382 300134
rect 257826 300218 258062 300454
rect 258146 300218 258382 300454
rect 257826 299898 258062 300134
rect 258146 299898 258382 300134
rect 293826 300218 294062 300454
rect 294146 300218 294382 300454
rect 293826 299898 294062 300134
rect 294146 299898 294382 300134
rect 329826 300218 330062 300454
rect 330146 300218 330382 300454
rect 329826 299898 330062 300134
rect 330146 299898 330382 300134
rect 365826 300218 366062 300454
rect 366146 300218 366382 300454
rect 365826 299898 366062 300134
rect 366146 299898 366382 300134
rect 401826 300218 402062 300454
rect 402146 300218 402382 300454
rect 401826 299898 402062 300134
rect 402146 299898 402382 300134
rect 568510 300218 568746 300454
rect 568830 300218 569066 300454
rect 568510 299898 568746 300134
rect 568830 299898 569066 300134
rect 577826 300218 578062 300454
rect 578146 300218 578382 300454
rect 577826 299898 578062 300134
rect 578146 299898 578382 300134
rect 9546 267938 9782 268174
rect 9866 267938 10102 268174
rect 9546 267618 9782 267854
rect 9866 267618 10102 267854
rect 189546 267938 189782 268174
rect 189866 267938 190102 268174
rect 189546 267618 189782 267854
rect 189866 267618 190102 267854
rect 225546 267938 225782 268174
rect 225866 267938 226102 268174
rect 225546 267618 225782 267854
rect 225866 267618 226102 267854
rect 261546 267938 261782 268174
rect 261866 267938 262102 268174
rect 261546 267618 261782 267854
rect 261866 267618 262102 267854
rect 297546 267938 297782 268174
rect 297866 267938 298102 268174
rect 297546 267618 297782 267854
rect 297866 267618 298102 267854
rect 333546 267938 333782 268174
rect 333866 267938 334102 268174
rect 333546 267618 333782 267854
rect 333866 267618 334102 267854
rect 369546 267938 369782 268174
rect 369866 267938 370102 268174
rect 369546 267618 369782 267854
rect 369866 267618 370102 267854
rect 405546 267938 405782 268174
rect 405866 267938 406102 268174
rect 405546 267618 405782 267854
rect 405866 267618 406102 267854
rect 572374 267938 572610 268174
rect 572694 267938 572930 268174
rect 572374 267618 572610 267854
rect 572694 267618 572930 267854
rect 1826 264218 2062 264454
rect 2146 264218 2382 264454
rect 1826 263898 2062 264134
rect 2146 263898 2382 264134
rect 5826 264218 6062 264454
rect 6146 264218 6382 264454
rect 5826 263898 6062 264134
rect 6146 263898 6382 264134
rect 185826 264218 186062 264454
rect 186146 264218 186382 264454
rect 185826 263898 186062 264134
rect 186146 263898 186382 264134
rect 221826 264218 222062 264454
rect 222146 264218 222382 264454
rect 221826 263898 222062 264134
rect 222146 263898 222382 264134
rect 257826 264218 258062 264454
rect 258146 264218 258382 264454
rect 257826 263898 258062 264134
rect 258146 263898 258382 264134
rect 293826 264218 294062 264454
rect 294146 264218 294382 264454
rect 293826 263898 294062 264134
rect 294146 263898 294382 264134
rect 329826 264218 330062 264454
rect 330146 264218 330382 264454
rect 329826 263898 330062 264134
rect 330146 263898 330382 264134
rect 365826 264218 366062 264454
rect 366146 264218 366382 264454
rect 365826 263898 366062 264134
rect 366146 263898 366382 264134
rect 401826 264218 402062 264454
rect 402146 264218 402382 264454
rect 401826 263898 402062 264134
rect 402146 263898 402382 264134
rect 568510 264218 568746 264454
rect 568830 264218 569066 264454
rect 568510 263898 568746 264134
rect 568830 263898 569066 264134
rect 577826 264218 578062 264454
rect 578146 264218 578382 264454
rect 577826 263898 578062 264134
rect 578146 263898 578382 264134
rect 9546 231938 9782 232174
rect 9866 231938 10102 232174
rect 9546 231618 9782 231854
rect 9866 231618 10102 231854
rect 45546 231938 45782 232174
rect 45866 231938 46102 232174
rect 45546 231618 45782 231854
rect 45866 231618 46102 231854
rect 81546 231938 81782 232174
rect 81866 231938 82102 232174
rect 81546 231618 81782 231854
rect 81866 231618 82102 231854
rect 117546 231938 117782 232174
rect 117866 231938 118102 232174
rect 117546 231618 117782 231854
rect 117866 231618 118102 231854
rect 153546 231938 153782 232174
rect 153866 231938 154102 232174
rect 153546 231618 153782 231854
rect 153866 231618 154102 231854
rect 189546 231938 189782 232174
rect 189866 231938 190102 232174
rect 189546 231618 189782 231854
rect 189866 231618 190102 231854
rect 225546 231938 225782 232174
rect 225866 231938 226102 232174
rect 225546 231618 225782 231854
rect 225866 231618 226102 231854
rect 261546 231938 261782 232174
rect 261866 231938 262102 232174
rect 261546 231618 261782 231854
rect 261866 231618 262102 231854
rect 297546 231938 297782 232174
rect 297866 231938 298102 232174
rect 297546 231618 297782 231854
rect 297866 231618 298102 231854
rect 333546 231938 333782 232174
rect 333866 231938 334102 232174
rect 333546 231618 333782 231854
rect 333866 231618 334102 231854
rect 369546 231938 369782 232174
rect 369866 231938 370102 232174
rect 369546 231618 369782 231854
rect 369866 231618 370102 231854
rect 405546 231938 405782 232174
rect 405866 231938 406102 232174
rect 405546 231618 405782 231854
rect 405866 231618 406102 231854
rect 441546 231938 441782 232174
rect 441866 231938 442102 232174
rect 441546 231618 441782 231854
rect 441866 231618 442102 231854
rect 477546 231938 477782 232174
rect 477866 231938 478102 232174
rect 477546 231618 477782 231854
rect 477866 231618 478102 231854
rect 513546 231938 513782 232174
rect 513866 231938 514102 232174
rect 513546 231618 513782 231854
rect 513866 231618 514102 231854
rect 549546 231938 549782 232174
rect 549866 231938 550102 232174
rect 549546 231618 549782 231854
rect 549866 231618 550102 231854
rect 1826 228218 2062 228454
rect 2146 228218 2382 228454
rect 1826 227898 2062 228134
rect 2146 227898 2382 228134
rect 5826 228218 6062 228454
rect 6146 228218 6382 228454
rect 5826 227898 6062 228134
rect 6146 227898 6382 228134
rect 41826 228218 42062 228454
rect 42146 228218 42382 228454
rect 41826 227898 42062 228134
rect 42146 227898 42382 228134
rect 77826 228218 78062 228454
rect 78146 228218 78382 228454
rect 77826 227898 78062 228134
rect 78146 227898 78382 228134
rect 113826 228218 114062 228454
rect 114146 228218 114382 228454
rect 113826 227898 114062 228134
rect 114146 227898 114382 228134
rect 149826 228218 150062 228454
rect 150146 228218 150382 228454
rect 149826 227898 150062 228134
rect 150146 227898 150382 228134
rect 185826 228218 186062 228454
rect 186146 228218 186382 228454
rect 185826 227898 186062 228134
rect 186146 227898 186382 228134
rect 221826 228218 222062 228454
rect 222146 228218 222382 228454
rect 221826 227898 222062 228134
rect 222146 227898 222382 228134
rect 257826 228218 258062 228454
rect 258146 228218 258382 228454
rect 257826 227898 258062 228134
rect 258146 227898 258382 228134
rect 293826 228218 294062 228454
rect 294146 228218 294382 228454
rect 293826 227898 294062 228134
rect 294146 227898 294382 228134
rect 329826 228218 330062 228454
rect 330146 228218 330382 228454
rect 329826 227898 330062 228134
rect 330146 227898 330382 228134
rect 365826 228218 366062 228454
rect 366146 228218 366382 228454
rect 365826 227898 366062 228134
rect 366146 227898 366382 228134
rect 401826 228218 402062 228454
rect 402146 228218 402382 228454
rect 401826 227898 402062 228134
rect 402146 227898 402382 228134
rect 437826 228218 438062 228454
rect 438146 228218 438382 228454
rect 437826 227898 438062 228134
rect 438146 227898 438382 228134
rect 473826 228218 474062 228454
rect 474146 228218 474382 228454
rect 473826 227898 474062 228134
rect 474146 227898 474382 228134
rect 509826 228218 510062 228454
rect 510146 228218 510382 228454
rect 509826 227898 510062 228134
rect 510146 227898 510382 228134
rect 545826 228218 546062 228454
rect 546146 228218 546382 228454
rect 577826 228218 578062 228454
rect 578146 228218 578382 228454
rect 545826 227898 546062 228134
rect 546146 227898 546382 228134
rect 568510 227903 568746 228139
rect 568830 227903 569066 228139
rect 577826 227898 578062 228134
rect 578146 227898 578382 228134
rect 9546 195938 9782 196174
rect 9866 195938 10102 196174
rect 9546 195618 9782 195854
rect 9866 195618 10102 195854
rect 189546 195938 189782 196174
rect 189866 195938 190102 196174
rect 189546 195618 189782 195854
rect 189866 195618 190102 195854
rect 225546 195938 225782 196174
rect 225866 195938 226102 196174
rect 225546 195618 225782 195854
rect 225866 195618 226102 195854
rect 261546 195938 261782 196174
rect 261866 195938 262102 196174
rect 261546 195618 261782 195854
rect 261866 195618 262102 195854
rect 297546 195938 297782 196174
rect 297866 195938 298102 196174
rect 297546 195618 297782 195854
rect 297866 195618 298102 195854
rect 333546 195938 333782 196174
rect 333866 195938 334102 196174
rect 333546 195618 333782 195854
rect 333866 195618 334102 195854
rect 369546 195938 369782 196174
rect 369866 195938 370102 196174
rect 369546 195618 369782 195854
rect 369866 195618 370102 195854
rect 405546 195938 405782 196174
rect 405866 195938 406102 196174
rect 405546 195618 405782 195854
rect 405866 195618 406102 195854
rect 572374 195938 572610 196174
rect 572694 195938 572930 196174
rect 572374 195618 572610 195854
rect 572694 195618 572930 195854
rect 1826 192218 2062 192454
rect 2146 192218 2382 192454
rect 1826 191898 2062 192134
rect 2146 191898 2382 192134
rect 5826 192218 6062 192454
rect 6146 192218 6382 192454
rect 5826 191898 6062 192134
rect 6146 191898 6382 192134
rect 185826 192218 186062 192454
rect 186146 192218 186382 192454
rect 185826 191898 186062 192134
rect 186146 191898 186382 192134
rect 221826 192218 222062 192454
rect 222146 192218 222382 192454
rect 221826 191898 222062 192134
rect 222146 191898 222382 192134
rect 257826 192218 258062 192454
rect 258146 192218 258382 192454
rect 257826 191898 258062 192134
rect 258146 191898 258382 192134
rect 293826 192218 294062 192454
rect 294146 192218 294382 192454
rect 293826 191898 294062 192134
rect 294146 191898 294382 192134
rect 329826 192218 330062 192454
rect 330146 192218 330382 192454
rect 329826 191898 330062 192134
rect 330146 191898 330382 192134
rect 365826 192218 366062 192454
rect 366146 192218 366382 192454
rect 365826 191898 366062 192134
rect 366146 191898 366382 192134
rect 401826 192218 402062 192454
rect 402146 192218 402382 192454
rect 401826 191898 402062 192134
rect 402146 191898 402382 192134
rect 568510 192218 568746 192454
rect 568830 192218 569066 192454
rect 568510 191898 568746 192134
rect 568830 191898 569066 192134
rect 577826 192218 578062 192454
rect 578146 192218 578382 192454
rect 577826 191898 578062 192134
rect 578146 191898 578382 192134
rect 9546 159938 9782 160174
rect 9866 159938 10102 160174
rect 9546 159618 9782 159854
rect 9866 159618 10102 159854
rect 189546 159938 189782 160174
rect 189866 159938 190102 160174
rect 189546 159618 189782 159854
rect 189866 159618 190102 159854
rect 225546 159938 225782 160174
rect 225866 159938 226102 160174
rect 225546 159618 225782 159854
rect 225866 159618 226102 159854
rect 261546 159938 261782 160174
rect 261866 159938 262102 160174
rect 261546 159618 261782 159854
rect 261866 159618 262102 159854
rect 297546 159938 297782 160174
rect 297866 159938 298102 160174
rect 297546 159618 297782 159854
rect 297866 159618 298102 159854
rect 333546 159938 333782 160174
rect 333866 159938 334102 160174
rect 333546 159618 333782 159854
rect 333866 159618 334102 159854
rect 369546 159938 369782 160174
rect 369866 159938 370102 160174
rect 369546 159618 369782 159854
rect 369866 159618 370102 159854
rect 405546 159938 405782 160174
rect 405866 159938 406102 160174
rect 405546 159618 405782 159854
rect 405866 159618 406102 159854
rect 572374 159938 572610 160174
rect 572694 159938 572930 160174
rect 572374 159618 572610 159854
rect 572694 159618 572930 159854
rect 1826 156218 2062 156454
rect 2146 156218 2382 156454
rect 1826 155898 2062 156134
rect 2146 155898 2382 156134
rect 5826 156218 6062 156454
rect 6146 156218 6382 156454
rect 5826 155898 6062 156134
rect 6146 155898 6382 156134
rect 185826 156218 186062 156454
rect 186146 156218 186382 156454
rect 185826 155898 186062 156134
rect 186146 155898 186382 156134
rect 221826 156218 222062 156454
rect 222146 156218 222382 156454
rect 221826 155898 222062 156134
rect 222146 155898 222382 156134
rect 257826 156218 258062 156454
rect 258146 156218 258382 156454
rect 257826 155898 258062 156134
rect 258146 155898 258382 156134
rect 293826 156218 294062 156454
rect 294146 156218 294382 156454
rect 293826 155898 294062 156134
rect 294146 155898 294382 156134
rect 329826 156218 330062 156454
rect 330146 156218 330382 156454
rect 329826 155898 330062 156134
rect 330146 155898 330382 156134
rect 365826 156218 366062 156454
rect 366146 156218 366382 156454
rect 365826 155898 366062 156134
rect 366146 155898 366382 156134
rect 401826 156218 402062 156454
rect 402146 156218 402382 156454
rect 401826 155898 402062 156134
rect 402146 155898 402382 156134
rect 568510 156218 568746 156454
rect 568830 156218 569066 156454
rect 568510 155898 568746 156134
rect 568830 155898 569066 156134
rect 577826 156218 578062 156454
rect 578146 156218 578382 156454
rect 577826 155898 578062 156134
rect 578146 155898 578382 156134
rect 9546 123938 9782 124174
rect 9866 123938 10102 124174
rect 9546 123618 9782 123854
rect 9866 123618 10102 123854
rect 45546 123938 45782 124174
rect 45866 123938 46102 124174
rect 45546 123618 45782 123854
rect 45866 123618 46102 123854
rect 81546 123938 81782 124174
rect 81866 123938 82102 124174
rect 81546 123618 81782 123854
rect 81866 123618 82102 123854
rect 117546 123938 117782 124174
rect 117866 123938 118102 124174
rect 117546 123618 117782 123854
rect 117866 123618 118102 123854
rect 153546 123938 153782 124174
rect 153866 123938 154102 124174
rect 153546 123618 153782 123854
rect 153866 123618 154102 123854
rect 189546 123938 189782 124174
rect 189866 123938 190102 124174
rect 189546 123618 189782 123854
rect 189866 123618 190102 123854
rect 225546 123938 225782 124174
rect 225866 123938 226102 124174
rect 225546 123618 225782 123854
rect 225866 123618 226102 123854
rect 261546 123938 261782 124174
rect 261866 123938 262102 124174
rect 261546 123618 261782 123854
rect 261866 123618 262102 123854
rect 297546 123938 297782 124174
rect 297866 123938 298102 124174
rect 297546 123618 297782 123854
rect 297866 123618 298102 123854
rect 333546 123938 333782 124174
rect 333866 123938 334102 124174
rect 333546 123618 333782 123854
rect 333866 123618 334102 123854
rect 369546 123938 369782 124174
rect 369866 123938 370102 124174
rect 369546 123618 369782 123854
rect 369866 123618 370102 123854
rect 405546 123938 405782 124174
rect 405866 123938 406102 124174
rect 405546 123618 405782 123854
rect 405866 123618 406102 123854
rect 441546 123938 441782 124174
rect 441866 123938 442102 124174
rect 441546 123618 441782 123854
rect 441866 123618 442102 123854
rect 477546 123938 477782 124174
rect 477866 123938 478102 124174
rect 477546 123618 477782 123854
rect 477866 123618 478102 123854
rect 513546 123938 513782 124174
rect 513866 123938 514102 124174
rect 513546 123618 513782 123854
rect 513866 123618 514102 123854
rect 549546 123938 549782 124174
rect 549866 123938 550102 124174
rect 549546 123618 549782 123854
rect 549866 123618 550102 123854
rect 1826 120218 2062 120454
rect 2146 120218 2382 120454
rect 1826 119898 2062 120134
rect 2146 119898 2382 120134
rect 5826 120218 6062 120454
rect 6146 120218 6382 120454
rect 5826 119898 6062 120134
rect 6146 119898 6382 120134
rect 41826 120218 42062 120454
rect 42146 120218 42382 120454
rect 41826 119898 42062 120134
rect 42146 119898 42382 120134
rect 77826 120218 78062 120454
rect 78146 120218 78382 120454
rect 77826 119898 78062 120134
rect 78146 119898 78382 120134
rect 113826 120218 114062 120454
rect 114146 120218 114382 120454
rect 113826 119898 114062 120134
rect 114146 119898 114382 120134
rect 149826 120218 150062 120454
rect 150146 120218 150382 120454
rect 149826 119898 150062 120134
rect 150146 119898 150382 120134
rect 185826 120218 186062 120454
rect 186146 120218 186382 120454
rect 185826 119898 186062 120134
rect 186146 119898 186382 120134
rect 221826 120218 222062 120454
rect 222146 120218 222382 120454
rect 221826 119898 222062 120134
rect 222146 119898 222382 120134
rect 257826 120218 258062 120454
rect 258146 120218 258382 120454
rect 257826 119898 258062 120134
rect 258146 119898 258382 120134
rect 293826 120218 294062 120454
rect 294146 120218 294382 120454
rect 293826 119898 294062 120134
rect 294146 119898 294382 120134
rect 329826 120218 330062 120454
rect 330146 120218 330382 120454
rect 329826 119898 330062 120134
rect 330146 119898 330382 120134
rect 365826 120218 366062 120454
rect 366146 120218 366382 120454
rect 365826 119898 366062 120134
rect 366146 119898 366382 120134
rect 401826 120218 402062 120454
rect 402146 120218 402382 120454
rect 401826 119898 402062 120134
rect 402146 119898 402382 120134
rect 437826 120218 438062 120454
rect 438146 120218 438382 120454
rect 437826 119898 438062 120134
rect 438146 119898 438382 120134
rect 473826 120218 474062 120454
rect 474146 120218 474382 120454
rect 473826 119898 474062 120134
rect 474146 119898 474382 120134
rect 509826 120218 510062 120454
rect 510146 120218 510382 120454
rect 509826 119898 510062 120134
rect 510146 119898 510382 120134
rect 545826 120218 546062 120454
rect 546146 120218 546382 120454
rect 545826 119898 546062 120134
rect 546146 119898 546382 120134
rect 577826 120218 578062 120454
rect 578146 120218 578382 120454
rect 577826 119898 578062 120134
rect 578146 119898 578382 120134
rect 9546 87938 9782 88174
rect 9866 87938 10102 88174
rect 9546 87618 9782 87854
rect 9866 87618 10102 87854
rect 189546 87938 189782 88174
rect 189866 87938 190102 88174
rect 189546 87618 189782 87854
rect 189866 87618 190102 87854
rect 369546 87938 369782 88174
rect 369866 87938 370102 88174
rect 369546 87618 369782 87854
rect 369866 87618 370102 87854
rect 405546 87938 405782 88174
rect 405866 87938 406102 88174
rect 405546 87618 405782 87854
rect 405866 87618 406102 87854
rect 572374 87938 572610 88174
rect 572694 87938 572930 88174
rect 572374 87618 572610 87854
rect 572694 87618 572930 87854
rect 1826 84218 2062 84454
rect 2146 84218 2382 84454
rect 1826 83898 2062 84134
rect 2146 83898 2382 84134
rect 5826 84218 6062 84454
rect 6146 84218 6382 84454
rect 5826 83898 6062 84134
rect 6146 83898 6382 84134
rect 185826 84218 186062 84454
rect 186146 84218 186382 84454
rect 185826 83898 186062 84134
rect 186146 83898 186382 84134
rect 365826 84218 366062 84454
rect 366146 84218 366382 84454
rect 365826 83898 366062 84134
rect 366146 83898 366382 84134
rect 401826 84218 402062 84454
rect 402146 84218 402382 84454
rect 401826 83898 402062 84134
rect 402146 83898 402382 84134
rect 568510 84218 568746 84454
rect 568830 84218 569066 84454
rect 568510 83898 568746 84134
rect 568830 83898 569066 84134
rect 577826 84218 578062 84454
rect 578146 84218 578382 84454
rect 577826 83898 578062 84134
rect 578146 83898 578382 84134
rect 9546 51938 9782 52174
rect 9866 51938 10102 52174
rect 9546 51618 9782 51854
rect 9866 51618 10102 51854
rect 189546 51938 189782 52174
rect 189866 51938 190102 52174
rect 189546 51618 189782 51854
rect 189866 51618 190102 51854
rect 369546 51938 369782 52174
rect 369866 51938 370102 52174
rect 369546 51618 369782 51854
rect 369866 51618 370102 51854
rect 405546 51938 405782 52174
rect 405866 51938 406102 52174
rect 405546 51618 405782 51854
rect 405866 51618 406102 51854
rect 572374 51938 572610 52174
rect 572694 51938 572930 52174
rect 572374 51618 572610 51854
rect 572694 51618 572930 51854
rect 1826 48218 2062 48454
rect 2146 48218 2382 48454
rect 1826 47898 2062 48134
rect 2146 47898 2382 48134
rect 5826 48218 6062 48454
rect 6146 48218 6382 48454
rect 5826 47898 6062 48134
rect 6146 47898 6382 48134
rect 185826 48218 186062 48454
rect 186146 48218 186382 48454
rect 185826 47898 186062 48134
rect 186146 47898 186382 48134
rect 365826 48218 366062 48454
rect 366146 48218 366382 48454
rect 365826 47898 366062 48134
rect 366146 47898 366382 48134
rect 401826 48218 402062 48454
rect 402146 48218 402382 48454
rect 401826 47898 402062 48134
rect 402146 47898 402382 48134
rect 568510 48218 568746 48454
rect 568830 48218 569066 48454
rect 568510 47898 568746 48134
rect 568830 47898 569066 48134
rect 577826 48218 578062 48454
rect 578146 48218 578382 48454
rect 577826 47898 578062 48134
rect 578146 47898 578382 48134
rect 9546 15938 9782 16174
rect 9866 15938 10102 16174
rect 9546 15618 9782 15854
rect 9866 15618 10102 15854
rect 45546 15938 45782 16174
rect 45866 15938 46102 16174
rect 45546 15618 45782 15854
rect 45866 15618 46102 15854
rect 81546 15938 81782 16174
rect 81866 15938 82102 16174
rect 81546 15618 81782 15854
rect 81866 15618 82102 15854
rect 117546 15938 117782 16174
rect 117866 15938 118102 16174
rect 117546 15618 117782 15854
rect 117866 15618 118102 15854
rect 153546 15938 153782 16174
rect 153866 15938 154102 16174
rect 153546 15618 153782 15854
rect 153866 15618 154102 15854
rect 189546 15938 189782 16174
rect 189866 15938 190102 16174
rect 189546 15618 189782 15854
rect 189866 15618 190102 15854
rect 225546 15938 225782 16174
rect 225866 15938 226102 16174
rect 225546 15618 225782 15854
rect 225866 15618 226102 15854
rect 261546 15938 261782 16174
rect 261866 15938 262102 16174
rect 261546 15618 261782 15854
rect 261866 15618 262102 15854
rect 297546 15938 297782 16174
rect 297866 15938 298102 16174
rect 297546 15618 297782 15854
rect 297866 15618 298102 15854
rect 333546 15938 333782 16174
rect 333866 15938 334102 16174
rect 333546 15618 333782 15854
rect 333866 15618 334102 15854
rect 369546 15938 369782 16174
rect 369866 15938 370102 16174
rect 369546 15618 369782 15854
rect 369866 15618 370102 15854
rect 405546 15938 405782 16174
rect 405866 15938 406102 16174
rect 405546 15618 405782 15854
rect 405866 15618 406102 15854
rect 441546 15938 441782 16174
rect 441866 15938 442102 16174
rect 441546 15618 441782 15854
rect 441866 15618 442102 15854
rect 477546 15938 477782 16174
rect 477866 15938 478102 16174
rect 477546 15618 477782 15854
rect 477866 15618 478102 15854
rect 513546 15938 513782 16174
rect 513866 15938 514102 16174
rect 513546 15618 513782 15854
rect 513866 15618 514102 15854
rect 549546 15938 549782 16174
rect 549866 15938 550102 16174
rect 549546 15618 549782 15854
rect 549866 15618 550102 15854
rect 1826 12218 2062 12454
rect 2146 12218 2382 12454
rect 1826 11898 2062 12134
rect 2146 11898 2382 12134
rect 5826 12218 6062 12454
rect 6146 12218 6382 12454
rect 5826 11898 6062 12134
rect 6146 11898 6382 12134
rect 41826 12218 42062 12454
rect 42146 12218 42382 12454
rect 41826 11898 42062 12134
rect 42146 11898 42382 12134
rect 77826 12218 78062 12454
rect 78146 12218 78382 12454
rect 77826 11898 78062 12134
rect 78146 11898 78382 12134
rect 113826 12218 114062 12454
rect 114146 12218 114382 12454
rect 113826 11898 114062 12134
rect 114146 11898 114382 12134
rect 149826 12218 150062 12454
rect 150146 12218 150382 12454
rect 149826 11898 150062 12134
rect 150146 11898 150382 12134
rect 185826 12218 186062 12454
rect 186146 12218 186382 12454
rect 185826 11898 186062 12134
rect 186146 11898 186382 12134
rect 221826 12218 222062 12454
rect 222146 12218 222382 12454
rect 221826 11898 222062 12134
rect 222146 11898 222382 12134
rect 257826 12218 258062 12454
rect 258146 12218 258382 12454
rect 257826 11898 258062 12134
rect 258146 11898 258382 12134
rect 293826 12218 294062 12454
rect 294146 12218 294382 12454
rect 293826 11898 294062 12134
rect 294146 11898 294382 12134
rect 329826 12218 330062 12454
rect 330146 12218 330382 12454
rect 329826 11898 330062 12134
rect 330146 11898 330382 12134
rect 365826 12218 366062 12454
rect 366146 12218 366382 12454
rect 365826 11898 366062 12134
rect 366146 11898 366382 12134
rect 401826 12218 402062 12454
rect 402146 12218 402382 12454
rect 401826 11898 402062 12134
rect 402146 11898 402382 12134
rect 437826 12218 438062 12454
rect 438146 12218 438382 12454
rect 437826 11898 438062 12134
rect 438146 11898 438382 12134
rect 473826 12218 474062 12454
rect 474146 12218 474382 12454
rect 473826 11898 474062 12134
rect 474146 11898 474382 12134
rect 509826 12218 510062 12454
rect 510146 12218 510382 12454
rect 509826 11898 510062 12134
rect 510146 11898 510382 12134
rect 545826 12218 546062 12454
rect 546146 12218 546382 12454
rect 545826 11898 546062 12134
rect 546146 11898 546382 12134
rect 577826 12218 578062 12454
rect 578146 12218 578382 12454
rect 577826 11898 578062 12134
rect 578146 11898 578382 12134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 699938 581782 700174
rect 581866 699938 582102 700174
rect 581546 699618 581782 699854
rect 581866 699618 582102 699854
rect 581546 663938 581782 664174
rect 581866 663938 582102 664174
rect 581546 663618 581782 663854
rect 581866 663618 582102 663854
rect 581546 627938 581782 628174
rect 581866 627938 582102 628174
rect 581546 627618 581782 627854
rect 581866 627618 582102 627854
rect 581546 591938 581782 592174
rect 581866 591938 582102 592174
rect 581546 591618 581782 591854
rect 581866 591618 582102 591854
rect 581546 555938 581782 556174
rect 581866 555938 582102 556174
rect 581546 555618 581782 555854
rect 581866 555618 582102 555854
rect 581546 519938 581782 520174
rect 581866 519938 582102 520174
rect 581546 519618 581782 519854
rect 581866 519618 582102 519854
rect 581546 483938 581782 484174
rect 581866 483938 582102 484174
rect 581546 483618 581782 483854
rect 581866 483618 582102 483854
rect 581546 447938 581782 448174
rect 581866 447938 582102 448174
rect 581546 447618 581782 447854
rect 581866 447618 582102 447854
rect 581546 411938 581782 412174
rect 581866 411938 582102 412174
rect 581546 411618 581782 411854
rect 581866 411618 582102 411854
rect 581546 375938 581782 376174
rect 581866 375938 582102 376174
rect 581546 375618 581782 375854
rect 581866 375618 582102 375854
rect 581546 339938 581782 340174
rect 581866 339938 582102 340174
rect 581546 339618 581782 339854
rect 581866 339618 582102 339854
rect 581546 303938 581782 304174
rect 581866 303938 582102 304174
rect 581546 303618 581782 303854
rect 581866 303618 582102 303854
rect 581546 267938 581782 268174
rect 581866 267938 582102 268174
rect 581546 267618 581782 267854
rect 581866 267618 582102 267854
rect 581546 231938 581782 232174
rect 581866 231938 582102 232174
rect 581546 231618 581782 231854
rect 581866 231618 582102 231854
rect 581546 195938 581782 196174
rect 581866 195938 582102 196174
rect 581546 195618 581782 195854
rect 581866 195618 582102 195854
rect 581546 159938 581782 160174
rect 581866 159938 582102 160174
rect 581546 159618 581782 159854
rect 581866 159618 582102 159854
rect 581546 123938 581782 124174
rect 581866 123938 582102 124174
rect 581546 123618 581782 123854
rect 581866 123618 582102 123854
rect 581546 87938 581782 88174
rect 581866 87938 582102 88174
rect 581546 87618 581782 87854
rect 581866 87618 582102 87854
rect 581546 51938 581782 52174
rect 581866 51938 582102 52174
rect 581546 51618 581782 51854
rect 581866 51618 582102 51854
rect 581546 15938 581782 16174
rect 581866 15938 582102 16174
rect 581546 15618 581782 15854
rect 581866 15618 582102 15854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 696218 585578 696454
rect 585662 696218 585898 696454
rect 585342 695898 585578 696134
rect 585662 695898 585898 696134
rect 585342 660218 585578 660454
rect 585662 660218 585898 660454
rect 585342 659898 585578 660134
rect 585662 659898 585898 660134
rect 585342 624218 585578 624454
rect 585662 624218 585898 624454
rect 585342 623898 585578 624134
rect 585662 623898 585898 624134
rect 585342 588218 585578 588454
rect 585662 588218 585898 588454
rect 585342 587898 585578 588134
rect 585662 587898 585898 588134
rect 585342 552218 585578 552454
rect 585662 552218 585898 552454
rect 585342 551898 585578 552134
rect 585662 551898 585898 552134
rect 585342 516218 585578 516454
rect 585662 516218 585898 516454
rect 585342 515898 585578 516134
rect 585662 515898 585898 516134
rect 585342 480218 585578 480454
rect 585662 480218 585898 480454
rect 585342 479898 585578 480134
rect 585662 479898 585898 480134
rect 585342 444218 585578 444454
rect 585662 444218 585898 444454
rect 585342 443898 585578 444134
rect 585662 443898 585898 444134
rect 585342 408218 585578 408454
rect 585662 408218 585898 408454
rect 585342 407898 585578 408134
rect 585662 407898 585898 408134
rect 585342 372218 585578 372454
rect 585662 372218 585898 372454
rect 585342 371898 585578 372134
rect 585662 371898 585898 372134
rect 585342 336218 585578 336454
rect 585662 336218 585898 336454
rect 585342 335898 585578 336134
rect 585662 335898 585898 336134
rect 585342 300218 585578 300454
rect 585662 300218 585898 300454
rect 585342 299898 585578 300134
rect 585662 299898 585898 300134
rect 585342 264218 585578 264454
rect 585662 264218 585898 264454
rect 585342 263898 585578 264134
rect 585662 263898 585898 264134
rect 585342 228218 585578 228454
rect 585662 228218 585898 228454
rect 585342 227898 585578 228134
rect 585662 227898 585898 228134
rect 585342 192218 585578 192454
rect 585662 192218 585898 192454
rect 585342 191898 585578 192134
rect 585662 191898 585898 192134
rect 585342 156218 585578 156454
rect 585662 156218 585898 156454
rect 585342 155898 585578 156134
rect 585662 155898 585898 156134
rect 585342 120218 585578 120454
rect 585662 120218 585898 120454
rect 585342 119898 585578 120134
rect 585662 119898 585898 120134
rect 585342 84218 585578 84454
rect 585662 84218 585898 84454
rect 585342 83898 585578 84134
rect 585662 83898 585898 84134
rect 585342 48218 585578 48454
rect 585662 48218 585898 48454
rect 585342 47898 585578 48134
rect 585662 47898 585898 48134
rect 585342 12218 585578 12454
rect 585662 12218 585898 12454
rect 585342 11898 585578 12134
rect 585662 11898 585898 12134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 699938 586538 700174
rect 586622 699938 586858 700174
rect 586302 699618 586538 699854
rect 586622 699618 586858 699854
rect 586302 663938 586538 664174
rect 586622 663938 586858 664174
rect 586302 663618 586538 663854
rect 586622 663618 586858 663854
rect 586302 627938 586538 628174
rect 586622 627938 586858 628174
rect 586302 627618 586538 627854
rect 586622 627618 586858 627854
rect 586302 591938 586538 592174
rect 586622 591938 586858 592174
rect 586302 591618 586538 591854
rect 586622 591618 586858 591854
rect 586302 555938 586538 556174
rect 586622 555938 586858 556174
rect 586302 555618 586538 555854
rect 586622 555618 586858 555854
rect 586302 519938 586538 520174
rect 586622 519938 586858 520174
rect 586302 519618 586538 519854
rect 586622 519618 586858 519854
rect 586302 483938 586538 484174
rect 586622 483938 586858 484174
rect 586302 483618 586538 483854
rect 586622 483618 586858 483854
rect 586302 447938 586538 448174
rect 586622 447938 586858 448174
rect 586302 447618 586538 447854
rect 586622 447618 586858 447854
rect 586302 411938 586538 412174
rect 586622 411938 586858 412174
rect 586302 411618 586538 411854
rect 586622 411618 586858 411854
rect 586302 375938 586538 376174
rect 586622 375938 586858 376174
rect 586302 375618 586538 375854
rect 586622 375618 586858 375854
rect 586302 339938 586538 340174
rect 586622 339938 586858 340174
rect 586302 339618 586538 339854
rect 586622 339618 586858 339854
rect 586302 303938 586538 304174
rect 586622 303938 586858 304174
rect 586302 303618 586538 303854
rect 586622 303618 586858 303854
rect 586302 267938 586538 268174
rect 586622 267938 586858 268174
rect 586302 267618 586538 267854
rect 586622 267618 586858 267854
rect 586302 231938 586538 232174
rect 586622 231938 586858 232174
rect 586302 231618 586538 231854
rect 586622 231618 586858 231854
rect 586302 195938 586538 196174
rect 586622 195938 586858 196174
rect 586302 195618 586538 195854
rect 586622 195618 586858 195854
rect 586302 159938 586538 160174
rect 586622 159938 586858 160174
rect 586302 159618 586538 159854
rect 586622 159618 586858 159854
rect 586302 123938 586538 124174
rect 586622 123938 586858 124174
rect 586302 123618 586538 123854
rect 586622 123618 586858 123854
rect 586302 87938 586538 88174
rect 586622 87938 586858 88174
rect 586302 87618 586538 87854
rect 586622 87618 586858 87854
rect 586302 51938 586538 52174
rect 586622 51938 586858 52174
rect 586302 51618 586538 51854
rect 586622 51618 586858 51854
rect 586302 15938 586538 16174
rect 586622 15938 586858 16174
rect 586302 15618 586538 15854
rect 586622 15618 586858 15854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700174 592650 700206
rect -8726 699938 -2934 700174
rect -2698 699938 -2614 700174
rect -2378 700085 581546 700174
rect -2378 699938 5546 700085
rect -8726 699854 5546 699938
rect -8726 699618 -2934 699854
rect -2698 699618 -2614 699854
rect -2378 699849 5546 699854
rect 5782 699849 5866 700085
rect 6102 699849 41546 700085
rect 41782 699849 41866 700085
rect 42102 699849 77546 700085
rect 77782 699849 77866 700085
rect 78102 699849 113546 700085
rect 113782 699849 113866 700085
rect 114102 699849 149546 700085
rect 149782 699849 149866 700085
rect 150102 699849 185546 700085
rect 185782 699849 185866 700085
rect 186102 699849 221546 700085
rect 221782 699849 221866 700085
rect 222102 699849 257546 700085
rect 257782 699849 257866 700085
rect 258102 699849 293546 700085
rect 293782 699849 293866 700085
rect 294102 699849 329546 700085
rect 329782 699849 329866 700085
rect 330102 699849 365546 700085
rect 365782 699849 365866 700085
rect 366102 699849 401546 700085
rect 401782 699849 401866 700085
rect 402102 699849 437546 700085
rect 437782 699849 437866 700085
rect 438102 699849 473546 700085
rect 473782 699849 473866 700085
rect 474102 699849 509546 700085
rect 509782 699849 509866 700085
rect 510102 699849 545546 700085
rect 545782 699849 545866 700085
rect 546102 699938 581546 700085
rect 581782 699938 581866 700174
rect 582102 699938 586302 700174
rect 586538 699938 586622 700174
rect 586858 699938 592650 700174
rect 546102 699854 592650 699938
rect 546102 699849 581546 699854
rect -2378 699618 581546 699849
rect 581782 699618 581866 699854
rect 582102 699618 586302 699854
rect 586538 699618 586622 699854
rect 586858 699618 592650 699854
rect -8726 699586 592650 699618
rect -8726 696454 592650 696486
rect -8726 696218 -1974 696454
rect -1738 696218 -1654 696454
rect -1418 696218 1826 696454
rect 2062 696218 2146 696454
rect 2382 696218 5826 696454
rect 6062 696218 6146 696454
rect 6382 696218 41826 696454
rect 42062 696218 42146 696454
rect 42382 696218 77826 696454
rect 78062 696218 78146 696454
rect 78382 696218 113826 696454
rect 114062 696218 114146 696454
rect 114382 696218 149826 696454
rect 150062 696218 150146 696454
rect 150382 696218 185826 696454
rect 186062 696218 186146 696454
rect 186382 696218 221826 696454
rect 222062 696218 222146 696454
rect 222382 696218 257826 696454
rect 258062 696218 258146 696454
rect 258382 696218 293826 696454
rect 294062 696218 294146 696454
rect 294382 696218 329826 696454
rect 330062 696218 330146 696454
rect 330382 696218 365826 696454
rect 366062 696218 366146 696454
rect 366382 696218 401826 696454
rect 402062 696218 402146 696454
rect 402382 696218 437826 696454
rect 438062 696218 438146 696454
rect 438382 696218 473826 696454
rect 474062 696218 474146 696454
rect 474382 696218 509826 696454
rect 510062 696218 510146 696454
rect 510382 696218 545826 696454
rect 546062 696218 546146 696454
rect 546382 696218 577826 696454
rect 578062 696218 578146 696454
rect 578382 696218 585342 696454
rect 585578 696218 585662 696454
rect 585898 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -1974 696134
rect -1738 695898 -1654 696134
rect -1418 695898 1826 696134
rect 2062 695898 2146 696134
rect 2382 695898 5826 696134
rect 6062 695898 6146 696134
rect 6382 695898 41826 696134
rect 42062 695898 42146 696134
rect 42382 695898 77826 696134
rect 78062 695898 78146 696134
rect 78382 695898 113826 696134
rect 114062 695898 114146 696134
rect 114382 695898 149826 696134
rect 150062 695898 150146 696134
rect 150382 695898 185826 696134
rect 186062 695898 186146 696134
rect 186382 695898 221826 696134
rect 222062 695898 222146 696134
rect 222382 695898 257826 696134
rect 258062 695898 258146 696134
rect 258382 695898 293826 696134
rect 294062 695898 294146 696134
rect 294382 695898 329826 696134
rect 330062 695898 330146 696134
rect 330382 695898 365826 696134
rect 366062 695898 366146 696134
rect 366382 695898 401826 696134
rect 402062 695898 402146 696134
rect 402382 695898 437826 696134
rect 438062 695898 438146 696134
rect 438382 695898 473826 696134
rect 474062 695898 474146 696134
rect 474382 695898 509826 696134
rect 510062 695898 510146 696134
rect 510382 695898 545826 696134
rect 546062 695898 546146 696134
rect 546382 695898 577826 696134
rect 578062 695898 578146 696134
rect 578382 695898 585342 696134
rect 585578 695898 585662 696134
rect 585898 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 664174 592650 664206
rect -8726 663938 -2934 664174
rect -2698 663938 -2614 664174
rect -2378 663938 9546 664174
rect 9782 663938 9866 664174
rect 10102 663938 189546 664174
rect 189782 663938 189866 664174
rect 190102 663938 369546 664174
rect 369782 663938 369866 664174
rect 370102 663938 405546 664174
rect 405782 663938 405866 664174
rect 406102 663938 572374 664174
rect 572610 663938 572694 664174
rect 572930 663938 581546 664174
rect 581782 663938 581866 664174
rect 582102 663938 586302 664174
rect 586538 663938 586622 664174
rect 586858 663938 592650 664174
rect -8726 663854 592650 663938
rect -8726 663618 -2934 663854
rect -2698 663618 -2614 663854
rect -2378 663618 9546 663854
rect 9782 663618 9866 663854
rect 10102 663618 189546 663854
rect 189782 663618 189866 663854
rect 190102 663618 369546 663854
rect 369782 663618 369866 663854
rect 370102 663618 405546 663854
rect 405782 663618 405866 663854
rect 406102 663618 572374 663854
rect 572610 663618 572694 663854
rect 572930 663618 581546 663854
rect 581782 663618 581866 663854
rect 582102 663618 586302 663854
rect 586538 663618 586622 663854
rect 586858 663618 592650 663854
rect -8726 663586 592650 663618
rect -8726 660454 592650 660486
rect -8726 660218 -1974 660454
rect -1738 660218 -1654 660454
rect -1418 660218 1826 660454
rect 2062 660218 2146 660454
rect 2382 660218 5826 660454
rect 6062 660218 6146 660454
rect 6382 660218 185826 660454
rect 186062 660218 186146 660454
rect 186382 660218 365826 660454
rect 366062 660218 366146 660454
rect 366382 660218 401826 660454
rect 402062 660218 402146 660454
rect 402382 660218 568510 660454
rect 568746 660218 568830 660454
rect 569066 660218 577826 660454
rect 578062 660218 578146 660454
rect 578382 660218 585342 660454
rect 585578 660218 585662 660454
rect 585898 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -1974 660134
rect -1738 659898 -1654 660134
rect -1418 659898 1826 660134
rect 2062 659898 2146 660134
rect 2382 659898 5826 660134
rect 6062 659898 6146 660134
rect 6382 659898 185826 660134
rect 186062 659898 186146 660134
rect 186382 659898 365826 660134
rect 366062 659898 366146 660134
rect 366382 659898 401826 660134
rect 402062 659898 402146 660134
rect 402382 659898 568510 660134
rect 568746 659898 568830 660134
rect 569066 659898 577826 660134
rect 578062 659898 578146 660134
rect 578382 659898 585342 660134
rect 585578 659898 585662 660134
rect 585898 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 628174 592650 628206
rect -8726 627938 -2934 628174
rect -2698 627938 -2614 628174
rect -2378 627938 9546 628174
rect 9782 627938 9866 628174
rect 10102 627938 189546 628174
rect 189782 627938 189866 628174
rect 190102 627938 369546 628174
rect 369782 627938 369866 628174
rect 370102 627938 405546 628174
rect 405782 627938 405866 628174
rect 406102 627938 572374 628174
rect 572610 627938 572694 628174
rect 572930 627938 581546 628174
rect 581782 627938 581866 628174
rect 582102 627938 586302 628174
rect 586538 627938 586622 628174
rect 586858 627938 592650 628174
rect -8726 627854 592650 627938
rect -8726 627618 -2934 627854
rect -2698 627618 -2614 627854
rect -2378 627618 9546 627854
rect 9782 627618 9866 627854
rect 10102 627618 189546 627854
rect 189782 627618 189866 627854
rect 190102 627618 369546 627854
rect 369782 627618 369866 627854
rect 370102 627618 405546 627854
rect 405782 627618 405866 627854
rect 406102 627618 572374 627854
rect 572610 627618 572694 627854
rect 572930 627618 581546 627854
rect 581782 627618 581866 627854
rect 582102 627618 586302 627854
rect 586538 627618 586622 627854
rect 586858 627618 592650 627854
rect -8726 627586 592650 627618
rect -8726 624454 592650 624486
rect -8726 624218 -1974 624454
rect -1738 624218 -1654 624454
rect -1418 624218 1826 624454
rect 2062 624218 2146 624454
rect 2382 624218 5826 624454
rect 6062 624218 6146 624454
rect 6382 624218 185826 624454
rect 186062 624218 186146 624454
rect 186382 624218 365826 624454
rect 366062 624218 366146 624454
rect 366382 624218 401826 624454
rect 402062 624218 402146 624454
rect 402382 624218 568510 624454
rect 568746 624218 568830 624454
rect 569066 624218 577826 624454
rect 578062 624218 578146 624454
rect 578382 624218 585342 624454
rect 585578 624218 585662 624454
rect 585898 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -1974 624134
rect -1738 623898 -1654 624134
rect -1418 623898 1826 624134
rect 2062 623898 2146 624134
rect 2382 623898 5826 624134
rect 6062 623898 6146 624134
rect 6382 623898 185826 624134
rect 186062 623898 186146 624134
rect 186382 623898 365826 624134
rect 366062 623898 366146 624134
rect 366382 623898 401826 624134
rect 402062 623898 402146 624134
rect 402382 623898 568510 624134
rect 568746 623898 568830 624134
rect 569066 623898 577826 624134
rect 578062 623898 578146 624134
rect 578382 623898 585342 624134
rect 585578 623898 585662 624134
rect 585898 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 592174 592650 592206
rect -8726 591938 -2934 592174
rect -2698 591938 -2614 592174
rect -2378 591938 9546 592174
rect 9782 591938 9866 592174
rect 10102 591938 45546 592174
rect 45782 591938 45866 592174
rect 46102 591938 81546 592174
rect 81782 591938 81866 592174
rect 82102 591938 117546 592174
rect 117782 591938 117866 592174
rect 118102 591938 153546 592174
rect 153782 591938 153866 592174
rect 154102 591938 189546 592174
rect 189782 591938 189866 592174
rect 190102 591938 225546 592174
rect 225782 591938 225866 592174
rect 226102 591938 261546 592174
rect 261782 591938 261866 592174
rect 262102 591938 297546 592174
rect 297782 591938 297866 592174
rect 298102 591938 333546 592174
rect 333782 591938 333866 592174
rect 334102 591938 369546 592174
rect 369782 591938 369866 592174
rect 370102 591938 405546 592174
rect 405782 591938 405866 592174
rect 406102 591938 441546 592174
rect 441782 591938 441866 592174
rect 442102 591938 477546 592174
rect 477782 591938 477866 592174
rect 478102 591938 513546 592174
rect 513782 591938 513866 592174
rect 514102 591938 549546 592174
rect 549782 591938 549866 592174
rect 550102 591938 581546 592174
rect 581782 591938 581866 592174
rect 582102 591938 586302 592174
rect 586538 591938 586622 592174
rect 586858 591938 592650 592174
rect -8726 591854 592650 591938
rect -8726 591618 -2934 591854
rect -2698 591618 -2614 591854
rect -2378 591618 9546 591854
rect 9782 591618 9866 591854
rect 10102 591618 45546 591854
rect 45782 591618 45866 591854
rect 46102 591618 81546 591854
rect 81782 591618 81866 591854
rect 82102 591618 117546 591854
rect 117782 591618 117866 591854
rect 118102 591618 153546 591854
rect 153782 591618 153866 591854
rect 154102 591618 189546 591854
rect 189782 591618 189866 591854
rect 190102 591618 225546 591854
rect 225782 591618 225866 591854
rect 226102 591618 261546 591854
rect 261782 591618 261866 591854
rect 262102 591618 297546 591854
rect 297782 591618 297866 591854
rect 298102 591618 333546 591854
rect 333782 591618 333866 591854
rect 334102 591618 369546 591854
rect 369782 591618 369866 591854
rect 370102 591618 405546 591854
rect 405782 591618 405866 591854
rect 406102 591618 441546 591854
rect 441782 591618 441866 591854
rect 442102 591618 477546 591854
rect 477782 591618 477866 591854
rect 478102 591618 513546 591854
rect 513782 591618 513866 591854
rect 514102 591618 549546 591854
rect 549782 591618 549866 591854
rect 550102 591618 581546 591854
rect 581782 591618 581866 591854
rect 582102 591618 586302 591854
rect 586538 591618 586622 591854
rect 586858 591618 592650 591854
rect -8726 591586 592650 591618
rect -8726 588454 592650 588486
rect -8726 588218 -1974 588454
rect -1738 588218 -1654 588454
rect -1418 588218 1826 588454
rect 2062 588218 2146 588454
rect 2382 588218 5826 588454
rect 6062 588218 6146 588454
rect 6382 588218 41826 588454
rect 42062 588218 42146 588454
rect 42382 588218 77826 588454
rect 78062 588218 78146 588454
rect 78382 588218 113826 588454
rect 114062 588218 114146 588454
rect 114382 588218 149826 588454
rect 150062 588218 150146 588454
rect 150382 588218 185826 588454
rect 186062 588218 186146 588454
rect 186382 588218 221826 588454
rect 222062 588218 222146 588454
rect 222382 588218 257826 588454
rect 258062 588218 258146 588454
rect 258382 588218 293826 588454
rect 294062 588218 294146 588454
rect 294382 588218 329826 588454
rect 330062 588218 330146 588454
rect 330382 588218 365826 588454
rect 366062 588218 366146 588454
rect 366382 588218 401826 588454
rect 402062 588218 402146 588454
rect 402382 588218 437826 588454
rect 438062 588218 438146 588454
rect 438382 588218 473826 588454
rect 474062 588218 474146 588454
rect 474382 588218 509826 588454
rect 510062 588218 510146 588454
rect 510382 588218 545826 588454
rect 546062 588218 546146 588454
rect 546382 588218 577826 588454
rect 578062 588218 578146 588454
rect 578382 588218 585342 588454
rect 585578 588218 585662 588454
rect 585898 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -1974 588134
rect -1738 587898 -1654 588134
rect -1418 587898 1826 588134
rect 2062 587898 2146 588134
rect 2382 587898 5826 588134
rect 6062 587898 6146 588134
rect 6382 587898 41826 588134
rect 42062 587898 42146 588134
rect 42382 587898 77826 588134
rect 78062 587898 78146 588134
rect 78382 587898 113826 588134
rect 114062 587898 114146 588134
rect 114382 587898 149826 588134
rect 150062 587898 150146 588134
rect 150382 587898 185826 588134
rect 186062 587898 186146 588134
rect 186382 587898 221826 588134
rect 222062 587898 222146 588134
rect 222382 587898 257826 588134
rect 258062 587898 258146 588134
rect 258382 587898 293826 588134
rect 294062 587898 294146 588134
rect 294382 587898 329826 588134
rect 330062 587898 330146 588134
rect 330382 587898 365826 588134
rect 366062 587898 366146 588134
rect 366382 587898 401826 588134
rect 402062 587898 402146 588134
rect 402382 587898 437826 588134
rect 438062 587898 438146 588134
rect 438382 587898 473826 588134
rect 474062 587898 474146 588134
rect 474382 587898 509826 588134
rect 510062 587898 510146 588134
rect 510382 587898 545826 588134
rect 546062 587898 546146 588134
rect 546382 587898 577826 588134
rect 578062 587898 578146 588134
rect 578382 587898 585342 588134
rect 585578 587898 585662 588134
rect 585898 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 556174 592650 556206
rect -8726 555938 -2934 556174
rect -2698 555938 -2614 556174
rect -2378 555938 9546 556174
rect 9782 555938 9866 556174
rect 10102 555938 189546 556174
rect 189782 555938 189866 556174
rect 190102 555938 225546 556174
rect 225782 555938 225866 556174
rect 226102 555938 261546 556174
rect 261782 555938 261866 556174
rect 262102 555938 297546 556174
rect 297782 555938 297866 556174
rect 298102 555938 333546 556174
rect 333782 555938 333866 556174
rect 334102 555938 369546 556174
rect 369782 555938 369866 556174
rect 370102 555938 405546 556174
rect 405782 555938 405866 556174
rect 406102 555938 572374 556174
rect 572610 555938 572694 556174
rect 572930 555938 581546 556174
rect 581782 555938 581866 556174
rect 582102 555938 586302 556174
rect 586538 555938 586622 556174
rect 586858 555938 592650 556174
rect -8726 555854 592650 555938
rect -8726 555618 -2934 555854
rect -2698 555618 -2614 555854
rect -2378 555618 9546 555854
rect 9782 555618 9866 555854
rect 10102 555618 189546 555854
rect 189782 555618 189866 555854
rect 190102 555618 225546 555854
rect 225782 555618 225866 555854
rect 226102 555618 261546 555854
rect 261782 555618 261866 555854
rect 262102 555618 297546 555854
rect 297782 555618 297866 555854
rect 298102 555618 333546 555854
rect 333782 555618 333866 555854
rect 334102 555618 369546 555854
rect 369782 555618 369866 555854
rect 370102 555618 405546 555854
rect 405782 555618 405866 555854
rect 406102 555618 572374 555854
rect 572610 555618 572694 555854
rect 572930 555618 581546 555854
rect 581782 555618 581866 555854
rect 582102 555618 586302 555854
rect 586538 555618 586622 555854
rect 586858 555618 592650 555854
rect -8726 555586 592650 555618
rect -8726 552454 592650 552486
rect -8726 552218 -1974 552454
rect -1738 552218 -1654 552454
rect -1418 552218 1826 552454
rect 2062 552218 2146 552454
rect 2382 552218 5826 552454
rect 6062 552218 6146 552454
rect 6382 552218 185826 552454
rect 186062 552218 186146 552454
rect 186382 552218 221826 552454
rect 222062 552218 222146 552454
rect 222382 552218 257826 552454
rect 258062 552218 258146 552454
rect 258382 552218 293826 552454
rect 294062 552218 294146 552454
rect 294382 552218 329826 552454
rect 330062 552218 330146 552454
rect 330382 552218 365826 552454
rect 366062 552218 366146 552454
rect 366382 552218 401826 552454
rect 402062 552218 402146 552454
rect 402382 552218 568510 552454
rect 568746 552218 568830 552454
rect 569066 552218 577826 552454
rect 578062 552218 578146 552454
rect 578382 552218 585342 552454
rect 585578 552218 585662 552454
rect 585898 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -1974 552134
rect -1738 551898 -1654 552134
rect -1418 551898 1826 552134
rect 2062 551898 2146 552134
rect 2382 551898 5826 552134
rect 6062 551898 6146 552134
rect 6382 551898 185826 552134
rect 186062 551898 186146 552134
rect 186382 551898 221826 552134
rect 222062 551898 222146 552134
rect 222382 551898 257826 552134
rect 258062 551898 258146 552134
rect 258382 551898 293826 552134
rect 294062 551898 294146 552134
rect 294382 551898 329826 552134
rect 330062 551898 330146 552134
rect 330382 551898 365826 552134
rect 366062 551898 366146 552134
rect 366382 551898 401826 552134
rect 402062 551898 402146 552134
rect 402382 551898 568510 552134
rect 568746 551898 568830 552134
rect 569066 551898 577826 552134
rect 578062 551898 578146 552134
rect 578382 551898 585342 552134
rect 585578 551898 585662 552134
rect 585898 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 520174 592650 520206
rect -8726 519938 -2934 520174
rect -2698 519938 -2614 520174
rect -2378 519938 9546 520174
rect 9782 519938 9866 520174
rect 10102 519938 189546 520174
rect 189782 519938 189866 520174
rect 190102 519938 225546 520174
rect 225782 519938 225866 520174
rect 226102 519938 261546 520174
rect 261782 519938 261866 520174
rect 262102 519938 297546 520174
rect 297782 519938 297866 520174
rect 298102 519938 333546 520174
rect 333782 519938 333866 520174
rect 334102 519938 369546 520174
rect 369782 519938 369866 520174
rect 370102 519938 405546 520174
rect 405782 519938 405866 520174
rect 406102 519938 572374 520174
rect 572610 519938 572694 520174
rect 572930 519938 581546 520174
rect 581782 519938 581866 520174
rect 582102 519938 586302 520174
rect 586538 519938 586622 520174
rect 586858 519938 592650 520174
rect -8726 519854 592650 519938
rect -8726 519618 -2934 519854
rect -2698 519618 -2614 519854
rect -2378 519618 9546 519854
rect 9782 519618 9866 519854
rect 10102 519618 189546 519854
rect 189782 519618 189866 519854
rect 190102 519618 225546 519854
rect 225782 519618 225866 519854
rect 226102 519618 261546 519854
rect 261782 519618 261866 519854
rect 262102 519618 297546 519854
rect 297782 519618 297866 519854
rect 298102 519618 333546 519854
rect 333782 519618 333866 519854
rect 334102 519618 369546 519854
rect 369782 519618 369866 519854
rect 370102 519618 405546 519854
rect 405782 519618 405866 519854
rect 406102 519618 572374 519854
rect 572610 519618 572694 519854
rect 572930 519618 581546 519854
rect 581782 519618 581866 519854
rect 582102 519618 586302 519854
rect 586538 519618 586622 519854
rect 586858 519618 592650 519854
rect -8726 519586 592650 519618
rect -8726 516454 592650 516486
rect -8726 516218 -1974 516454
rect -1738 516218 -1654 516454
rect -1418 516218 1826 516454
rect 2062 516218 2146 516454
rect 2382 516218 5826 516454
rect 6062 516218 6146 516454
rect 6382 516218 185826 516454
rect 186062 516218 186146 516454
rect 186382 516218 221826 516454
rect 222062 516218 222146 516454
rect 222382 516218 257826 516454
rect 258062 516218 258146 516454
rect 258382 516218 293826 516454
rect 294062 516218 294146 516454
rect 294382 516218 329826 516454
rect 330062 516218 330146 516454
rect 330382 516218 365826 516454
rect 366062 516218 366146 516454
rect 366382 516218 401826 516454
rect 402062 516218 402146 516454
rect 402382 516218 568510 516454
rect 568746 516218 568830 516454
rect 569066 516218 577826 516454
rect 578062 516218 578146 516454
rect 578382 516218 585342 516454
rect 585578 516218 585662 516454
rect 585898 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -1974 516134
rect -1738 515898 -1654 516134
rect -1418 515898 1826 516134
rect 2062 515898 2146 516134
rect 2382 515898 5826 516134
rect 6062 515898 6146 516134
rect 6382 515898 185826 516134
rect 186062 515898 186146 516134
rect 186382 515898 221826 516134
rect 222062 515898 222146 516134
rect 222382 515898 257826 516134
rect 258062 515898 258146 516134
rect 258382 515898 293826 516134
rect 294062 515898 294146 516134
rect 294382 515898 329826 516134
rect 330062 515898 330146 516134
rect 330382 515898 365826 516134
rect 366062 515898 366146 516134
rect 366382 515898 401826 516134
rect 402062 515898 402146 516134
rect 402382 515898 568510 516134
rect 568746 515898 568830 516134
rect 569066 515898 577826 516134
rect 578062 515898 578146 516134
rect 578382 515898 585342 516134
rect 585578 515898 585662 516134
rect 585898 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 484174 592650 484206
rect -8726 483938 -2934 484174
rect -2698 483938 -2614 484174
rect -2378 483938 9546 484174
rect 9782 483938 9866 484174
rect 10102 483938 45546 484174
rect 45782 483938 45866 484174
rect 46102 483938 81546 484174
rect 81782 483938 81866 484174
rect 82102 483938 117546 484174
rect 117782 483938 117866 484174
rect 118102 483938 153546 484174
rect 153782 483938 153866 484174
rect 154102 483938 189546 484174
rect 189782 483938 189866 484174
rect 190102 483938 225546 484174
rect 225782 483938 225866 484174
rect 226102 483938 261546 484174
rect 261782 483938 261866 484174
rect 262102 483938 297546 484174
rect 297782 483938 297866 484174
rect 298102 483938 333546 484174
rect 333782 483938 333866 484174
rect 334102 483938 369546 484174
rect 369782 483938 369866 484174
rect 370102 483938 405546 484174
rect 405782 483938 405866 484174
rect 406102 483938 441546 484174
rect 441782 483938 441866 484174
rect 442102 483938 477546 484174
rect 477782 483938 477866 484174
rect 478102 483938 513546 484174
rect 513782 483938 513866 484174
rect 514102 483938 549546 484174
rect 549782 483938 549866 484174
rect 550102 483938 581546 484174
rect 581782 483938 581866 484174
rect 582102 483938 586302 484174
rect 586538 483938 586622 484174
rect 586858 483938 592650 484174
rect -8726 483854 592650 483938
rect -8726 483618 -2934 483854
rect -2698 483618 -2614 483854
rect -2378 483618 9546 483854
rect 9782 483618 9866 483854
rect 10102 483618 45546 483854
rect 45782 483618 45866 483854
rect 46102 483618 81546 483854
rect 81782 483618 81866 483854
rect 82102 483618 117546 483854
rect 117782 483618 117866 483854
rect 118102 483618 153546 483854
rect 153782 483618 153866 483854
rect 154102 483618 189546 483854
rect 189782 483618 189866 483854
rect 190102 483618 225546 483854
rect 225782 483618 225866 483854
rect 226102 483618 261546 483854
rect 261782 483618 261866 483854
rect 262102 483618 297546 483854
rect 297782 483618 297866 483854
rect 298102 483618 333546 483854
rect 333782 483618 333866 483854
rect 334102 483618 369546 483854
rect 369782 483618 369866 483854
rect 370102 483618 405546 483854
rect 405782 483618 405866 483854
rect 406102 483618 441546 483854
rect 441782 483618 441866 483854
rect 442102 483618 477546 483854
rect 477782 483618 477866 483854
rect 478102 483618 513546 483854
rect 513782 483618 513866 483854
rect 514102 483618 549546 483854
rect 549782 483618 549866 483854
rect 550102 483618 581546 483854
rect 581782 483618 581866 483854
rect 582102 483618 586302 483854
rect 586538 483618 586622 483854
rect 586858 483618 592650 483854
rect -8726 483586 592650 483618
rect -8726 480454 592650 480486
rect -8726 480218 -1974 480454
rect -1738 480218 -1654 480454
rect -1418 480218 1826 480454
rect 2062 480218 2146 480454
rect 2382 480218 5826 480454
rect 6062 480218 6146 480454
rect 6382 480218 41826 480454
rect 42062 480218 42146 480454
rect 42382 480218 77826 480454
rect 78062 480218 78146 480454
rect 78382 480218 113826 480454
rect 114062 480218 114146 480454
rect 114382 480218 149826 480454
rect 150062 480218 150146 480454
rect 150382 480218 185826 480454
rect 186062 480218 186146 480454
rect 186382 480218 221826 480454
rect 222062 480218 222146 480454
rect 222382 480218 257826 480454
rect 258062 480218 258146 480454
rect 258382 480218 293826 480454
rect 294062 480218 294146 480454
rect 294382 480218 329826 480454
rect 330062 480218 330146 480454
rect 330382 480218 365826 480454
rect 366062 480218 366146 480454
rect 366382 480218 401826 480454
rect 402062 480218 402146 480454
rect 402382 480218 437826 480454
rect 438062 480218 438146 480454
rect 438382 480218 473826 480454
rect 474062 480218 474146 480454
rect 474382 480218 509826 480454
rect 510062 480218 510146 480454
rect 510382 480218 545826 480454
rect 546062 480218 546146 480454
rect 546382 480218 577826 480454
rect 578062 480218 578146 480454
rect 578382 480218 585342 480454
rect 585578 480218 585662 480454
rect 585898 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -1974 480134
rect -1738 479898 -1654 480134
rect -1418 479898 1826 480134
rect 2062 479898 2146 480134
rect 2382 479898 5826 480134
rect 6062 479898 6146 480134
rect 6382 479898 41826 480134
rect 42062 479898 42146 480134
rect 42382 479898 77826 480134
rect 78062 479898 78146 480134
rect 78382 479898 113826 480134
rect 114062 479898 114146 480134
rect 114382 479898 149826 480134
rect 150062 479898 150146 480134
rect 150382 479898 185826 480134
rect 186062 479898 186146 480134
rect 186382 479898 221826 480134
rect 222062 479898 222146 480134
rect 222382 479898 257826 480134
rect 258062 479898 258146 480134
rect 258382 479898 293826 480134
rect 294062 479898 294146 480134
rect 294382 479898 329826 480134
rect 330062 479898 330146 480134
rect 330382 479898 365826 480134
rect 366062 479898 366146 480134
rect 366382 479898 401826 480134
rect 402062 479898 402146 480134
rect 402382 479898 437826 480134
rect 438062 479898 438146 480134
rect 438382 479898 473826 480134
rect 474062 479898 474146 480134
rect 474382 479898 509826 480134
rect 510062 479898 510146 480134
rect 510382 479898 545826 480134
rect 546062 479898 546146 480134
rect 546382 479898 577826 480134
rect 578062 479898 578146 480134
rect 578382 479898 585342 480134
rect 585578 479898 585662 480134
rect 585898 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 448174 592650 448206
rect -8726 447938 -2934 448174
rect -2698 447938 -2614 448174
rect -2378 447938 9546 448174
rect 9782 447938 9866 448174
rect 10102 447938 189546 448174
rect 189782 447938 189866 448174
rect 190102 447938 225546 448174
rect 225782 447938 225866 448174
rect 226102 447938 261546 448174
rect 261782 447938 261866 448174
rect 262102 447938 297546 448174
rect 297782 447938 297866 448174
rect 298102 447938 333546 448174
rect 333782 447938 333866 448174
rect 334102 447938 369546 448174
rect 369782 447938 369866 448174
rect 370102 447938 405546 448174
rect 405782 447938 405866 448174
rect 406102 447938 572374 448174
rect 572610 447938 572694 448174
rect 572930 447938 581546 448174
rect 581782 447938 581866 448174
rect 582102 447938 586302 448174
rect 586538 447938 586622 448174
rect 586858 447938 592650 448174
rect -8726 447854 592650 447938
rect -8726 447618 -2934 447854
rect -2698 447618 -2614 447854
rect -2378 447618 9546 447854
rect 9782 447618 9866 447854
rect 10102 447618 189546 447854
rect 189782 447618 189866 447854
rect 190102 447618 225546 447854
rect 225782 447618 225866 447854
rect 226102 447618 261546 447854
rect 261782 447618 261866 447854
rect 262102 447618 297546 447854
rect 297782 447618 297866 447854
rect 298102 447618 333546 447854
rect 333782 447618 333866 447854
rect 334102 447618 369546 447854
rect 369782 447618 369866 447854
rect 370102 447618 405546 447854
rect 405782 447618 405866 447854
rect 406102 447618 572374 447854
rect 572610 447618 572694 447854
rect 572930 447618 581546 447854
rect 581782 447618 581866 447854
rect 582102 447618 586302 447854
rect 586538 447618 586622 447854
rect 586858 447618 592650 447854
rect -8726 447586 592650 447618
rect -8726 444454 592650 444486
rect -8726 444218 -1974 444454
rect -1738 444218 -1654 444454
rect -1418 444218 1826 444454
rect 2062 444218 2146 444454
rect 2382 444218 5826 444454
rect 6062 444218 6146 444454
rect 6382 444218 185826 444454
rect 186062 444218 186146 444454
rect 186382 444218 221826 444454
rect 222062 444218 222146 444454
rect 222382 444218 257826 444454
rect 258062 444218 258146 444454
rect 258382 444218 293826 444454
rect 294062 444218 294146 444454
rect 294382 444218 329826 444454
rect 330062 444218 330146 444454
rect 330382 444218 365826 444454
rect 366062 444218 366146 444454
rect 366382 444218 401826 444454
rect 402062 444218 402146 444454
rect 402382 444218 568510 444454
rect 568746 444218 568830 444454
rect 569066 444218 577826 444454
rect 578062 444218 578146 444454
rect 578382 444218 585342 444454
rect 585578 444218 585662 444454
rect 585898 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -1974 444134
rect -1738 443898 -1654 444134
rect -1418 443898 1826 444134
rect 2062 443898 2146 444134
rect 2382 443898 5826 444134
rect 6062 443898 6146 444134
rect 6382 443898 185826 444134
rect 186062 443898 186146 444134
rect 186382 443898 221826 444134
rect 222062 443898 222146 444134
rect 222382 443898 257826 444134
rect 258062 443898 258146 444134
rect 258382 443898 293826 444134
rect 294062 443898 294146 444134
rect 294382 443898 329826 444134
rect 330062 443898 330146 444134
rect 330382 443898 365826 444134
rect 366062 443898 366146 444134
rect 366382 443898 401826 444134
rect 402062 443898 402146 444134
rect 402382 443898 568510 444134
rect 568746 443898 568830 444134
rect 569066 443898 577826 444134
rect 578062 443898 578146 444134
rect 578382 443898 585342 444134
rect 585578 443898 585662 444134
rect 585898 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 412174 592650 412206
rect -8726 411938 -2934 412174
rect -2698 411938 -2614 412174
rect -2378 411938 9546 412174
rect 9782 411938 9866 412174
rect 10102 411938 189546 412174
rect 189782 411938 189866 412174
rect 190102 411938 225546 412174
rect 225782 411938 225866 412174
rect 226102 411938 261546 412174
rect 261782 411938 261866 412174
rect 262102 411938 297546 412174
rect 297782 411938 297866 412174
rect 298102 411938 333546 412174
rect 333782 411938 333866 412174
rect 334102 411938 369546 412174
rect 369782 411938 369866 412174
rect 370102 411938 405546 412174
rect 405782 411938 405866 412174
rect 406102 411938 572374 412174
rect 572610 411938 572694 412174
rect 572930 411938 581546 412174
rect 581782 411938 581866 412174
rect 582102 411938 586302 412174
rect 586538 411938 586622 412174
rect 586858 411938 592650 412174
rect -8726 411854 592650 411938
rect -8726 411618 -2934 411854
rect -2698 411618 -2614 411854
rect -2378 411618 9546 411854
rect 9782 411618 9866 411854
rect 10102 411618 189546 411854
rect 189782 411618 189866 411854
rect 190102 411618 225546 411854
rect 225782 411618 225866 411854
rect 226102 411618 261546 411854
rect 261782 411618 261866 411854
rect 262102 411618 297546 411854
rect 297782 411618 297866 411854
rect 298102 411618 333546 411854
rect 333782 411618 333866 411854
rect 334102 411618 369546 411854
rect 369782 411618 369866 411854
rect 370102 411618 405546 411854
rect 405782 411618 405866 411854
rect 406102 411618 572374 411854
rect 572610 411618 572694 411854
rect 572930 411618 581546 411854
rect 581782 411618 581866 411854
rect 582102 411618 586302 411854
rect 586538 411618 586622 411854
rect 586858 411618 592650 411854
rect -8726 411586 592650 411618
rect -8726 408454 592650 408486
rect -8726 408218 -1974 408454
rect -1738 408218 -1654 408454
rect -1418 408218 1826 408454
rect 2062 408218 2146 408454
rect 2382 408218 5826 408454
rect 6062 408218 6146 408454
rect 6382 408218 185826 408454
rect 186062 408218 186146 408454
rect 186382 408218 221826 408454
rect 222062 408218 222146 408454
rect 222382 408218 257826 408454
rect 258062 408218 258146 408454
rect 258382 408218 293826 408454
rect 294062 408218 294146 408454
rect 294382 408218 329826 408454
rect 330062 408218 330146 408454
rect 330382 408218 365826 408454
rect 366062 408218 366146 408454
rect 366382 408218 401826 408454
rect 402062 408218 402146 408454
rect 402382 408218 568510 408454
rect 568746 408218 568830 408454
rect 569066 408218 577826 408454
rect 578062 408218 578146 408454
rect 578382 408218 585342 408454
rect 585578 408218 585662 408454
rect 585898 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -1974 408134
rect -1738 407898 -1654 408134
rect -1418 407898 1826 408134
rect 2062 407898 2146 408134
rect 2382 407898 5826 408134
rect 6062 407898 6146 408134
rect 6382 407898 185826 408134
rect 186062 407898 186146 408134
rect 186382 407898 221826 408134
rect 222062 407898 222146 408134
rect 222382 407898 257826 408134
rect 258062 407898 258146 408134
rect 258382 407898 293826 408134
rect 294062 407898 294146 408134
rect 294382 407898 329826 408134
rect 330062 407898 330146 408134
rect 330382 407898 365826 408134
rect 366062 407898 366146 408134
rect 366382 407898 401826 408134
rect 402062 407898 402146 408134
rect 402382 407898 568510 408134
rect 568746 407898 568830 408134
rect 569066 407898 577826 408134
rect 578062 407898 578146 408134
rect 578382 407898 585342 408134
rect 585578 407898 585662 408134
rect 585898 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 376174 592650 376206
rect -8726 375938 -2934 376174
rect -2698 375938 -2614 376174
rect -2378 375938 9546 376174
rect 9782 375938 9866 376174
rect 10102 375938 189546 376174
rect 189782 375938 189866 376174
rect 190102 375938 225546 376174
rect 225782 375938 225866 376174
rect 226102 375938 261546 376174
rect 261782 375938 261866 376174
rect 262102 375938 297546 376174
rect 297782 375938 297866 376174
rect 298102 375938 333546 376174
rect 333782 375938 333866 376174
rect 334102 375938 369546 376174
rect 369782 375938 369866 376174
rect 370102 375938 405546 376174
rect 405782 375938 405866 376174
rect 406102 375938 572374 376174
rect 572610 375938 572694 376174
rect 572930 375938 581546 376174
rect 581782 375938 581866 376174
rect 582102 375938 586302 376174
rect 586538 375938 586622 376174
rect 586858 375938 592650 376174
rect -8726 375854 592650 375938
rect -8726 375618 -2934 375854
rect -2698 375618 -2614 375854
rect -2378 375618 9546 375854
rect 9782 375618 9866 375854
rect 10102 375618 189546 375854
rect 189782 375618 189866 375854
rect 190102 375618 225546 375854
rect 225782 375618 225866 375854
rect 226102 375618 261546 375854
rect 261782 375618 261866 375854
rect 262102 375618 297546 375854
rect 297782 375618 297866 375854
rect 298102 375618 333546 375854
rect 333782 375618 333866 375854
rect 334102 375618 369546 375854
rect 369782 375618 369866 375854
rect 370102 375618 405546 375854
rect 405782 375618 405866 375854
rect 406102 375618 572374 375854
rect 572610 375618 572694 375854
rect 572930 375618 581546 375854
rect 581782 375618 581866 375854
rect 582102 375618 586302 375854
rect 586538 375618 586622 375854
rect 586858 375618 592650 375854
rect -8726 375586 592650 375618
rect -8726 372454 592650 372486
rect -8726 372218 -1974 372454
rect -1738 372218 -1654 372454
rect -1418 372218 1826 372454
rect 2062 372218 2146 372454
rect 2382 372218 5826 372454
rect 6062 372218 6146 372454
rect 6382 372218 185826 372454
rect 186062 372218 186146 372454
rect 186382 372218 221826 372454
rect 222062 372218 222146 372454
rect 222382 372218 257826 372454
rect 258062 372218 258146 372454
rect 258382 372218 293826 372454
rect 294062 372218 294146 372454
rect 294382 372218 329826 372454
rect 330062 372218 330146 372454
rect 330382 372218 365826 372454
rect 366062 372218 366146 372454
rect 366382 372218 401826 372454
rect 402062 372218 402146 372454
rect 402382 372218 568510 372454
rect 568746 372218 568830 372454
rect 569066 372218 577826 372454
rect 578062 372218 578146 372454
rect 578382 372218 585342 372454
rect 585578 372218 585662 372454
rect 585898 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -1974 372134
rect -1738 371898 -1654 372134
rect -1418 371898 1826 372134
rect 2062 371898 2146 372134
rect 2382 371898 5826 372134
rect 6062 371898 6146 372134
rect 6382 371898 185826 372134
rect 186062 371898 186146 372134
rect 186382 371898 221826 372134
rect 222062 371898 222146 372134
rect 222382 371898 257826 372134
rect 258062 371898 258146 372134
rect 258382 371898 293826 372134
rect 294062 371898 294146 372134
rect 294382 371898 329826 372134
rect 330062 371898 330146 372134
rect 330382 371898 365826 372134
rect 366062 371898 366146 372134
rect 366382 371898 401826 372134
rect 402062 371898 402146 372134
rect 402382 371898 568510 372134
rect 568746 371898 568830 372134
rect 569066 371898 577826 372134
rect 578062 371898 578146 372134
rect 578382 371898 585342 372134
rect 585578 371898 585662 372134
rect 585898 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 340174 592650 340206
rect -8726 339938 -2934 340174
rect -2698 339938 -2614 340174
rect -2378 339938 9546 340174
rect 9782 339938 9866 340174
rect 10102 339938 189546 340174
rect 189782 339938 189866 340174
rect 190102 339938 225546 340174
rect 225782 339938 225866 340174
rect 226102 339938 261546 340174
rect 261782 339938 261866 340174
rect 262102 339938 297546 340174
rect 297782 339938 297866 340174
rect 298102 339938 333546 340174
rect 333782 339938 333866 340174
rect 334102 339938 369546 340174
rect 369782 339938 369866 340174
rect 370102 339938 405546 340174
rect 405782 339938 405866 340174
rect 406102 339938 572374 340174
rect 572610 339938 572694 340174
rect 572930 339938 581546 340174
rect 581782 339938 581866 340174
rect 582102 339938 586302 340174
rect 586538 339938 586622 340174
rect 586858 339938 592650 340174
rect -8726 339854 592650 339938
rect -8726 339618 -2934 339854
rect -2698 339618 -2614 339854
rect -2378 339618 9546 339854
rect 9782 339618 9866 339854
rect 10102 339618 189546 339854
rect 189782 339618 189866 339854
rect 190102 339618 225546 339854
rect 225782 339618 225866 339854
rect 226102 339618 261546 339854
rect 261782 339618 261866 339854
rect 262102 339618 297546 339854
rect 297782 339618 297866 339854
rect 298102 339618 333546 339854
rect 333782 339618 333866 339854
rect 334102 339618 369546 339854
rect 369782 339618 369866 339854
rect 370102 339618 405546 339854
rect 405782 339618 405866 339854
rect 406102 339618 572374 339854
rect 572610 339618 572694 339854
rect 572930 339618 581546 339854
rect 581782 339618 581866 339854
rect 582102 339618 586302 339854
rect 586538 339618 586622 339854
rect 586858 339618 592650 339854
rect -8726 339586 592650 339618
rect -8726 336454 592650 336486
rect -8726 336218 -1974 336454
rect -1738 336218 -1654 336454
rect -1418 336218 1826 336454
rect 2062 336218 2146 336454
rect 2382 336218 5826 336454
rect 6062 336218 6146 336454
rect 6382 336218 185826 336454
rect 186062 336218 186146 336454
rect 186382 336218 221826 336454
rect 222062 336218 222146 336454
rect 222382 336218 257826 336454
rect 258062 336218 258146 336454
rect 258382 336218 293826 336454
rect 294062 336218 294146 336454
rect 294382 336218 329826 336454
rect 330062 336218 330146 336454
rect 330382 336218 365826 336454
rect 366062 336218 366146 336454
rect 366382 336218 401826 336454
rect 402062 336218 402146 336454
rect 402382 336218 568510 336454
rect 568746 336218 568830 336454
rect 569066 336218 577826 336454
rect 578062 336218 578146 336454
rect 578382 336218 585342 336454
rect 585578 336218 585662 336454
rect 585898 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -1974 336134
rect -1738 335898 -1654 336134
rect -1418 335898 1826 336134
rect 2062 335898 2146 336134
rect 2382 335898 5826 336134
rect 6062 335898 6146 336134
rect 6382 335898 185826 336134
rect 186062 335898 186146 336134
rect 186382 335898 221826 336134
rect 222062 335898 222146 336134
rect 222382 335898 257826 336134
rect 258062 335898 258146 336134
rect 258382 335898 293826 336134
rect 294062 335898 294146 336134
rect 294382 335898 329826 336134
rect 330062 335898 330146 336134
rect 330382 335898 365826 336134
rect 366062 335898 366146 336134
rect 366382 335898 401826 336134
rect 402062 335898 402146 336134
rect 402382 335898 568510 336134
rect 568746 335898 568830 336134
rect 569066 335898 577826 336134
rect 578062 335898 578146 336134
rect 578382 335898 585342 336134
rect 585578 335898 585662 336134
rect 585898 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 304174 592650 304206
rect -8726 303938 -2934 304174
rect -2698 303938 -2614 304174
rect -2378 303938 9546 304174
rect 9782 303938 9866 304174
rect 10102 303938 189546 304174
rect 189782 303938 189866 304174
rect 190102 303938 225546 304174
rect 225782 303938 225866 304174
rect 226102 303938 261546 304174
rect 261782 303938 261866 304174
rect 262102 303938 297546 304174
rect 297782 303938 297866 304174
rect 298102 303938 333546 304174
rect 333782 303938 333866 304174
rect 334102 303938 369546 304174
rect 369782 303938 369866 304174
rect 370102 303938 405546 304174
rect 405782 303938 405866 304174
rect 406102 303938 572374 304174
rect 572610 303938 572694 304174
rect 572930 303938 581546 304174
rect 581782 303938 581866 304174
rect 582102 303938 586302 304174
rect 586538 303938 586622 304174
rect 586858 303938 592650 304174
rect -8726 303854 592650 303938
rect -8726 303618 -2934 303854
rect -2698 303618 -2614 303854
rect -2378 303618 9546 303854
rect 9782 303618 9866 303854
rect 10102 303618 189546 303854
rect 189782 303618 189866 303854
rect 190102 303618 225546 303854
rect 225782 303618 225866 303854
rect 226102 303618 261546 303854
rect 261782 303618 261866 303854
rect 262102 303618 297546 303854
rect 297782 303618 297866 303854
rect 298102 303618 333546 303854
rect 333782 303618 333866 303854
rect 334102 303618 369546 303854
rect 369782 303618 369866 303854
rect 370102 303618 405546 303854
rect 405782 303618 405866 303854
rect 406102 303618 572374 303854
rect 572610 303618 572694 303854
rect 572930 303618 581546 303854
rect 581782 303618 581866 303854
rect 582102 303618 586302 303854
rect 586538 303618 586622 303854
rect 586858 303618 592650 303854
rect -8726 303586 592650 303618
rect -8726 300454 592650 300486
rect -8726 300218 -1974 300454
rect -1738 300218 -1654 300454
rect -1418 300218 1826 300454
rect 2062 300218 2146 300454
rect 2382 300218 5826 300454
rect 6062 300218 6146 300454
rect 6382 300218 185826 300454
rect 186062 300218 186146 300454
rect 186382 300218 221826 300454
rect 222062 300218 222146 300454
rect 222382 300218 257826 300454
rect 258062 300218 258146 300454
rect 258382 300218 293826 300454
rect 294062 300218 294146 300454
rect 294382 300218 329826 300454
rect 330062 300218 330146 300454
rect 330382 300218 365826 300454
rect 366062 300218 366146 300454
rect 366382 300218 401826 300454
rect 402062 300218 402146 300454
rect 402382 300218 568510 300454
rect 568746 300218 568830 300454
rect 569066 300218 577826 300454
rect 578062 300218 578146 300454
rect 578382 300218 585342 300454
rect 585578 300218 585662 300454
rect 585898 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -1974 300134
rect -1738 299898 -1654 300134
rect -1418 299898 1826 300134
rect 2062 299898 2146 300134
rect 2382 299898 5826 300134
rect 6062 299898 6146 300134
rect 6382 299898 185826 300134
rect 186062 299898 186146 300134
rect 186382 299898 221826 300134
rect 222062 299898 222146 300134
rect 222382 299898 257826 300134
rect 258062 299898 258146 300134
rect 258382 299898 293826 300134
rect 294062 299898 294146 300134
rect 294382 299898 329826 300134
rect 330062 299898 330146 300134
rect 330382 299898 365826 300134
rect 366062 299898 366146 300134
rect 366382 299898 401826 300134
rect 402062 299898 402146 300134
rect 402382 299898 568510 300134
rect 568746 299898 568830 300134
rect 569066 299898 577826 300134
rect 578062 299898 578146 300134
rect 578382 299898 585342 300134
rect 585578 299898 585662 300134
rect 585898 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 268174 592650 268206
rect -8726 267938 -2934 268174
rect -2698 267938 -2614 268174
rect -2378 267938 9546 268174
rect 9782 267938 9866 268174
rect 10102 267938 189546 268174
rect 189782 267938 189866 268174
rect 190102 267938 225546 268174
rect 225782 267938 225866 268174
rect 226102 267938 261546 268174
rect 261782 267938 261866 268174
rect 262102 267938 297546 268174
rect 297782 267938 297866 268174
rect 298102 267938 333546 268174
rect 333782 267938 333866 268174
rect 334102 267938 369546 268174
rect 369782 267938 369866 268174
rect 370102 267938 405546 268174
rect 405782 267938 405866 268174
rect 406102 267938 572374 268174
rect 572610 267938 572694 268174
rect 572930 267938 581546 268174
rect 581782 267938 581866 268174
rect 582102 267938 586302 268174
rect 586538 267938 586622 268174
rect 586858 267938 592650 268174
rect -8726 267854 592650 267938
rect -8726 267618 -2934 267854
rect -2698 267618 -2614 267854
rect -2378 267618 9546 267854
rect 9782 267618 9866 267854
rect 10102 267618 189546 267854
rect 189782 267618 189866 267854
rect 190102 267618 225546 267854
rect 225782 267618 225866 267854
rect 226102 267618 261546 267854
rect 261782 267618 261866 267854
rect 262102 267618 297546 267854
rect 297782 267618 297866 267854
rect 298102 267618 333546 267854
rect 333782 267618 333866 267854
rect 334102 267618 369546 267854
rect 369782 267618 369866 267854
rect 370102 267618 405546 267854
rect 405782 267618 405866 267854
rect 406102 267618 572374 267854
rect 572610 267618 572694 267854
rect 572930 267618 581546 267854
rect 581782 267618 581866 267854
rect 582102 267618 586302 267854
rect 586538 267618 586622 267854
rect 586858 267618 592650 267854
rect -8726 267586 592650 267618
rect -8726 264454 592650 264486
rect -8726 264218 -1974 264454
rect -1738 264218 -1654 264454
rect -1418 264218 1826 264454
rect 2062 264218 2146 264454
rect 2382 264218 5826 264454
rect 6062 264218 6146 264454
rect 6382 264218 185826 264454
rect 186062 264218 186146 264454
rect 186382 264218 221826 264454
rect 222062 264218 222146 264454
rect 222382 264218 257826 264454
rect 258062 264218 258146 264454
rect 258382 264218 293826 264454
rect 294062 264218 294146 264454
rect 294382 264218 329826 264454
rect 330062 264218 330146 264454
rect 330382 264218 365826 264454
rect 366062 264218 366146 264454
rect 366382 264218 401826 264454
rect 402062 264218 402146 264454
rect 402382 264218 568510 264454
rect 568746 264218 568830 264454
rect 569066 264218 577826 264454
rect 578062 264218 578146 264454
rect 578382 264218 585342 264454
rect 585578 264218 585662 264454
rect 585898 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -1974 264134
rect -1738 263898 -1654 264134
rect -1418 263898 1826 264134
rect 2062 263898 2146 264134
rect 2382 263898 5826 264134
rect 6062 263898 6146 264134
rect 6382 263898 185826 264134
rect 186062 263898 186146 264134
rect 186382 263898 221826 264134
rect 222062 263898 222146 264134
rect 222382 263898 257826 264134
rect 258062 263898 258146 264134
rect 258382 263898 293826 264134
rect 294062 263898 294146 264134
rect 294382 263898 329826 264134
rect 330062 263898 330146 264134
rect 330382 263898 365826 264134
rect 366062 263898 366146 264134
rect 366382 263898 401826 264134
rect 402062 263898 402146 264134
rect 402382 263898 568510 264134
rect 568746 263898 568830 264134
rect 569066 263898 577826 264134
rect 578062 263898 578146 264134
rect 578382 263898 585342 264134
rect 585578 263898 585662 264134
rect 585898 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 232174 592650 232206
rect -8726 231938 -2934 232174
rect -2698 231938 -2614 232174
rect -2378 231938 9546 232174
rect 9782 231938 9866 232174
rect 10102 231938 45546 232174
rect 45782 231938 45866 232174
rect 46102 231938 81546 232174
rect 81782 231938 81866 232174
rect 82102 231938 117546 232174
rect 117782 231938 117866 232174
rect 118102 231938 153546 232174
rect 153782 231938 153866 232174
rect 154102 231938 189546 232174
rect 189782 231938 189866 232174
rect 190102 231938 225546 232174
rect 225782 231938 225866 232174
rect 226102 231938 261546 232174
rect 261782 231938 261866 232174
rect 262102 231938 297546 232174
rect 297782 231938 297866 232174
rect 298102 231938 333546 232174
rect 333782 231938 333866 232174
rect 334102 231938 369546 232174
rect 369782 231938 369866 232174
rect 370102 231938 405546 232174
rect 405782 231938 405866 232174
rect 406102 231938 441546 232174
rect 441782 231938 441866 232174
rect 442102 231938 477546 232174
rect 477782 231938 477866 232174
rect 478102 231938 513546 232174
rect 513782 231938 513866 232174
rect 514102 231938 549546 232174
rect 549782 231938 549866 232174
rect 550102 231938 581546 232174
rect 581782 231938 581866 232174
rect 582102 231938 586302 232174
rect 586538 231938 586622 232174
rect 586858 231938 592650 232174
rect -8726 231854 592650 231938
rect -8726 231618 -2934 231854
rect -2698 231618 -2614 231854
rect -2378 231618 9546 231854
rect 9782 231618 9866 231854
rect 10102 231618 45546 231854
rect 45782 231618 45866 231854
rect 46102 231618 81546 231854
rect 81782 231618 81866 231854
rect 82102 231618 117546 231854
rect 117782 231618 117866 231854
rect 118102 231618 153546 231854
rect 153782 231618 153866 231854
rect 154102 231618 189546 231854
rect 189782 231618 189866 231854
rect 190102 231618 225546 231854
rect 225782 231618 225866 231854
rect 226102 231618 261546 231854
rect 261782 231618 261866 231854
rect 262102 231618 297546 231854
rect 297782 231618 297866 231854
rect 298102 231618 333546 231854
rect 333782 231618 333866 231854
rect 334102 231618 369546 231854
rect 369782 231618 369866 231854
rect 370102 231618 405546 231854
rect 405782 231618 405866 231854
rect 406102 231618 441546 231854
rect 441782 231618 441866 231854
rect 442102 231618 477546 231854
rect 477782 231618 477866 231854
rect 478102 231618 513546 231854
rect 513782 231618 513866 231854
rect 514102 231618 549546 231854
rect 549782 231618 549866 231854
rect 550102 231618 581546 231854
rect 581782 231618 581866 231854
rect 582102 231618 586302 231854
rect 586538 231618 586622 231854
rect 586858 231618 592650 231854
rect -8726 231586 592650 231618
rect -8726 228454 592650 228486
rect -8726 228218 -1974 228454
rect -1738 228218 -1654 228454
rect -1418 228218 1826 228454
rect 2062 228218 2146 228454
rect 2382 228218 5826 228454
rect 6062 228218 6146 228454
rect 6382 228218 41826 228454
rect 42062 228218 42146 228454
rect 42382 228218 77826 228454
rect 78062 228218 78146 228454
rect 78382 228218 113826 228454
rect 114062 228218 114146 228454
rect 114382 228218 149826 228454
rect 150062 228218 150146 228454
rect 150382 228218 185826 228454
rect 186062 228218 186146 228454
rect 186382 228218 221826 228454
rect 222062 228218 222146 228454
rect 222382 228218 257826 228454
rect 258062 228218 258146 228454
rect 258382 228218 293826 228454
rect 294062 228218 294146 228454
rect 294382 228218 329826 228454
rect 330062 228218 330146 228454
rect 330382 228218 365826 228454
rect 366062 228218 366146 228454
rect 366382 228218 401826 228454
rect 402062 228218 402146 228454
rect 402382 228218 437826 228454
rect 438062 228218 438146 228454
rect 438382 228218 473826 228454
rect 474062 228218 474146 228454
rect 474382 228218 509826 228454
rect 510062 228218 510146 228454
rect 510382 228218 545826 228454
rect 546062 228218 546146 228454
rect 546382 228218 577826 228454
rect 578062 228218 578146 228454
rect 578382 228218 585342 228454
rect 585578 228218 585662 228454
rect 585898 228218 592650 228454
rect -8726 228139 592650 228218
rect -8726 228134 568510 228139
rect -8726 227898 -1974 228134
rect -1738 227898 -1654 228134
rect -1418 227898 1826 228134
rect 2062 227898 2146 228134
rect 2382 227898 5826 228134
rect 6062 227898 6146 228134
rect 6382 227898 41826 228134
rect 42062 227898 42146 228134
rect 42382 227898 77826 228134
rect 78062 227898 78146 228134
rect 78382 227898 113826 228134
rect 114062 227898 114146 228134
rect 114382 227898 149826 228134
rect 150062 227898 150146 228134
rect 150382 227898 185826 228134
rect 186062 227898 186146 228134
rect 186382 227898 221826 228134
rect 222062 227898 222146 228134
rect 222382 227898 257826 228134
rect 258062 227898 258146 228134
rect 258382 227898 293826 228134
rect 294062 227898 294146 228134
rect 294382 227898 329826 228134
rect 330062 227898 330146 228134
rect 330382 227898 365826 228134
rect 366062 227898 366146 228134
rect 366382 227898 401826 228134
rect 402062 227898 402146 228134
rect 402382 227898 437826 228134
rect 438062 227898 438146 228134
rect 438382 227898 473826 228134
rect 474062 227898 474146 228134
rect 474382 227898 509826 228134
rect 510062 227898 510146 228134
rect 510382 227898 545826 228134
rect 546062 227898 546146 228134
rect 546382 227903 568510 228134
rect 568746 227903 568830 228139
rect 569066 228134 592650 228139
rect 569066 227903 577826 228134
rect 546382 227898 577826 227903
rect 578062 227898 578146 228134
rect 578382 227898 585342 228134
rect 585578 227898 585662 228134
rect 585898 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 196174 592650 196206
rect -8726 195938 -2934 196174
rect -2698 195938 -2614 196174
rect -2378 195938 9546 196174
rect 9782 195938 9866 196174
rect 10102 195938 189546 196174
rect 189782 195938 189866 196174
rect 190102 195938 225546 196174
rect 225782 195938 225866 196174
rect 226102 195938 261546 196174
rect 261782 195938 261866 196174
rect 262102 195938 297546 196174
rect 297782 195938 297866 196174
rect 298102 195938 333546 196174
rect 333782 195938 333866 196174
rect 334102 195938 369546 196174
rect 369782 195938 369866 196174
rect 370102 195938 405546 196174
rect 405782 195938 405866 196174
rect 406102 195938 572374 196174
rect 572610 195938 572694 196174
rect 572930 195938 581546 196174
rect 581782 195938 581866 196174
rect 582102 195938 586302 196174
rect 586538 195938 586622 196174
rect 586858 195938 592650 196174
rect -8726 195854 592650 195938
rect -8726 195618 -2934 195854
rect -2698 195618 -2614 195854
rect -2378 195618 9546 195854
rect 9782 195618 9866 195854
rect 10102 195618 189546 195854
rect 189782 195618 189866 195854
rect 190102 195618 225546 195854
rect 225782 195618 225866 195854
rect 226102 195618 261546 195854
rect 261782 195618 261866 195854
rect 262102 195618 297546 195854
rect 297782 195618 297866 195854
rect 298102 195618 333546 195854
rect 333782 195618 333866 195854
rect 334102 195618 369546 195854
rect 369782 195618 369866 195854
rect 370102 195618 405546 195854
rect 405782 195618 405866 195854
rect 406102 195618 572374 195854
rect 572610 195618 572694 195854
rect 572930 195618 581546 195854
rect 581782 195618 581866 195854
rect 582102 195618 586302 195854
rect 586538 195618 586622 195854
rect 586858 195618 592650 195854
rect -8726 195586 592650 195618
rect -8726 192454 592650 192486
rect -8726 192218 -1974 192454
rect -1738 192218 -1654 192454
rect -1418 192218 1826 192454
rect 2062 192218 2146 192454
rect 2382 192218 5826 192454
rect 6062 192218 6146 192454
rect 6382 192218 185826 192454
rect 186062 192218 186146 192454
rect 186382 192218 221826 192454
rect 222062 192218 222146 192454
rect 222382 192218 257826 192454
rect 258062 192218 258146 192454
rect 258382 192218 293826 192454
rect 294062 192218 294146 192454
rect 294382 192218 329826 192454
rect 330062 192218 330146 192454
rect 330382 192218 365826 192454
rect 366062 192218 366146 192454
rect 366382 192218 401826 192454
rect 402062 192218 402146 192454
rect 402382 192218 568510 192454
rect 568746 192218 568830 192454
rect 569066 192218 577826 192454
rect 578062 192218 578146 192454
rect 578382 192218 585342 192454
rect 585578 192218 585662 192454
rect 585898 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -1974 192134
rect -1738 191898 -1654 192134
rect -1418 191898 1826 192134
rect 2062 191898 2146 192134
rect 2382 191898 5826 192134
rect 6062 191898 6146 192134
rect 6382 191898 185826 192134
rect 186062 191898 186146 192134
rect 186382 191898 221826 192134
rect 222062 191898 222146 192134
rect 222382 191898 257826 192134
rect 258062 191898 258146 192134
rect 258382 191898 293826 192134
rect 294062 191898 294146 192134
rect 294382 191898 329826 192134
rect 330062 191898 330146 192134
rect 330382 191898 365826 192134
rect 366062 191898 366146 192134
rect 366382 191898 401826 192134
rect 402062 191898 402146 192134
rect 402382 191898 568510 192134
rect 568746 191898 568830 192134
rect 569066 191898 577826 192134
rect 578062 191898 578146 192134
rect 578382 191898 585342 192134
rect 585578 191898 585662 192134
rect 585898 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 160174 592650 160206
rect -8726 159938 -2934 160174
rect -2698 159938 -2614 160174
rect -2378 159938 9546 160174
rect 9782 159938 9866 160174
rect 10102 159938 189546 160174
rect 189782 159938 189866 160174
rect 190102 159938 225546 160174
rect 225782 159938 225866 160174
rect 226102 159938 261546 160174
rect 261782 159938 261866 160174
rect 262102 159938 297546 160174
rect 297782 159938 297866 160174
rect 298102 159938 333546 160174
rect 333782 159938 333866 160174
rect 334102 159938 369546 160174
rect 369782 159938 369866 160174
rect 370102 159938 405546 160174
rect 405782 159938 405866 160174
rect 406102 159938 572374 160174
rect 572610 159938 572694 160174
rect 572930 159938 581546 160174
rect 581782 159938 581866 160174
rect 582102 159938 586302 160174
rect 586538 159938 586622 160174
rect 586858 159938 592650 160174
rect -8726 159854 592650 159938
rect -8726 159618 -2934 159854
rect -2698 159618 -2614 159854
rect -2378 159618 9546 159854
rect 9782 159618 9866 159854
rect 10102 159618 189546 159854
rect 189782 159618 189866 159854
rect 190102 159618 225546 159854
rect 225782 159618 225866 159854
rect 226102 159618 261546 159854
rect 261782 159618 261866 159854
rect 262102 159618 297546 159854
rect 297782 159618 297866 159854
rect 298102 159618 333546 159854
rect 333782 159618 333866 159854
rect 334102 159618 369546 159854
rect 369782 159618 369866 159854
rect 370102 159618 405546 159854
rect 405782 159618 405866 159854
rect 406102 159618 572374 159854
rect 572610 159618 572694 159854
rect 572930 159618 581546 159854
rect 581782 159618 581866 159854
rect 582102 159618 586302 159854
rect 586538 159618 586622 159854
rect 586858 159618 592650 159854
rect -8726 159586 592650 159618
rect -8726 156454 592650 156486
rect -8726 156218 -1974 156454
rect -1738 156218 -1654 156454
rect -1418 156218 1826 156454
rect 2062 156218 2146 156454
rect 2382 156218 5826 156454
rect 6062 156218 6146 156454
rect 6382 156218 185826 156454
rect 186062 156218 186146 156454
rect 186382 156218 221826 156454
rect 222062 156218 222146 156454
rect 222382 156218 257826 156454
rect 258062 156218 258146 156454
rect 258382 156218 293826 156454
rect 294062 156218 294146 156454
rect 294382 156218 329826 156454
rect 330062 156218 330146 156454
rect 330382 156218 365826 156454
rect 366062 156218 366146 156454
rect 366382 156218 401826 156454
rect 402062 156218 402146 156454
rect 402382 156218 568510 156454
rect 568746 156218 568830 156454
rect 569066 156218 577826 156454
rect 578062 156218 578146 156454
rect 578382 156218 585342 156454
rect 585578 156218 585662 156454
rect 585898 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -1974 156134
rect -1738 155898 -1654 156134
rect -1418 155898 1826 156134
rect 2062 155898 2146 156134
rect 2382 155898 5826 156134
rect 6062 155898 6146 156134
rect 6382 155898 185826 156134
rect 186062 155898 186146 156134
rect 186382 155898 221826 156134
rect 222062 155898 222146 156134
rect 222382 155898 257826 156134
rect 258062 155898 258146 156134
rect 258382 155898 293826 156134
rect 294062 155898 294146 156134
rect 294382 155898 329826 156134
rect 330062 155898 330146 156134
rect 330382 155898 365826 156134
rect 366062 155898 366146 156134
rect 366382 155898 401826 156134
rect 402062 155898 402146 156134
rect 402382 155898 568510 156134
rect 568746 155898 568830 156134
rect 569066 155898 577826 156134
rect 578062 155898 578146 156134
rect 578382 155898 585342 156134
rect 585578 155898 585662 156134
rect 585898 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 124174 592650 124206
rect -8726 123938 -2934 124174
rect -2698 123938 -2614 124174
rect -2378 123938 9546 124174
rect 9782 123938 9866 124174
rect 10102 123938 45546 124174
rect 45782 123938 45866 124174
rect 46102 123938 81546 124174
rect 81782 123938 81866 124174
rect 82102 123938 117546 124174
rect 117782 123938 117866 124174
rect 118102 123938 153546 124174
rect 153782 123938 153866 124174
rect 154102 123938 189546 124174
rect 189782 123938 189866 124174
rect 190102 123938 225546 124174
rect 225782 123938 225866 124174
rect 226102 123938 261546 124174
rect 261782 123938 261866 124174
rect 262102 123938 297546 124174
rect 297782 123938 297866 124174
rect 298102 123938 333546 124174
rect 333782 123938 333866 124174
rect 334102 123938 369546 124174
rect 369782 123938 369866 124174
rect 370102 123938 405546 124174
rect 405782 123938 405866 124174
rect 406102 123938 441546 124174
rect 441782 123938 441866 124174
rect 442102 123938 477546 124174
rect 477782 123938 477866 124174
rect 478102 123938 513546 124174
rect 513782 123938 513866 124174
rect 514102 123938 549546 124174
rect 549782 123938 549866 124174
rect 550102 123938 581546 124174
rect 581782 123938 581866 124174
rect 582102 123938 586302 124174
rect 586538 123938 586622 124174
rect 586858 123938 592650 124174
rect -8726 123854 592650 123938
rect -8726 123618 -2934 123854
rect -2698 123618 -2614 123854
rect -2378 123618 9546 123854
rect 9782 123618 9866 123854
rect 10102 123618 45546 123854
rect 45782 123618 45866 123854
rect 46102 123618 81546 123854
rect 81782 123618 81866 123854
rect 82102 123618 117546 123854
rect 117782 123618 117866 123854
rect 118102 123618 153546 123854
rect 153782 123618 153866 123854
rect 154102 123618 189546 123854
rect 189782 123618 189866 123854
rect 190102 123618 225546 123854
rect 225782 123618 225866 123854
rect 226102 123618 261546 123854
rect 261782 123618 261866 123854
rect 262102 123618 297546 123854
rect 297782 123618 297866 123854
rect 298102 123618 333546 123854
rect 333782 123618 333866 123854
rect 334102 123618 369546 123854
rect 369782 123618 369866 123854
rect 370102 123618 405546 123854
rect 405782 123618 405866 123854
rect 406102 123618 441546 123854
rect 441782 123618 441866 123854
rect 442102 123618 477546 123854
rect 477782 123618 477866 123854
rect 478102 123618 513546 123854
rect 513782 123618 513866 123854
rect 514102 123618 549546 123854
rect 549782 123618 549866 123854
rect 550102 123618 581546 123854
rect 581782 123618 581866 123854
rect 582102 123618 586302 123854
rect 586538 123618 586622 123854
rect 586858 123618 592650 123854
rect -8726 123586 592650 123618
rect -8726 120454 592650 120486
rect -8726 120218 -1974 120454
rect -1738 120218 -1654 120454
rect -1418 120218 1826 120454
rect 2062 120218 2146 120454
rect 2382 120218 5826 120454
rect 6062 120218 6146 120454
rect 6382 120218 41826 120454
rect 42062 120218 42146 120454
rect 42382 120218 77826 120454
rect 78062 120218 78146 120454
rect 78382 120218 113826 120454
rect 114062 120218 114146 120454
rect 114382 120218 149826 120454
rect 150062 120218 150146 120454
rect 150382 120218 185826 120454
rect 186062 120218 186146 120454
rect 186382 120218 221826 120454
rect 222062 120218 222146 120454
rect 222382 120218 257826 120454
rect 258062 120218 258146 120454
rect 258382 120218 293826 120454
rect 294062 120218 294146 120454
rect 294382 120218 329826 120454
rect 330062 120218 330146 120454
rect 330382 120218 365826 120454
rect 366062 120218 366146 120454
rect 366382 120218 401826 120454
rect 402062 120218 402146 120454
rect 402382 120218 437826 120454
rect 438062 120218 438146 120454
rect 438382 120218 473826 120454
rect 474062 120218 474146 120454
rect 474382 120218 509826 120454
rect 510062 120218 510146 120454
rect 510382 120218 545826 120454
rect 546062 120218 546146 120454
rect 546382 120218 577826 120454
rect 578062 120218 578146 120454
rect 578382 120218 585342 120454
rect 585578 120218 585662 120454
rect 585898 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -1974 120134
rect -1738 119898 -1654 120134
rect -1418 119898 1826 120134
rect 2062 119898 2146 120134
rect 2382 119898 5826 120134
rect 6062 119898 6146 120134
rect 6382 119898 41826 120134
rect 42062 119898 42146 120134
rect 42382 119898 77826 120134
rect 78062 119898 78146 120134
rect 78382 119898 113826 120134
rect 114062 119898 114146 120134
rect 114382 119898 149826 120134
rect 150062 119898 150146 120134
rect 150382 119898 185826 120134
rect 186062 119898 186146 120134
rect 186382 119898 221826 120134
rect 222062 119898 222146 120134
rect 222382 119898 257826 120134
rect 258062 119898 258146 120134
rect 258382 119898 293826 120134
rect 294062 119898 294146 120134
rect 294382 119898 329826 120134
rect 330062 119898 330146 120134
rect 330382 119898 365826 120134
rect 366062 119898 366146 120134
rect 366382 119898 401826 120134
rect 402062 119898 402146 120134
rect 402382 119898 437826 120134
rect 438062 119898 438146 120134
rect 438382 119898 473826 120134
rect 474062 119898 474146 120134
rect 474382 119898 509826 120134
rect 510062 119898 510146 120134
rect 510382 119898 545826 120134
rect 546062 119898 546146 120134
rect 546382 119898 577826 120134
rect 578062 119898 578146 120134
rect 578382 119898 585342 120134
rect 585578 119898 585662 120134
rect 585898 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 88174 592650 88206
rect -8726 87938 -2934 88174
rect -2698 87938 -2614 88174
rect -2378 87938 9546 88174
rect 9782 87938 9866 88174
rect 10102 87938 189546 88174
rect 189782 87938 189866 88174
rect 190102 87938 369546 88174
rect 369782 87938 369866 88174
rect 370102 87938 405546 88174
rect 405782 87938 405866 88174
rect 406102 87938 572374 88174
rect 572610 87938 572694 88174
rect 572930 87938 581546 88174
rect 581782 87938 581866 88174
rect 582102 87938 586302 88174
rect 586538 87938 586622 88174
rect 586858 87938 592650 88174
rect -8726 87854 592650 87938
rect -8726 87618 -2934 87854
rect -2698 87618 -2614 87854
rect -2378 87618 9546 87854
rect 9782 87618 9866 87854
rect 10102 87618 189546 87854
rect 189782 87618 189866 87854
rect 190102 87618 369546 87854
rect 369782 87618 369866 87854
rect 370102 87618 405546 87854
rect 405782 87618 405866 87854
rect 406102 87618 572374 87854
rect 572610 87618 572694 87854
rect 572930 87618 581546 87854
rect 581782 87618 581866 87854
rect 582102 87618 586302 87854
rect 586538 87618 586622 87854
rect 586858 87618 592650 87854
rect -8726 87586 592650 87618
rect -8726 84454 592650 84486
rect -8726 84218 -1974 84454
rect -1738 84218 -1654 84454
rect -1418 84218 1826 84454
rect 2062 84218 2146 84454
rect 2382 84218 5826 84454
rect 6062 84218 6146 84454
rect 6382 84218 185826 84454
rect 186062 84218 186146 84454
rect 186382 84218 365826 84454
rect 366062 84218 366146 84454
rect 366382 84218 401826 84454
rect 402062 84218 402146 84454
rect 402382 84218 568510 84454
rect 568746 84218 568830 84454
rect 569066 84218 577826 84454
rect 578062 84218 578146 84454
rect 578382 84218 585342 84454
rect 585578 84218 585662 84454
rect 585898 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -1974 84134
rect -1738 83898 -1654 84134
rect -1418 83898 1826 84134
rect 2062 83898 2146 84134
rect 2382 83898 5826 84134
rect 6062 83898 6146 84134
rect 6382 83898 185826 84134
rect 186062 83898 186146 84134
rect 186382 83898 365826 84134
rect 366062 83898 366146 84134
rect 366382 83898 401826 84134
rect 402062 83898 402146 84134
rect 402382 83898 568510 84134
rect 568746 83898 568830 84134
rect 569066 83898 577826 84134
rect 578062 83898 578146 84134
rect 578382 83898 585342 84134
rect 585578 83898 585662 84134
rect 585898 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 52174 592650 52206
rect -8726 51938 -2934 52174
rect -2698 51938 -2614 52174
rect -2378 51938 9546 52174
rect 9782 51938 9866 52174
rect 10102 51938 189546 52174
rect 189782 51938 189866 52174
rect 190102 51938 369546 52174
rect 369782 51938 369866 52174
rect 370102 51938 405546 52174
rect 405782 51938 405866 52174
rect 406102 51938 572374 52174
rect 572610 51938 572694 52174
rect 572930 51938 581546 52174
rect 581782 51938 581866 52174
rect 582102 51938 586302 52174
rect 586538 51938 586622 52174
rect 586858 51938 592650 52174
rect -8726 51854 592650 51938
rect -8726 51618 -2934 51854
rect -2698 51618 -2614 51854
rect -2378 51618 9546 51854
rect 9782 51618 9866 51854
rect 10102 51618 189546 51854
rect 189782 51618 189866 51854
rect 190102 51618 369546 51854
rect 369782 51618 369866 51854
rect 370102 51618 405546 51854
rect 405782 51618 405866 51854
rect 406102 51618 572374 51854
rect 572610 51618 572694 51854
rect 572930 51618 581546 51854
rect 581782 51618 581866 51854
rect 582102 51618 586302 51854
rect 586538 51618 586622 51854
rect 586858 51618 592650 51854
rect -8726 51586 592650 51618
rect -8726 48454 592650 48486
rect -8726 48218 -1974 48454
rect -1738 48218 -1654 48454
rect -1418 48218 1826 48454
rect 2062 48218 2146 48454
rect 2382 48218 5826 48454
rect 6062 48218 6146 48454
rect 6382 48218 185826 48454
rect 186062 48218 186146 48454
rect 186382 48218 365826 48454
rect 366062 48218 366146 48454
rect 366382 48218 401826 48454
rect 402062 48218 402146 48454
rect 402382 48218 568510 48454
rect 568746 48218 568830 48454
rect 569066 48218 577826 48454
rect 578062 48218 578146 48454
rect 578382 48218 585342 48454
rect 585578 48218 585662 48454
rect 585898 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -1974 48134
rect -1738 47898 -1654 48134
rect -1418 47898 1826 48134
rect 2062 47898 2146 48134
rect 2382 47898 5826 48134
rect 6062 47898 6146 48134
rect 6382 47898 185826 48134
rect 186062 47898 186146 48134
rect 186382 47898 365826 48134
rect 366062 47898 366146 48134
rect 366382 47898 401826 48134
rect 402062 47898 402146 48134
rect 402382 47898 568510 48134
rect 568746 47898 568830 48134
rect 569066 47898 577826 48134
rect 578062 47898 578146 48134
rect 578382 47898 585342 48134
rect 585578 47898 585662 48134
rect 585898 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 16174 592650 16206
rect -8726 15938 -2934 16174
rect -2698 15938 -2614 16174
rect -2378 15938 9546 16174
rect 9782 15938 9866 16174
rect 10102 15938 45546 16174
rect 45782 15938 45866 16174
rect 46102 15938 81546 16174
rect 81782 15938 81866 16174
rect 82102 15938 117546 16174
rect 117782 15938 117866 16174
rect 118102 15938 153546 16174
rect 153782 15938 153866 16174
rect 154102 15938 189546 16174
rect 189782 15938 189866 16174
rect 190102 15938 225546 16174
rect 225782 15938 225866 16174
rect 226102 15938 261546 16174
rect 261782 15938 261866 16174
rect 262102 15938 297546 16174
rect 297782 15938 297866 16174
rect 298102 15938 333546 16174
rect 333782 15938 333866 16174
rect 334102 15938 369546 16174
rect 369782 15938 369866 16174
rect 370102 15938 405546 16174
rect 405782 15938 405866 16174
rect 406102 15938 441546 16174
rect 441782 15938 441866 16174
rect 442102 15938 477546 16174
rect 477782 15938 477866 16174
rect 478102 15938 513546 16174
rect 513782 15938 513866 16174
rect 514102 15938 549546 16174
rect 549782 15938 549866 16174
rect 550102 15938 581546 16174
rect 581782 15938 581866 16174
rect 582102 15938 586302 16174
rect 586538 15938 586622 16174
rect 586858 15938 592650 16174
rect -8726 15854 592650 15938
rect -8726 15618 -2934 15854
rect -2698 15618 -2614 15854
rect -2378 15618 9546 15854
rect 9782 15618 9866 15854
rect 10102 15618 45546 15854
rect 45782 15618 45866 15854
rect 46102 15618 81546 15854
rect 81782 15618 81866 15854
rect 82102 15618 117546 15854
rect 117782 15618 117866 15854
rect 118102 15618 153546 15854
rect 153782 15618 153866 15854
rect 154102 15618 189546 15854
rect 189782 15618 189866 15854
rect 190102 15618 225546 15854
rect 225782 15618 225866 15854
rect 226102 15618 261546 15854
rect 261782 15618 261866 15854
rect 262102 15618 297546 15854
rect 297782 15618 297866 15854
rect 298102 15618 333546 15854
rect 333782 15618 333866 15854
rect 334102 15618 369546 15854
rect 369782 15618 369866 15854
rect 370102 15618 405546 15854
rect 405782 15618 405866 15854
rect 406102 15618 441546 15854
rect 441782 15618 441866 15854
rect 442102 15618 477546 15854
rect 477782 15618 477866 15854
rect 478102 15618 513546 15854
rect 513782 15618 513866 15854
rect 514102 15618 549546 15854
rect 549782 15618 549866 15854
rect 550102 15618 581546 15854
rect 581782 15618 581866 15854
rect 582102 15618 586302 15854
rect 586538 15618 586622 15854
rect 586858 15618 592650 15854
rect -8726 15586 592650 15618
rect -8726 12454 592650 12486
rect -8726 12218 -1974 12454
rect -1738 12218 -1654 12454
rect -1418 12218 1826 12454
rect 2062 12218 2146 12454
rect 2382 12218 5826 12454
rect 6062 12218 6146 12454
rect 6382 12218 41826 12454
rect 42062 12218 42146 12454
rect 42382 12218 77826 12454
rect 78062 12218 78146 12454
rect 78382 12218 113826 12454
rect 114062 12218 114146 12454
rect 114382 12218 149826 12454
rect 150062 12218 150146 12454
rect 150382 12218 185826 12454
rect 186062 12218 186146 12454
rect 186382 12218 221826 12454
rect 222062 12218 222146 12454
rect 222382 12218 257826 12454
rect 258062 12218 258146 12454
rect 258382 12218 293826 12454
rect 294062 12218 294146 12454
rect 294382 12218 329826 12454
rect 330062 12218 330146 12454
rect 330382 12218 365826 12454
rect 366062 12218 366146 12454
rect 366382 12218 401826 12454
rect 402062 12218 402146 12454
rect 402382 12218 437826 12454
rect 438062 12218 438146 12454
rect 438382 12218 473826 12454
rect 474062 12218 474146 12454
rect 474382 12218 509826 12454
rect 510062 12218 510146 12454
rect 510382 12218 545826 12454
rect 546062 12218 546146 12454
rect 546382 12218 577826 12454
rect 578062 12218 578146 12454
rect 578382 12218 585342 12454
rect 585578 12218 585662 12454
rect 585898 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -1974 12134
rect -1738 11898 -1654 12134
rect -1418 11898 1826 12134
rect 2062 11898 2146 12134
rect 2382 11898 5826 12134
rect 6062 11898 6146 12134
rect 6382 11898 41826 12134
rect 42062 11898 42146 12134
rect 42382 11898 77826 12134
rect 78062 11898 78146 12134
rect 78382 11898 113826 12134
rect 114062 11898 114146 12134
rect 114382 11898 149826 12134
rect 150062 11898 150146 12134
rect 150382 11898 185826 12134
rect 186062 11898 186146 12134
rect 186382 11898 221826 12134
rect 222062 11898 222146 12134
rect 222382 11898 257826 12134
rect 258062 11898 258146 12134
rect 258382 11898 293826 12134
rect 294062 11898 294146 12134
rect 294382 11898 329826 12134
rect 330062 11898 330146 12134
rect 330382 11898 365826 12134
rect 366062 11898 366146 12134
rect 366382 11898 401826 12134
rect 402062 11898 402146 12134
rect 402382 11898 437826 12134
rect 438062 11898 438146 12134
rect 438382 11898 473826 12134
rect 474062 11898 474146 12134
rect 474382 11898 509826 12134
rect 510062 11898 510146 12134
rect 510382 11898 545826 12134
rect 546062 11898 546146 12134
rect 546382 11898 577826 12134
rect 578062 11898 578146 12134
rect 578382 11898 585342 12134
rect 585578 11898 585662 12134
rect 585898 11898 592650 12134
rect -8726 11866 592650 11898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use j202_soc_core_wrapper  j202_soc_core_wrapper
timestamp 0
transform 1 0 4000 0 1 4000
box -960 -960 576960 696960
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 699728 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 699728 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 699728 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 699728 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 699728 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 699728 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 699728 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 699728 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 699728 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 699728 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 699728 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 699728 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 699728 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 699728 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 699728 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 699728 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 15586 592650 16206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 51586 592650 52206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 87586 592650 88206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 123586 592650 124206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 159586 592650 160206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 195586 592650 196206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 231586 592650 232206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 267586 592650 268206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 303586 592650 304206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 339586 592650 340206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 375586 592650 376206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 411586 592650 412206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 447586 592650 448206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 483586 592650 484206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 519586 592650 520206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 555586 592650 556206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 591586 592650 592206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 627586 592650 628206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 663586 592650 664206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 699586 592650 700206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 578264 696336 578264 696336 0 vccd1
rlabel metal4 587540 351968 587540 351968 0 vccd2
rlabel metal4 589460 351968 589460 351968 0 vdda1
rlabel metal4 591380 351968 591380 351968 0 vdda2
rlabel metal4 590420 351968 590420 351968 0 vssa1
rlabel metal4 592340 351968 592340 351968 0 vssa2
rlabel via4 572812 664056 572812 664056 0 vssd1
rlabel metal4 588500 351968 588500 351968 0 vssd2
rlabel metal3 580796 286265 580796 286265 0 analog_io[0]
rlabel metal2 443401 700876 443401 700876 0 analog_io[10]
rlabel metal2 379401 700876 379401 700876 0 analog_io[11]
rlabel metal2 315981 700876 315981 700876 0 analog_io[12]
rlabel metal2 251981 700876 251981 700876 0 analog_io[13]
rlabel metal1 187496 703018 187496 703018 0 analog_io[14]
rlabel metal2 121670 702280 121670 702280 0 analog_io[15]
rlabel metal1 58788 700978 58788 700978 0 analog_io[16]
rlabel metal3 1188 697340 1188 697340 0 analog_io[17]
rlabel metal3 2262 639676 2262 639676 0 analog_io[18]
rlabel metal3 1556 593028 1556 593028 0 analog_io[19]
rlabel metal3 580796 338693 580796 338693 0 analog_io[1]
rlabel metal3 866 540804 866 540804 0 analog_io[20]
rlabel metal3 958 488716 958 488716 0 analog_io[21]
rlabel metal3 1556 436628 1556 436628 0 analog_io[22]
rlabel metal3 1763 384404 1763 384404 0 analog_io[23]
rlabel metal3 1763 332316 1763 332316 0 analog_io[24]
rlabel metal3 1556 280092 1556 280092 0 analog_io[25]
rlabel metal3 2998 230588 2998 230588 0 analog_io[26]
rlabel metal3 1556 175916 1556 175916 0 analog_io[27]
rlabel metal3 544 123692 544 123692 0 analog_io[28]
rlabel metal3 580796 391491 580796 391491 0 analog_io[2]
rlabel metal3 580796 443783 580796 443783 0 analog_io[3]
rlabel metal3 581248 495652 581248 495652 0 analog_io[4]
rlabel metal3 581248 547740 581248 547740 0 analog_io[5]
rlabel metal3 581248 600100 581248 600100 0 analog_io[6]
rlabel metal3 582966 657356 582966 657356 0 analog_io[7]
rlabel metal1 573206 703018 573206 703018 0 analog_io[8]
rlabel metal2 506874 701682 506874 701682 0 analog_io[9]
rlabel metal3 581724 6596 581724 6596 0 io_in[0]
rlabel metal3 581248 456484 581248 456484 0 io_in[10]
rlabel metal3 581616 508708 581616 508708 0 io_in[11]
rlabel metal3 581616 560932 581616 560932 0 io_in[12]
rlabel metal3 582598 617508 582598 617508 0 io_in[13]
rlabel metal3 581616 665380 581616 665380 0 io_in[14]
rlabel metal2 559682 703028 559682 703028 0 io_in[15]
rlabel metal1 492890 702746 492890 702746 0 io_in[16]
rlabel metal2 427439 700876 427439 700876 0 io_in[17]
rlabel metal2 365010 702280 365010 702280 0 io_in[18]
rlabel metal2 300065 700876 300065 700876 0 io_in[19]
rlabel metal3 580796 51325 580796 51325 0 io_in[1]
rlabel metal1 235704 703018 235704 703018 0 io_in[20]
rlabel metal2 172454 700927 172454 700927 0 io_in[21]
rlabel metal1 107042 700978 107042 700978 0 io_in[22]
rlabel metal1 42734 700978 42734 700978 0 io_in[23]
rlabel metal3 2124 678028 2124 678028 0 io_in[24]
rlabel metal3 820 632060 820 632060 0 io_in[25]
rlabel metal3 1556 579972 1556 579972 0 io_in[26]
rlabel metal3 912 527884 912 527884 0 io_in[27]
rlabel metal3 1556 475660 1556 475660 0 io_in[28]
rlabel metal3 1556 423572 1556 423572 0 io_in[29]
rlabel metal3 580796 90493 580796 90493 0 io_in[2]
rlabel metal3 1763 371348 1763 371348 0 io_in[30]
rlabel metal3 1763 319260 1763 319260 0 io_in[31]
rlabel metal3 2262 268804 2262 268804 0 io_in[32]
rlabel metal3 1556 214948 1556 214948 0 io_in[33]
rlabel metal3 1556 162860 1556 162860 0 io_in[34]
rlabel metal3 2262 115396 2262 115396 0 io_in[35]
rlabel metal3 2400 77044 2400 77044 0 io_in[36]
rlabel metal3 2998 38692 2998 38692 0 io_in[37]
rlabel metal3 580796 130167 580796 130167 0 io_in[3]
rlabel metal3 580796 168829 580796 168829 0 io_in[4]
rlabel metal3 581616 208284 581616 208284 0 io_in[5]
rlabel metal3 580796 247233 580796 247233 0 io_in[6]
rlabel metal3 580796 299457 580796 299457 0 io_in[7]
rlabel metal3 582176 351900 582176 351900 0 io_in[8]
rlabel metal3 580796 404615 580796 404615 0 io_in[9]
rlabel metal3 580865 38012 580865 38012 0 io_oeb[0]
rlabel metal3 581616 482596 581616 482596 0 io_oeb[10]
rlabel metal3 581616 534820 581616 534820 0 io_oeb[11]
rlabel metal3 581248 587044 581248 587044 0 io_oeb[12]
rlabel metal3 581248 639268 581248 639268 0 io_oeb[13]
rlabel metal3 582598 697204 582598 697204 0 io_oeb[14]
rlabel metal1 524952 703018 524952 703018 0 io_oeb[15]
rlabel metal2 462346 703028 462346 703028 0 io_oeb[16]
rlabel metal2 395607 700876 395607 700876 0 io_oeb[17]
rlabel metal2 331989 700876 331989 700876 0 io_oeb[18]
rlabel metal2 267851 700876 267851 700876 0 io_oeb[19]
rlabel metal3 579991 77316 579991 77316 0 io_oeb[1]
rlabel metal1 203550 700978 203550 700978 0 io_oeb[20]
rlabel metal1 139150 700978 139150 700978 0 io_oeb[21]
rlabel metal2 76774 700927 76774 700927 0 io_oeb[22]
rlabel metal1 10626 700978 10626 700978 0 io_oeb[23]
rlabel via2 69 657628 69 657628 0 io_oeb[24]
rlabel metal3 2032 601324 2032 601324 0 io_oeb[25]
rlabel metal3 1556 553860 1556 553860 0 io_oeb[26]
rlabel metal3 958 501772 958 501772 0 io_oeb[27]
rlabel metal3 1556 449548 1556 449548 0 io_oeb[28]
rlabel metal3 1763 397460 1763 397460 0 io_oeb[29]
rlabel metal3 579991 116348 579991 116348 0 io_oeb[2]
rlabel metal3 935 345372 935 345372 0 io_oeb[30]
rlabel metal3 820 293148 820 293148 0 io_oeb[31]
rlabel metal3 1556 241060 1556 241060 0 io_oeb[32]
rlabel metal3 2262 192100 2262 192100 0 io_oeb[33]
rlabel metal3 452 136748 452 136748 0 io_oeb[34]
rlabel metal3 958 84660 958 84660 0 io_oeb[35]
rlabel metal3 1556 45492 1556 45492 0 io_oeb[36]
rlabel metal3 1556 6460 1556 6460 0 io_oeb[37]
rlabel metal3 580796 156279 580796 156279 0 io_oeb[3]
rlabel metal3 580796 194941 580796 194941 0 io_oeb[4]
rlabel metal3 581616 234396 581616 234396 0 io_oeb[5]
rlabel metal3 580796 273209 580796 273209 0 io_oeb[6]
rlabel metal3 582161 325244 582161 325244 0 io_oeb[7]
rlabel metal3 580796 378299 580796 378299 0 io_oeb[8]
rlabel metal3 580796 430727 580796 430727 0 io_oeb[9]
rlabel metal3 580796 25213 580796 25213 0 io_out[0]
rlabel metal3 581248 469540 581248 469540 0 io_out[10]
rlabel metal3 581616 521764 581616 521764 0 io_out[11]
rlabel metal3 582598 577660 582598 577660 0 io_out[12]
rlabel metal3 581616 626212 581616 626212 0 io_out[13]
rlabel metal3 581616 678436 581616 678436 0 io_out[14]
rlabel metal1 541098 702746 541098 702746 0 io_out[15]
rlabel metal2 475233 700876 475233 700876 0 io_out[16]
rlabel metal2 411569 700876 411569 700876 0 io_out[17]
rlabel metal2 347905 700876 347905 700876 0 io_out[18]
rlabel metal2 283905 700876 283905 700876 0 io_out[19]
rlabel metal3 580796 64381 580796 64381 0 io_out[1]
rlabel metal2 219006 703028 219006 703028 0 io_out[20]
rlabel metal1 155204 700978 155204 700978 0 io_out[21]
rlabel metal1 90896 700978 90896 700978 0 io_out[22]
rlabel metal2 24334 703028 24334 703028 0 io_out[23]
rlabel metal3 682 671228 682 671228 0 io_out[24]
rlabel via2 69 618596 69 618596 0 io_out[25]
rlabel metal3 1556 566916 1556 566916 0 io_out[26]
rlabel metal3 1556 514828 1556 514828 0 io_out[27]
rlabel metal3 958 462604 958 462604 0 io_out[28]
rlabel metal3 1763 410516 1763 410516 0 io_out[29]
rlabel metal3 582230 99484 582230 99484 0 io_out[2]
rlabel metal3 1748 358428 1748 358428 0 io_out[30]
rlabel metal3 1763 306204 1763 306204 0 io_out[31]
rlabel metal3 820 254116 820 254116 0 io_out[32]
rlabel metal3 1556 201892 1556 201892 0 io_out[33]
rlabel metal3 2262 153748 2262 153748 0 io_out[34]
rlabel metal3 958 97580 958 97580 0 io_out[35]
rlabel metal3 912 58548 912 58548 0 io_out[36]
rlabel metal3 912 19380 912 19380 0 io_out[37]
rlabel metal3 582230 139332 582230 139332 0 io_out[3]
rlabel metal3 582230 179180 582230 179180 0 io_out[4]
rlabel metal3 582230 219028 582230 219028 0 io_out[5]
rlabel metal3 581616 260508 581616 260508 0 io_out[6]
rlabel metal3 580796 312377 580796 312377 0 io_out[7]
rlabel metal3 582176 365092 582176 365092 0 io_out[8]
rlabel metal3 580796 417535 580796 417535 0 io_out[9]
rlabel via1 136666 3757 136666 3757 0 la_data_in[0]
rlabel metal2 468142 1846 468142 1846 0 la_data_in[100]
rlabel via1 484242 187 484242 187 0 la_data_in[101]
rlabel metal2 487455 340 487455 340 0 la_data_in[102]
rlabel metal2 478354 1649 478354 1649 0 la_data_in[103]
rlabel metal2 481574 1853 481574 1853 0 la_data_in[104]
rlabel metal2 484702 1540 484702 1540 0 la_data_in[105]
rlabel metal2 488014 1880 488014 1880 0 la_data_in[106]
rlabel metal2 505402 500 505402 500 0 la_data_in[107]
rlabel metal2 508898 636 508898 636 0 la_data_in[108]
rlabel metal2 500434 884 500434 884 0 la_data_in[109]
rlabel metal2 161322 1792 161322 1792 0 la_data_in[10]
rlabel metal2 501262 1778 501262 1778 0 la_data_in[110]
rlabel metal1 506874 680 506874 680 0 la_data_in[111]
rlabel metal2 507886 527 507886 527 0 la_data_in[112]
rlabel metal2 526463 340 526463 340 0 la_data_in[113]
rlabel metal2 514510 1710 514510 1710 0 la_data_in[114]
rlabel metal2 517822 2118 517822 2118 0 la_data_in[115]
rlabel metal2 521134 1676 521134 1676 0 la_data_in[116]
rlabel metal2 524354 1880 524354 1880 0 la_data_in[117]
rlabel metal2 527758 1914 527758 1914 0 la_data_in[118]
rlabel metal2 531070 1574 531070 1574 0 la_data_in[119]
rlabel via1 173006 3315 173006 3315 0 la_data_in[11]
rlabel metal2 534382 2016 534382 2016 0 la_data_in[120]
rlabel metal2 537694 1608 537694 1608 0 la_data_in[121]
rlabel metal2 540914 1880 540914 1880 0 la_data_in[122]
rlabel metal2 544594 1785 544594 1785 0 la_data_in[123]
rlabel metal2 547630 1914 547630 1914 0 la_data_in[124]
rlabel metal2 550942 1948 550942 1948 0 la_data_in[125]
rlabel metal2 554254 1642 554254 1642 0 la_data_in[126]
rlabel metal2 557198 1683 557198 1683 0 la_data_in[127]
rlabel metal2 176594 2968 176594 2968 0 la_data_in[12]
rlabel metal2 171994 1690 171994 1690 0 la_data_in[13]
rlabel metal2 175490 1588 175490 1588 0 la_data_in[14]
rlabel metal2 179078 1758 179078 1758 0 la_data_in[15]
rlabel metal2 182574 1792 182574 1792 0 la_data_in[16]
rlabel metal2 193154 3002 193154 3002 0 la_data_in[17]
rlabel via1 196190 3315 196190 3315 0 la_data_in[18]
rlabel metal2 193246 1554 193246 1554 0 la_data_in[19]
rlabel via1 139886 3485 139886 3485 0 la_data_in[1]
rlabel metal2 196834 1724 196834 1724 0 la_data_in[20]
rlabel metal2 200330 1792 200330 1792 0 la_data_in[21]
rlabel metal2 203918 1656 203918 1656 0 la_data_in[22]
rlabel metal2 213026 2186 213026 2186 0 la_data_in[23]
rlabel metal2 211002 1588 211002 1588 0 la_data_in[24]
rlabel metal2 214498 1758 214498 1758 0 la_data_in[25]
rlabel metal2 218086 1690 218086 1690 0 la_data_in[26]
rlabel metal2 221582 1724 221582 1724 0 la_data_in[27]
rlabel via1 229310 3043 229310 3043 0 la_data_in[28]
rlabel metal2 232898 2934 232898 2934 0 la_data_in[29]
rlabel metal2 132986 1962 132986 1962 0 la_data_in[2]
rlabel metal2 232254 1622 232254 1622 0 la_data_in[30]
rlabel metal2 235842 1588 235842 1588 0 la_data_in[31]
rlabel metal2 239338 1656 239338 1656 0 la_data_in[32]
rlabel metal2 242926 1656 242926 1656 0 la_data_in[33]
rlabel metal2 249458 3002 249458 3002 0 la_data_in[34]
rlabel metal2 250010 1622 250010 1622 0 la_data_in[35]
rlabel metal2 253506 1656 253506 1656 0 la_data_in[36]
rlabel metal2 257094 840 257094 840 0 la_data_in[37]
rlabel metal2 260682 1588 260682 1588 0 la_data_in[38]
rlabel metal2 264178 806 264178 806 0 la_data_in[39]
rlabel metal2 136482 1588 136482 1588 0 la_data_in[3]
rlabel metal2 267766 840 267766 840 0 la_data_in[40]
rlabel metal2 271262 840 271262 840 0 la_data_in[41]
rlabel metal2 275087 340 275087 340 0 la_data_in[42]
rlabel metal2 278583 340 278583 340 0 la_data_in[43]
rlabel metal2 281934 1707 281934 1707 0 la_data_in[44]
rlabel metal2 285430 1707 285430 1707 0 la_data_in[45]
rlabel metal2 289018 1707 289018 1707 0 la_data_in[46]
rlabel metal2 292606 1700 292606 1700 0 la_data_in[47]
rlabel metal2 296102 1707 296102 1707 0 la_data_in[48]
rlabel metal2 299690 1707 299690 1707 0 la_data_in[49]
rlabel metal2 140070 1690 140070 1690 0 la_data_in[4]
rlabel metal2 303186 1707 303186 1707 0 la_data_in[50]
rlabel metal2 306314 1700 306314 1700 0 la_data_in[51]
rlabel metal2 310270 1588 310270 1588 0 la_data_in[52]
rlabel metal2 313858 1622 313858 1622 0 la_data_in[53]
rlabel metal2 315790 2934 315790 2934 0 la_data_in[54]
rlabel metal2 320942 1622 320942 1622 0 la_data_in[55]
rlabel metal2 324438 1588 324438 1588 0 la_data_in[56]
rlabel metal2 328026 1656 328026 1656 0 la_data_in[57]
rlabel metal2 331614 1656 331614 1656 0 la_data_in[58]
rlabel metal2 335110 1656 335110 1656 0 la_data_in[59]
rlabel via1 153226 3315 153226 3315 0 la_data_in[5]
rlabel metal2 338698 1588 338698 1588 0 la_data_in[60]
rlabel metal2 342194 755 342194 755 0 la_data_in[61]
rlabel metal2 345782 840 345782 840 0 la_data_in[62]
rlabel metal2 349278 670 349278 670 0 la_data_in[63]
rlabel metal2 352866 840 352866 840 0 la_data_in[64]
rlabel metal2 352222 2084 352222 2084 0 la_data_in[65]
rlabel metal2 359950 704 359950 704 0 la_data_in[66]
rlabel metal2 363538 636 363538 636 0 la_data_in[67]
rlabel metal2 367034 670 367034 670 0 la_data_in[68]
rlabel metal2 370431 340 370431 340 0 la_data_in[69]
rlabel via1 156446 3179 156446 3179 0 la_data_in[6]
rlabel metal2 373934 765 373934 765 0 la_data_in[70]
rlabel metal2 372370 2941 372370 2941 0 la_data_in[71]
rlabel metal2 381202 738 381202 738 0 la_data_in[72]
rlabel metal2 384599 340 384599 340 0 la_data_in[73]
rlabel via1 387918 323 387918 323 0 la_data_in[74]
rlabel metal2 391874 738 391874 738 0 la_data_in[75]
rlabel metal2 388654 1812 388654 1812 0 la_data_in[76]
rlabel metal2 391690 1615 391690 1615 0 la_data_in[77]
rlabel metal2 402546 772 402546 772 0 la_data_in[78]
rlabel via1 406226 85 406226 85 0 la_data_in[79]
rlabel via1 159758 3213 159758 3213 0 la_data_in[7]
rlabel metal2 409439 340 409439 340 0 la_data_in[80]
rlabel metal2 405214 1608 405214 1608 0 la_data_in[81]
rlabel metal2 408434 1880 408434 1880 0 la_data_in[82]
rlabel metal2 412114 1581 412114 1581 0 la_data_in[83]
rlabel via1 423614 221 423614 221 0 la_data_in[84]
rlabel metal2 427294 500 427294 500 0 la_data_in[85]
rlabel via1 431066 51 431066 51 0 la_data_in[86]
rlabel metal2 424810 1751 424810 1751 0 la_data_in[87]
rlabel metal2 428674 1717 428674 1717 0 la_data_in[88]
rlabel metal2 431710 1608 431710 1608 0 la_data_in[89]
rlabel metal2 154238 1826 154238 1826 0 la_data_in[8]
rlabel metal2 445149 340 445149 340 0 la_data_in[90]
rlabel metal2 448447 340 448447 340 0 la_data_in[91]
rlabel metal2 441554 1948 441554 1948 0 la_data_in[92]
rlabel metal2 444958 1982 444958 1982 0 la_data_in[93]
rlabel metal2 448270 2016 448270 2016 0 la_data_in[94]
rlabel metal2 462615 340 462615 340 0 la_data_in[95]
rlabel metal2 466111 340 466111 340 0 la_data_in[96]
rlabel metal2 469989 340 469989 340 0 la_data_in[97]
rlabel metal2 461794 1785 461794 1785 0 la_data_in[98]
rlabel metal2 464830 1812 464830 1812 0 la_data_in[99]
rlabel metal2 157826 1656 157826 1656 0 la_data_in[9]
rlabel via1 137678 3349 137678 3349 0 la_data_out[0]
rlabel metal2 469154 2118 469154 2118 0 la_data_out[100]
rlabel metal2 485063 340 485063 340 0 la_data_out[101]
rlabel metal2 488842 840 488842 840 0 la_data_out[102]
rlabel metal2 479550 1683 479550 1683 0 la_data_out[103]
rlabel metal2 482494 2016 482494 2016 0 la_data_out[104]
rlabel metal2 485714 2084 485714 2084 0 la_data_out[105]
rlabel metal2 489118 2050 489118 2050 0 la_data_out[106]
rlabel metal2 506506 602 506506 602 0 la_data_out[107]
rlabel metal2 495742 2016 495742 2016 0 la_data_out[108]
rlabel metal2 499054 2152 499054 2152 0 la_data_out[109]
rlabel metal2 162518 1758 162518 1758 0 la_data_out[10]
rlabel metal1 506966 748 506966 748 0 la_data_out[110]
rlabel metal2 505678 1676 505678 1676 0 la_data_out[111]
rlabel metal2 508990 1948 508990 1948 0 la_data_out[112]
rlabel metal2 527850 806 527850 806 0 la_data_out[113]
rlabel metal2 515522 1642 515522 1642 0 la_data_out[114]
rlabel metal2 518834 1778 518834 1778 0 la_data_out[115]
rlabel metal2 522238 1812 522238 1812 0 la_data_out[116]
rlabel metal2 525550 1846 525550 1846 0 la_data_out[117]
rlabel metal2 545613 340 545613 340 0 la_data_out[118]
rlabel metal2 532174 1982 532174 1982 0 la_data_out[119]
rlabel metal2 174386 3002 174386 3002 0 la_data_out[11]
rlabel metal2 535394 1642 535394 1642 0 la_data_out[120]
rlabel metal2 538798 1676 538798 1676 0 la_data_out[121]
rlabel metal2 542110 1812 542110 1812 0 la_data_out[122]
rlabel metal2 545422 1846 545422 1846 0 la_data_out[123]
rlabel metal2 566957 340 566957 340 0 la_data_out[124]
rlabel metal2 551954 1574 551954 1574 0 la_data_out[125]
rlabel metal2 555358 1710 555358 1710 0 la_data_out[126]
rlabel metal2 558854 1615 558854 1615 0 la_data_out[127]
rlabel via1 177422 3451 177422 3451 0 la_data_out[12]
rlabel metal2 173190 1792 173190 1792 0 la_data_out[13]
rlabel metal2 176686 959 176686 959 0 la_data_out[14]
rlabel metal2 180274 1860 180274 1860 0 la_data_out[15]
rlabel via1 190670 3451 190670 3451 0 la_data_out[16]
rlabel via1 193982 3043 193982 3043 0 la_data_out[17]
rlabel metal2 190854 1792 190854 1792 0 la_data_out[18]
rlabel metal2 194442 1690 194442 1690 0 la_data_out[19]
rlabel via1 140990 3315 140990 3315 0 la_data_out[1]
rlabel metal2 198129 340 198129 340 0 la_data_out[20]
rlabel metal2 201526 1758 201526 1758 0 la_data_out[21]
rlabel metal2 210542 2941 210542 2941 0 la_data_out[22]
rlabel via1 213854 3077 213854 3077 0 la_data_out[23]
rlabel metal2 212198 1656 212198 1656 0 la_data_out[24]
rlabel metal2 215694 1724 215694 1724 0 la_data_out[25]
rlabel metal2 219282 1622 219282 1622 0 la_data_out[26]
rlabel metal2 222778 1656 222778 1656 0 la_data_out[27]
rlabel metal2 230690 2968 230690 2968 0 la_data_out[28]
rlabel metal2 229862 1758 229862 1758 0 la_data_out[29]
rlabel metal2 134182 1724 134182 1724 0 la_data_out[2]
rlabel metal2 233450 1690 233450 1690 0 la_data_out[30]
rlabel metal2 237038 1622 237038 1622 0 la_data_out[31]
rlabel metal2 240534 1588 240534 1588 0 la_data_out[32]
rlabel metal2 244122 1588 244122 1588 0 la_data_out[33]
rlabel metal2 250562 2934 250562 2934 0 la_data_out[34]
rlabel metal2 251206 568 251206 568 0 la_data_out[35]
rlabel metal2 254702 1622 254702 1622 0 la_data_out[36]
rlabel metal2 258290 806 258290 806 0 la_data_out[37]
rlabel metal2 261786 1622 261786 1622 0 la_data_out[38]
rlabel metal2 265374 840 265374 840 0 la_data_out[39]
rlabel metal2 137579 204 137579 204 0 la_data_out[3]
rlabel metal2 268870 772 268870 772 0 la_data_out[40]
rlabel metal2 272458 806 272458 806 0 la_data_out[41]
rlabel metal2 276046 959 276046 959 0 la_data_out[42]
rlabel metal2 279542 840 279542 840 0 la_data_out[43]
rlabel metal2 283275 340 283275 340 0 la_data_out[44]
rlabel metal2 286817 340 286817 340 0 la_data_out[45]
rlabel metal2 290214 1707 290214 1707 0 la_data_out[46]
rlabel metal2 293710 1700 293710 1700 0 la_data_out[47]
rlabel metal2 297298 1707 297298 1707 0 la_data_out[48]
rlabel metal2 300794 1707 300794 1707 0 la_data_out[49]
rlabel metal2 141266 1622 141266 1622 0 la_data_out[4]
rlabel metal2 304145 340 304145 340 0 la_data_out[50]
rlabel metal2 307970 1588 307970 1588 0 la_data_out[51]
rlabel metal2 311466 1656 311466 1656 0 la_data_out[52]
rlabel metal2 315054 1588 315054 1588 0 la_data_out[53]
rlabel metal2 318550 1622 318550 1622 0 la_data_out[54]
rlabel metal2 322138 1588 322138 1588 0 la_data_out[55]
rlabel metal2 325634 1622 325634 1622 0 la_data_out[56]
rlabel metal2 329222 1588 329222 1588 0 la_data_out[57]
rlabel metal2 332718 1588 332718 1588 0 la_data_out[58]
rlabel metal2 333454 2968 333454 2968 0 la_data_out[59]
rlabel via1 154238 3621 154238 3621 0 la_data_out[5]
rlabel metal2 339894 840 339894 840 0 la_data_out[60]
rlabel metal2 343199 340 343199 340 0 la_data_out[61]
rlabel metal2 346978 806 346978 806 0 la_data_out[62]
rlabel metal2 350474 1588 350474 1588 0 la_data_out[63]
rlabel metal2 354062 806 354062 806 0 la_data_out[64]
rlabel metal2 353234 2934 353234 2934 0 la_data_out[65]
rlabel metal2 361146 840 361146 840 0 la_data_out[66]
rlabel metal2 364642 772 364642 772 0 la_data_out[67]
rlabel via1 367862 51 367862 51 0 la_data_out[68]
rlabel metal2 371535 340 371535 340 0 la_data_out[69]
rlabel via1 157550 3587 157550 3587 0 la_data_out[6]
rlabel metal2 369794 2186 369794 2186 0 la_data_out[70]
rlabel metal2 373198 2016 373198 2016 0 la_data_out[71]
rlabel metal2 382398 840 382398 840 0 la_data_out[72]
rlabel metal2 385986 772 385986 772 0 la_data_out[73]
rlabel via1 389666 85 389666 85 0 la_data_out[74]
rlabel metal2 392879 340 392879 340 0 la_data_out[75]
rlabel metal2 389758 1676 389758 1676 0 la_data_out[76]
rlabel metal2 393070 1846 393070 1846 0 la_data_out[77]
rlabel metal2 403650 806 403650 806 0 la_data_out[78]
rlabel via1 407054 51 407054 51 0 la_data_out[79]
rlabel metal2 151846 1724 151846 1724 0 la_data_out[7]
rlabel via1 411010 221 411010 221 0 la_data_out[80]
rlabel metal2 406318 2186 406318 2186 0 la_data_out[81]
rlabel metal2 409630 1846 409630 1846 0 la_data_out[82]
rlabel metal2 421406 738 421406 738 0 la_data_out[83]
rlabel metal2 424994 670 424994 670 0 la_data_out[84]
rlabel via1 428674 187 428674 187 0 la_data_out[85]
rlabel via1 431894 85 431894 85 0 la_data_out[86]
rlabel metal2 426190 1812 426190 1812 0 la_data_out[87]
rlabel metal2 429502 1778 429502 1778 0 la_data_out[88]
rlabel via1 442842 221 442842 221 0 la_data_out[89]
rlabel metal2 155434 1860 155434 1860 0 la_data_out[8]
rlabel metal2 446055 340 446055 340 0 la_data_out[90]
rlabel via1 450018 51 450018 51 0 la_data_out[91]
rlabel metal2 442750 1846 442750 1846 0 la_data_out[92]
rlabel metal2 446062 1880 446062 1880 0 la_data_out[93]
rlabel metal2 449374 1914 449374 1914 0 la_data_out[94]
rlabel via1 464186 51 464186 51 0 la_data_out[95]
rlabel metal2 467498 636 467498 636 0 la_data_out[96]
rlabel metal2 459494 1717 459494 1717 0 la_data_out[97]
rlabel metal2 462622 2186 462622 2186 0 la_data_out[98]
rlabel metal2 465842 1540 465842 1540 0 la_data_out[99]
rlabel metal2 158930 1622 158930 1622 0 la_data_out[9]
rlabel via1 138782 3043 138782 3043 0 la_oenb[0]
rlabel metal2 470350 1744 470350 1744 0 la_oenb[100]
rlabel metal2 486450 466 486450 466 0 la_oenb[101]
rlabel metal2 477250 1581 477250 1581 0 la_oenb[102]
rlabel metal2 480194 1982 480194 1982 0 la_oenb[103]
rlabel metal2 483598 1914 483598 1914 0 la_oenb[104]
rlabel metal2 486910 1778 486910 1778 0 la_oenb[105]
rlabel metal2 504015 340 504015 340 0 la_oenb[106]
rlabel metal2 507511 340 507511 340 0 la_oenb[107]
rlabel metal2 496754 1710 496754 1710 0 la_oenb[108]
rlabel metal2 507058 1054 507058 1054 0 la_oenb[109]
rlabel via1 171902 3485 171902 3485 0 la_oenb[10]
rlabel metal2 503470 2050 503470 2050 0 la_oenb[110]
rlabel metal2 506782 1540 506782 1540 0 la_oenb[111]
rlabel metal2 525458 636 525458 636 0 la_oenb[112]
rlabel metal2 513314 1574 513314 1574 0 la_oenb[113]
rlabel metal2 516718 2186 516718 2186 0 la_oenb[114]
rlabel metal2 520030 1608 520030 1608 0 la_oenb[115]
rlabel metal2 523342 1540 523342 1540 0 la_oenb[116]
rlabel metal2 526654 2968 526654 2968 0 la_oenb[117]
rlabel metal2 546710 1724 546710 1724 0 la_oenb[118]
rlabel metal2 533278 1710 533278 1710 0 la_oenb[119]
rlabel via1 175306 3349 175306 3349 0 la_oenb[11]
rlabel metal2 536590 3002 536590 3002 0 la_oenb[120]
rlabel metal2 546526 2074 546526 2074 0 la_oenb[121]
rlabel via1 543490 3043 543490 3043 0 la_oenb[122]
rlabel metal2 546434 1540 546434 1540 0 la_oenb[123]
rlabel metal2 549838 2968 549838 2968 0 la_oenb[124]
rlabel via1 553334 3213 553334 3213 0 la_oenb[125]
rlabel via1 556738 3179 556738 3179 0 la_oenb[126]
rlabel via1 560050 3315 560050 3315 0 la_oenb[127]
rlabel via1 178526 3179 178526 3179 0 la_oenb[12]
rlabel metal2 174294 1826 174294 1826 0 la_oenb[13]
rlabel metal2 177882 1656 177882 1656 0 la_oenb[14]
rlabel metal2 181470 1622 181470 1622 0 la_oenb[15]
rlabel metal2 192050 2934 192050 2934 0 la_oenb[16]
rlabel metal2 195362 2968 195362 2968 0 la_oenb[17]
rlabel metal2 192241 340 192241 340 0 la_oenb[18]
rlabel metal2 195638 1656 195638 1656 0 la_oenb[19]
rlabel metal2 131790 1656 131790 1656 0 la_oenb[1]
rlabel metal2 199134 1622 199134 1622 0 la_oenb[20]
rlabel metal2 202722 1690 202722 1690 0 la_oenb[21]
rlabel metal2 211646 2975 211646 2975 0 la_oenb[22]
rlabel metal2 209806 1656 209806 1656 0 la_oenb[23]
rlabel metal2 213394 1622 213394 1622 0 la_oenb[24]
rlabel metal2 216890 1588 216890 1588 0 la_oenb[25]
rlabel metal2 220379 204 220379 204 0 la_oenb[26]
rlabel metal2 223974 1588 223974 1588 0 la_oenb[27]
rlabel metal2 231794 3002 231794 3002 0 la_oenb[28]
rlabel metal2 231058 1724 231058 1724 0 la_oenb[29]
rlabel metal2 135286 1758 135286 1758 0 la_oenb[2]
rlabel metal2 234646 1656 234646 1656 0 la_oenb[30]
rlabel metal2 238142 1690 238142 1690 0 la_oenb[31]
rlabel metal2 241921 340 241921 340 0 la_oenb[32]
rlabel metal2 245226 1622 245226 1622 0 la_oenb[33]
rlabel metal2 248814 1690 248814 1690 0 la_oenb[34]
rlabel metal2 252402 1588 252402 1588 0 la_oenb[35]
rlabel metal2 255898 1588 255898 1588 0 la_oenb[36]
rlabel metal2 259486 840 259486 840 0 la_oenb[37]
rlabel metal2 262982 840 262982 840 0 la_oenb[38]
rlabel metal2 268226 2152 268226 2152 0 la_oenb[39]
rlabel metal2 139065 340 139065 340 0 la_oenb[3]
rlabel metal2 270066 806 270066 806 0 la_oenb[40]
rlabel metal2 273654 840 273654 840 0 la_oenb[41]
rlabel metal2 277150 840 277150 840 0 la_oenb[42]
rlabel metal2 280975 340 280975 340 0 la_oenb[43]
rlabel metal2 284326 1707 284326 1707 0 la_oenb[44]
rlabel metal2 287822 1707 287822 1707 0 la_oenb[45]
rlabel metal2 291410 1700 291410 1700 0 la_oenb[46]
rlabel metal2 294906 1707 294906 1707 0 la_oenb[47]
rlabel metal2 298303 340 298303 340 0 la_oenb[48]
rlabel metal2 301845 340 301845 340 0 la_oenb[49]
rlabel via1 152030 3485 152030 3485 0 la_oenb[4]
rlabel metal2 305578 1588 305578 1588 0 la_oenb[50]
rlabel metal2 309074 959 309074 959 0 la_oenb[51]
rlabel metal2 312662 1588 312662 1588 0 la_oenb[52]
rlabel metal2 314594 2968 314594 2968 0 la_oenb[53]
rlabel metal2 319746 1588 319746 1588 0 la_oenb[54]
rlabel metal2 323334 1622 323334 1622 0 la_oenb[55]
rlabel metal2 326830 1588 326830 1588 0 la_oenb[56]
rlabel metal2 330418 1622 330418 1622 0 la_oenb[57]
rlabel metal2 333914 1690 333914 1690 0 la_oenb[58]
rlabel via1 334834 3043 334834 3043 0 la_oenb[59]
rlabel metal2 155618 3002 155618 3002 0 la_oenb[5]
rlabel metal2 340998 602 340998 602 0 la_oenb[60]
rlabel metal2 344586 1656 344586 1656 0 la_oenb[61]
rlabel via1 348266 85 348266 85 0 la_oenb[62]
rlabel metal2 351670 602 351670 602 0 la_oenb[63]
rlabel metal2 351118 2016 351118 2016 0 la_oenb[64]
rlabel metal2 354430 1574 354430 1574 0 la_oenb[65]
rlabel metal2 362342 806 362342 806 0 la_oenb[66]
rlabel metal2 365647 340 365647 340 0 la_oenb[67]
rlabel metal2 369426 840 369426 840 0 la_oenb[68]
rlabel metal2 372922 704 372922 704 0 la_oenb[69]
rlabel metal2 158746 2941 158746 2941 0 la_oenb[6]
rlabel metal2 370990 2152 370990 2152 0 la_oenb[70]
rlabel metal2 379815 340 379815 340 0 la_oenb[71]
rlabel metal2 383594 704 383594 704 0 la_oenb[72]
rlabel via1 386814 187 386814 187 0 la_oenb[73]
rlabel metal2 390678 840 390678 840 0 la_oenb[74]
rlabel metal2 387550 2152 387550 2152 0 la_oenb[75]
rlabel metal2 390862 1642 390862 1642 0 la_oenb[76]
rlabel metal2 401350 840 401350 840 0 la_oenb[77]
rlabel metal2 404846 738 404846 738 0 la_oenb[78]
rlabel metal2 408434 466 408434 466 0 la_oenb[79]
rlabel metal2 153042 1894 153042 1894 0 la_oenb[7]
rlabel metal2 411930 806 411930 806 0 la_oenb[80]
rlabel metal2 407422 1710 407422 1710 0 la_oenb[81]
rlabel metal2 410642 1540 410642 1540 0 la_oenb[82]
rlabel via1 422786 323 422786 323 0 la_oenb[83]
rlabel metal2 425999 340 425999 340 0 la_oenb[84]
rlabel metal2 429495 340 429495 340 0 la_oenb[85]
rlabel metal2 423982 1880 423982 1880 0 la_oenb[86]
rlabel metal2 427570 1683 427570 1683 0 la_oenb[87]
rlabel metal2 430514 2152 430514 2152 0 la_oenb[88]
rlabel via1 443486 85 443486 85 0 la_oenb[89]
rlabel metal2 156630 1690 156630 1690 0 la_oenb[8]
rlabel metal2 447442 738 447442 738 0 la_oenb[90]
rlabel via1 451122 323 451122 323 0 la_oenb[91]
rlabel metal2 443854 2118 443854 2118 0 la_oenb[92]
rlabel metal2 447074 2152 447074 2152 0 la_oenb[93]
rlabel metal2 450478 2186 450478 2186 0 la_oenb[94]
rlabel via1 465014 187 465014 187 0 la_oenb[95]
rlabel metal2 468503 340 468503 340 0 la_oenb[96]
rlabel metal2 460598 1649 460598 1649 0 la_oenb[97]
rlabel metal2 463634 1574 463634 1574 0 la_oenb[98]
rlabel metal2 467038 1676 467038 1676 0 la_oenb[99]
rlabel metal2 160126 1588 160126 1588 0 la_oenb[9]
rlabel metal2 560878 3002 560878 3002 0 user_clock2
rlabel via1 562258 3043 562258 3043 0 user_irq[0]
rlabel metal2 562994 2934 562994 2934 0 user_irq[1]
rlabel via1 564374 3077 564374 3077 0 user_irq[2]
rlabel via1 414 51 414 51 0 wb_clk_i
rlabel via1 1518 187 1518 187 0 wb_rst_i
rlabel metal2 3089 340 3089 340 0 wbs_ack_o
rlabel via1 8050 85 8050 85 0 wbs_adr_i[0]
rlabel via1 63710 3043 63710 3043 0 wbs_adr_i[10]
rlabel metal2 51382 1758 51382 1758 0 wbs_adr_i[11]
rlabel metal2 54970 1656 54970 1656 0 wbs_adr_i[12]
rlabel metal2 58657 340 58657 340 0 wbs_adr_i[13]
rlabel metal2 62054 1826 62054 1826 0 wbs_adr_i[14]
rlabel metal2 79994 2941 79994 2941 0 wbs_adr_i[15]
rlabel metal2 83858 3002 83858 3002 0 wbs_adr_i[16]
rlabel metal2 72634 1962 72634 1962 0 wbs_adr_i[17]
rlabel metal2 76222 959 76222 959 0 wbs_adr_i[18]
rlabel metal2 79718 1996 79718 1996 0 wbs_adr_i[19]
rlabel metal2 12275 340 12275 340 0 wbs_adr_i[1]
rlabel metal2 83306 2030 83306 2030 0 wbs_adr_i[20]
rlabel metal2 86894 1588 86894 1588 0 wbs_adr_i[21]
rlabel metal2 90245 340 90245 340 0 wbs_adr_i[22]
rlabel metal2 93978 1894 93978 1894 0 wbs_adr_i[23]
rlabel metal2 97474 1758 97474 1758 0 wbs_adr_i[24]
rlabel via1 113114 3213 113114 3213 0 wbs_adr_i[25]
rlabel metal2 116978 2152 116978 2152 0 wbs_adr_i[26]
rlabel via1 120014 3043 120014 3043 0 wbs_adr_i[27]
rlabel metal2 111642 1588 111642 1588 0 wbs_adr_i[28]
rlabel metal2 115230 1724 115230 1724 0 wbs_adr_i[29]
rlabel via1 17434 323 17434 323 0 wbs_adr_i[2]
rlabel metal2 118818 2030 118818 2030 0 wbs_adr_i[30]
rlabel metal2 122314 1792 122314 1792 0 wbs_adr_i[31]
rlabel metal2 21850 670 21850 670 0 wbs_adr_i[3]
rlabel metal2 43838 2975 43838 2975 0 wbs_adr_i[4]
rlabel via1 30314 51 30314 51 0 wbs_adr_i[5]
rlabel metal2 33626 1656 33626 1656 0 wbs_adr_i[6]
rlabel metal2 37115 68 37115 68 0 wbs_adr_i[7]
rlabel metal2 40565 340 40565 340 0 wbs_adr_i[8]
rlabel metal2 44298 1622 44298 1622 0 wbs_adr_i[9]
rlabel via1 3910 221 3910 221 0 wbs_cyc_i
rlabel metal2 8977 340 8977 340 0 wbs_dat_i[0]
rlabel metal1 60030 3264 60030 3264 0 wbs_dat_i[10]
rlabel metal2 52578 1860 52578 1860 0 wbs_dat_i[11]
rlabel metal2 56074 1724 56074 1724 0 wbs_dat_i[12]
rlabel metal2 59662 1027 59662 1027 0 wbs_dat_i[13]
rlabel metal2 63250 2030 63250 2030 0 wbs_dat_i[14]
rlabel via1 81374 3179 81374 3179 0 wbs_dat_i[15]
rlabel metal2 70235 204 70235 204 0 wbs_dat_i[16]
rlabel metal2 73685 340 73685 340 0 wbs_dat_i[17]
rlabel metal2 77418 2064 77418 2064 0 wbs_dat_i[18]
rlabel metal2 80914 1792 80914 1792 0 wbs_dat_i[19]
rlabel metal2 13669 340 13669 340 0 wbs_dat_i[1]
rlabel metal2 98210 3002 98210 3002 0 wbs_dat_i[20]
rlabel metal2 87998 1724 87998 1724 0 wbs_dat_i[21]
rlabel metal2 91777 340 91777 340 0 wbs_dat_i[22]
rlabel metal2 95174 1996 95174 1996 0 wbs_dat_i[23]
rlabel metal2 98670 1928 98670 1928 0 wbs_dat_i[24]
rlabel via1 114586 3077 114586 3077 0 wbs_dat_i[25]
rlabel via1 117806 3757 117806 3757 0 wbs_dat_i[26]
rlabel via1 121118 3315 121118 3315 0 wbs_dat_i[27]
rlabel metal2 112838 1622 112838 1622 0 wbs_dat_i[28]
rlabel metal2 116426 1894 116426 1894 0 wbs_dat_i[29]
rlabel metal2 18262 500 18262 500 0 wbs_dat_i[2]
rlabel metal2 119922 1656 119922 1656 0 wbs_dat_i[30]
rlabel metal2 134642 2934 134642 2934 0 wbs_dat_i[31]
rlabel metal2 22947 340 22947 340 0 wbs_dat_i[3]
rlabel metal2 44942 2941 44942 2941 0 wbs_dat_i[4]
rlabel via1 31142 85 31142 85 0 wbs_dat_i[5]
rlabel metal2 34822 466 34822 466 0 wbs_dat_i[6]
rlabel via1 38594 323 38594 323 0 wbs_dat_i[7]
rlabel via1 42274 221 42274 221 0 wbs_dat_i[8]
rlabel metal2 45395 340 45395 340 0 wbs_dat_i[9]
rlabel metal2 9883 340 9883 340 0 wbs_dat_o[0]
rlabel metal2 50186 1588 50186 1588 0 wbs_dat_o[10]
rlabel via1 53590 51 53590 51 0 wbs_dat_o[11]
rlabel metal2 57125 340 57125 340 0 wbs_dat_o[12]
rlabel metal2 60858 1996 60858 1996 0 wbs_dat_o[13]
rlabel metal2 64354 2132 64354 2132 0 wbs_dat_o[14]
rlabel via1 82478 3349 82478 3349 0 wbs_dat_o[15]
rlabel metal2 71530 1095 71530 1095 0 wbs_dat_o[16]
rlabel metal2 75217 340 75217 340 0 wbs_dat_o[17]
rlabel metal2 78614 1622 78614 1622 0 wbs_dat_o[18]
rlabel metal2 82110 1758 82110 1758 0 wbs_dat_o[19]
rlabel metal2 14766 534 14766 534 0 wbs_dat_o[1]
rlabel via1 99038 3315 99038 3315 0 wbs_dat_o[20]
rlabel metal2 89385 340 89385 340 0 wbs_dat_o[21]
rlabel metal2 92782 1622 92782 1622 0 wbs_dat_o[22]
rlabel metal2 96278 1792 96278 1792 0 wbs_dat_o[23]
rlabel via1 112286 3859 112286 3859 0 wbs_dat_o[24]
rlabel via1 115598 3587 115598 3587 0 wbs_dat_o[25]
rlabel metal2 119186 3002 119186 3002 0 wbs_dat_o[26]
rlabel metal2 122222 3247 122222 3247 0 wbs_dat_o[27]
rlabel metal2 114034 1860 114034 1860 0 wbs_dat_o[28]
rlabel metal2 117622 1996 117622 1996 0 wbs_dat_o[29]
rlabel metal2 19458 636 19458 636 0 wbs_dat_o[2]
rlabel metal2 121019 204 121019 204 0 wbs_dat_o[30]
rlabel metal2 135746 2968 135746 2968 0 wbs_dat_o[31]
rlabel via1 24610 187 24610 187 0 wbs_dat_o[3]
rlabel metal2 28934 483 28934 483 0 wbs_dat_o[4]
rlabel metal2 32331 340 32331 340 0 wbs_dat_o[5]
rlabel metal2 36018 500 36018 500 0 wbs_dat_o[6]
rlabel metal2 39507 340 39507 340 0 wbs_dat_o[7]
rlabel via1 42918 187 42918 187 0 wbs_dat_o[8]
rlabel metal2 62882 1625 62882 1625 0 wbs_dat_o[9]
rlabel metal2 11178 602 11178 602 0 wbs_sel_i[0]
rlabel metal2 15962 466 15962 466 0 wbs_sel_i[1]
rlabel metal2 20654 568 20654 568 0 wbs_sel_i[2]
rlabel metal2 25537 204 25537 204 0 wbs_sel_i[3]
rlabel metal2 5389 204 5389 204 0 wbs_stb_i
rlabel metal2 6387 68 6387 68 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
