// SPDX-FileCopyrightText: 2022 SH CONSULTING K.K.
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

module j202_soc_core_wrapper ( wb_clk_i, wb_rst_i, wbs_stb_i, wbs_cyc_i, 
        wbs_we_i, wbs_sel_i, wbs_dat_i, wbs_adr_i, wbs_ack_o, wbs_dat_o, 
        la_data_in, la_data_out, la_oenb, io_in, io_out, io_oeb, analog_io, 
        user_clock2, user_irq );
  input [3:0] wbs_sel_i;
  input [31:0] wbs_dat_i;
  input [31:0] wbs_adr_i;
  output [31:0] wbs_dat_o;
  input [127:0] la_data_in;
  output [127:0] la_data_out;
  input [127:0] la_oenb;
  input [37:0] io_in;
  output [37:0] io_out;
  output [37:0] io_oeb;
  inout [28:0] analog_io;
  output [2:0] user_irq;
  input wb_clk_i, wb_rst_i, wbs_stb_i, wbs_cyc_i, wbs_we_i, user_clock2;
  output wbs_ack_o;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n220, n230, n240, n250, n260, n270, n280, n290, n300,
         n310, n320, n330, n340, n350, n360, n370, n380, n390,
         j202_soc_core_qspi_wb_we, j202_soc_core_qspi_wb_cyc,
         j202_soc_core_qspi_wb_ack, j202_soc_core_aquc_STB_,
         j202_soc_core_aquc_ADR__0_, j202_soc_core_aquc_ADR__1_,
         j202_soc_core_aquc_ADR__2_, j202_soc_core_aquc_ADR__3_,
         j202_soc_core_aquc_ADR__4_, j202_soc_core_aquc_ADR__5_,
         j202_soc_core_aquc_ADR__6_, j202_soc_core_aquc_ADR__7_,
         j202_soc_core_aquc_SEL__0_, j202_soc_core_aquc_SEL__2_,
         j202_soc_core_aquc_SEL__3_, j202_soc_core_aquc_WE_,
         j202_soc_core_aquc_CE__0_, j202_soc_core_aquc_CE__1_,
         j202_soc_core_bldc_int, j202_soc_core_qspi_int,
         j202_soc_core_ahbcs_6__HREADY_, j202_soc_core_intr_vec__0_,
         j202_soc_core_intr_vec__1_, j202_soc_core_intr_vec__2_,
         j202_soc_core_intr_vec__3_, j202_soc_core_intr_vec__4_,
         j202_soc_core_intr_vec__6_, j202_soc_core_intr_level__0_,
         j202_soc_core_intr_level__1_, j202_soc_core_intr_level__2_,
         j202_soc_core_intr_level__3_, j202_soc_core_intr_level__4_,
         j202_soc_core_intr_req_, j202_soc_core_rst, j202_soc_core_rst1,
         j202_soc_core_rst0, j202_soc_core_j22_cpu_regop_M_Wm__0_,
         j202_soc_core_j22_cpu_regop_M_Wm__1_,
         j202_soc_core_j22_cpu_regop_M_Wm__2_,
         j202_soc_core_j22_cpu_regop_M_Wm__3_,
         j202_soc_core_j22_cpu_regop_M_Rn__0_,
         j202_soc_core_j22_cpu_regop_M_Rn__1_,
         j202_soc_core_j22_cpu_regop_M_Rn__2_,
         j202_soc_core_j22_cpu_regop_M_Rn__3_,
         j202_soc_core_j22_cpu_regop_Wm__0_,
         j202_soc_core_j22_cpu_regop_Wm__1_,
         j202_soc_core_j22_cpu_regop_Wm__2_,
         j202_soc_core_j22_cpu_regop_Wm__3_,
         j202_soc_core_j22_cpu_regop_We__0_,
         j202_soc_core_j22_cpu_regop_We__1_,
         j202_soc_core_j22_cpu_regop_We__2_,
         j202_soc_core_j22_cpu_regop_We__3_,
         j202_soc_core_j22_cpu_regop_Rs__0_,
         j202_soc_core_j22_cpu_regop_Rs__1_,
         j202_soc_core_j22_cpu_regop_Rb__0_,
         j202_soc_core_j22_cpu_regop_Rb__1_,
         j202_soc_core_j22_cpu_regop_Ra__0_,
         j202_soc_core_j22_cpu_regop_Ra__1_,
         j202_soc_core_j22_cpu_regop_other__0_,
         j202_soc_core_j22_cpu_regop_other__1_,
         j202_soc_core_j22_cpu_regop_other__2_,
         j202_soc_core_j22_cpu_regop_imm__0_,
         j202_soc_core_j22_cpu_regop_imm__1_,
         j202_soc_core_j22_cpu_regop_imm__2_,
         j202_soc_core_j22_cpu_regop_imm__3_,
         j202_soc_core_j22_cpu_regop_imm__4_,
         j202_soc_core_j22_cpu_regop_imm__5_,
         j202_soc_core_j22_cpu_regop_imm__6_,
         j202_soc_core_j22_cpu_regop_imm__7_,
         j202_soc_core_j22_cpu_regop_imm__8_,
         j202_soc_core_j22_cpu_regop_imm__9_,
         j202_soc_core_j22_cpu_regop_imm__10_,
         j202_soc_core_j22_cpu_regop_imm__11_,
         j202_soc_core_j22_cpu_regop_imm__12_,
         j202_soc_core_j22_cpu_regop_Rm__0_,
         j202_soc_core_j22_cpu_regop_Rm__1_,
         j202_soc_core_j22_cpu_regop_Rm__2_,
         j202_soc_core_j22_cpu_regop_Rm__3_,
         j202_soc_core_j22_cpu_regop_Rn__0_,
         j202_soc_core_j22_cpu_regop_Rn__1_,
         j202_soc_core_j22_cpu_regop_Rn__2_,
         j202_soc_core_j22_cpu_regop_Rn__3_, j202_soc_core_j22_cpu_ifetch,
         j202_soc_core_j22_cpu_memop_Ma__0_,
         j202_soc_core_j22_cpu_memop_Ma__1_,
         j202_soc_core_j22_cpu_memop_MEM__0_,
         j202_soc_core_j22_cpu_memop_MEM__1_,
         j202_soc_core_j22_cpu_memop_MEM__2_,
         j202_soc_core_j22_cpu_memop_MEM__3_, j202_soc_core_j22_cpu_pc_hold,
         j202_soc_core_j22_cpu_istall, j202_soc_core_j22_cpu_intack,
         j202_soc_core_j22_cpu_N8, j202_soc_core_j22_cpu_rte4,
         j202_soc_core_j22_cpu_rfuo_sr__t_, j202_soc_core_j22_cpu_rfuo_sr__s_,
         j202_soc_core_j22_cpu_rfuo_sr__i__0_,
         j202_soc_core_j22_cpu_rfuo_sr__i__1_,
         j202_soc_core_j22_cpu_rfuo_sr__i__2_,
         j202_soc_core_j22_cpu_rfuo_sr__i__3_,
         j202_soc_core_j22_cpu_rfuo_sr__q_, j202_soc_core_j22_cpu_rfuo_sr__m_,
         j202_soc_core_j22_cpu_ifetchl, j202_soc_core_j22_cpu_id_opn_v_,
         j202_soc_core_j22_cpu_id_opn_inst__0_,
         j202_soc_core_j22_cpu_id_opn_inst__1_,
         j202_soc_core_j22_cpu_id_opn_inst__2_,
         j202_soc_core_j22_cpu_id_opn_inst__3_,
         j202_soc_core_j22_cpu_id_opn_inst__4_,
         j202_soc_core_j22_cpu_id_opn_inst__5_,
         j202_soc_core_j22_cpu_id_opn_inst__6_,
         j202_soc_core_j22_cpu_id_opn_inst__7_,
         j202_soc_core_j22_cpu_id_opn_inst__8_,
         j202_soc_core_j22_cpu_id_opn_inst__9_,
         j202_soc_core_j22_cpu_id_opn_inst__10_,
         j202_soc_core_j22_cpu_id_opn_inst__11_,
         j202_soc_core_j22_cpu_id_opn_inst__12_,
         j202_soc_core_j22_cpu_id_opn_inst__13_,
         j202_soc_core_j22_cpu_id_opn_inst__14_,
         j202_soc_core_j22_cpu_id_opn_inst__15_, j202_soc_core_j22_cpu_id_N7,
         j202_soc_core_j22_cpu_id_op2_v_,
         j202_soc_core_j22_cpu_id_op2_inst__0_,
         j202_soc_core_j22_cpu_id_op2_inst__1_,
         j202_soc_core_j22_cpu_id_op2_inst__2_,
         j202_soc_core_j22_cpu_id_op2_inst__3_,
         j202_soc_core_j22_cpu_id_op2_inst__4_,
         j202_soc_core_j22_cpu_id_op2_inst__5_,
         j202_soc_core_j22_cpu_id_op2_inst__6_,
         j202_soc_core_j22_cpu_id_op2_inst__7_,
         j202_soc_core_j22_cpu_id_op2_inst__8_,
         j202_soc_core_j22_cpu_id_op2_inst__9_,
         j202_soc_core_j22_cpu_id_op2_inst__10_,
         j202_soc_core_j22_cpu_id_op2_inst__11_,
         j202_soc_core_j22_cpu_id_op2_inst__12_,
         j202_soc_core_j22_cpu_id_op2_inst__13_,
         j202_soc_core_j22_cpu_id_op2_inst__14_,
         j202_soc_core_j22_cpu_id_op2_inst__15_,
         j202_soc_core_j22_cpu_id_idec_N960,
         j202_soc_core_j22_cpu_id_idec_N959,
         j202_soc_core_j22_cpu_id_idec_N958,
         j202_soc_core_j22_cpu_id_idec_N957,
         j202_soc_core_j22_cpu_id_idec_N956,
         j202_soc_core_j22_cpu_id_idec_N937,
         j202_soc_core_j22_cpu_id_idec_N917,
         j202_soc_core_j22_cpu_id_idec_N900,
         j202_soc_core_j22_cpu_id_idec_N894,
         j202_soc_core_j22_cpu_id_idec_N857,
         j202_soc_core_j22_cpu_id_idec_N822, j202_soc_core_j22_cpu_rf_N3392,
         j202_soc_core_j22_cpu_rf_N3391, j202_soc_core_j22_cpu_rf_N3390,
         j202_soc_core_j22_cpu_rf_N3388, j202_soc_core_j22_cpu_rf_N3386,
         j202_soc_core_j22_cpu_rf_N3379, j202_soc_core_j22_cpu_rf_N3378,
         j202_soc_core_j22_cpu_rf_N3377, j202_soc_core_j22_cpu_rf_N3376,
         j202_soc_core_j22_cpu_rf_N3375, j202_soc_core_j22_cpu_rf_N3374,
         j202_soc_core_j22_cpu_rf_N3373, j202_soc_core_j22_cpu_rf_N3372,
         j202_soc_core_j22_cpu_rf_N3371, j202_soc_core_j22_cpu_rf_N3370,
         j202_soc_core_j22_cpu_rf_N3369, j202_soc_core_j22_cpu_rf_N3368,
         j202_soc_core_j22_cpu_rf_N3367, j202_soc_core_j22_cpu_rf_N3366,
         j202_soc_core_j22_cpu_rf_N3365, j202_soc_core_j22_cpu_rf_N3364,
         j202_soc_core_j22_cpu_rf_N3363, j202_soc_core_j22_cpu_rf_N3361,
         j202_soc_core_j22_cpu_rf_N3360, j202_soc_core_j22_cpu_rf_N3359,
         j202_soc_core_j22_cpu_rf_N3358, j202_soc_core_j22_cpu_rf_N3357,
         j202_soc_core_j22_cpu_rf_N3356, j202_soc_core_j22_cpu_rf_N3355,
         j202_soc_core_j22_cpu_rf_N3354, j202_soc_core_j22_cpu_rf_N3352,
         j202_soc_core_j22_cpu_rf_N3351, j202_soc_core_j22_cpu_rf_N3350,
         j202_soc_core_j22_cpu_rf_N3349, j202_soc_core_j22_cpu_rf_N3348,
         j202_soc_core_j22_cpu_rf_N3347, j202_soc_core_j22_cpu_rf_N3346,
         j202_soc_core_j22_cpu_rf_N3345, j202_soc_core_j22_cpu_rf_N3343,
         j202_soc_core_j22_cpu_rf_N3342, j202_soc_core_j22_cpu_rf_N3341,
         j202_soc_core_j22_cpu_rf_N3340, j202_soc_core_j22_cpu_rf_N3339,
         j202_soc_core_j22_cpu_rf_N3338, j202_soc_core_j22_cpu_rf_N3337,
         j202_soc_core_j22_cpu_rf_N3336, j202_soc_core_j22_cpu_rf_N3335,
         j202_soc_core_j22_cpu_rf_N3334, j202_soc_core_j22_cpu_rf_N3333,
         j202_soc_core_j22_cpu_rf_N3331, j202_soc_core_j22_cpu_rf_N3330,
         j202_soc_core_j22_cpu_rf_N3329, j202_soc_core_j22_cpu_rf_N3328,
         j202_soc_core_j22_cpu_rf_N3327, j202_soc_core_j22_cpu_rf_N3326,
         j202_soc_core_j22_cpu_rf_N3325, j202_soc_core_j22_cpu_rf_N3324,
         j202_soc_core_j22_cpu_rf_N3323, j202_soc_core_j22_cpu_rf_N3322,
         j202_soc_core_j22_cpu_rf_N3321, j202_soc_core_j22_cpu_rf_N3319,
         j202_soc_core_j22_cpu_rf_N3318, j202_soc_core_j22_cpu_rf_N3317,
         j202_soc_core_j22_cpu_rf_N3316, j202_soc_core_j22_cpu_rf_N3315,
         j202_soc_core_j22_cpu_rf_N3314, j202_soc_core_j22_cpu_rf_N3313,
         j202_soc_core_j22_cpu_rf_N3311, j202_soc_core_j22_cpu_rf_N3309,
         j202_soc_core_j22_cpu_rf_N3307, j202_soc_core_j22_cpu_rf_N3305,
         j202_soc_core_j22_cpu_rf_N3304, j202_soc_core_j22_cpu_rf_N3303,
         j202_soc_core_j22_cpu_rf_N3302, j202_soc_core_j22_cpu_rf_N3301,
         j202_soc_core_j22_cpu_rf_N3300, j202_soc_core_j22_cpu_rf_N3299,
         j202_soc_core_j22_cpu_rf_N3298, j202_soc_core_j22_cpu_rf_N3297,
         j202_soc_core_j22_cpu_rf_N3296, j202_soc_core_j22_cpu_rf_N3295,
         j202_soc_core_j22_cpu_rf_N3294, j202_soc_core_j22_cpu_rf_N3292,
         j202_soc_core_j22_cpu_rf_N3291, j202_soc_core_j22_cpu_rf_N3290,
         j202_soc_core_j22_cpu_rf_N3289, j202_soc_core_j22_cpu_rf_N3288,
         j202_soc_core_j22_cpu_rf_N3287, j202_soc_core_j22_cpu_rf_N3286,
         j202_soc_core_j22_cpu_rf_N3284, j202_soc_core_j22_cpu_rf_N3283,
         j202_soc_core_j22_cpu_rf_N3282, j202_soc_core_j22_cpu_rf_N3281,
         j202_soc_core_j22_cpu_rf_N3280, j202_soc_core_j22_cpu_rf_N3279,
         j202_soc_core_j22_cpu_rf_N3278, j202_soc_core_j22_cpu_rf_N3276,
         j202_soc_core_j22_cpu_rf_N3275, j202_soc_core_j22_cpu_rf_N3274,
         j202_soc_core_j22_cpu_rf_N3273, j202_soc_core_j22_cpu_rf_N3272,
         j202_soc_core_j22_cpu_rf_N3271, j202_soc_core_j22_cpu_rf_N3270,
         j202_soc_core_j22_cpu_rf_N3268, j202_soc_core_j22_cpu_rf_N3267,
         j202_soc_core_j22_cpu_rf_N3266, j202_soc_core_j22_cpu_rf_N3265,
         j202_soc_core_j22_cpu_rf_N3264, j202_soc_core_j22_cpu_rf_N3263,
         j202_soc_core_j22_cpu_rf_N3262, j202_soc_core_j22_cpu_rf_N3261,
         j202_soc_core_j22_cpu_rf_N3260, j202_soc_core_j22_cpu_rf_N3259,
         j202_soc_core_j22_cpu_rf_N3258, j202_soc_core_j22_cpu_rf_N3257,
         j202_soc_core_j22_cpu_rf_N3255, j202_soc_core_j22_cpu_rf_N3254,
         j202_soc_core_j22_cpu_rf_N3253, j202_soc_core_j22_cpu_rf_N3252,
         j202_soc_core_j22_cpu_rf_N3251, j202_soc_core_j22_cpu_rf_N3250,
         j202_soc_core_j22_cpu_rf_N3249, j202_soc_core_j22_cpu_rf_N3247,
         j202_soc_core_j22_cpu_rf_N3246, j202_soc_core_j22_cpu_rf_N3245,
         j202_soc_core_j22_cpu_rf_N3244, j202_soc_core_j22_cpu_rf_N3243,
         j202_soc_core_j22_cpu_rf_N3242, j202_soc_core_j22_cpu_rf_N3241,
         j202_soc_core_j22_cpu_rf_N3239, j202_soc_core_j22_cpu_rf_N3238,
         j202_soc_core_j22_cpu_rf_N3237, j202_soc_core_j22_cpu_rf_N3236,
         j202_soc_core_j22_cpu_rf_N3235, j202_soc_core_j22_cpu_rf_N3234,
         j202_soc_core_j22_cpu_rf_N3233, j202_soc_core_j22_cpu_rf_N3231,
         j202_soc_core_j22_cpu_rf_N3230, j202_soc_core_j22_cpu_rf_N3229,
         j202_soc_core_j22_cpu_rf_N3228, j202_soc_core_j22_cpu_rf_N3227,
         j202_soc_core_j22_cpu_rf_N3226, j202_soc_core_j22_cpu_rf_N3225,
         j202_soc_core_j22_cpu_rf_N3224, j202_soc_core_j22_cpu_rf_N3223,
         j202_soc_core_j22_cpu_rf_N3222, j202_soc_core_j22_cpu_rf_N3221,
         j202_soc_core_j22_cpu_rf_N3220, j202_soc_core_j22_cpu_rf_N3218,
         j202_soc_core_j22_cpu_rf_N3217, j202_soc_core_j22_cpu_rf_N3216,
         j202_soc_core_j22_cpu_rf_N3215, j202_soc_core_j22_cpu_rf_N3214,
         j202_soc_core_j22_cpu_rf_N3213, j202_soc_core_j22_cpu_rf_N3212,
         j202_soc_core_j22_cpu_rf_N3210, j202_soc_core_j22_cpu_rf_N3209,
         j202_soc_core_j22_cpu_rf_N3208, j202_soc_core_j22_cpu_rf_N3207,
         j202_soc_core_j22_cpu_rf_N3206, j202_soc_core_j22_cpu_rf_N3205,
         j202_soc_core_j22_cpu_rf_N3204, j202_soc_core_j22_cpu_rf_N3202,
         j202_soc_core_j22_cpu_rf_N3201, j202_soc_core_j22_cpu_rf_N3200,
         j202_soc_core_j22_cpu_rf_N3199, j202_soc_core_j22_cpu_rf_N3198,
         j202_soc_core_j22_cpu_rf_N3197, j202_soc_core_j22_cpu_rf_N3196,
         j202_soc_core_j22_cpu_rf_N3194, j202_soc_core_j22_cpu_rf_N3193,
         j202_soc_core_j22_cpu_rf_N3192, j202_soc_core_j22_cpu_rf_N3191,
         j202_soc_core_j22_cpu_rf_N3190, j202_soc_core_j22_cpu_rf_N3189,
         j202_soc_core_j22_cpu_rf_N3188, j202_soc_core_j22_cpu_rf_N3187,
         j202_soc_core_j22_cpu_rf_N3186, j202_soc_core_j22_cpu_rf_N3185,
         j202_soc_core_j22_cpu_rf_N3184, j202_soc_core_j22_cpu_rf_N3183,
         j202_soc_core_j22_cpu_rf_N3181, j202_soc_core_j22_cpu_rf_N3180,
         j202_soc_core_j22_cpu_rf_N3179, j202_soc_core_j22_cpu_rf_N3178,
         j202_soc_core_j22_cpu_rf_N3177, j202_soc_core_j22_cpu_rf_N3176,
         j202_soc_core_j22_cpu_rf_N3175, j202_soc_core_j22_cpu_rf_N3173,
         j202_soc_core_j22_cpu_rf_N3172, j202_soc_core_j22_cpu_rf_N3171,
         j202_soc_core_j22_cpu_rf_N3170, j202_soc_core_j22_cpu_rf_N3169,
         j202_soc_core_j22_cpu_rf_N3168, j202_soc_core_j22_cpu_rf_N3167,
         j202_soc_core_j22_cpu_rf_N3165, j202_soc_core_j22_cpu_rf_N3164,
         j202_soc_core_j22_cpu_rf_N3163, j202_soc_core_j22_cpu_rf_N3162,
         j202_soc_core_j22_cpu_rf_N3161, j202_soc_core_j22_cpu_rf_N3160,
         j202_soc_core_j22_cpu_rf_N3159, j202_soc_core_j22_cpu_rf_N3157,
         j202_soc_core_j22_cpu_rf_N3156, j202_soc_core_j22_cpu_rf_N3155,
         j202_soc_core_j22_cpu_rf_N3154, j202_soc_core_j22_cpu_rf_N3153,
         j202_soc_core_j22_cpu_rf_N3152, j202_soc_core_j22_cpu_rf_N3151,
         j202_soc_core_j22_cpu_rf_N3150, j202_soc_core_j22_cpu_rf_N3149,
         j202_soc_core_j22_cpu_rf_N3148, j202_soc_core_j22_cpu_rf_N3147,
         j202_soc_core_j22_cpu_rf_N3146, j202_soc_core_j22_cpu_rf_N3144,
         j202_soc_core_j22_cpu_rf_N3143, j202_soc_core_j22_cpu_rf_N3142,
         j202_soc_core_j22_cpu_rf_N3141, j202_soc_core_j22_cpu_rf_N3140,
         j202_soc_core_j22_cpu_rf_N3139, j202_soc_core_j22_cpu_rf_N3138,
         j202_soc_core_j22_cpu_rf_N3136, j202_soc_core_j22_cpu_rf_N3135,
         j202_soc_core_j22_cpu_rf_N3134, j202_soc_core_j22_cpu_rf_N3133,
         j202_soc_core_j22_cpu_rf_N3132, j202_soc_core_j22_cpu_rf_N3131,
         j202_soc_core_j22_cpu_rf_N3130, j202_soc_core_j22_cpu_rf_N3128,
         j202_soc_core_j22_cpu_rf_N3127, j202_soc_core_j22_cpu_rf_N3126,
         j202_soc_core_j22_cpu_rf_N3125, j202_soc_core_j22_cpu_rf_N3124,
         j202_soc_core_j22_cpu_rf_N3123, j202_soc_core_j22_cpu_rf_N3122,
         j202_soc_core_j22_cpu_rf_N3120, j202_soc_core_j22_cpu_rf_N3119,
         j202_soc_core_j22_cpu_rf_N3118, j202_soc_core_j22_cpu_rf_N3117,
         j202_soc_core_j22_cpu_rf_N3116, j202_soc_core_j22_cpu_rf_N3115,
         j202_soc_core_j22_cpu_rf_N3114, j202_soc_core_j22_cpu_rf_N3113,
         j202_soc_core_j22_cpu_rf_N3112, j202_soc_core_j22_cpu_rf_N3111,
         j202_soc_core_j22_cpu_rf_N3110, j202_soc_core_j22_cpu_rf_N3109,
         j202_soc_core_j22_cpu_rf_N3107, j202_soc_core_j22_cpu_rf_N3106,
         j202_soc_core_j22_cpu_rf_N3105, j202_soc_core_j22_cpu_rf_N3104,
         j202_soc_core_j22_cpu_rf_N3103, j202_soc_core_j22_cpu_rf_N3102,
         j202_soc_core_j22_cpu_rf_N3101, j202_soc_core_j22_cpu_rf_N3099,
         j202_soc_core_j22_cpu_rf_N3098, j202_soc_core_j22_cpu_rf_N3097,
         j202_soc_core_j22_cpu_rf_N3096, j202_soc_core_j22_cpu_rf_N3095,
         j202_soc_core_j22_cpu_rf_N3094, j202_soc_core_j22_cpu_rf_N3093,
         j202_soc_core_j22_cpu_rf_N3091, j202_soc_core_j22_cpu_rf_N3090,
         j202_soc_core_j22_cpu_rf_N3089, j202_soc_core_j22_cpu_rf_N3088,
         j202_soc_core_j22_cpu_rf_N3087, j202_soc_core_j22_cpu_rf_N3086,
         j202_soc_core_j22_cpu_rf_N3085, j202_soc_core_j22_cpu_rf_N3083,
         j202_soc_core_j22_cpu_rf_N3082, j202_soc_core_j22_cpu_rf_N3081,
         j202_soc_core_j22_cpu_rf_N3080, j202_soc_core_j22_cpu_rf_N3079,
         j202_soc_core_j22_cpu_rf_N3078, j202_soc_core_j22_cpu_rf_N3077,
         j202_soc_core_j22_cpu_rf_N3076, j202_soc_core_j22_cpu_rf_N3075,
         j202_soc_core_j22_cpu_rf_N3074, j202_soc_core_j22_cpu_rf_N3073,
         j202_soc_core_j22_cpu_rf_N3072, j202_soc_core_j22_cpu_rf_N3070,
         j202_soc_core_j22_cpu_rf_N3069, j202_soc_core_j22_cpu_rf_N3068,
         j202_soc_core_j22_cpu_rf_N3067, j202_soc_core_j22_cpu_rf_N3066,
         j202_soc_core_j22_cpu_rf_N3065, j202_soc_core_j22_cpu_rf_N3064,
         j202_soc_core_j22_cpu_rf_N3062, j202_soc_core_j22_cpu_rf_N3061,
         j202_soc_core_j22_cpu_rf_N3060, j202_soc_core_j22_cpu_rf_N3059,
         j202_soc_core_j22_cpu_rf_N3058, j202_soc_core_j22_cpu_rf_N3057,
         j202_soc_core_j22_cpu_rf_N3056, j202_soc_core_j22_cpu_rf_N3054,
         j202_soc_core_j22_cpu_rf_N3053, j202_soc_core_j22_cpu_rf_N3052,
         j202_soc_core_j22_cpu_rf_N3051, j202_soc_core_j22_cpu_rf_N3050,
         j202_soc_core_j22_cpu_rf_N3049, j202_soc_core_j22_cpu_rf_N3048,
         j202_soc_core_j22_cpu_rf_N3046, j202_soc_core_j22_cpu_rf_N3045,
         j202_soc_core_j22_cpu_rf_N3044, j202_soc_core_j22_cpu_rf_N3043,
         j202_soc_core_j22_cpu_rf_N3042, j202_soc_core_j22_cpu_rf_N3041,
         j202_soc_core_j22_cpu_rf_N3040, j202_soc_core_j22_cpu_rf_N3039,
         j202_soc_core_j22_cpu_rf_N3038, j202_soc_core_j22_cpu_rf_N3037,
         j202_soc_core_j22_cpu_rf_N3036, j202_soc_core_j22_cpu_rf_N3035,
         j202_soc_core_j22_cpu_rf_N3033, j202_soc_core_j22_cpu_rf_N3032,
         j202_soc_core_j22_cpu_rf_N3031, j202_soc_core_j22_cpu_rf_N3030,
         j202_soc_core_j22_cpu_rf_N3029, j202_soc_core_j22_cpu_rf_N3028,
         j202_soc_core_j22_cpu_rf_N3027, j202_soc_core_j22_cpu_rf_N3025,
         j202_soc_core_j22_cpu_rf_N3024, j202_soc_core_j22_cpu_rf_N3023,
         j202_soc_core_j22_cpu_rf_N3022, j202_soc_core_j22_cpu_rf_N3021,
         j202_soc_core_j22_cpu_rf_N3020, j202_soc_core_j22_cpu_rf_N3019,
         j202_soc_core_j22_cpu_rf_N3017, j202_soc_core_j22_cpu_rf_N3016,
         j202_soc_core_j22_cpu_rf_N3015, j202_soc_core_j22_cpu_rf_N3014,
         j202_soc_core_j22_cpu_rf_N3013, j202_soc_core_j22_cpu_rf_N3012,
         j202_soc_core_j22_cpu_rf_N3011, j202_soc_core_j22_cpu_rf_N3009,
         j202_soc_core_j22_cpu_rf_N3008, j202_soc_core_j22_cpu_rf_N3007,
         j202_soc_core_j22_cpu_rf_N3006, j202_soc_core_j22_cpu_rf_N3005,
         j202_soc_core_j22_cpu_rf_N3004, j202_soc_core_j22_cpu_rf_N3003,
         j202_soc_core_j22_cpu_rf_N3002, j202_soc_core_j22_cpu_rf_N3001,
         j202_soc_core_j22_cpu_rf_N3000, j202_soc_core_j22_cpu_rf_N2999,
         j202_soc_core_j22_cpu_rf_N2998, j202_soc_core_j22_cpu_rf_N2996,
         j202_soc_core_j22_cpu_rf_N2995, j202_soc_core_j22_cpu_rf_N2994,
         j202_soc_core_j22_cpu_rf_N2993, j202_soc_core_j22_cpu_rf_N2992,
         j202_soc_core_j22_cpu_rf_N2991, j202_soc_core_j22_cpu_rf_N2990,
         j202_soc_core_j22_cpu_rf_N2988, j202_soc_core_j22_cpu_rf_N2987,
         j202_soc_core_j22_cpu_rf_N2986, j202_soc_core_j22_cpu_rf_N2985,
         j202_soc_core_j22_cpu_rf_N2984, j202_soc_core_j22_cpu_rf_N2983,
         j202_soc_core_j22_cpu_rf_N2982, j202_soc_core_j22_cpu_rf_N2980,
         j202_soc_core_j22_cpu_rf_N2979, j202_soc_core_j22_cpu_rf_N2978,
         j202_soc_core_j22_cpu_rf_N2977, j202_soc_core_j22_cpu_rf_N2976,
         j202_soc_core_j22_cpu_rf_N2975, j202_soc_core_j22_cpu_rf_N2974,
         j202_soc_core_j22_cpu_rf_N2972, j202_soc_core_j22_cpu_rf_N2971,
         j202_soc_core_j22_cpu_rf_N2970, j202_soc_core_j22_cpu_rf_N2969,
         j202_soc_core_j22_cpu_rf_N2968, j202_soc_core_j22_cpu_rf_N2967,
         j202_soc_core_j22_cpu_rf_N2966, j202_soc_core_j22_cpu_rf_N2965,
         j202_soc_core_j22_cpu_rf_N2964, j202_soc_core_j22_cpu_rf_N2963,
         j202_soc_core_j22_cpu_rf_N2962, j202_soc_core_j22_cpu_rf_N2961,
         j202_soc_core_j22_cpu_rf_N2959, j202_soc_core_j22_cpu_rf_N2958,
         j202_soc_core_j22_cpu_rf_N2957, j202_soc_core_j22_cpu_rf_N2956,
         j202_soc_core_j22_cpu_rf_N2955, j202_soc_core_j22_cpu_rf_N2954,
         j202_soc_core_j22_cpu_rf_N2953, j202_soc_core_j22_cpu_rf_N2951,
         j202_soc_core_j22_cpu_rf_N2950, j202_soc_core_j22_cpu_rf_N2949,
         j202_soc_core_j22_cpu_rf_N2948, j202_soc_core_j22_cpu_rf_N2947,
         j202_soc_core_j22_cpu_rf_N2946, j202_soc_core_j22_cpu_rf_N2945,
         j202_soc_core_j22_cpu_rf_N2943, j202_soc_core_j22_cpu_rf_N2942,
         j202_soc_core_j22_cpu_rf_N2941, j202_soc_core_j22_cpu_rf_N2940,
         j202_soc_core_j22_cpu_rf_N2939, j202_soc_core_j22_cpu_rf_N2938,
         j202_soc_core_j22_cpu_rf_N2937, j202_soc_core_j22_cpu_rf_N2935,
         j202_soc_core_j22_cpu_rf_N2934, j202_soc_core_j22_cpu_rf_N2933,
         j202_soc_core_j22_cpu_rf_N2932, j202_soc_core_j22_cpu_rf_N2931,
         j202_soc_core_j22_cpu_rf_N2930, j202_soc_core_j22_cpu_rf_N2929,
         j202_soc_core_j22_cpu_rf_N2928, j202_soc_core_j22_cpu_rf_N2927,
         j202_soc_core_j22_cpu_rf_N2926, j202_soc_core_j22_cpu_rf_N2925,
         j202_soc_core_j22_cpu_rf_N2924, j202_soc_core_j22_cpu_rf_N2922,
         j202_soc_core_j22_cpu_rf_N2921, j202_soc_core_j22_cpu_rf_N2920,
         j202_soc_core_j22_cpu_rf_N2919, j202_soc_core_j22_cpu_rf_N2918,
         j202_soc_core_j22_cpu_rf_N2917, j202_soc_core_j22_cpu_rf_N2916,
         j202_soc_core_j22_cpu_rf_N2914, j202_soc_core_j22_cpu_rf_N2913,
         j202_soc_core_j22_cpu_rf_N2912, j202_soc_core_j22_cpu_rf_N2911,
         j202_soc_core_j22_cpu_rf_N2910, j202_soc_core_j22_cpu_rf_N2909,
         j202_soc_core_j22_cpu_rf_N2908, j202_soc_core_j22_cpu_rf_N2906,
         j202_soc_core_j22_cpu_rf_N2905, j202_soc_core_j22_cpu_rf_N2904,
         j202_soc_core_j22_cpu_rf_N2903, j202_soc_core_j22_cpu_rf_N2902,
         j202_soc_core_j22_cpu_rf_N2901, j202_soc_core_j22_cpu_rf_N2900,
         j202_soc_core_j22_cpu_rf_N2898, j202_soc_core_j22_cpu_rf_N2897,
         j202_soc_core_j22_cpu_rf_N2896, j202_soc_core_j22_cpu_rf_N2895,
         j202_soc_core_j22_cpu_rf_N2894, j202_soc_core_j22_cpu_rf_N2893,
         j202_soc_core_j22_cpu_rf_N2892, j202_soc_core_j22_cpu_rf_N2891,
         j202_soc_core_j22_cpu_rf_N2890, j202_soc_core_j22_cpu_rf_N2889,
         j202_soc_core_j22_cpu_rf_N2888, j202_soc_core_j22_cpu_rf_N2887,
         j202_soc_core_j22_cpu_rf_N2885, j202_soc_core_j22_cpu_rf_N2884,
         j202_soc_core_j22_cpu_rf_N2883, j202_soc_core_j22_cpu_rf_N2882,
         j202_soc_core_j22_cpu_rf_N2881, j202_soc_core_j22_cpu_rf_N2880,
         j202_soc_core_j22_cpu_rf_N2879, j202_soc_core_j22_cpu_rf_N2877,
         j202_soc_core_j22_cpu_rf_N2876, j202_soc_core_j22_cpu_rf_N2875,
         j202_soc_core_j22_cpu_rf_N2874, j202_soc_core_j22_cpu_rf_N2873,
         j202_soc_core_j22_cpu_rf_N2872, j202_soc_core_j22_cpu_rf_N2871,
         j202_soc_core_j22_cpu_rf_N2869, j202_soc_core_j22_cpu_rf_N2868,
         j202_soc_core_j22_cpu_rf_N2867, j202_soc_core_j22_cpu_rf_N2866,
         j202_soc_core_j22_cpu_rf_N2865, j202_soc_core_j22_cpu_rf_N2864,
         j202_soc_core_j22_cpu_rf_N2863, j202_soc_core_j22_cpu_rf_N2861,
         j202_soc_core_j22_cpu_rf_N2860, j202_soc_core_j22_cpu_rf_N2859,
         j202_soc_core_j22_cpu_rf_N2858, j202_soc_core_j22_cpu_rf_N2857,
         j202_soc_core_j22_cpu_rf_N2856, j202_soc_core_j22_cpu_rf_N2855,
         j202_soc_core_j22_cpu_rf_N2854, j202_soc_core_j22_cpu_rf_N2853,
         j202_soc_core_j22_cpu_rf_N2852, j202_soc_core_j22_cpu_rf_N2851,
         j202_soc_core_j22_cpu_rf_N2850, j202_soc_core_j22_cpu_rf_N2848,
         j202_soc_core_j22_cpu_rf_N2847, j202_soc_core_j22_cpu_rf_N2846,
         j202_soc_core_j22_cpu_rf_N2845, j202_soc_core_j22_cpu_rf_N2844,
         j202_soc_core_j22_cpu_rf_N2843, j202_soc_core_j22_cpu_rf_N2842,
         j202_soc_core_j22_cpu_rf_N2840, j202_soc_core_j22_cpu_rf_N2839,
         j202_soc_core_j22_cpu_rf_N2838, j202_soc_core_j22_cpu_rf_N2837,
         j202_soc_core_j22_cpu_rf_N2836, j202_soc_core_j22_cpu_rf_N2835,
         j202_soc_core_j22_cpu_rf_N2834, j202_soc_core_j22_cpu_rf_N2832,
         j202_soc_core_j22_cpu_rf_N2831, j202_soc_core_j22_cpu_rf_N2830,
         j202_soc_core_j22_cpu_rf_N2829, j202_soc_core_j22_cpu_rf_N2828,
         j202_soc_core_j22_cpu_rf_N2827, j202_soc_core_j22_cpu_rf_N2826,
         j202_soc_core_j22_cpu_rf_N2824, j202_soc_core_j22_cpu_rf_N2823,
         j202_soc_core_j22_cpu_rf_N2822, j202_soc_core_j22_cpu_rf_N2821,
         j202_soc_core_j22_cpu_rf_N2820, j202_soc_core_j22_cpu_rf_N2819,
         j202_soc_core_j22_cpu_rf_N2818, j202_soc_core_j22_cpu_rf_N2817,
         j202_soc_core_j22_cpu_rf_N2816, j202_soc_core_j22_cpu_rf_N2815,
         j202_soc_core_j22_cpu_rf_N2814, j202_soc_core_j22_cpu_rf_N2813,
         j202_soc_core_j22_cpu_rf_N2811, j202_soc_core_j22_cpu_rf_N2810,
         j202_soc_core_j22_cpu_rf_N2809, j202_soc_core_j22_cpu_rf_N2808,
         j202_soc_core_j22_cpu_rf_N2807, j202_soc_core_j22_cpu_rf_N2806,
         j202_soc_core_j22_cpu_rf_N2805, j202_soc_core_j22_cpu_rf_N2803,
         j202_soc_core_j22_cpu_rf_N2802, j202_soc_core_j22_cpu_rf_N2801,
         j202_soc_core_j22_cpu_rf_N2800, j202_soc_core_j22_cpu_rf_N2799,
         j202_soc_core_j22_cpu_rf_N2798, j202_soc_core_j22_cpu_rf_N2797,
         j202_soc_core_j22_cpu_rf_N2795, j202_soc_core_j22_cpu_rf_N2794,
         j202_soc_core_j22_cpu_rf_N2793, j202_soc_core_j22_cpu_rf_N2792,
         j202_soc_core_j22_cpu_rf_N2791, j202_soc_core_j22_cpu_rf_N2790,
         j202_soc_core_j22_cpu_rf_N2789, j202_soc_core_j22_cpu_rf_N2787,
         j202_soc_core_j22_cpu_rf_N2786, j202_soc_core_j22_cpu_rf_N2785,
         j202_soc_core_j22_cpu_rf_N2784, j202_soc_core_j22_cpu_rf_N2783,
         j202_soc_core_j22_cpu_rf_N2782, j202_soc_core_j22_cpu_rf_N2781,
         j202_soc_core_j22_cpu_rf_N2780, j202_soc_core_j22_cpu_rf_N2779,
         j202_soc_core_j22_cpu_rf_N2778, j202_soc_core_j22_cpu_rf_N2777,
         j202_soc_core_j22_cpu_rf_N2776, j202_soc_core_j22_cpu_rf_N2774,
         j202_soc_core_j22_cpu_rf_N2773, j202_soc_core_j22_cpu_rf_N2772,
         j202_soc_core_j22_cpu_rf_N2771, j202_soc_core_j22_cpu_rf_N2770,
         j202_soc_core_j22_cpu_rf_N2769, j202_soc_core_j22_cpu_rf_N2768,
         j202_soc_core_j22_cpu_rf_N2766, j202_soc_core_j22_cpu_rf_N2765,
         j202_soc_core_j22_cpu_rf_N2764, j202_soc_core_j22_cpu_rf_N2763,
         j202_soc_core_j22_cpu_rf_N2762, j202_soc_core_j22_cpu_rf_N2761,
         j202_soc_core_j22_cpu_rf_N2760, j202_soc_core_j22_cpu_rf_N2758,
         j202_soc_core_j22_cpu_rf_N2757, j202_soc_core_j22_cpu_rf_N2756,
         j202_soc_core_j22_cpu_rf_N2755, j202_soc_core_j22_cpu_rf_N2754,
         j202_soc_core_j22_cpu_rf_N2753, j202_soc_core_j22_cpu_rf_N2752,
         j202_soc_core_j22_cpu_rf_N2750, j202_soc_core_j22_cpu_rf_N2749,
         j202_soc_core_j22_cpu_rf_N2748, j202_soc_core_j22_cpu_rf_N2747,
         j202_soc_core_j22_cpu_rf_N2746, j202_soc_core_j22_cpu_rf_N2745,
         j202_soc_core_j22_cpu_rf_N2744, j202_soc_core_j22_cpu_rf_N2743,
         j202_soc_core_j22_cpu_rf_N2742, j202_soc_core_j22_cpu_rf_N2741,
         j202_soc_core_j22_cpu_rf_N2740, j202_soc_core_j22_cpu_rf_N2739,
         j202_soc_core_j22_cpu_rf_N2737, j202_soc_core_j22_cpu_rf_N2736,
         j202_soc_core_j22_cpu_rf_N2735, j202_soc_core_j22_cpu_rf_N2734,
         j202_soc_core_j22_cpu_rf_N2733, j202_soc_core_j22_cpu_rf_N2732,
         j202_soc_core_j22_cpu_rf_N2731, j202_soc_core_j22_cpu_rf_N2729,
         j202_soc_core_j22_cpu_rf_N2728, j202_soc_core_j22_cpu_rf_N2727,
         j202_soc_core_j22_cpu_rf_N2726, j202_soc_core_j22_cpu_rf_N2725,
         j202_soc_core_j22_cpu_rf_N2724, j202_soc_core_j22_cpu_rf_N2723,
         j202_soc_core_j22_cpu_rf_N2721, j202_soc_core_j22_cpu_rf_N2720,
         j202_soc_core_j22_cpu_rf_N2719, j202_soc_core_j22_cpu_rf_N2718,
         j202_soc_core_j22_cpu_rf_N2717, j202_soc_core_j22_cpu_rf_N2716,
         j202_soc_core_j22_cpu_rf_N2715, j202_soc_core_j22_cpu_rf_N2713,
         j202_soc_core_j22_cpu_rf_N2712, j202_soc_core_j22_cpu_rf_N2711,
         j202_soc_core_j22_cpu_rf_N2710, j202_soc_core_j22_cpu_rf_N2709,
         j202_soc_core_j22_cpu_rf_N2708, j202_soc_core_j22_cpu_rf_N2707,
         j202_soc_core_j22_cpu_rf_N2706, j202_soc_core_j22_cpu_rf_N2705,
         j202_soc_core_j22_cpu_rf_N2704, j202_soc_core_j22_cpu_rf_N2703,
         j202_soc_core_j22_cpu_rf_N2702, j202_soc_core_j22_cpu_rf_N2700,
         j202_soc_core_j22_cpu_rf_N2699, j202_soc_core_j22_cpu_rf_N2698,
         j202_soc_core_j22_cpu_rf_N2697, j202_soc_core_j22_cpu_rf_N2696,
         j202_soc_core_j22_cpu_rf_N2695, j202_soc_core_j22_cpu_rf_N2694,
         j202_soc_core_j22_cpu_rf_N2692, j202_soc_core_j22_cpu_rf_N2691,
         j202_soc_core_j22_cpu_rf_N2690, j202_soc_core_j22_cpu_rf_N2689,
         j202_soc_core_j22_cpu_rf_N2688, j202_soc_core_j22_cpu_rf_N2687,
         j202_soc_core_j22_cpu_rf_N2686, j202_soc_core_j22_cpu_rf_N2684,
         j202_soc_core_j22_cpu_rf_N2683, j202_soc_core_j22_cpu_rf_N2682,
         j202_soc_core_j22_cpu_rf_N2681, j202_soc_core_j22_cpu_rf_N2680,
         j202_soc_core_j22_cpu_rf_N2679, j202_soc_core_j22_cpu_rf_N2678,
         j202_soc_core_j22_cpu_rf_N2676, j202_soc_core_j22_cpu_rf_N2675,
         j202_soc_core_j22_cpu_rf_N2660, j202_soc_core_j22_cpu_rf_N2656,
         j202_soc_core_j22_cpu_rf_N2655, j202_soc_core_j22_cpu_rf_N2653,
         j202_soc_core_j22_cpu_rf_N2652, j202_soc_core_j22_cpu_rf_N2646,
         j202_soc_core_j22_cpu_rf_N2645, j202_soc_core_j22_cpu_rf_N2640,
         j202_soc_core_j22_cpu_rf_N2639, j202_soc_core_j22_cpu_rf_N2638,
         j202_soc_core_j22_cpu_rf_N2637, j202_soc_core_j22_cpu_rf_N2628,
         j202_soc_core_j22_cpu_rf_N2627, j202_soc_core_j22_cpu_rf_N2626,
         j202_soc_core_j22_cpu_rf_N2625, j202_soc_core_j22_cpu_rf_N329,
         j202_soc_core_j22_cpu_rf_N328, j202_soc_core_j22_cpu_rf_N327,
         j202_soc_core_j22_cpu_rf_N326, j202_soc_core_j22_cpu_rf_N325,
         j202_soc_core_j22_cpu_rf_N324, j202_soc_core_j22_cpu_rf_N323,
         j202_soc_core_j22_cpu_rf_N322, j202_soc_core_j22_cpu_rf_N321,
         j202_soc_core_j22_cpu_rf_N320, j202_soc_core_j22_cpu_rf_N319,
         j202_soc_core_j22_cpu_rf_N318, j202_soc_core_j22_cpu_rf_N317,
         j202_soc_core_j22_cpu_rf_N316, j202_soc_core_j22_cpu_rf_N315,
         j202_soc_core_j22_cpu_rf_N314, j202_soc_core_j22_cpu_rf_N313,
         j202_soc_core_j22_cpu_rf_N312, j202_soc_core_j22_cpu_rf_N311,
         j202_soc_core_j22_cpu_rf_N310, j202_soc_core_j22_cpu_rf_N309,
         j202_soc_core_j22_cpu_rf_N308, j202_soc_core_j22_cpu_rf_N307,
         j202_soc_core_j22_cpu_rf_N306, j202_soc_core_j22_cpu_rf_N305,
         j202_soc_core_j22_cpu_rf_N304, j202_soc_core_j22_cpu_rf_N303,
         j202_soc_core_j22_cpu_rf_N302, j202_soc_core_j22_cpu_rf_N301,
         j202_soc_core_j22_cpu_rf_N300, j202_soc_core_j22_cpu_rf_N299,
         j202_soc_core_j22_cpu_rf_N298, j202_soc_core_j22_cpu_ma_N56,
         j202_soc_core_j22_cpu_ma_N55, j202_soc_core_j22_cpu_ma_N54,
         j202_soc_core_j22_cpu_ma_N53, j202_soc_core_j22_cpu_ml_N429,
         j202_soc_core_j22_cpu_ml_N427, j202_soc_core_j22_cpu_ml_N426,
         j202_soc_core_j22_cpu_ml_N425, j202_soc_core_j22_cpu_ml_N424,
         j202_soc_core_j22_cpu_ml_N423, j202_soc_core_j22_cpu_ml_N422,
         j202_soc_core_j22_cpu_ml_N421, j202_soc_core_j22_cpu_ml_N420,
         j202_soc_core_j22_cpu_ml_N419, j202_soc_core_j22_cpu_ml_N418,
         j202_soc_core_j22_cpu_ml_N417, j202_soc_core_j22_cpu_ml_N416,
         j202_soc_core_j22_cpu_ml_N415, j202_soc_core_j22_cpu_ml_N414,
         j202_soc_core_j22_cpu_ml_N413, j202_soc_core_j22_cpu_ml_N412,
         j202_soc_core_j22_cpu_ml_N370, j202_soc_core_j22_cpu_ml_N369,
         j202_soc_core_j22_cpu_ml_N368, j202_soc_core_j22_cpu_ml_N367,
         j202_soc_core_j22_cpu_ml_N366, j202_soc_core_j22_cpu_ml_N365,
         j202_soc_core_j22_cpu_ml_N364, j202_soc_core_j22_cpu_ml_N363,
         j202_soc_core_j22_cpu_ml_N362, j202_soc_core_j22_cpu_ml_N361,
         j202_soc_core_j22_cpu_ml_N360, j202_soc_core_j22_cpu_ml_N359,
         j202_soc_core_j22_cpu_ml_N357, j202_soc_core_j22_cpu_ml_N356,
         j202_soc_core_j22_cpu_ml_N355, j202_soc_core_j22_cpu_ml_N354,
         j202_soc_core_j22_cpu_ml_N336, j202_soc_core_j22_cpu_ml_N335,
         j202_soc_core_j22_cpu_ml_N334, j202_soc_core_j22_cpu_ml_N333,
         j202_soc_core_j22_cpu_ml_N332, j202_soc_core_j22_cpu_ml_N331,
         j202_soc_core_j22_cpu_ml_N330, j202_soc_core_j22_cpu_ml_N329,
         j202_soc_core_j22_cpu_ml_N328, j202_soc_core_j22_cpu_ml_N327,
         j202_soc_core_j22_cpu_ml_N326, j202_soc_core_j22_cpu_ml_N325,
         j202_soc_core_j22_cpu_ml_N324, j202_soc_core_j22_cpu_ml_N323,
         j202_soc_core_j22_cpu_ml_N322, j202_soc_core_j22_cpu_ml_N321,
         j202_soc_core_j22_cpu_ml_N320, j202_soc_core_j22_cpu_ml_N319,
         j202_soc_core_j22_cpu_ml_N318, j202_soc_core_j22_cpu_ml_N317,
         j202_soc_core_j22_cpu_ml_N316, j202_soc_core_j22_cpu_ml_N315,
         j202_soc_core_j22_cpu_ml_N314, j202_soc_core_j22_cpu_ml_N313,
         j202_soc_core_j22_cpu_ml_N312, j202_soc_core_j22_cpu_ml_N311,
         j202_soc_core_j22_cpu_ml_N310, j202_soc_core_j22_cpu_ml_N309,
         j202_soc_core_j22_cpu_ml_N308, j202_soc_core_j22_cpu_ml_N307,
         j202_soc_core_j22_cpu_ml_N306, j202_soc_core_j22_cpu_ml_N305,
         j202_soc_core_j22_cpu_ml_N304, j202_soc_core_j22_cpu_ml_N303,
         j202_soc_core_j22_cpu_ml_N195, j202_soc_core_j22_cpu_ml_N194,
         j202_soc_core_j22_cpu_ml_N193, j202_soc_core_j22_cpu_ml_N192,
         j202_soc_core_j22_cpu_ml_N191, j202_soc_core_j22_cpu_ml_N156,
         j202_soc_core_j22_cpu_ml_N155, j202_soc_core_j22_cpu_ml_N154,
         j202_soc_core_j22_cpu_ml_N153, j202_soc_core_j22_cpu_ml_N152,
         j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_N497,
         j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_N487,
         j202_soc_core_ahb2apb_00_N143, j202_soc_core_ahb2apb_00_N142,
         j202_soc_core_ahb2apb_00_N141, j202_soc_core_ahb2apb_00_N140,
         j202_soc_core_ahb2apb_00_N139, j202_soc_core_ahb2apb_00_N138,
         j202_soc_core_ahb2apb_00_N137, j202_soc_core_ahb2apb_00_N136,
         j202_soc_core_ahb2apb_00_N135, j202_soc_core_ahb2apb_00_N134,
         j202_soc_core_ahb2apb_00_N133, j202_soc_core_ahb2apb_00_N132,
         j202_soc_core_ahb2apb_00_N131, j202_soc_core_ahb2apb_00_N130,
         j202_soc_core_ahb2apb_00_N129, j202_soc_core_ahb2apb_00_N128,
         j202_soc_core_ahb2apb_00_N127, j202_soc_core_ahb2apb_00_N91,
         j202_soc_core_ahb2apb_00_N90, j202_soc_core_ahb2apb_00_N89,
         j202_soc_core_ahb2apb_00_N55, j202_soc_core_ahb2apb_00_N30,
         j202_soc_core_ahb2apb_00_N29, j202_soc_core_ahb2apb_00_N28,
         j202_soc_core_ahb2apb_00_N27, j202_soc_core_ahb2apb_00_N26,
         j202_soc_core_ahb2apb_00_N25, j202_soc_core_ahb2apb_00_N24,
         j202_soc_core_ahb2apb_00_N23, j202_soc_core_ahb2apb_00_N22,
         j202_soc_core_cmt_core_00_cmf1, j202_soc_core_cmt_core_00_cmf0,
         j202_soc_core_cmt_core_00_str1, j202_soc_core_cmt_core_00_str0,
         j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_2,
         j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_1,
         j202_soc_core_cmt_core_00_cmt_apb_00_nxt_state_0_,
         j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen,
         j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_nxt_latch_status_0_,
         j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_0_,
         j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_nxt_latch_status_0_,
         j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_0_,
         j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt1_to1,
         j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt0_to1,
         j202_soc_core_ahb2apb_01_N159, j202_soc_core_ahb2apb_01_N158,
         j202_soc_core_ahb2apb_01_N157, j202_soc_core_ahb2apb_01_N156,
         j202_soc_core_ahb2apb_01_N155, j202_soc_core_ahb2apb_01_N154,
         j202_soc_core_ahb2apb_01_N153, j202_soc_core_ahb2apb_01_N152,
         j202_soc_core_ahb2apb_01_N151, j202_soc_core_ahb2apb_01_N150,
         j202_soc_core_ahb2apb_01_N149, j202_soc_core_ahb2apb_01_N148,
         j202_soc_core_ahb2apb_01_N147, j202_soc_core_ahb2apb_01_N146,
         j202_soc_core_ahb2apb_01_N145, j202_soc_core_ahb2apb_01_N144,
         j202_soc_core_ahb2apb_01_N143, j202_soc_core_ahb2apb_01_N142,
         j202_soc_core_ahb2apb_01_N141, j202_soc_core_ahb2apb_01_N140,
         j202_soc_core_ahb2apb_01_N139, j202_soc_core_ahb2apb_01_N138,
         j202_soc_core_ahb2apb_01_N137, j202_soc_core_ahb2apb_01_N136,
         j202_soc_core_ahb2apb_01_N135, j202_soc_core_ahb2apb_01_N134,
         j202_soc_core_ahb2apb_01_N133, j202_soc_core_ahb2apb_01_N132,
         j202_soc_core_ahb2apb_01_N131, j202_soc_core_ahb2apb_01_N130,
         j202_soc_core_ahb2apb_01_N129, j202_soc_core_ahb2apb_01_N128,
         j202_soc_core_ahb2apb_01_N123, j202_soc_core_ahb2apb_01_N22,
         j202_soc_core_intc_core_00_cp_intack_all_0_,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_0__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_1__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_2__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_3__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_4__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_5__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_6__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_7__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_8__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_9__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_10__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_11__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_12__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_13__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_14__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_sint_label_15__rg_sint_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N23,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N22,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N21,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N20,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N19,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N18,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N17,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N16,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N15,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N14,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N13,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N12,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N11,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N10,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N9,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N8,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N7,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N6,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N5,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N4,
         j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N3,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N34,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N33,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N32,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N31,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N30,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N29,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N28,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N27,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N26,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N25,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N24,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N23,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N22,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N21,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N20,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N19,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N18,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N17,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N16,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N15,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N14,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N13,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N12,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N11,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N10,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N9,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N8,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N7,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N6,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N5,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N4,
         j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N3,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N23,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N22,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N21,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N20,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N19,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N18,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N17,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N16,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N15,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N14,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N13,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N12,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N11,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N10,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N9,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N8,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N7,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N6,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N5,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N4,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N3,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N23,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N22,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N21,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N20,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N19,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N18,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N17,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N16,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N15,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N14,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N13,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N12,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N11,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N10,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N9,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N8,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N7,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N6,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N5,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N4,
         j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N3,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_req_N3,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N6,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N5,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N4,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N3,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N6,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N5,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N4,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N3,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N9,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N7,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N6,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N5,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N4,
         j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N3,
         j202_soc_core_ahb2apb_02_N159, j202_soc_core_ahb2apb_02_N158,
         j202_soc_core_ahb2apb_02_N157, j202_soc_core_ahb2apb_02_N156,
         j202_soc_core_ahb2apb_02_N155, j202_soc_core_ahb2apb_02_N154,
         j202_soc_core_ahb2apb_02_N153, j202_soc_core_ahb2apb_02_N152,
         j202_soc_core_ahb2apb_02_N151, j202_soc_core_ahb2apb_02_N150,
         j202_soc_core_ahb2apb_02_N149, j202_soc_core_ahb2apb_02_N148,
         j202_soc_core_ahb2apb_02_N147, j202_soc_core_ahb2apb_02_N146,
         j202_soc_core_ahb2apb_02_N145, j202_soc_core_ahb2apb_02_N144,
         j202_soc_core_ahb2apb_02_N143, j202_soc_core_ahb2apb_02_N142,
         j202_soc_core_ahb2apb_02_N141, j202_soc_core_ahb2apb_02_N140,
         j202_soc_core_ahb2apb_02_N139, j202_soc_core_ahb2apb_02_N138,
         j202_soc_core_ahb2apb_02_N137, j202_soc_core_ahb2apb_02_N136,
         j202_soc_core_ahb2apb_02_N135, j202_soc_core_ahb2apb_02_N134,
         j202_soc_core_ahb2apb_02_N133, j202_soc_core_ahb2apb_02_N132,
         j202_soc_core_ahb2apb_02_N131, j202_soc_core_ahb2apb_02_N130,
         j202_soc_core_ahb2apb_02_N129, j202_soc_core_ahb2apb_02_N128,
         j202_soc_core_ahb2apb_02_N123, j202_soc_core_ahb2apb_02_N22,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N34,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N33,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N32,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N31,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N30,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N29,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N28,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N27,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N26,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N25,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N24,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N23,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N22,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N21,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N20,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N19,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N18,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N17,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N16,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N15,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N14,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N13,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N12,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N11,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N10,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N9,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N8,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N7,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N6,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N5,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N4,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N3,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N34,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N33,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N32,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N31,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N30,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N29,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N28,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N27,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N26,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N25,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N24,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N23,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N22,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N21,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N20,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N19,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N18,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N17,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N16,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N15,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N14,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N13,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N12,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N11,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N10,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N9,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N8,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N7,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N6,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N5,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N4,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N3,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N71,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N70,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N69,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N68,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N67,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N66,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N65,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N64,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N63,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N62,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N61,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N60,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N59,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N58,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N57,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N56,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N55,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N54,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N53,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N52,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N51,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N50,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N49,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N48,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N47,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N46,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N45,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N44,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N43,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N42,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N41,
         j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N40,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N34,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N33,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N32,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N31,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N30,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N29,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N28,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N27,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N26,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N25,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N24,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N23,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N22,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N21,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N20,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N19,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N18,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N17,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N16,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N15,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N14,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N13,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N12,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N11,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N10,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N9,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N8,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N7,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N6,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N5,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N4,
         j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N3,
         j202_soc_core_ahb2aqu_00_N164, j202_soc_core_ahb2aqu_00_N163,
         j202_soc_core_ahb2aqu_00_N161, j202_soc_core_ahb2aqu_00_N136,
         j202_soc_core_ahb2aqu_00_N135, j202_soc_core_ahb2aqu_00_N134,
         j202_soc_core_ahb2aqu_00_N133, j202_soc_core_ahb2aqu_00_N132,
         j202_soc_core_ahb2aqu_00_N131, j202_soc_core_ahb2aqu_00_N130,
         j202_soc_core_ahb2aqu_00_N129, j202_soc_core_ahb2aqu_00_N128,
         j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N98,
         j202_soc_core_ahb2aqu_00_N97, j202_soc_core_ahb2aqu_00_N95,
         j202_soc_core_ahb2aqu_00_N93, j202_soc_core_ahb2aqu_00_aqu_st_0_,
         j202_soc_core_uart_sio_ce_x4, j202_soc_core_uart_sio_ce,
         j202_soc_core_uart_RDRXD1, j202_soc_core_uart_WRTXD1,
         j202_soc_core_uart_N5, j202_soc_core_uart_TOP_N137,
         j202_soc_core_uart_TOP_N128, j202_soc_core_uart_TOP_N123,
         j202_soc_core_uart_TOP_N118, j202_soc_core_uart_TOP_rx_sio_ce_r2,
         j202_soc_core_uart_TOP_rx_sio_ce_r1, j202_soc_core_uart_TOP_N102,
         j202_soc_core_uart_TOP_N101, j202_soc_core_uart_TOP_change,
         j202_soc_core_uart_TOP_N95, j202_soc_core_uart_TOP_rx_valid_r,
         j202_soc_core_uart_TOP_rx_valid, j202_soc_core_uart_TOP_N89,
         j202_soc_core_uart_TOP_N88, j202_soc_core_uart_TOP_N87,
         j202_soc_core_uart_TOP_N86, j202_soc_core_uart_TOP_N85,
         j202_soc_core_uart_TOP_rx_sio_ce, j202_soc_core_uart_TOP_rx_go,
         j202_soc_core_uart_TOP_rxd_r, j202_soc_core_uart_TOP_rxd_s,
         j202_soc_core_uart_TOP_N61, j202_soc_core_uart_TOP_N60,
         j202_soc_core_uart_TOP_N59, j202_soc_core_uart_TOP_N58,
         j202_soc_core_uart_TOP_N57, j202_soc_core_uart_TOP_N43,
         j202_soc_core_uart_TOP_shift_en_r, j202_soc_core_uart_TOP_N33,
         j202_soc_core_uart_TOP_N32, j202_soc_core_uart_TOP_N31,
         j202_soc_core_uart_TOP_N30, j202_soc_core_uart_TOP_N29,
         j202_soc_core_uart_TOP_N28, j202_soc_core_uart_TOP_N27,
         j202_soc_core_uart_TOP_N26, j202_soc_core_uart_TOP_N25,
         j202_soc_core_uart_TOP_N24, j202_soc_core_uart_TOP_load,
         j202_soc_core_uart_TOP_shift_en, j202_soc_core_uart_TOP_N16,
         j202_soc_core_uart_TOP_txf_empty_r,
         j202_soc_core_uart_TOP_tx_fifo_N42,
         j202_soc_core_uart_TOP_tx_fifo_N41, j202_soc_core_uart_TOP_tx_fifo_gb,
         j202_soc_core_uart_TOP_tx_fifo_N32,
         j202_soc_core_uart_TOP_tx_fifo_N31,
         j202_soc_core_uart_TOP_tx_fifo_N30,
         j202_soc_core_uart_TOP_tx_fifo_N29,
         j202_soc_core_uart_TOP_rx_fifo_N42,
         j202_soc_core_uart_TOP_rx_fifo_N41, j202_soc_core_uart_TOP_rx_fifo_gb,
         j202_soc_core_uart_TOP_rx_fifo_N32,
         j202_soc_core_uart_TOP_rx_fifo_N31,
         j202_soc_core_uart_TOP_rx_fifo_N30,
         j202_soc_core_uart_TOP_rx_fifo_N29, j202_soc_core_uart_BRG_N59,
         j202_soc_core_uart_BRG_sio_ce_r, j202_soc_core_uart_BRG_N57,
         j202_soc_core_uart_BRG_N56, j202_soc_core_uart_BRG_N55,
         j202_soc_core_uart_BRG_sio_ce_x4_t,
         j202_soc_core_uart_BRG_sio_ce_x4_r, j202_soc_core_uart_BRG_N47,
         j202_soc_core_uart_BRG_N42, j202_soc_core_uart_BRG_N41,
         j202_soc_core_uart_BRG_N40, j202_soc_core_uart_BRG_N39,
         j202_soc_core_uart_BRG_N38, j202_soc_core_uart_BRG_N37,
         j202_soc_core_uart_BRG_N36, j202_soc_core_uart_BRG_N35,
         j202_soc_core_uart_BRG_br_clr, j202_soc_core_uart_BRG_N21,
         j202_soc_core_uart_BRG_N19, j202_soc_core_uart_BRG_N18,
         j202_soc_core_uart_BRG_N17, j202_soc_core_uart_BRG_N16,
         j202_soc_core_uart_BRG_N15, j202_soc_core_uart_BRG_N14,
         j202_soc_core_uart_BRG_N13, j202_soc_core_uart_BRG_N12,
         j202_soc_core_uart_BRG_ps_clr, j202_soc_core_bldc_core_00_adc_en,
         j202_soc_core_bldc_core_00_pwm_en,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_nxt_bldc_int,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_0_,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_wen,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_nxt_latch_status_0_,
         j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_0_,
         j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_2,
         j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1,
         j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posc,
         j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_negb,
         j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posb,
         j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posa,
         j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld,
         j202_soc_core_ahb2wbqspi_00_stb_o, j202_soc_core_wbqspiflash_00_N755,
         j202_soc_core_wbqspiflash_00_N752, j202_soc_core_wbqspiflash_00_N751,
         j202_soc_core_wbqspiflash_00_N750, j202_soc_core_wbqspiflash_00_N749,
         j202_soc_core_wbqspiflash_00_N748, j202_soc_core_wbqspiflash_00_N747,
         j202_soc_core_wbqspiflash_00_N746, j202_soc_core_wbqspiflash_00_N745,
         j202_soc_core_wbqspiflash_00_N744, j202_soc_core_wbqspiflash_00_N743,
         j202_soc_core_wbqspiflash_00_N742, j202_soc_core_wbqspiflash_00_N741,
         j202_soc_core_wbqspiflash_00_N740, j202_soc_core_wbqspiflash_00_N739,
         j202_soc_core_wbqspiflash_00_N738, j202_soc_core_wbqspiflash_00_N737,
         j202_soc_core_wbqspiflash_00_N736, j202_soc_core_wbqspiflash_00_N735,
         j202_soc_core_wbqspiflash_00_N734, j202_soc_core_wbqspiflash_00_N733,
         j202_soc_core_wbqspiflash_00_N730, j202_soc_core_wbqspiflash_00_N729,
         j202_soc_core_wbqspiflash_00_N728, j202_soc_core_wbqspiflash_00_N727,
         j202_soc_core_wbqspiflash_00_N726, j202_soc_core_wbqspiflash_00_N725,
         j202_soc_core_wbqspiflash_00_N724, j202_soc_core_wbqspiflash_00_N723,
         j202_soc_core_wbqspiflash_00_N722, j202_soc_core_wbqspiflash_00_N721,
         j202_soc_core_wbqspiflash_00_N720, j202_soc_core_wbqspiflash_00_N719,
         j202_soc_core_wbqspiflash_00_N718, j202_soc_core_wbqspiflash_00_N717,
         j202_soc_core_wbqspiflash_00_N716, j202_soc_core_wbqspiflash_00_N715,
         j202_soc_core_wbqspiflash_00_N714, j202_soc_core_wbqspiflash_00_N713,
         j202_soc_core_wbqspiflash_00_N712, j202_soc_core_wbqspiflash_00_N711,
         j202_soc_core_wbqspiflash_00_N710, j202_soc_core_wbqspiflash_00_N709,
         j202_soc_core_wbqspiflash_00_N708, j202_soc_core_wbqspiflash_00_N698,
         j202_soc_core_wbqspiflash_00_N697, j202_soc_core_wbqspiflash_00_N696,
         j202_soc_core_wbqspiflash_00_N695, j202_soc_core_wbqspiflash_00_N694,
         j202_soc_core_wbqspiflash_00_N693, j202_soc_core_wbqspiflash_00_N692,
         j202_soc_core_wbqspiflash_00_N691, j202_soc_core_wbqspiflash_00_N690,
         j202_soc_core_wbqspiflash_00_N689, j202_soc_core_wbqspiflash_00_N688,
         j202_soc_core_wbqspiflash_00_N687, j202_soc_core_wbqspiflash_00_N686,
         j202_soc_core_wbqspiflash_00_N685, j202_soc_core_wbqspiflash_00_N684,
         j202_soc_core_wbqspiflash_00_N683, j202_soc_core_wbqspiflash_00_N682,
         j202_soc_core_wbqspiflash_00_N681, j202_soc_core_wbqspiflash_00_N680,
         j202_soc_core_wbqspiflash_00_N679, j202_soc_core_wbqspiflash_00_N678,
         j202_soc_core_wbqspiflash_00_N677, j202_soc_core_wbqspiflash_00_N676,
         j202_soc_core_wbqspiflash_00_N675, j202_soc_core_wbqspiflash_00_N674,
         j202_soc_core_wbqspiflash_00_N673, j202_soc_core_wbqspiflash_00_N672,
         j202_soc_core_wbqspiflash_00_N671, j202_soc_core_wbqspiflash_00_N670,
         j202_soc_core_wbqspiflash_00_N669, j202_soc_core_wbqspiflash_00_N668,
         j202_soc_core_wbqspiflash_00_N667, j202_soc_core_wbqspiflash_00_N663,
         j202_soc_core_wbqspiflash_00_N629, j202_soc_core_wbqspiflash_00_N628,
         j202_soc_core_wbqspiflash_00_N623, j202_soc_core_wbqspiflash_00_N622,
         j202_soc_core_wbqspiflash_00_N621, j202_soc_core_wbqspiflash_00_N620,
         j202_soc_core_wbqspiflash_00_N619, j202_soc_core_wbqspiflash_00_N618,
         j202_soc_core_wbqspiflash_00_N617, j202_soc_core_wbqspiflash_00_N616,
         j202_soc_core_wbqspiflash_00_N615, j202_soc_core_wbqspiflash_00_N614,
         j202_soc_core_wbqspiflash_00_N613, j202_soc_core_wbqspiflash_00_N612,
         j202_soc_core_wbqspiflash_00_N611, j202_soc_core_wbqspiflash_00_N609,
         j202_soc_core_wbqspiflash_00_N608, j202_soc_core_wbqspiflash_00_N607,
         j202_soc_core_wbqspiflash_00_N606, j202_soc_core_wbqspiflash_00_N605,
         j202_soc_core_wbqspiflash_00_N594, j202_soc_core_wbqspiflash_00_N592,
         j202_soc_core_wbqspiflash_00_N590,
         j202_soc_core_wbqspiflash_00_spif_cmd,
         j202_soc_core_wbqspiflash_00_spif_req,
         j202_soc_core_wbqspiflash_00_N86,
         j202_soc_core_wbqspiflash_00_alt_ctrl,
         j202_soc_core_wbqspiflash_00_N85,
         j202_soc_core_wbqspiflash_00_alt_cmd,
         j202_soc_core_wbqspiflash_00_spif_ctrl,
         j202_soc_core_wbqspiflash_00_spif_override,
         j202_soc_core_wbqspiflash_00_quad_mode_enabled,
         j202_soc_core_wbqspiflash_00_write_protect,
         j202_soc_core_wbqspiflash_00_dirty_sector,
         j202_soc_core_wbqspiflash_00_write_in_progress,
         j202_soc_core_wbqspiflash_00_w_qspi_cs_n,
         j202_soc_core_wbqspiflash_00_w_qspi_sck,
         j202_soc_core_wbqspiflash_00_spi_busy,
         j202_soc_core_wbqspiflash_00_spi_valid,
         j202_soc_core_wbqspiflash_00_spi_dir,
         j202_soc_core_wbqspiflash_00_spi_spd,
         j202_soc_core_wbqspiflash_00_spi_hold,
         j202_soc_core_wbqspiflash_00_spi_wr,
         j202_soc_core_wbqspiflash_00_lldriver_N430,
         j202_soc_core_wbqspiflash_00_lldriver_N429,
         j202_soc_core_wbqspiflash_00_lldriver_N428,
         j202_soc_core_wbqspiflash_00_lldriver_N427,
         j202_soc_core_wbqspiflash_00_lldriver_N426,
         j202_soc_core_wbqspiflash_00_lldriver_N425,
         j202_soc_core_wbqspiflash_00_lldriver_N424,
         j202_soc_core_wbqspiflash_00_lldriver_N423,
         j202_soc_core_wbqspiflash_00_lldriver_N422,
         j202_soc_core_wbqspiflash_00_lldriver_N421,
         j202_soc_core_wbqspiflash_00_lldriver_N420,
         j202_soc_core_wbqspiflash_00_lldriver_N419,
         j202_soc_core_wbqspiflash_00_lldriver_N418,
         j202_soc_core_wbqspiflash_00_lldriver_N417,
         j202_soc_core_wbqspiflash_00_lldriver_N416,
         j202_soc_core_wbqspiflash_00_lldriver_N415,
         j202_soc_core_wbqspiflash_00_lldriver_N414,
         j202_soc_core_wbqspiflash_00_lldriver_N413,
         j202_soc_core_wbqspiflash_00_lldriver_N412,
         j202_soc_core_wbqspiflash_00_lldriver_N411,
         j202_soc_core_wbqspiflash_00_lldriver_N410,
         j202_soc_core_wbqspiflash_00_lldriver_N409,
         j202_soc_core_wbqspiflash_00_lldriver_N408,
         j202_soc_core_wbqspiflash_00_lldriver_N407,
         j202_soc_core_wbqspiflash_00_lldriver_N406,
         j202_soc_core_wbqspiflash_00_lldriver_N405,
         j202_soc_core_wbqspiflash_00_lldriver_N404,
         j202_soc_core_wbqspiflash_00_lldriver_N403,
         j202_soc_core_wbqspiflash_00_lldriver_N402,
         j202_soc_core_wbqspiflash_00_lldriver_N401,
         j202_soc_core_wbqspiflash_00_lldriver_N400,
         j202_soc_core_wbqspiflash_00_lldriver_N399,
         j202_soc_core_wbqspiflash_00_lldriver_N398,
         j202_soc_core_wbqspiflash_00_lldriver_N397,
         j202_soc_core_wbqspiflash_00_lldriver_N396,
         j202_soc_core_wbqspiflash_00_lldriver_N395,
         j202_soc_core_wbqspiflash_00_lldriver_N394,
         j202_soc_core_wbqspiflash_00_lldriver_N393,
         j202_soc_core_wbqspiflash_00_lldriver_N392,
         j202_soc_core_wbqspiflash_00_lldriver_N391,
         j202_soc_core_wbqspiflash_00_lldriver_N389,
         j202_soc_core_wbqspiflash_00_lldriver_N388,
         j202_soc_core_wbqspiflash_00_lldriver_N387,
         j202_soc_core_wbqspiflash_00_lldriver_N386,
         j202_soc_core_wbqspiflash_00_lldriver_N385,
         j202_soc_core_wbqspiflash_00_lldriver_N384,
         j202_soc_core_wbqspiflash_00_lldriver_N383,
         j202_soc_core_wbqspiflash_00_lldriver_N382,
         j202_soc_core_wbqspiflash_00_lldriver_N381,
         j202_soc_core_wbqspiflash_00_lldriver_N380,
         j202_soc_core_wbqspiflash_00_lldriver_N379,
         j202_soc_core_wbqspiflash_00_lldriver_N378,
         j202_soc_core_wbqspiflash_00_lldriver_N377,
         j202_soc_core_wbqspiflash_00_lldriver_N376,
         j202_soc_core_wbqspiflash_00_lldriver_N375,
         j202_soc_core_wbqspiflash_00_lldriver_N374,
         j202_soc_core_wbqspiflash_00_lldriver_N373,
         j202_soc_core_wbqspiflash_00_lldriver_N372,
         j202_soc_core_wbqspiflash_00_lldriver_N371,
         j202_soc_core_wbqspiflash_00_lldriver_N370,
         j202_soc_core_wbqspiflash_00_lldriver_N369,
         j202_soc_core_wbqspiflash_00_lldriver_N368,
         j202_soc_core_wbqspiflash_00_lldriver_N367,
         j202_soc_core_wbqspiflash_00_lldriver_N366,
         j202_soc_core_wbqspiflash_00_lldriver_N365,
         j202_soc_core_wbqspiflash_00_lldriver_N364,
         j202_soc_core_wbqspiflash_00_lldriver_N363,
         j202_soc_core_wbqspiflash_00_lldriver_N362,
         j202_soc_core_wbqspiflash_00_lldriver_N361,
         j202_soc_core_wbqspiflash_00_lldriver_N360,
         j202_soc_core_wbqspiflash_00_lldriver_N359,
         j202_soc_core_wbqspiflash_00_lldriver_N358,
         j202_soc_core_wbqspiflash_00_lldriver_N356,
         j202_soc_core_wbqspiflash_00_lldriver_N355,
         j202_soc_core_wbqspiflash_00_lldriver_N354,
         j202_soc_core_wbqspiflash_00_lldriver_N353,
         j202_soc_core_wbqspiflash_00_lldriver_N352,
         j202_soc_core_wbqspiflash_00_lldriver_N351,
         j202_soc_core_wbqspiflash_00_lldriver_N350,
         j202_soc_core_wbqspiflash_00_lldriver_N349,
         j202_soc_core_wbqspiflash_00_lldriver_N348,
         j202_soc_core_wbqspiflash_00_lldriver_N347,
         j202_soc_core_wbqspiflash_00_lldriver_N346,
         j202_soc_core_wbqspiflash_00_lldriver_N345,
         j202_soc_core_wbqspiflash_00_lldriver_N344,
         j202_soc_core_wbqspiflash_00_lldriver_N343,
         j202_soc_core_wbqspiflash_00_lldriver_N342,
         j202_soc_core_wbqspiflash_00_lldriver_N341,
         j202_soc_core_wbqspiflash_00_lldriver_N340,
         j202_soc_core_wbqspiflash_00_lldriver_N339,
         j202_soc_core_wbqspiflash_00_lldriver_N338,
         j202_soc_core_wbqspiflash_00_lldriver_N337,
         j202_soc_core_wbqspiflash_00_lldriver_N336,
         j202_soc_core_wbqspiflash_00_lldriver_N335,
         j202_soc_core_wbqspiflash_00_lldriver_N334,
         j202_soc_core_wbqspiflash_00_lldriver_N333,
         j202_soc_core_wbqspiflash_00_lldriver_N332,
         j202_soc_core_wbqspiflash_00_lldriver_N331,
         j202_soc_core_wbqspiflash_00_lldriver_N330,
         j202_soc_core_wbqspiflash_00_lldriver_N329,
         j202_soc_core_wbqspiflash_00_lldriver_N328,
         j202_soc_core_wbqspiflash_00_lldriver_N327,
         j202_soc_core_wbqspiflash_00_lldriver_N326,
         j202_soc_core_wbqspiflash_00_lldriver_N325,
         j202_soc_core_wbqspiflash_00_lldriver_N324,
         j202_soc_core_wbqspiflash_00_lldriver_N323,
         j202_soc_core_wbqspiflash_00_lldriver_N321,
         j202_soc_core_wbqspiflash_00_lldriver_N319,
         j202_soc_core_wbqspiflash_00_lldriver_N318,
         j202_soc_core_wbqspiflash_00_lldriver_N317,
         j202_soc_core_wbqspiflash_00_lldriver_N316,
         j202_soc_core_wbqspiflash_00_lldriver_N315,
         j202_soc_core_wbqspiflash_00_lldriver_N314,
         j202_soc_core_wbqspiflash_00_lldriver_N313,
         j202_soc_core_wbqspiflash_00_lldriver_N312,
         j202_soc_core_wbqspiflash_00_lldriver_N311,
         j202_soc_core_wbqspiflash_00_lldriver_N310,
         j202_soc_core_wbqspiflash_00_lldriver_N308,
         j202_soc_core_wbqspiflash_00_lldriver_N307,
         j202_soc_core_wbqspiflash_00_lldriver_r_dir,
         j202_soc_core_wbqspiflash_00_lldriver_r_spd,
         j202_soc_core_bootrom_00_sel_w, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10558, n10559, n10560, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10602, n10603, n10604, n10605,
         n10670, n10671, n10672, n10673, n10675, n10676, n10742, n10743,
         n10744, n10745, n10901, n10902, n10903, n10904, n10908,
         DP_OP_1501J1_126_8405_n3, DP_OP_1501J1_126_8405_n4,
         U7_RSOP_1488_C3_DATA3_2, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10974, n10976, n10978, n10979, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10999, n11000, n11001, n11002, n11004, n11005, n11006, n11007,
         n11009, n11010, n11011, n11012, n11014, n11015, n11016, n11017,
         n11019, n11020, n11021, n11022, n11024, n11025, n11026, n11027,
         n11029, n11030, n11031, n11032, n11034, n11035, n11036, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
         n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183,
         n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191,
         n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
         n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207,
         n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
         n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
         n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231,
         n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
         n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
         n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255,
         n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
         n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279,
         n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287,
         n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295,
         n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303,
         n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311,
         n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319,
         n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327,
         n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335,
         n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
         n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351,
         n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359,
         n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
         n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
         n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383,
         n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
         n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399,
         n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
         n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
         n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423,
         n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
         n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
         n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447,
         n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455,
         n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463,
         n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471,
         n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479,
         n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
         n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495,
         n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503,
         n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
         n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519,
         n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527,
         n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535,
         n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543,
         n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551,
         n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
         n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
         n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
         n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
         n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591,
         n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
         n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607,
         n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615,
         n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
         n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
         n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639,
         n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647,
         n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655,
         n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663,
         n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
         n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
         n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
         n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
         n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
         n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711,
         n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719,
         n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
         n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
         n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
         n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
         n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759,
         n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
         n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
         n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
         n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
         n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
         n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807,
         n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
         n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
         n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831,
         n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
         n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
         n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855,
         n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863,
         n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
         n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879,
         n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
         n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
         n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
         n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
         n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
         n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
         n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
         n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
         n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
         n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
         n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999,
         n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
         n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
         n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
         n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
         n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
         n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
         n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
         n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
         n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071,
         n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
         n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
         n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095,
         n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
         n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111,
         n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119,
         n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
         n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
         n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143,
         n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151,
         n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
         n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167,
         n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
         n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183,
         n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
         n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
         n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
         n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215,
         n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223,
         n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
         n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239,
         n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247,
         n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255,
         n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263,
         n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271,
         n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
         n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287,
         n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295,
         n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
         n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311,
         n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
         n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
         n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
         n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343,
         n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
         n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359,
         n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367,
         n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375,
         n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383,
         n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391,
         n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399,
         n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
         n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415,
         n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423,
         n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431,
         n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439,
         n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
         n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455,
         n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463,
         n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
         n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479,
         n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487,
         n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495,
         n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503,
         n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511,
         n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519,
         n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527,
         n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535,
         n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543,
         n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551,
         n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559,
         n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567,
         n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575,
         n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583,
         n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591,
         n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599,
         n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607,
         n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615,
         n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623,
         n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631,
         n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639,
         n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647,
         n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655,
         n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663,
         n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671,
         n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679,
         n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687,
         n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695,
         n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703,
         n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711,
         n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719,
         n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727,
         n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735,
         n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743,
         n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751,
         n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759,
         n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767,
         n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775,
         n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783,
         n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791,
         n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799,
         n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807,
         n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815,
         n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823,
         n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831,
         n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839,
         n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847,
         n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855,
         n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863,
         n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871,
         n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879,
         n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887,
         n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895,
         n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903,
         n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911,
         n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919,
         n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927,
         n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935,
         n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943,
         n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951,
         n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959,
         n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967,
         n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975,
         n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983,
         n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991,
         n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999,
         n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007,
         n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015,
         n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023,
         n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031,
         n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039,
         n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047,
         n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055,
         n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063,
         n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071,
         n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079,
         n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087,
         n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095,
         n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103,
         n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111,
         n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119,
         n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127,
         n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135,
         n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143,
         n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151,
         n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159,
         n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167,
         n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175,
         n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183,
         n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191,
         n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199,
         n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207,
         n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215,
         n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223,
         n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231,
         n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239,
         n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247,
         n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255,
         n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263,
         n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271,
         n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279,
         n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287,
         n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295,
         n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303,
         n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311,
         n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319,
         n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327,
         n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335,
         n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343,
         n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351,
         n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359,
         n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367,
         n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375,
         n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383,
         n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391,
         n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399,
         n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407,
         n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415,
         n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423,
         n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431,
         n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439,
         n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447,
         n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455,
         n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463,
         n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471,
         n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479,
         n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487,
         n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495,
         n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503,
         n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511,
         n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519,
         n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527,
         n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535,
         n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543,
         n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551,
         n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559,
         n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567,
         n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575,
         n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583,
         n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591,
         n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599,
         n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607,
         n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615,
         n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623,
         n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631,
         n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639,
         n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647,
         n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655,
         n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663,
         n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671,
         n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679,
         n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687,
         n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695,
         n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703,
         n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711,
         n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719,
         n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727,
         n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735,
         n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743,
         n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751,
         n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759,
         n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767,
         n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775,
         n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783,
         n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791,
         n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799,
         n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807,
         n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815,
         n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823,
         n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831,
         n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839,
         n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847,
         n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855,
         n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863,
         n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871,
         n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879,
         n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887,
         n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895,
         n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903,
         n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911,
         n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919,
         n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927,
         n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935,
         n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943,
         n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951,
         n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959,
         n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967,
         n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975,
         n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983,
         n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991,
         n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999,
         n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007,
         n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015,
         n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023,
         n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031,
         n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039,
         n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047,
         n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055,
         n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063,
         n24064, n24065, n24067, n24068, n24069, n24070, n24071, n24072,
         n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080,
         n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088,
         n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096,
         n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104,
         n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112,
         n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120,
         n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128,
         n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136,
         n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144,
         n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152,
         n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160,
         n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168,
         n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176,
         n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184,
         n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192,
         n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200,
         n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208,
         n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216,
         n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224,
         n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232,
         n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240,
         n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248,
         n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256,
         n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264,
         n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272,
         n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280,
         n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288,
         n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296,
         n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304,
         n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312,
         n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320,
         n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328,
         n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336,
         n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344,
         n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352,
         n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360,
         n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368,
         n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376,
         n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384,
         n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392,
         n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400,
         n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408,
         n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416,
         n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424,
         n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432,
         n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440,
         n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448,
         n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456,
         n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464,
         n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472,
         n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480,
         n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488,
         n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496,
         n24497, n24498, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24823, n24824, n24825, n24826,
         n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834,
         n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842,
         n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850,
         n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858,
         n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866,
         n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874,
         n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882,
         n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890,
         n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898,
         n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906,
         n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914,
         n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922,
         n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930,
         n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938,
         n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946,
         n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954,
         n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962,
         n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970,
         n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978,
         n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986,
         n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994,
         n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002,
         n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010,
         n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018,
         n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026,
         n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034,
         n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042,
         n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050,
         n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058,
         n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066,
         n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074,
         n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082,
         n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090,
         n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098,
         n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106,
         n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114,
         n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122,
         n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130,
         n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138,
         n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146,
         n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154,
         n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162,
         n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170,
         n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178,
         n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186,
         n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194,
         n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202,
         n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
         n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218,
         n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226,
         n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
         n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242,
         n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
         n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
         n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
         n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274,
         n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
         n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290,
         n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
         n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
         n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314,
         n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322,
         n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
         n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338,
         n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346,
         n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
         n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362,
         n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
         n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378,
         n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386,
         n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394,
         n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
         n25403, n25404, n25405, n25406, n25427, n25428, n25429, n25430,
         n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438,
         n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446,
         n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454,
         n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462,
         n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470,
         n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478,
         n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486,
         n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494,
         n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502,
         n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510,
         n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518,
         n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526,
         n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534,
         n25535, n25536, n25537, n25541, n25542, n25543, n25544, n25545,
         n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675,
         n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683,
         n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
         n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
         n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
         n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
         n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
         n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731,
         n25732, n25733, n25734, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45,
         SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53,
         SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55,
         SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57,
         SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59,
         SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61,
         SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63,
         SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65,
         SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67,
         SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69,
         SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71,
         SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73,
         SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75,
         SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77,
         SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79,
         SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81,
         SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83,
         SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85,
         SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87,
         SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89,
         SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91,
         SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93,
         SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95,
         SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97,
         SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99,
         SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101,
         SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103,
         SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105,
         SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107,
         SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109,
         SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111,
         SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113,
         SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115,
         SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117,
         SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119,
         SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121,
         SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123,
         SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125,
         SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127,
         SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129,
         SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131,
         SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133,
         SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135,
         SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137,
         SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139,
         SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141,
         SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143,
         SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145,
         SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147,
         SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149,
         SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151,
         SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153,
         SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155,
         SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157,
         SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159,
         SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161,
         SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163,
         SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165,
         SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167,
         SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169,
         SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171,
         SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173,
         SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175,
         SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177,
         SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179,
         SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181,
         SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183,
         SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185,
         SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187,
         SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189,
         SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191,
         SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193,
         SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195,
         SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197,
         SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199,
         SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201,
         SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203,
         SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205,
         SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207,
         SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209,
         SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211,
         SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213,
         SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215,
         SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217,
         SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219,
         SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221,
         SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223,
         SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225,
         SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227,
         SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229,
         SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231,
         SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233,
         SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235,
         SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237,
         SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239,
         SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241,
         SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243,
         SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245,
         SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247,
         SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249,
         SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251,
         SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253,
         SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255,
         SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257,
         SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259,
         SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261,
         SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263,
         SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265,
         SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267,
         SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269,
         SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271,
         SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273,
         SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275,
         SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277,
         SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279,
         SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281,
         SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283,
         SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285,
         SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287,
         SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289,
         SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291,
         SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293,
         SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295,
         SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297,
         SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299,
         SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301,
         SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303,
         SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305,
         SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307,
         SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309,
         SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311,
         SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313,
         SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315,
         SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317,
         SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319,
         SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321,
         SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323,
         SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325,
         SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327,
         SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329,
         SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331,
         SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333,
         SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335,
         SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337,
         SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339,
         SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341,
         SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343,
         SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345,
         SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347,
         SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349,
         SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351,
         SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353,
         SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355,
         SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357,
         SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359,
         SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361,
         SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363,
         SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365,
         SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367,
         SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369,
         SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371,
         SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373,
         SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375,
         SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377,
         SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379,
         SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381,
         SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383,
         SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385,
         SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387,
         SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389,
         SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391,
         SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393,
         SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395,
         SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397,
         SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399,
         SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401,
         SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403,
         SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405,
         SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407,
         SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409,
         SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411,
         SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413,
         SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415,
         SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417,
         SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419,
         SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421,
         SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423,
         SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425,
         SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427,
         SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429,
         SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431,
         SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433,
         SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435,
         SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437,
         SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439,
         SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441,
         SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443,
         SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445,
         SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447,
         SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449,
         SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451,
         SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453,
         SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455,
         SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457,
         SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459,
         SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461,
         SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463,
         SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465,
         SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467,
         SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469,
         SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471,
         SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473,
         SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475,
         SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477,
         SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479,
         SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481,
         SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483,
         SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485,
         SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487,
         SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489,
         SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491,
         SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493,
         SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495,
         SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497,
         SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499,
         SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501,
         SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503,
         SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505,
         SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507,
         SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509,
         SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511,
         SYNOPSYS_UNCONNECTED_512;
  wire   [31:0] gpio_en_o;
  wire   [31:0] j202_soc_core_qspi_wb_wdat;
  wire   [24:2] j202_soc_core_qspi_wb_addr;
  wire   [15:0] j202_soc_core_prdata;
  wire   [7:0] j202_soc_core_paddr;
  wire   [7:0] j202_soc_core_pstrb;
  wire   [0:2] j202_soc_core_pwrite;
  wire   [5:0] j202_soc_core_j22_cpu_exuop_EXU_;
  wire   [4:0] j202_soc_core_j22_cpu_macop_MAC_;
  wire   [31:0] j202_soc_core_j22_cpu_pc;
  wire   [4:0] j202_soc_core_j22_cpu_opst;
  wire   [31:0] j202_soc_core_j22_cpu_rf_tmp;
  wire   [31:0] j202_soc_core_j22_cpu_rf_vbr;
  wire   [31:0] j202_soc_core_j22_cpu_rf_gbr;
  wire   [31:0] j202_soc_core_j22_cpu_rf_pr;
  wire   [511:0] j202_soc_core_j22_cpu_rf_gpr;
  wire   [1:0] j202_soc_core_j22_cpu_ma_M_address;
  wire   [1:0] j202_soc_core_j22_cpu_ma_M_area;
  wire   [3:0] j202_soc_core_j22_cpu_ma_M_MEM;
  wire   [31:0] j202_soc_core_j22_cpu_ml_maclj;
  wire   [31:0] j202_soc_core_j22_cpu_ml_machj;
  wire   [31:0] j202_soc_core_j22_cpu_ml_mach;
  wire   [31:0] j202_soc_core_j22_cpu_ml_macl;
  wire   [32:0] j202_soc_core_j22_cpu_ml_bufb;
  wire   [32:0] j202_soc_core_j22_cpu_ml_bufa;
  wire   [4:0] j202_soc_core_j22_cpu_ml_X_macop_MAC_;
  wire   [4:0] j202_soc_core_j22_cpu_ml_M_macop_MAC_;
  wire   [511:0] j202_soc_core_memory0_ram_dout0;
  wire   [15:0] j202_soc_core_memory0_ram_dout0_sel;
  wire   [111:0] j202_soc_core_ahblite_interconnect_s_hrdata;
  wire  
         [0:6] j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel
;
  wire   [2:0] j202_soc_core_ahb2apb_00_state;
  wire   [15:0] j202_soc_core_cmt_core_00_cnt1;
  wire   [15:0] j202_soc_core_cmt_core_00_cnt0;
  wire   [15:0] j202_soc_core_cmt_core_00_const1;
  wire   [15:0] j202_soc_core_cmt_core_00_const0;
  wire   [15:0] j202_soc_core_cmt_core_00_wdata_cnt0;
  wire   [1:0] j202_soc_core_cmt_core_00_cks1;
  wire   [1:0] j202_soc_core_cmt_core_00_cks0;
  wire   [7:0] j202_soc_core_cmt_core_00_reg_addr;
  wire   [1:0] j202_soc_core_cmt_core_00_cmt_apb_00_state;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata;
  wire   [6:2] j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1;
  wire   [6:2] j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1;
  wire   [9:0] j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1;
  wire   [9:0] j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1;
  wire   [15:0] j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0;
  wire   [9:0] j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0;
  wire   [9:0] j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0;
  wire   [2:0] j202_soc_core_ahb2apb_01_state;
  wire   [1:0] j202_soc_core_ahb2apb_01_hsize_buf;
  wire   [20:0] j202_soc_core_intc_core_00_in_intreq;
  wire   [127:0] j202_soc_core_intc_core_00_rg_ipr;
  wire   [127:0] j202_soc_core_intc_core_00_rg_itgt;
  wire   [20:0] j202_soc_core_intc_core_00_rg_irqc;
  wire   [31:0] j202_soc_core_intc_core_00_rg_ie;
  wire   [7:0] j202_soc_core_intc_core_00_rg_eimk;
  wire   [15:0] j202_soc_core_intc_core_00_rg_sint;
  wire   [11:0] j202_soc_core_intc_core_00_bs_addr;
  wire  
         [20:0] j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int
;
  wire  
         [6:0] j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch
;
  wire   [2:0] j202_soc_core_ahb2apb_02_state;
  wire   [1:0] j202_soc_core_ahb2apb_02_hsize_buf;
  wire   [7:0] j202_soc_core_gpio_core_00_reg_addr;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_dtr;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_isr;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_ier;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2;
  wire   [31:0] j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1;
  wire   [7:0] j202_soc_core_uart_din_i;
  wire   [7:0] j202_soc_core_uart_div1;
  wire   [7:0] j202_soc_core_uart_div0;
  wire   [1:0] j202_soc_core_uart_TOP_dpll_state;
  wire   [3:0] j202_soc_core_uart_TOP_rx_bit_cnt;
  wire   [3:0] j202_soc_core_uart_TOP_tx_bit_cnt;
  wire   [8:0] j202_soc_core_uart_TOP_hold_reg;
  wire   [9:2] j202_soc_core_uart_TOP_rxr;
  wire   [31:0] j202_soc_core_uart_TOP_tx_fifo_mem;
  wire   [1:0] j202_soc_core_uart_TOP_tx_fifo_rp;
  wire   [1:0] j202_soc_core_uart_TOP_tx_fifo_wp;
  wire   [31:0] j202_soc_core_uart_TOP_rx_fifo_mem;
  wire   [1:0] j202_soc_core_uart_TOP_rx_fifo_rp;
  wire   [1:0] j202_soc_core_uart_TOP_rx_fifo_wp;
  wire   [1:0] j202_soc_core_uart_BRG_cnt;
  wire   [7:0] j202_soc_core_uart_BRG_br_cnt;
  wire   [7:0] j202_soc_core_uart_BRG_ps;
  wire   [2:0] j202_soc_core_bldc_core_00_hall_value;
  wire   [2:0] j202_soc_core_bldc_core_00_comm;
  wire   [11:0] j202_soc_core_bldc_core_00_pwm_period;
  wire   [11:0] j202_soc_core_bldc_core_00_pwm_duty;
  wire   [23:0] j202_soc_core_bldc_core_00_wdata;
  wire   [7:0] j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1;
  wire   [1:0] j202_soc_core_bldc_core_00_bldc_wb_slave_00_state;
  wire  
         [2:0] j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status
;
  wire   [2:0] j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3;
  wire   [2:0] j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2;
  wire   [2:0] j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1;
  wire   [11:0] j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt;
  wire   [11:0] j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt;
  wire   [31:0] j202_soc_core_wbqspiflash_00_spif_data;
  wire   [7:0] j202_soc_core_wbqspiflash_00_last_status;
  wire   [9:0] j202_soc_core_wbqspiflash_00_reset_counter;
  wire   [4:0] j202_soc_core_wbqspiflash_00_state;
  wire   [7:0] j202_soc_core_wbqspiflash_00_erased_sector;
  wire   [23:2] j202_soc_core_wbqspiflash_00_w_spif_addr;
  wire   [3:0] j202_soc_core_wbqspiflash_00_w_qspi_dat;
  wire   [1:0] j202_soc_core_wbqspiflash_00_w_qspi_mod;
  wire   [31:0] j202_soc_core_wbqspiflash_00_spi_out;
  wire   [1:0] j202_soc_core_wbqspiflash_00_spi_len;
  wire   [31:0] j202_soc_core_wbqspiflash_00_spi_in;
  wire   [5:0] j202_soc_core_wbqspiflash_00_lldriver_spi_len;
  wire   [31:0] j202_soc_core_wbqspiflash_00_lldriver_r_word;
  wire   [30:0] j202_soc_core_wbqspiflash_00_lldriver_r_input;
  wire   [2:0] j202_soc_core_wbqspiflash_00_lldriver_state;
  wire   [17:2] j202_soc_core_bootrom_00_address_w;

/*sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_15__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[511:480]), .addr0({n25694, n25715, 
        n10938, n25706, n10940, n25709, n25700, n25697, n25712}), .wmask0({
        n11168, n10976, n25703, n25722}), .dout1({SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_1}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10555), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );*/

  assign j202_soc_core_memory0_ram_dout0[511:480] = 32'd0;

  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_14__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[479:448]), .addr0({n11032, n10997, 
        n10983, n11012, n10988, n11007, n11022, n11027, n11002}), .wmask0({
        n10966, n10958, n11017, n10969}), .dout1({SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_33}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10554), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_13__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[447:416]), .addr0({n25693, n25714, 
        n10938, n25705, n10940, n25708, n25699, n25696, n25711}), .wmask0({
        n10962, n10959, n25702, n25723}), .dout1({SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_96, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_90, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_65}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10553), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_12__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[415:384]), .addr0({n25694, n25715, 
        n25729, n25706, n25727, n25709, n25700, n25697, n25712}), .wmask0({
        n11168, n10960, n25703, n25725}), .dout1({SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_118, 
        SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_116, 
        SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_114, 
        SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_112, 
        SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_110, 
        SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_128, 
        SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_126, 
        SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_124, 
        SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_122, 
        SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_108, 
        SYNOPSYS_UNCONNECTED_97}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10552), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_11__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[383:352]), .addr0({n10956, n10942, 
        n10938, n10948, n10940, n10946, n10952, n10954, n10944}), .wmask0({
        n10963, n10960, n10950, n10993}), .dout1({SYNOPSYS_UNCONNECTED_153, 
        SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_140, 
        SYNOPSYS_UNCONNECTED_129}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10551), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_10__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[351:320]), .addr0({n25670, n25691, 
        n25721, n25682, n25720, n25685, n25676, n25673, n25688}), .wmask0({
        n10978, n10976, n25679, n10969}), .dout1({SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_178, 
        SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_176, 
        SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_174, 
        SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_171, 
        SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_169, 
        SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_167, 
        SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_165, 
        SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_163, 
        SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_192, 
        SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_190, 
        SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_188, 
        SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_186, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_172, 
        SYNOPSYS_UNCONNECTED_161}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10550), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_9__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[319:288]), .addr0({n25670, n25691, 
        n10918, n25682, n10920, n25685, n25676, n25673, n25688}), .wmask0({
        n10963, n10974, n25679, n10968}), .dout1({SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_214, 
        SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_212, 
        SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_210, 
        SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_208, 
        SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_206, 
        SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_224, 
        SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_222, 
        SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_220, 
        SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_218, 
        SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_204, 
        SYNOPSYS_UNCONNECTED_193}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10549), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_8__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[287:256]), .addr0({n10936, n10922, 
        n10983, n10928, n10988, n10926, n10932, n10934, n10924}), .wmask0({
        n10979, n25718, n10930, n10968}), .dout1({SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_246, 
        SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_244, 
        SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_242, 
        SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_240, 
        SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_238, 
        SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_256, 
        SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_254, 
        SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_252, 
        SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_250, 
        SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_236, 
        SYNOPSYS_UNCONNECTED_225}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10548), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
/*sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_7__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[255:224]), .addr0({n11032, n10997, 
        n10983, n11012, n10988, n11007, n11022, n11027, n11002}), .wmask0({
        n10979, n25717, n11017, n10969}), .dout1({SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_278, 
        SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_276, 
        SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_274, 
        SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_272, 
        SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_270, 
        SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_288, 
        SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_286, 
        SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_284, 
        SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_282, 
        SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_268, 
        SYNOPSYS_UNCONNECTED_257}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10547), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );*/

  assign j202_soc_core_memory0_ram_dout0[255:224] = 32'd0;

  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_6__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[223:192]), .addr0({n11035, n11000, 
        n25729, n11015, n25727, n11010, n11025, n11030, n11005}), .wmask0({
        n10971, n10976, n11020, n10993}), .dout1({SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_299, 
        SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_297, 
        SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_295, 
        SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_293, 
        SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_291, 
        SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_320, 
        SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_318, 
        SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_316, 
        SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_314, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_289}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10546), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_5__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[191:160]), .addr0({n11032, n10997, 
        n25721, n11012, n25720, n11007, n11022, n11027, n11002}), .wmask0({
        n10962, n10974, n11017, n25724}), .dout1({SYNOPSYS_UNCONNECTED_345, 
        SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_338, 
        SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_336, 
        SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_334, 
        SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_331, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_352, 
        SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_350, 
        SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_348, 
        SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_346, 
        SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_332, 
        SYNOPSYS_UNCONNECTED_321}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10545), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_4__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[159:128]), .addr0({n11032, n10997, 
        n10918, n11012, n10920, n11007, n11022, n11027, n11002}), .wmask0({
        n10965, n10974, n11017, n10995}), .dout1({SYNOPSYS_UNCONNECTED_377, 
        SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_374, 
        SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_372, 
        SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_370, 
        SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_368, 
        SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_366, 
        SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_363, 
        SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_361, 
        SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_359, 
        SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_357, 
        SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_355, 
        SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_384, 
        SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_382, 
        SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_380, 
        SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_378, 
        SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_364, 
        SYNOPSYS_UNCONNECTED_353}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10544), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_3__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[127:96]), .addr0({n25669, n25690, 
        n10918, n25681, n10920, n25684, n25675, n25672, n25687}), .wmask0({
        n10971, n10974, n25678, n10995}), .dout1({SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_406, 
        SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_404, 
        SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_402, 
        SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_400, 
        SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_398, 
        SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_389, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_416, 
        SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_414, 
        SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_412, 
        SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_410, 
        SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_396, 
        SYNOPSYS_UNCONNECTED_385}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10543), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_2__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[95:64]), .addr0({n11032, n10997, 
        n10983, n11012, n10988, n11007, n11022, n11027, n11002}), .wmask0({
        n10966, n10959, n11017, n10995}), .dout1({SYNOPSYS_UNCONNECTED_441, 
        SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_438, 
        SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_436, 
        SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_434, 
        SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_432, 
        SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_430, 
        SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_427, 
        SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_425, 
        SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_423, 
        SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_421, 
        SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_419, 
        SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_448, 
        SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_446, 
        SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_444, 
        SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_442, 
        SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_428, 
        SYNOPSYS_UNCONNECTED_417}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10542), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_1__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[63:32]), .addr0({n25693, n25714, 
        n10938, n25705, n10940, n25708, n25699, n25696, n25711}), .wmask0({
        n10965, n25718, n25702, n10993}), .dout1({SYNOPSYS_UNCONNECTED_473, 
        SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_470, 
        SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_468, 
        SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_466, 
        SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_464, 
        SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_462, 
        SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_459, 
        SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_457, 
        SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_455, 
        SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_453, 
        SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_451, 
        SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_480, 
        SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_478, 
        SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_476, 
        SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_474, 
        SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_460, 
        SYNOPSYS_UNCONNECTED_449}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10541), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_sram_2kbyte_1rw1r_32x512_8 j202_soc_core_memory0_g_ram_0__ram ( 
        .din0({n25519, n25518, n25516, n25515, n25514, n25513, n25512, n25511, 
        n25510, n25509, n25508, n25507, n25505, n25504, n25503, n25502, n25501, 
        n25500, n25499, n25498, n25497, n25496, n25526, n25525, n25524, n25523, 
        n25522, n25521, n25520, n25517, n25506, n25495}), .dout0(
        j202_soc_core_memory0_ram_dout0[31:0]), .addr0({n25669, n25690, n10918, 
        n25681, n10920, n25684, n25675, n25672, n25687}), .wmask0({n10971, 
        n25717, n25678, n10968}), .dout1({SYNOPSYS_UNCONNECTED_505, 
        SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_502, 
        SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_500, 
        SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_498, 
        SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_496, 
        SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_494, 
        SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_491, 
        SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_489, 
        SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_487, 
        SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_485, 
        SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_483, 
        SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_512, 
        SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_510, 
        SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_508, 
        SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_506, 
        SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_492, 
        SYNOPSYS_UNCONNECTED_481}), .addr1({j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127, 
        j202_soc_core_ahb2aqu_00_N127, j202_soc_core_ahb2aqu_00_N127}), .csb0(
        n10540), .web0(n10539), .clk0(wb_clk_i), .csb1(
        j202_soc_core_ahb2aqu_00_N127), .clk1(wb_clk_i) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_31_ ( .D(n390), .DE(n310), .CLK(
        wb_clk_i), .Q(wbs_dat_o[31]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_30_ ( .D(n380), .DE(n310), .CLK(
        wb_clk_i), .Q(wbs_dat_o[30]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_29_ ( .D(n370), .DE(n310), .CLK(
        wb_clk_i), .Q(wbs_dat_o[29]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_28_ ( .D(n360), .DE(n310), .CLK(
        wb_clk_i), .Q(wbs_dat_o[28]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_27_ ( .D(n350), .DE(n310), .CLK(
        wb_clk_i), .Q(wbs_dat_o[27]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_26_ ( .D(n340), .DE(n310), .CLK(
        wb_clk_i), .Q(wbs_dat_o[26]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_25_ ( .D(n330), .DE(n310), .CLK(
        wb_clk_i), .Q(wbs_dat_o[25]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_24_ ( .D(n320), .DE(n310), .CLK(
        wb_clk_i), .Q(wbs_dat_o[24]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_23_ ( .D(n300), .DE(n220), .CLK(
        wb_clk_i), .Q(wbs_dat_o[23]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_22_ ( .D(n290), .DE(n220), .CLK(
        wb_clk_i), .Q(wbs_dat_o[22]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_21_ ( .D(n280), .DE(n220), .CLK(
        wb_clk_i), .Q(wbs_dat_o[21]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_20_ ( .D(n270), .DE(n220), .CLK(
        wb_clk_i), .Q(wbs_dat_o[20]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_19_ ( .D(n260), .DE(n220), .CLK(
        wb_clk_i), .Q(wbs_dat_o[19]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_18_ ( .D(n250), .DE(n220), .CLK(
        wb_clk_i), .Q(wbs_dat_o[18]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_17_ ( .D(n240), .DE(n220), .CLK(
        wb_clk_i), .Q(wbs_dat_o[17]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_16_ ( .D(n230), .DE(n220), .CLK(
        wb_clk_i), .Q(wbs_dat_o[16]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_15_ ( .D(n21), .DE(n13), .CLK(wb_clk_i), .Q(wbs_dat_o[15]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_14_ ( .D(n20), .DE(n13), .CLK(wb_clk_i), .Q(wbs_dat_o[14]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_13_ ( .D(n19), .DE(n13), .CLK(wb_clk_i), .Q(wbs_dat_o[13]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_12_ ( .D(n18), .DE(n13), .CLK(wb_clk_i), .Q(wbs_dat_o[12]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_11_ ( .D(n17), .DE(n13), .CLK(wb_clk_i), .Q(wbs_dat_o[11]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_10_ ( .D(n16), .DE(n13), .CLK(wb_clk_i), .Q(wbs_dat_o[10]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_9_ ( .D(n15), .DE(n13), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[9]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_8_ ( .D(n14), .DE(n13), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[8]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_7_ ( .D(n12), .DE(n4), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[7]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_6_ ( .D(n11), .DE(n4), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[6]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_5_ ( .D(n10), .DE(n4), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[5]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_4_ ( .D(n9), .DE(n4), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[4]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_3_ ( .D(n8), .DE(n4), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[3]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_2_ ( .D(n7), .DE(n4), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[2]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_1_ ( .D(n6), .DE(n4), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[1]) );
  sky130_fd_sc_hd__edfxtp_1 reg_val_reg_0_ ( .D(n5), .DE(n4), .CLK(wb_clk_i), 
        .Q(wbs_dat_o[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_rst0_reg ( .D(n10484), .CLK(wb_clk_i), 
        .Q(j202_soc_core_rst0) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_rst1_reg ( .D(j202_soc_core_rst0), 
        .CLK(wb_clk_i), .Q(j202_soc_core_rst1) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_0_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N3), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_1_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N4), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_2_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N5), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_3_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N6), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_4_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N7), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_5_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N8), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_6_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N9), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_7_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N10), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_8_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N11), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_9_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N12), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_10_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N13), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[10])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_11_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N14), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[11])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_12_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N15), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[12])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_13_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N16), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[13])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_14_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N17), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[14])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_15_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N18), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[15])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_16_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N19), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[16])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_17_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N20), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[17])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_18_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N21), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[18])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_19_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N22), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[19])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_20_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N23), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[20])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_21_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[21])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_22_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N25), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[22])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_23_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N26), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[23])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_24_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N27), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[24])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_25_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N28), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[25])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_26_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N29), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[26])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_27_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N30), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[27])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_28_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N31), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[28])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_29_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N32), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[29])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_30_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N33), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[30])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_dout_reg_31_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N34), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[31])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_0_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N3), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_1_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N4), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_2_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N5), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_3_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N6), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_4_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N7), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_5_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N8), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_6_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N9), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_7_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N10), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_8_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N11), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_9_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N12), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_10_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N13), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[10])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_11_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N14), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[11])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_12_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N15), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[12])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_13_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N16), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_14_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N17), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_15_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N18), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_16_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N19), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_17_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N20), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[17])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_18_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N21), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[18])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_19_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N22), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[19])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_20_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N23), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[20])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_21_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[21])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_22_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N25), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[22])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_23_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N26), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[23])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_24_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N27), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[24])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_25_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N28), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[25])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_26_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N29), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[26])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_27_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N30), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[27])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_28_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N31), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[28])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_29_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N32), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[29])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_30_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N33), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[30])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_dout_reg_31_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N34), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[31])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_0_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N3), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_1_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N4), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_2_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N5), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_3_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N6), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_4_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N7), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_5_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N8), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_6_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N9), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_7_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N10), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_8_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N11), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_9_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N12), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_10_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N13), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[10])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_11_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N14), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[11])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_12_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N15), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[12])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_13_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N16), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[13])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_14_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N17), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[14])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_15_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N18), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[15])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_16_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N19), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[16])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_17_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N20), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[17])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_18_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N21), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[18])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_19_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N22), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[19])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_20_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N23), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[20])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_21_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[21])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_22_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N25), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[22])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_23_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N26), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[23])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_24_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N27), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[24])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_25_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N28), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[25])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_26_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N29), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[26])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_27_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N30), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[27])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_28_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N31), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[28])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_29_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N32), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[29])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_30_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N33), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[30])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_dout_reg_31_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N34), .CLK(
        wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[31])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rxd_s_reg ( .D(io_in[5]), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rxd_s) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rxd_r_reg ( .D(
        j202_soc_core_uart_TOP_rxd_s), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rxd_r) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1_reg_0_ ( 
        .D(io_in[22]), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2_reg_0_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[0]), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3_reg_0_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[0]), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1_reg_1_ ( 
        .D(io_in[23]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2_reg_1_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[1]), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3_reg_1_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[1]), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1_reg_2_ ( 
        .D(io_in[24]), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2_reg_2_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[2]), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3_reg_2_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_2[2]), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1_reg ( 
        .D(n25406), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_2_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_2) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_o_reg_2_ ( 
        .D(n138), .CLK(wb_clk_i), .RESET_B(n25732), .Q(
        j202_soc_core_bldc_core_00_hall_value[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status_reg_2_ ( 
        .D(j202_soc_core_bldc_core_00_hall_value[2]), .CLK(wb_clk_i), 
        .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_o_reg_0_ ( 
        .D(n137), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_hall_value[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status_reg_0_ ( 
        .D(j202_soc_core_bldc_core_00_hall_value[0]), .CLK(wb_clk_i), 
        .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_o_reg_1_ ( 
        .D(n136), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_hall_value[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status_reg_1_ ( 
        .D(j202_soc_core_bldc_core_00_hall_value[1]), .CLK(wb_clk_i), 
        .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_0_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[0]), .CLK(
        wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_1_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[1]), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_2_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[2]), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_3_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[3]), .CLK(
        wb_clk_i), .RESET_B(n25732), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_4_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[4]), .CLK(
        wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_5_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[5]), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_6_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[6]), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_7_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[7]), .CLK(
        wb_clk_i), .RESET_B(n25732), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_8_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[8]), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_9_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[9]), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_10_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[10]), .CLK(
        wb_clk_i), .RESET_B(n25732), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt_reg_11_ ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[11]), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_bootrom_00_sel_w_reg ( .D(n25542), 
        .CLK(wb_clk_i), .Q(j202_soc_core_bootrom_00_sel_w) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_other__2_ ( 
        .D(n10485), .DE(n10581), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_other__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_ifetchl_reg ( .D(
        j202_soc_core_j22_cpu_ifetch), .DE(j202_soc_core_ahbcs_6__HREADY_), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ifetchl) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_area_reg_0_ ( .D(n10538), .DE(n10559), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ma_M_area[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aqu_st_reg_0_ ( .D(
        j202_soc_core_ahb2aqu_00_N93), .DE(j202_soc_core_ahb2aqu_00_N95), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2aqu_00_aqu_st_0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_STB_ ( .D(
        j202_soc_core_ahb2aqu_00_N128), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_STB_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_area_reg_1_ ( .D(n10537), .DE(n10559), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ma_M_area[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_WE_ ( .D(n25248), .DE(j202_soc_core_ahb2aqu_00_N95), .CLK(wb_clk_i), .Q(j202_soc_core_aquc_WE_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_state_reg_0_ ( 
        .D(n25245), .CLK(wb_clk_i), .RESET_B(n25732), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_1_ ( .D(
        n10564), .DE(n10560), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_opst[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rb__1_ ( 
        .D(n10579), .DE(n10568), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rb__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__2_ ( 
        .D(n10498), .DE(n10582), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__2_ ( .D(
        j202_soc_core_ahb2aqu_00_N131), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_ADR__2_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_2_ ( 
        .D(j202_soc_core_aquc_ADR__2_), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_2_ ( .D(
        n25333), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_other__0_ ( 
        .D(n10487), .DE(n10581), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_other__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__15_ ( 
        .D(n25345), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_15_ ( 
        .D(j202_soc_core_qspi_wb_wdat[15]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_bldc_core_00_wdata[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_15_ ( 
        .D(j202_soc_core_qspi_wb_wdat[15]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_15_ ( 
        .D(n25262), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_15_ ( .D(
        j202_soc_core_ahb2apb_02_N143), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[47]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__7_ ( 
        .D(n10493), .DE(n10582), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__7_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__7_ ( .D(
        j202_soc_core_ahb2aqu_00_N136), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_ADR__7_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_7_ ( 
        .D(j202_soc_core_aquc_ADR__7_), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_7_ ( .D(
        n25338), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rn__3_ ( 
        .D(n10574), .DE(n10569), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rn__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__10_ ( 
        .D(n25342), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_10_ ( 
        .D(j202_soc_core_qspi_wb_wdat[10]), .CLK(wb_clk_i), .RESET_B(n25732), 
        .Q(j202_soc_core_bldc_core_00_wdata[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_10_ ( 
        .D(j202_soc_core_qspi_wb_wdat[10]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_10_ ( 
        .D(n25263), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_10_ ( .D(
        j202_soc_core_ahb2apb_02_N138), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[42]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__0_ ( 
        .D(n10583), .DE(n10560), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__4_ ( .D(
        j202_soc_core_j22_cpu_ml_N195), .DE(j202_soc_core_ahbcs_6__HREADY_), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_M_macop_MAC_[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__4_ ( .D(
        j202_soc_core_j22_cpu_ml_N156), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_Ma__1_ ( 
        .D(n10500), .DE(n10570), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_memop_Ma__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_4_ ( 
        .D(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_N487), .DE(n10559), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_other__1_ ( 
        .D(n10486), .DE(n10581), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_other__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_20_ ( .D(
        j202_soc_core_j22_cpu_rf_N318), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__12_ ( 
        .D(n10488), .DE(n10582), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__12_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__12_ ( 
        .D(n25302), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_12_ ( 
        .D(j202_soc_core_qspi_wb_wdat[12]), .CLK(wb_clk_i), .RESET_B(n25732), 
        .Q(j202_soc_core_bldc_core_00_wdata[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_12_ ( 
        .D(j202_soc_core_qspi_wb_wdat[12]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__0_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__3_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_4_ ( 
        .D(n25370), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__4_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_6_ ( 
        .D(n25544), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__6_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__2_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_4_ ( 
        .D(n25390), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__4_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__1_ ( .D(
        n25274), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__2_ ( .D(
        n25246), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__3_ ( .D(
        n25253), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__7_ ( .D(
        n25247), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__7_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__10_ ( .D(
        n25314), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__10_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__11_ ( .D(
        n25311), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__11_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__12_ ( .D(
        n25312), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__12_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__15_ ( .D(
        n25388), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__15_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__0_ ( .D(
        n25259), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_v_ ( .D(n25434), 
        .DE(n10533), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_id_opn_v_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_We__0_ ( 
        .D(n10575), .DE(n10604), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_We__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Wm__3_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N900), .DE(n10604), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_Wm__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_2_ ( .D(
        n10563), .DE(n10560), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_opst[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__4_ ( 
        .D(n10587), .DE(n10560), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__1_ ( 
        .D(n10499), .DE(n10582), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_address_reg_1_ ( .D(
        n25391), .DE(n25543), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_address[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__1_ ( .D(
        j202_soc_core_ahb2aqu_00_N130), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_ADR__1_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_1_ ( 
        .D(j202_soc_core_aquc_ADR__1_), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_SEL__3_ ( .D(
        j202_soc_core_ahb2aqu_00_N164), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_SEL__3_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_1_ ( .D(n135), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_uart_div0[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__3_ ( 
        .D(n10497), .DE(n10582), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__3_ ( .D(
        j202_soc_core_ahb2aqu_00_N132), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_ADR__3_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_3_ ( 
        .D(j202_soc_core_aquc_ADR__3_), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_3_ ( .D(
        n25334), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__8_ ( .D(
        n25308), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__8_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__0_ ( 
        .D(n10591), .DE(n10568), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_istall_reg ( .D(n10556), 
        .DE(n10605), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_istall) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_v_ ( .D(n25299), 
        .DE(j202_soc_core_ahbcs_6__HREADY_), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_v_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__0_ ( .D(
        n25372), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__1_ ( .D(
        n25377), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__2_ ( .D(
        n25381), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__3_ ( .D(
        n25380), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__6_ ( .D(
        n25384), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__6_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__7_ ( .D(
        n25383), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__7_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__8_ ( .D(
        n25387), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__8_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__9_ ( .D(
        n25385), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__9_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__10_ ( .D(
        n25369), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__10_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__11_ ( .D(
        n25258), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__11_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__12_ ( .D(
        n25315), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__12_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__15_ ( .D(
        n25316), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__15_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_30_ ( .D(
        j202_soc_core_j22_cpu_rf_N328), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_5_ ( 
        .D(n25249), .DE(n10559), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_2_ ( .D(
        n25333), .DE(n11200), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_3_ ( .D(
        n25334), .DE(n11200), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_7_ ( .D(
        n25338), .DE(n11200), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_18_ ( 
        .D(n25251), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_20_ ( 
        .D(n25250), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_hwrite_temp_reg ( .D(
        n25248), .DE(n11200), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_we) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_req_reg ( .D(
        n10502), .DE(j202_soc_core_wbqspiflash_00_N748), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_req) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_ack_reg ( .D(
        j202_soc_core_wbqspiflash_00_N730), .DE(
        j202_soc_core_wbqspiflash_00_N729), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_ack) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_stb_o_reg ( .D(n11200), 
        .DE(n10536), .CLK(wb_clk_i), .Q(j202_soc_core_ahb2wbqspi_00_stb_o) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_cyc_o_reg ( .D(n11200), 
        .DE(n10536), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_cyc) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_1_ ( .D(
        j202_soc_core_wbqspiflash_00_N725), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_hold_reg ( .D(
        j202_soc_core_wbqspiflash_00_N590), .DE(
        j202_soc_core_wbqspiflash_00_N745), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_hold) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_state_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N308), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N307), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_state[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_write_in_progress_reg ( 
        .D(j202_soc_core_wbqspiflash_00_N709), .DE(
        j202_soc_core_wbqspiflash_00_N708), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_write_in_progress) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_31_ ( .D(
        n10503), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_2_ ( .D(
        j202_soc_core_wbqspiflash_00_N726), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_0_ ( .D(
        j202_soc_core_wbqspiflash_00_N724), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_len_reg_1_ ( .D(
        j202_soc_core_wbqspiflash_00_N737), .DE(
        j202_soc_core_wbqspiflash_00_N735), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_len[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N429), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_state_reg_1_ ( 
        .D(n25396), .DE(j202_soc_core_wbqspiflash_00_lldriver_N307), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_state_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N310), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N307), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_state[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_sck_reg ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N312), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_sck) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_cs_n_reg ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N314), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N313), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_cs_n) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_write_protect_reg ( 
        .D(j202_soc_core_wbqspiflash_00_N722), .DE(
        j202_soc_core_wbqspiflash_00_N721), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_write_protect) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_28_ ( 
        .D(j202_soc_core_wbqspiflash_00_N695), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_0_ ( 
        .D(n25541), .DE(n10559), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_00_state_reg_0_ ( .D(
        j202_soc_core_ahb2apb_00_N89), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_00_state[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_00_state_reg_2_ ( .D(
        j202_soc_core_ahb2apb_00_N91), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_00_state[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_00_state_reg_1_ ( .D(
        j202_soc_core_ahb2apb_00_N90), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_00_state[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_state_reg_1_ ( 
        .D(n25403), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_state_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_apb_00_nxt_state_0_), .CLK(wb_clk_i), 
        .RESET_B(n25734), .Q(j202_soc_core_cmt_core_00_cmt_apb_00_state[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_hwrite_buf_reg ( .D(
        j202_soc_core_ahb2apb_00_N55), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_pwrite[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_1_reg ( 
        .D(j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen), .CLK(wb_clk_i), 
        .RESET_B(n25730), .Q(j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_1)
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_2_reg ( 
        .D(j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_1), .CLK(wb_clk_i), 
        .RESET_B(n25733), .Q(j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_2)
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_7_ ( .D(
        j202_soc_core_ahb2apb_00_N30), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_7_ ( 
        .D(j202_soc_core_paddr[7]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_reg_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_3_ ( .D(
        j202_soc_core_ahb2apb_00_N26), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_3_ ( 
        .D(j202_soc_core_paddr[3]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_reg_addr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_2_ ( .D(
        j202_soc_core_ahb2apb_00_N25), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_2_ ( 
        .D(j202_soc_core_paddr[2]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_reg_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_00_N24), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_1_ ( 
        .D(j202_soc_core_paddr[1]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_reg_addr[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_6_ ( 
        .D(n134), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N19), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[16])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_16_ ( .D(
        j202_soc_core_ahb2apb_01_N144), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[80]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_16_ ( 
        .D(n25260), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_3_ ( 
        .D(n25376), .DE(n10559), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_CE__1_ ( .D(
        j202_soc_core_ahb2aqu_00_N98), .DE(j202_soc_core_ahb2aqu_00_N95), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_CE__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_19_ ( 
        .D(n25252), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_17_ ( 
        .D(j202_soc_core_qspi_wb_addr[19]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_dirty_sector_reg ( 
        .D(j202_soc_core_wbqspiflash_00_N720), .DE(
        j202_soc_core_wbqspiflash_00_N719), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_dirty_sector) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_30_ ( 
        .D(j202_soc_core_wbqspiflash_00_N697), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__14_ ( .D(
        n25304), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__14_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rb__0_ ( 
        .D(n10578), .DE(n10568), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rb__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_21_ ( .D(
        j202_soc_core_j22_cpu_rf_N319), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__13_ ( .D(
        n25309), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__13_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__13_ ( .D(
        n25303), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__13_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rm__2_ ( 
        .D(n25384), .DE(j202_soc_core_j22_cpu_id_idec_N857), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_Rm__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rm__3_ ( 
        .D(n25383), .DE(j202_soc_core_j22_cpu_id_idec_N857), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_Rm__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__14_ ( .D(
        n25310), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__14_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_14_ ( 
        .D(n25273), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_0_ ( .D(
        n25321), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__t_ ( .D(
        j202_soc_core_j22_cpu_rf_N2626), .DE(j202_soc_core_j22_cpu_rf_N2625), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__t_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_19_ ( .D(
        j202_soc_core_j22_cpu_rf_N317), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__11_ ( 
        .D(n25343), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_11_ ( 
        .D(j202_soc_core_qspi_wb_wdat[11]), .CLK(wb_clk_i), .RESET_B(n25732), 
        .Q(j202_soc_core_bldc_core_00_wdata[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_11_ ( 
        .D(j202_soc_core_qspi_wb_wdat[11]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[11]), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_cmt_core_00_cnt1[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[11]), .CLK(wb_clk_i), .RESET_B(
        n25732), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmf1_o_reg ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt1_to1), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_cmt_core_00_cmf1) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[9]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_cmt_core_00_cnt1[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[9]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[9]), .CLK(wb_clk_i), 
        .RESET_B(n25733), .Q(j202_soc_core_prdata[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_9_ ( .D(
        j202_soc_core_ahb2apb_00_N137), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[105])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__9_ ( .D(
        n25313), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__9_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_9_ ( .D(
        n25375), .DE(n11200), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_9_ ( .D(
        n25375), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3204), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[455]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__14_ ( 
        .D(n25301), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_14_ ( 
        .D(j202_soc_core_qspi_wb_wdat[14]), .CLK(wb_clk_i), .RESET_B(n25730), 
        .Q(j202_soc_core_bldc_core_00_wdata[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_14_ ( 
        .D(j202_soc_core_qspi_wb_wdat[14]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__i__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3390), .DE(j202_soc_core_j22_cpu_rf_N3391), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__i__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_6_ ( .D(
        j202_soc_core_ahb2apb_00_N29), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_6_ ( 
        .D(j202_soc_core_paddr[6]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_reg_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__6_ ( .D(
        j202_soc_core_ahb2aqu_00_N135), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_ADR__6_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_6_ ( 
        .D(j202_soc_core_aquc_ADR__6_), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_6_ ( .D(
        n25337), .DE(n11200), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_6_ ( .D(
        n25337), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_17_ ( 
        .D(n25254), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_17_ ( .D(
        n25254), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__5_ ( .D(
        n25382), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__5_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rm__1_ ( 
        .D(n25382), .DE(j202_soc_core_j22_cpu_id_idec_N857), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_Rm__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__5_ ( 
        .D(n10495), .DE(n10582), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__5_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_5_ ( .D(
        j202_soc_core_ahb2apb_00_N28), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_5_ ( 
        .D(j202_soc_core_paddr[5]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_reg_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__5_ ( .D(
        j202_soc_core_ahb2aqu_00_N134), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_ADR__5_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_5_ ( 
        .D(j202_soc_core_aquc_ADR__5_), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_5_ ( .D(
        n25336), .DE(n11200), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_5_ ( .D(
        n25336), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__4_ ( .D(
        n25256), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__4_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_op2_reg_inst__4_ ( .D(
        n25386), .DE(j202_soc_core_j22_cpu_id_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_op2_inst__4_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rm__0_ ( 
        .D(n25386), .DE(j202_soc_core_j22_cpu_id_idec_N857), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_Rm__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__0_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N917), .DE(n10582), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_imm__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_MEM__1_ ( 
        .D(n10588), .DE(n10560), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_memop_MEM__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_MEM_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ma_N54), .DE(n10559), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_MEM[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_SEL__2_ ( .D(
        j202_soc_core_ahb2aqu_00_N163), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_SEL__2_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_1_ ( .D(n133), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_uart_div1[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_br_clr_reg ( .D(
        j202_soc_core_uart_BRG_N47), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_clr) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_x4_r_reg ( .D(
        j202_soc_core_uart_BRG_br_clr), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_sio_ce_x4_r) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_x4_t_reg ( .D(n25400), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_BRG_sio_ce_x4_t) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_x4_reg ( .D(
        j202_soc_core_uart_BRG_sio_ce_x4_t), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_sio_ce_x4) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_change_reg ( .D(
        j202_soc_core_uart_TOP_N102), .DE(j202_soc_core_uart_TOP_N101), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_change) );
  sky130_fd_sc_hd__dfstp_1 j202_soc_core_uart_TOP_dpll_state_reg_0_ ( .D(n132), 
        .CLK(wb_clk_i), .SET_B(n25733), .Q(
        j202_soc_core_uart_TOP_dpll_state[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_sio_ce_r1_reg ( .D(n25405), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_sio_ce_r1) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_sio_ce_r2_reg ( .D(
        j202_soc_core_uart_TOP_rx_sio_ce_r1), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_sio_ce_r2) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_sio_ce_reg ( .D(
        j202_soc_core_uart_TOP_N118), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_sio_ce) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_9_ ( .D(
        j202_soc_core_uart_TOP_rxd_s), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_8_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_7_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_6_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_5_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_4_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_3_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rxr_reg_2_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(j202_soc_core_uart_TOP_N95), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rxr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_bit_cnt_reg_0_ ( .D(
        j202_soc_core_uart_TOP_N86), .DE(j202_soc_core_uart_TOP_N85), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_bit_cnt[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_bit_cnt_reg_1_ ( .D(
        j202_soc_core_uart_TOP_N87), .DE(j202_soc_core_uart_TOP_N85), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_bit_cnt[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_bit_cnt_reg_2_ ( .D(
        j202_soc_core_uart_TOP_N88), .DE(j202_soc_core_uart_TOP_N85), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_bit_cnt[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_bit_cnt_reg_3_ ( .D(
        j202_soc_core_uart_TOP_N89), .DE(j202_soc_core_uart_TOP_N85), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_bit_cnt[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_go_reg ( .D(
        j202_soc_core_uart_TOP_N128), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_go) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_valid_reg ( .D(n10908), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_valid) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_rx_valid_r_reg ( .D(
        j202_soc_core_uart_TOP_rx_valid), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_valid_r) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_rx_fifo_wp_reg_0_ ( .D(n131), 
        .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_uart_TOP_rx_fifo_wp[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_rx_fifo_wp_reg_1_ ( .D(n130), 
        .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_uart_TOP_rx_fifo_wp[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__0_ ( .D(
        j202_soc_core_uart_TOP_rxr[2]), .DE(j202_soc_core_uart_TOP_rx_fifo_N29), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__7_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(j202_soc_core_uart_TOP_rx_fifo_N29), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__6_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(j202_soc_core_uart_TOP_rx_fifo_N29), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__5_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(j202_soc_core_uart_TOP_rx_fifo_N29), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__4_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(j202_soc_core_uart_TOP_rx_fifo_N29), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__3_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(j202_soc_core_uart_TOP_rx_fifo_N29), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__2_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(j202_soc_core_uart_TOP_rx_fifo_N29), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_3__1_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(j202_soc_core_uart_TOP_rx_fifo_N29), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__0_ ( .D(
        j202_soc_core_uart_TOP_rxr[2]), .DE(j202_soc_core_uart_TOP_rx_fifo_N30), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__7_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(j202_soc_core_uart_TOP_rx_fifo_N30), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__6_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(j202_soc_core_uart_TOP_rx_fifo_N30), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__5_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(j202_soc_core_uart_TOP_rx_fifo_N30), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__4_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(j202_soc_core_uart_TOP_rx_fifo_N30), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__3_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(j202_soc_core_uart_TOP_rx_fifo_N30), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__2_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(j202_soc_core_uart_TOP_rx_fifo_N30), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_2__1_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(j202_soc_core_uart_TOP_rx_fifo_N30), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__0_ ( .D(
        j202_soc_core_uart_TOP_rxr[2]), .DE(j202_soc_core_uart_TOP_rx_fifo_N31), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__7_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(j202_soc_core_uart_TOP_rx_fifo_N31), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__6_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(j202_soc_core_uart_TOP_rx_fifo_N31), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__5_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(j202_soc_core_uart_TOP_rx_fifo_N31), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__4_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(j202_soc_core_uart_TOP_rx_fifo_N31), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__3_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(j202_soc_core_uart_TOP_rx_fifo_N31), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__2_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(j202_soc_core_uart_TOP_rx_fifo_N31), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_1__1_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(j202_soc_core_uart_TOP_rx_fifo_N31), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__0_ ( .D(
        j202_soc_core_uart_TOP_rxr[2]), .DE(j202_soc_core_uart_TOP_rx_fifo_N32), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__7_ ( .D(
        j202_soc_core_uart_TOP_rxr[9]), .DE(j202_soc_core_uart_TOP_rx_fifo_N32), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__6_ ( .D(
        j202_soc_core_uart_TOP_rxr[8]), .DE(j202_soc_core_uart_TOP_rx_fifo_N32), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__5_ ( .D(
        j202_soc_core_uart_TOP_rxr[7]), .DE(j202_soc_core_uart_TOP_rx_fifo_N32), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__5_ ( .D(
        n25255), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__5_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__13_ ( 
        .D(n25344), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_13_ ( 
        .D(j202_soc_core_qspi_wb_wdat[13]), .CLK(wb_clk_i), .RESET_B(n25732), 
        .Q(j202_soc_core_bldc_core_00_wdata[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_13_ ( 
        .D(j202_soc_core_qspi_wb_wdat[13]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__i__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3388), .DE(j202_soc_core_j22_cpu_rf_N3391), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__i__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N302), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_4_ ( .D(
        j202_soc_core_ahb2apb_00_N27), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_4_ ( 
        .D(j202_soc_core_paddr[4]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_reg_addr[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_14_ ( 
        .D(n129), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const0[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_13_ ( 
        .D(n128), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const0[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_12_ ( 
        .D(n127), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const0[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_11_ ( 
        .D(n126), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const0[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_10_ ( 
        .D(n125), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const0[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_15_ ( 
        .D(n124), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const0[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_14_ ( 
        .D(n123), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const1[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_13_ ( 
        .D(n122), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const1[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_12_ ( 
        .D(n121), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const1[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_11_ ( 
        .D(n120), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const1[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_10_ ( 
        .D(n119), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const1[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_15_ ( 
        .D(n118), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const1[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__4_ ( .D(
        j202_soc_core_ahb2aqu_00_N133), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_ADR__4_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_4_ ( 
        .D(j202_soc_core_aquc_ADR__4_), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_4_ ( .D(
        n25335), .DE(n11200), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_4_ ( .D(
        n25335), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_31_ ( .D(
        j202_soc_core_j22_cpu_rf_N329), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2676), .DE(n25489), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__8_ ( .D(
        n25367), .DE(n25488), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_8_ ( 
        .D(j202_soc_core_qspi_wb_wdat[8]), .CLK(wb_clk_i), .RESET_B(n25732), 
        .Q(j202_soc_core_bldc_core_00_wdata[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_8_ ( 
        .D(j202_soc_core_qspi_wb_wdat[8]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_8_ ( 
        .D(n117), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_cmt_core_00_const1[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_8_ ( 
        .D(n116), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const0[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intr_level__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__i__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3386), .DE(j202_soc_core_j22_cpu_rf_N3391), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__i__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_6_ ( .D(
        j202_soc_core_j22_cpu_ml_N309), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_24_ ( 
        .D(n25257), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_len_reg_0_ ( .D(
        j202_soc_core_wbqspiflash_00_N736), .DE(
        j202_soc_core_wbqspiflash_00_N735), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_len[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_26_ ( 
        .D(j202_soc_core_wbqspiflash_00_N693), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_26_ ( .D(
        j202_soc_core_j22_cpu_rf_N324), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_26_ ( .D(n25448), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_28_ ( .D(n25432), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2675), .DE(n25489), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_29_ ( .D(n25477), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_16_ ( .D(
        n25260), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_14_ ( .D(
        n25273), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_6_ ( 
        .D(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_N497), .DE(n10559), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_29_ ( .D(
        j202_soc_core_j22_cpu_rf_N327), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2656), .DE(n25489), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_13_ ( 
        .D(n25271), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_13_ ( .D(
        n25271), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_1_ ( .D(
        n25324), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N301), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__3_ ( .D(
        n25363), .DE(n25488), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_3_ ( 
        .D(j202_soc_core_qspi_wb_wdat[3]), .CLK(wb_clk_i), .RESET_B(n25732), 
        .Q(j202_soc_core_bldc_core_00_wdata[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_3_ ( 
        .D(j202_soc_core_qspi_wb_wdat[3]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_3_ ( 
        .D(n115), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_cmt_core_00_const1[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_3_ ( 
        .D(n114), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_cmt_core_00_const0[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_3_ ( 
        .D(n113), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_3_ ( 
        .D(n112), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intr_vec__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_3_ ( .D(
        j202_soc_core_j22_cpu_id_idec_N894), .DE(n10560), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_opst[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_MEM__2_ ( 
        .D(n10589), .DE(n10560), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_memop_MEM__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_MEM_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ma_N55), .DE(n10559), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_MEM[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__5_ ( 
        .D(n10596), .DE(n10568), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__1_ ( 
        .D(n10592), .DE(n10568), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_4_ ( .D(
        n10565), .DE(n10560), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_opst[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rs__0_ ( 
        .D(n25371), .DE(n10568), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rs__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_We__1_ ( 
        .D(n10600), .DE(n10604), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_We__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Wm__1_ ( 
        .D(n10598), .DE(n10604), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Wm__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_opst_reg_0_ ( .D(
        n10567), .DE(n10560), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_opst[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_MEM__3_ ( 
        .D(n10590), .DE(n10560), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_memop_MEM__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_MEM_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ma_N56), .DE(n10559), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_MEM[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_intack_reg ( .D(
        j202_soc_core_j22_cpu_id_idec_N822), .DE(n10562), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_intack) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intack_all_dout_reg_0_ ( 
        .D(n25393), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_cp_intack_all_0_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N4), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N5), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N6), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N9), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rte4_reg ( .D(
        j202_soc_core_j22_cpu_N8), .DE(n10562), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rte4) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Wm__2_ ( 
        .D(n10599), .DE(n10604), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Wm__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Wm__0_ ( 
        .D(n10597), .DE(n10604), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Wm__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_MEM__0_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N937), .DE(n10560), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_memop_MEM__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_MEM_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ma_N53), .DE(n10559), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_MEM[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Rn__3_ ( 
        .D(j202_soc_core_j22_cpu_regop_Rn__3_), .DE(
        j202_soc_core_j22_cpu_id_idec_N960), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_M_Rn__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Wm__0_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N956), .DE(n10558), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Wm__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Wm__3_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N959), .DE(n10558), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Wm__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Wm__2_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N958), .DE(n10558), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Wm__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Wm__1_ ( 
        .D(j202_soc_core_j22_cpu_id_idec_N957), .DE(n10558), .CLK(wb_clk_i), 
        .Q(j202_soc_core_j22_cpu_regop_M_Wm__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__23_ ( 
        .D(n25353), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[23]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_23_ ( 
        .D(j202_soc_core_qspi_wb_wdat[23]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_bldc_core_00_wdata[23]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_7_ ( .D(n111), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_uart_div1[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__21_ ( 
        .D(n25351), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[21]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_21_ ( 
        .D(j202_soc_core_qspi_wb_wdat[21]), .CLK(wb_clk_i), .RESET_B(n25731), 
        .Q(j202_soc_core_bldc_core_00_wdata[21]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_5_ ( .D(n110), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_uart_div1[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__20_ ( 
        .D(n25350), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[20]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_20_ ( 
        .D(j202_soc_core_qspi_wb_wdat[20]), .CLK(wb_clk_i), .RESET_B(n25731), 
        .Q(j202_soc_core_bldc_core_00_wdata[20]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_4_ ( .D(n109), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_uart_div1[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__18_ ( 
        .D(n25348), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[18]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_18_ ( 
        .D(j202_soc_core_qspi_wb_wdat[18]), .CLK(wb_clk_i), .RESET_B(n25730), 
        .Q(j202_soc_core_bldc_core_00_wdata[18]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_2_ ( .D(n108), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_uart_div1[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__7_ ( .D(
        n25366), .DE(n25488), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_7_ ( 
        .D(j202_soc_core_qspi_wb_wdat[7]), .CLK(wb_clk_i), .RESET_B(n25732), 
        .Q(j202_soc_core_bldc_core_00_wdata[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_7_ ( 
        .D(j202_soc_core_qspi_wb_wdat[7]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_7_ ( 
        .D(n107), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_cmt_core_00_const1[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_7_ ( 
        .D(n106), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const0[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_nxt_latch_status_0_), 
        .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__6_ ( .D(
        n25300), .DE(n25488), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_6_ ( 
        .D(j202_soc_core_qspi_wb_wdat[6]), .CLK(wb_clk_i), .RESET_B(n25732), 
        .Q(j202_soc_core_bldc_core_00_wdata[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_6_ ( 
        .D(j202_soc_core_qspi_wb_wdat[6]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_6_ ( 
        .D(n105), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_cmt_core_00_const1[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_6_ ( 
        .D(n104), .CLK(wb_clk_i), .RESET_B(n25732), .Q(
        j202_soc_core_cmt_core_00_const0[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_6_ ( 
        .D(n103), .CLK(wb_clk_i), .RESET_B(n25732), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N20), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[17])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__5_ ( .D(
        n25365), .DE(n25488), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_5_ ( 
        .D(j202_soc_core_qspi_wb_wdat[5]), .CLK(wb_clk_i), .RESET_B(n25732), 
        .Q(j202_soc_core_bldc_core_00_wdata[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_5_ ( 
        .D(j202_soc_core_qspi_wb_wdat[5]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_5_ ( 
        .D(n102), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_cmt_core_00_const1[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_5_ ( 
        .D(n101), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_const0[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_5_ ( 
        .D(n100), .CLK(wb_clk_i), .RESET_B(n25732), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_5_ ( 
        .D(n99), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__4_ ( .D(
        n25364), .DE(n25488), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_4_ ( 
        .D(j202_soc_core_qspi_wb_wdat[4]), .CLK(wb_clk_i), .RESET_B(n25732), 
        .Q(j202_soc_core_bldc_core_00_wdata[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_4_ ( 
        .D(j202_soc_core_qspi_wb_wdat[4]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_4_ ( 
        .D(n98), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_cmt_core_00_const1[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_4_ ( 
        .D(n97), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_cmt_core_00_const0[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_4_ ( 
        .D(n96), .CLK(wb_clk_i), .RESET_B(n25734), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_4_ ( 
        .D(n95), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_pc_hold_reg ( .D(
        n10566), .DE(n10560), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_pc_hold) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_memop_reg_Ma__0_ ( 
        .D(n10501), .DE(n10570), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_memop_Ma__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_We__2_ ( 
        .D(n10576), .DE(n10604), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_We__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rn__2_ ( 
        .D(n10573), .DE(n10569), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rn__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Rn__2_ ( 
        .D(j202_soc_core_j22_cpu_regop_Rn__2_), .DE(
        j202_soc_core_j22_cpu_id_idec_N960), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_M_Rn__2_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rn__1_ ( 
        .D(n10572), .DE(n10569), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rn__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Rn__1_ ( 
        .D(j202_soc_core_j22_cpu_regop_Rn__1_), .DE(
        j202_soc_core_j22_cpu_id_idec_N960), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_M_Rn__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rn__0_ ( 
        .D(n10571), .DE(n10569), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rn__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_M_Rn__0_ ( 
        .D(j202_soc_core_j22_cpu_regop_Rn__0_), .DE(
        j202_soc_core_j22_cpu_id_idec_N960), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_M_Rn__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__4_ ( 
        .D(n10496), .DE(n10582), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__4_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__6_ ( 
        .D(n10494), .DE(n10582), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__6_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__8_ ( 
        .D(n10492), .DE(n10582), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__8_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__9_ ( 
        .D(n10491), .DE(n10582), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__9_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__10_ ( 
        .D(n10490), .DE(n10582), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__10_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_imm__11_ ( 
        .D(n10489), .DE(n10582), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_imm__11_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__4_ ( 
        .D(n10595), .DE(n10568), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__3_ ( 
        .D(n10594), .DE(n10568), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_exuop_reg_EXU__2_ ( 
        .D(n10593), .DE(n10568), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_exuop_EXU_[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_We__3_ ( 
        .D(n25305), .DE(n10604), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_We__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3324), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3313), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3314), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3315), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3316), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3317), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3311), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3338), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3340), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3341), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3342), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3343), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_2_ ( .D(n25480), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2645), .DE(n25489), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2646), .DE(n25489), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_5_ ( .D(n25479), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_6_ ( .D(n25476), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_7_ ( .D(n25431), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_0_ ( .D(n25478), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3302), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3303), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3304), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3305), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3299), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3284), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3278), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3276), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3275), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3274), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3273), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3272), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3347), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3348), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3349), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3350), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3351), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3352), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3359), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3374), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3376), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3377), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3378), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3379), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2710), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2713), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2712), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2711), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2707), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2692), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2686), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2680), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2681), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2682), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2683), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2684), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2747), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[60]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2750), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[63]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2749), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[62]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2748), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[61]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2744), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[58]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2729), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[45]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2723), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[39]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2717), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[34]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2718), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[35]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2719), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[36]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2720), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[37]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2721), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[38]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2784), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[92]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2787), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[95]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2786), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[94]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2785), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[93]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2781), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[90]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2766), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[77]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2760), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[71]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2754), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[66]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2755), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[67]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2756), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[68]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2757), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[69]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2758), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[70]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2821), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[124]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2824), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[127]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2823), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[126]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2822), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[125]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2818), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[122]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2803), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[109]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2797), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[103]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2791), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[98]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2792), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[99]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2793), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[100]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2794), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[101]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2795), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[102]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2858), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[156]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2861), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[159]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2860), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[158]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2859), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[157]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2855), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[154]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2840), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[141]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2834), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[135]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2828), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[130]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2829), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[131]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2830), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[132]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2831), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[133]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2832), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[134]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2895), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[188]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2898), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[191]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2897), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[190]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2896), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[189]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2892), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[186]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2877), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[173]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2871), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[167]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2865), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[162]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2866), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[163]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2867), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[164]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2868), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[165]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2869), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[166]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2932), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[220]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2935), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[223]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2934), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[222]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2933), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[221]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2929), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[218]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2914), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[205]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2908), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[199]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2902), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[194]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2903), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[195]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2904), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[196]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2905), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[197]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2906), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[198]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N2969), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[252]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N2972), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[255]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N2971), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[254]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N2970), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[253]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N2966), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[250]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2951), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[237]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2945), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[231]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2939), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[226]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2940), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[227]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2941), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[228]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2942), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[229]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2943), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[230]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3006), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[284]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3009), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[287]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3008), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[286]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3007), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[285]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3003), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[282]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N2988), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[269]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N2982), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[263]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N2976), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[258]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N2977), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[259]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N2978), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[260]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N2979), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[261]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N2980), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[262]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3043), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[316]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3046), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[319]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3045), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[318]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3044), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[317]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3040), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[314]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3025), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[301]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3019), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[295]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3013), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[290]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3014), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[291]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3015), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[292]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3016), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[293]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3017), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[294]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3080), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[348]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3083), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[351]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3082), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[350]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3081), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[349]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3077), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[346]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3062), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[333]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3056), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[327]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3050), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[322]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3051), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[323]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3052), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[324]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3053), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[325]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3054), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[326]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3117), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[380]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3120), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[383]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3119), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[382]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3118), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[381]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3114), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[378]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3099), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[365]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3093), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[359]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3087), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[354]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3088), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[355]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3089), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[356]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3090), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[357]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3091), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[358]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3154), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[412]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3157), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[415]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3156), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[414]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3155), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[413]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3151), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[410]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3136), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[397]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3130), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[391]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3124), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[386]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3125), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[387]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3126), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[388]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3127), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[389]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3128), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[390]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3191), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[444]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3194), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[447]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3193), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[446]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3192), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[445]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3188), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[442]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3173), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[429]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3167), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[423]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3161), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[418]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3162), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[419]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3163), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[420]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3164), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[421]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3165), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[422]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3228), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[476]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3231), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[479]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3230), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[478]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3229), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[477]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3225), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[474]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3210), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[461]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3198), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[450]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3199), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[451]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3200), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[452]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3201), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[453]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3202), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[454]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__28_ ( .D(
        j202_soc_core_j22_cpu_rf_N3265), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[508]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__31_ ( .D(
        j202_soc_core_j22_cpu_rf_N3268), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[511]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__30_ ( .D(
        j202_soc_core_j22_cpu_rf_N3267), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[510]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__29_ ( .D(
        j202_soc_core_j22_cpu_rf_N3266), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[509]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__26_ ( .D(
        j202_soc_core_j22_cpu_rf_N3262), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[506]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__13_ ( .D(
        j202_soc_core_j22_cpu_rf_N3247), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[493]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__7_ ( .D(
        j202_soc_core_j22_cpu_rf_N3241), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[487]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__2_ ( .D(
        j202_soc_core_j22_cpu_rf_N3235), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[482]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3236), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[483]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__4_ ( .D(
        j202_soc_core_j22_cpu_rf_N3237), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[484]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__5_ ( .D(
        j202_soc_core_j22_cpu_rf_N3238), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[485]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__6_ ( .D(
        j202_soc_core_j22_cpu_rf_N3239), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[486]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__3_ ( 
        .D(n10586), .DE(n10560), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__2_ ( 
        .D(n10585), .DE(n10560), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_macop_reg_MAC__1_ ( 
        .D(n10584), .DE(n10560), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_macop_MAC_[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_2_ ( .D(
        j202_soc_core_j22_cpu_rf_N300), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_5_ ( .D(
        j202_soc_core_j22_cpu_rf_N303), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_6_ ( .D(
        j202_soc_core_j22_cpu_rf_N304), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_13_ ( .D(
        j202_soc_core_j22_cpu_rf_N311), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_28_ ( .D(
        j202_soc_core_j22_cpu_rf_N326), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Ra__1_ ( 
        .D(n10580), .DE(n10568), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Ra__1_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Ra__0_ ( 
        .D(n10603), .DE(n10568), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Ra__0_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_idec_regop_reg_Rs__1_ ( 
        .D(n10602), .DE(n10568), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_regop_Rs__1_) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_req_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_req_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intr_req_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_haddr_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_00_N23), .DE(j202_soc_core_ahb2apb_00_N22), 
        .CLK(wb_clk_i), .Q(j202_soc_core_paddr[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_reg_addr_o_reg_0_ ( 
        .D(j202_soc_core_paddr[0]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_cmt_core_00_reg_addr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_ADR__0_ ( .D(
        j202_soc_core_ahb2aqu_00_N129), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_ADR__0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1_reg_0_ ( 
        .D(j202_soc_core_aquc_ADR__0_), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_SEL__0_ ( .D(
        j202_soc_core_ahb2aqu_00_N161), .DE(j202_soc_core_ahb2aqu_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_SEL__0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_RDRXD1_reg ( .D(n25394), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_uart_RDRXD1) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_rx_fifo_rp_reg_0_ ( .D(n94), 
        .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_uart_TOP_rx_fifo_rp[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_rx_fifo_rp_reg_1_ ( .D(n93), 
        .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_uart_TOP_rx_fifo_rp[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_gb_reg ( .D(
        j202_soc_core_uart_TOP_rx_fifo_N42), .DE(
        j202_soc_core_uart_TOP_rx_fifo_N41), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_rx_fifo_gb) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_3_ ( .D(n92), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_uart_din_i[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_4_ ( .D(n91), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_uart_din_i[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_5_ ( .D(n90), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_uart_din_i[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_6_ ( .D(n89), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_uart_din_i[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_7_ ( .D(n88), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_uart_din_i[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_WRTXD1_reg ( .D(
        j202_soc_core_uart_N5), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_uart_WRTXD1) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_tx_fifo_wp_reg_0_ ( .D(n87), 
        .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_uart_TOP_tx_fifo_wp[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_tx_fifo_wp_reg_1_ ( .D(n86), 
        .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_uart_TOP_tx_fifo_wp[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__7_ ( .D(
        j202_soc_core_uart_din_i[7]), .DE(j202_soc_core_uart_TOP_tx_fifo_N29), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__6_ ( .D(
        j202_soc_core_uart_din_i[6]), .DE(j202_soc_core_uart_TOP_tx_fifo_N29), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__5_ ( .D(
        j202_soc_core_uart_din_i[5]), .DE(j202_soc_core_uart_TOP_tx_fifo_N29), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__4_ ( .D(
        j202_soc_core_uart_din_i[4]), .DE(j202_soc_core_uart_TOP_tx_fifo_N29), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__3_ ( .D(
        j202_soc_core_uart_din_i[3]), .DE(j202_soc_core_uart_TOP_tx_fifo_N29), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__7_ ( .D(
        j202_soc_core_uart_din_i[7]), .DE(j202_soc_core_uart_TOP_tx_fifo_N30), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__6_ ( .D(
        j202_soc_core_uart_din_i[6]), .DE(j202_soc_core_uart_TOP_tx_fifo_N30), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__5_ ( .D(
        j202_soc_core_uart_din_i[5]), .DE(j202_soc_core_uart_TOP_tx_fifo_N30), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__4_ ( .D(
        j202_soc_core_uart_din_i[4]), .DE(j202_soc_core_uart_TOP_tx_fifo_N30), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__3_ ( .D(
        j202_soc_core_uart_din_i[3]), .DE(j202_soc_core_uart_TOP_tx_fifo_N30), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__7_ ( .D(
        j202_soc_core_uart_din_i[7]), .DE(j202_soc_core_uart_TOP_tx_fifo_N31), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__6_ ( .D(
        j202_soc_core_uart_din_i[6]), .DE(j202_soc_core_uart_TOP_tx_fifo_N31), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__5_ ( .D(
        j202_soc_core_uart_din_i[5]), .DE(j202_soc_core_uart_TOP_tx_fifo_N31), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__4_ ( .D(
        j202_soc_core_uart_din_i[4]), .DE(j202_soc_core_uart_TOP_tx_fifo_N31), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__3_ ( .D(
        j202_soc_core_uart_din_i[3]), .DE(j202_soc_core_uart_TOP_tx_fifo_N31), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__7_ ( .D(
        j202_soc_core_uart_din_i[7]), .DE(j202_soc_core_uart_TOP_tx_fifo_N32), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__6_ ( .D(
        j202_soc_core_uart_din_i[6]), .DE(j202_soc_core_uart_TOP_tx_fifo_N32), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__5_ ( .D(
        j202_soc_core_uart_din_i[5]), .DE(j202_soc_core_uart_TOP_tx_fifo_N32), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__4_ ( .D(
        j202_soc_core_uart_din_i[4]), .DE(j202_soc_core_uart_TOP_tx_fifo_N32), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__3_ ( .D(
        j202_soc_core_uart_din_i[3]), .DE(j202_soc_core_uart_TOP_tx_fifo_N32), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_M_address_reg_0_ ( .D(
        n25379), .DE(n25543), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ma_M_address[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3307), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3270), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2678), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3233), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[480]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2715), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[32]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2752), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[64]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2789), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[96]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2826), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[128]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2863), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[160]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2900), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[192]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2937), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[224]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N2974), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[256]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3011), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[288]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3048), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[320]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3085), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[352]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3122), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[384]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3159), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[416]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3196), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[448]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_0_ ( .D(
        j202_soc_core_j22_cpu_rf_N298), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_0_ ( .D(
        j202_soc_core_j22_cpu_rf_N3345), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3370), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3335), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3296), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2704), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2741), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[55]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2778), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[87]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2815), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[119]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2852), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[151]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2889), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[183]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2926), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[215]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N2963), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[247]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3000), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[279]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3037), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[311]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3074), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[343]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3111), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[375]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3148), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[407]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3185), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[439]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3222), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[471]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__23_ ( .D(
        j202_soc_core_j22_cpu_rf_N3259), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[503]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_23_ ( .D(n25475), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_23_ ( .D(
        j202_soc_core_j22_cpu_rf_N321), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3373), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3337), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3298), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2706), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2743), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[57]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2780), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[89]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2817), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[121]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2854), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[153]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2891), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[185]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2928), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[217]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N2965), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[249]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3002), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[281]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3039), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[313]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3076), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[345]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3113), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[377]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3150), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[409]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3187), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[441]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3224), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[473]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__25_ ( .D(
        j202_soc_core_j22_cpu_rf_N3261), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[505]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_25_ ( .D(n25427), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_25_ ( .D(
        j202_soc_core_j22_cpu_rf_N323), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3355), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3319), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3280), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2688), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2725), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[41]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2762), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[73]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2799), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[105]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2836), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[137]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2873), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[169]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2910), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[201]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2947), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[233]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2984), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[265]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3021), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[297]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3058), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[329]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3095), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[361]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3132), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[393]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3169), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[425]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3206), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[457]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__9_ ( .D(
        j202_soc_core_j22_cpu_rf_N3243), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[489]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_9_ ( .D(
        j202_soc_core_j22_cpu_rf_N2652), .DE(n25489), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__m_ ( .D(
        j202_soc_core_j22_cpu_rf_N2640), .DE(j202_soc_core_j22_cpu_rf_N2639), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__m_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3309), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3271), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2679), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2716), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[33]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2753), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[65]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2790), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[97]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2827), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[129]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2864), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[161]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2901), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[193]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2938), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[225]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N2975), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[257]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3012), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[289]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3049), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[321]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3086), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[353]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3123), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[385]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3160), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[417]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3197), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[449]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3234), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[481]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_1_ ( .D(n25474), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__s_ ( .D(
        j202_soc_core_j22_cpu_rf_N2628), .DE(j202_soc_core_j22_cpu_rf_N2627), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__s_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__0_ ( .D(
        j202_soc_core_j22_cpu_ml_N191), .DE(j202_soc_core_ahbcs_6__HREADY_), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__2_ ( .D(
        j202_soc_core_j22_cpu_ml_N193), .DE(j202_soc_core_ahbcs_6__HREADY_), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_M_macop_MAC_[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__3_ ( .D(
        j202_soc_core_j22_cpu_ml_N194), .DE(j202_soc_core_ahbcs_6__HREADY_), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_M_macop_MAC_[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_M_macop_reg_MAC__1_ ( .D(
        j202_soc_core_j22_cpu_ml_N192), .DE(j202_soc_core_ahbcs_6__HREADY_), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__1_ ( .D(
        j202_soc_core_j22_cpu_ml_N153), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__2_ ( .D(
        j202_soc_core_j22_cpu_ml_N154), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__0_ ( .D(
        j202_soc_core_j22_cpu_ml_N152), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_X_macop_reg_MAC__3_ ( .D(
        j202_soc_core_j22_cpu_ml_N155), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_6_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[6]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_7_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[7]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_6_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[6]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ml_N303), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[0]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[0]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__0_ ( .D(
        n25341), .DE(n25488), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_0_ ( 
        .D(j202_soc_core_qspi_wb_wdat[0]), .CLK(wb_clk_i), .RESET_B(n25732), 
        .Q(j202_soc_core_bldc_core_00_wdata[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_0_ ( .D(n85), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_uart_din_i[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__0_ ( .D(
        j202_soc_core_uart_din_i[0]), .DE(j202_soc_core_uart_TOP_tx_fifo_N32), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__0_ ( .D(
        j202_soc_core_uart_din_i[0]), .DE(j202_soc_core_uart_TOP_tx_fifo_N31), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__0_ ( .D(
        j202_soc_core_uart_din_i[0]), .DE(j202_soc_core_uart_TOP_tx_fifo_N30), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__0_ ( .D(
        j202_soc_core_uart_din_i[0]), .DE(j202_soc_core_uart_TOP_tx_fifo_N29), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_0_ ( 
        .D(j202_soc_core_qspi_wb_wdat[0]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_0_ ( 
        .D(n84), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_cmt_core_00_const1[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_0_ ( 
        .D(n83), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_cmt_core_00_const0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_0_ ( 
        .D(n82), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_cmt_core_00_cks1[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_0_ ( 
        .D(n81), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_cmt_core_00_cks0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmstr_reg_reg_o_reg_0_ ( 
        .D(n80), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_cmt_core_00_str0) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ml_N304), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[1]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[1]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ml_N305), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[2]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[2]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__2_ ( .D(
        n25360), .DE(n25488), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_2_ ( 
        .D(j202_soc_core_qspi_wb_wdat[2]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_bldc_core_00_wdata[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_2_ ( .D(n79), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_uart_din_i[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__2_ ( .D(
        j202_soc_core_uart_din_i[2]), .DE(j202_soc_core_uart_TOP_tx_fifo_N32), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__2_ ( .D(
        j202_soc_core_uart_din_i[2]), .DE(j202_soc_core_uart_TOP_tx_fifo_N31), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__2_ ( .D(
        j202_soc_core_uart_din_i[2]), .DE(j202_soc_core_uart_TOP_tx_fifo_N30), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__2_ ( .D(
        j202_soc_core_uart_din_i[2]), .DE(j202_soc_core_uart_TOP_tx_fifo_N29), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_2_ ( 
        .D(j202_soc_core_qspi_wb_wdat[2]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_2_ ( 
        .D(n78), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_cmt_core_00_const1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_2_ ( 
        .D(n77), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_cmt_core_00_const0[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_2_ ( 
        .D(n76), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_2_ ( 
        .D(n75), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ml_N306), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[3]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[3]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_4_ ( .D(
        j202_soc_core_j22_cpu_ml_N307), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_4_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[4]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_4_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[4]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_5_ ( .D(
        j202_soc_core_j22_cpu_ml_N308), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_5_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[5]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_5_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[5]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_7_ ( .D(
        j202_soc_core_j22_cpu_ml_N310), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_7_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[7]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_9_ ( .D(
        j202_soc_core_j22_cpu_ml_N312), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_9_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[9]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_9_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[9]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_13_ ( .D(
        j202_soc_core_j22_cpu_ml_N316), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_13_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[13]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_13_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[13]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_20_ ( .D(
        j202_soc_core_j22_cpu_ml_N359), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_4_ ( .D(
        j202_soc_core_j22_cpu_ml_N416), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_21_ ( .D(
        j202_soc_core_j22_cpu_ml_N360), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_5_ ( .D(
        j202_soc_core_j22_cpu_ml_N417), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_23_ ( .D(
        j202_soc_core_j22_cpu_ml_N362), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_7_ ( .D(
        j202_soc_core_j22_cpu_ml_N419), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_25_ ( .D(
        j202_soc_core_j22_cpu_ml_N364), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_9_ ( .D(
        j202_soc_core_j22_cpu_ml_N421), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_26_ ( .D(
        j202_soc_core_j22_cpu_ml_N365), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_28_ ( .D(
        j202_soc_core_j22_cpu_ml_N367), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_30_ ( .D(
        j202_soc_core_j22_cpu_ml_N369), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_19_ ( .D(
        j202_soc_core_j22_cpu_ml_N357), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_3_ ( .D(
        j202_soc_core_j22_cpu_ml_N415), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_18_ ( .D(
        j202_soc_core_j22_cpu_ml_N356), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_2_ ( .D(
        j202_soc_core_j22_cpu_ml_N414), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3364), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3328), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3289), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2697), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2734), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[49]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2771), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[81]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2808), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[113]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2845), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[145]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2882), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[177]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2919), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[209]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2956), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[241]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N2993), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[273]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3030), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[305]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3067), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[337]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3104), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[369]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3141), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[401]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3178), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[433]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3215), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[465]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__17_ ( .D(
        j202_soc_core_j22_cpu_rf_N3252), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[497]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_17_ ( .D(n25430), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3366), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3330), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3291), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2699), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2736), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[51]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2773), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[83]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2810), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[115]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2847), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[147]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2884), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[179]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2921), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[211]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2958), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[243]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N2995), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[275]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3032), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[307]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3069), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[339]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3106), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[371]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3143), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[403]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3180), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[435]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3217), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[467]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__19_ ( .D(
        j202_soc_core_j22_cpu_rf_N3254), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[499]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_19_ ( .D(n25473), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3375), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3339), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3300), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2708), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2745), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[59]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2782), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[91]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2819), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[123]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2856), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[155]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2893), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[187]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2930), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[219]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N2967), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[251]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3004), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[283]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3041), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[315]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3078), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[347]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3115), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[379]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3152), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[411]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3189), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[443]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3226), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[475]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__27_ ( .D(
        j202_soc_core_j22_cpu_rf_N3263), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[507]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_27_ ( .D(n25447), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_27_ ( .D(
        j202_soc_core_j22_cpu_ml_N366), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_27_ ( .D(
        j202_soc_core_j22_cpu_rf_N325), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3357), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3322), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3282), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2690), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2727), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[43]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2764), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[75]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2801), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[107]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2838), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[139]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2875), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[171]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2912), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[203]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2949), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[235]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N2986), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[267]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3023), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[299]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3060), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[331]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3097), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[363]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3134), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[395]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3171), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[427]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3208), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[459]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__11_ ( .D(
        j202_soc_core_j22_cpu_rf_N3245), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[491]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_11_ ( .D(n25472), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3358), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3323), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3283), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2691), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2728), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[44]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2765), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[76]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2802), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[108]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2839), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[140]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2876), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[172]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2913), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[204]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2950), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[236]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2987), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[268]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3024), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[300]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3061), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[332]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3098), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[364]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3135), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[396]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3172), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[428]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3209), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[460]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__12_ ( .D(
        j202_soc_core_j22_cpu_rf_N3246), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[492]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_12_ ( .D(
        j202_soc_core_j22_cpu_rf_N2655), .DE(n25489), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3360), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3325), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3286), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2694), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2731), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[46]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2768), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[78]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2805), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[110]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2842), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[142]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2879), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[174]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2916), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[206]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2953), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[238]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N2990), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[270]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3027), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[302]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3064), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[334]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3101), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[366]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3138), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[398]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3175), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[430]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3212), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[462]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__14_ ( .D(
        j202_soc_core_j22_cpu_rf_N3249), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[494]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_14_ ( .D(n25471), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3369), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3334), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3295), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2703), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2740), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[54]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2777), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[86]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2814), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[118]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2851), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[150]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2888), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[182]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2925), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[214]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2962), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[246]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N2999), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[278]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3036), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[310]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3073), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[342]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3110), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[374]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3147), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[406]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3184), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[438]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3221), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[470]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__22_ ( .D(
        j202_soc_core_j22_cpu_rf_N3258), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[502]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_22_ ( .D(n25470), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_22_ ( .D(
        j202_soc_core_j22_cpu_ml_N361), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_22_ ( .D(
        j202_soc_core_j22_cpu_rf_N320), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3372), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3336), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3297), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2705), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2742), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[56]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2779), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[88]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2816), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[120]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2853), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[152]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2890), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[184]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2927), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[216]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N2964), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[248]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3001), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[280]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3038), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[312]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3075), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[344]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3112), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[376]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3149), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[408]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3186), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[440]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3223), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[472]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__24_ ( .D(
        j202_soc_core_j22_cpu_rf_N3260), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[504]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_24_ ( .D(n25469), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_24_ ( .D(
        j202_soc_core_j22_cpu_ml_N363), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_24_ ( .D(
        j202_soc_core_j22_cpu_rf_N322), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3354), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3318), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3279), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2687), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2724), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[40]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2761), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[72]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2798), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[104]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2835), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[136]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2872), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[168]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2909), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[200]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2946), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[232]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N2983), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[264]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3020), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[296]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3057), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[328]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3094), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[360]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3131), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[392]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3168), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[424]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3205), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[456]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__8_ ( .D(
        j202_soc_core_j22_cpu_rf_N3242), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[488]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_8_ ( .D(n25468), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3356), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3321), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3281), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2689), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2726), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[42]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2763), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[74]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2800), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[106]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2837), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[138]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2874), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[170]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2911), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[202]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2948), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[234]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2985), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[266]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3022), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[298]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3059), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[330]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3096), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[362]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3133), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[394]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3170), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[426]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3207), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[458]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__10_ ( .D(
        j202_soc_core_j22_cpu_rf_N3244), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[490]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N2653), .DE(n25489), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_10_ ( .D(
        j202_soc_core_j22_cpu_ml_N313), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_10_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[10]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_10_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[10]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_10_ ( .D(
        j202_soc_core_j22_cpu_ml_N422), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_10_ ( .D(
        j202_soc_core_j22_cpu_rf_N308), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_10_ ( 
        .D(n25373), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_10_ ( .D(
        n25373), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3363), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3327), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3288), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2696), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2733), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[48]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2770), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[80]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2807), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[112]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2844), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[144]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2881), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[176]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2918), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[208]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2955), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[240]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2992), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[272]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3029), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[304]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3066), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[336]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3103), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[368]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3140), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[400]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3177), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[432]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3214), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[464]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__16_ ( .D(
        j202_soc_core_j22_cpu_rf_N3251), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[496]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_16_ ( .D(
        j202_soc_core_j22_cpu_rf_N2660), .DE(n25489), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_tmp[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3361), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3326), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3287), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2695), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2732), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[47]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2769), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[79]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2806), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[111]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2843), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[143]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2880), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[175]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2917), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[207]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2954), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[239]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N2991), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[271]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3028), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[303]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3065), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[335]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3102), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[367]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3139), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[399]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3176), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[431]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3213), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[463]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__15_ ( .D(
        j202_soc_core_j22_cpu_rf_N3250), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[495]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_15_ ( .D(n25467), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_15_ ( .D(
        j202_soc_core_j22_cpu_ml_N318), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_15_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[15]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_15_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[15]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_18_ ( .D(
        j202_soc_core_j22_cpu_ml_N321), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_18_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[18]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_18_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[18]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_19_ ( .D(
        j202_soc_core_j22_cpu_ml_N322), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_19_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[19]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_19_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[19]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_20_ ( .D(
        j202_soc_core_j22_cpu_ml_N324), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_20_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[20]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_20_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[20]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_21_ ( .D(
        j202_soc_core_j22_cpu_ml_N325), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_21_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[21]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_21_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[21]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_22_ ( .D(
        j202_soc_core_j22_cpu_ml_N326), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_22_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[22]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_22_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[22]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__22_ ( 
        .D(n25352), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[22]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_22_ ( 
        .D(j202_soc_core_qspi_wb_wdat[22]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_bldc_core_00_wdata[22]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_6_ ( .D(n74), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_uart_div1[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_23_ ( .D(
        j202_soc_core_j22_cpu_ml_N327), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_23_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[23]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_23_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[23]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_24_ ( .D(
        j202_soc_core_j22_cpu_ml_N328), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_24_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[24]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_24_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[24]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_25_ ( .D(
        j202_soc_core_j22_cpu_ml_N329), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_25_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[25]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_25_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[25]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_26_ ( .D(
        j202_soc_core_j22_cpu_ml_N330), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_26_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[26]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_26_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[26]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__26_ ( 
        .D(n25356), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[26]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_2_ ( .D(n73), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_uart_div0[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_27_ ( .D(
        j202_soc_core_j22_cpu_ml_N331), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_27_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[27]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_27_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[27]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_28_ ( .D(
        j202_soc_core_j22_cpu_ml_N332), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_28_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[28]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_28_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[28]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_29_ ( .D(
        j202_soc_core_j22_cpu_ml_N333), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_29_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[29]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_29_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[29]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__29_ ( 
        .D(n25359), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[29]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_5_ ( .D(n72), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_uart_div0[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_30_ ( .D(
        j202_soc_core_j22_cpu_ml_N334), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_30_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[30]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_30_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[30]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_31_ ( .D(
        j202_soc_core_j22_cpu_ml_N335), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_31_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[31]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_31_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[31]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_32_ ( .D(
        j202_soc_core_j22_cpu_ml_N336), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[32]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_15_ ( .D(
        j202_soc_core_j22_cpu_rf_N313), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__31_ ( 
        .D(n25362), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[31]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_7_ ( .D(n71), .CLK(
        wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_uart_div0[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_3_ ( .D(
        j202_soc_core_wbqspiflash_00_N727), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_9_ ( 
        .D(j202_soc_core_wbqspiflash_00_N623), .DE(
        j202_soc_core_wbqspiflash_00_N751), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_reset_counter[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_N614), .DE(
        j202_soc_core_wbqspiflash_00_N751), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_reset_counter[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_8_ ( 
        .D(j202_soc_core_wbqspiflash_00_N622), .DE(
        j202_soc_core_wbqspiflash_00_N751), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_reset_counter[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_N621), .DE(
        j202_soc_core_wbqspiflash_00_N751), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_reset_counter[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_N620), .DE(
        j202_soc_core_wbqspiflash_00_N751), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_reset_counter[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_N619), .DE(
        j202_soc_core_wbqspiflash_00_N751), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_reset_counter[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_N618), .DE(
        j202_soc_core_wbqspiflash_00_N751), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_reset_counter[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_N617), .DE(
        j202_soc_core_wbqspiflash_00_N751), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_reset_counter[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_N616), .DE(
        j202_soc_core_wbqspiflash_00_N751), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_reset_counter[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_reset_counter_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_N615), .DE(
        j202_soc_core_wbqspiflash_00_N751), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_reset_counter[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_alt_ctrl_reg ( .D(
        j202_soc_core_wbqspiflash_00_N86), .DE(n25734), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_alt_ctrl) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_alt_cmd_reg ( .D(
        j202_soc_core_wbqspiflash_00_N85), .DE(n25734), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_alt_cmd) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_ctrl_reg ( .D(
        j202_soc_core_wbqspiflash_00_N744), .DE(
        j202_soc_core_wbqspiflash_00_N743), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_ctrl) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_wr_reg ( .D(
        j202_soc_core_wbqspiflash_00_N734), .DE(
        j202_soc_core_wbqspiflash_00_N733), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_wr) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_0_ ( 
        .D(j202_soc_core_qspi_wb_addr[2]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_18_ ( 
        .D(j202_soc_core_qspi_wb_addr[20]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_16_ ( 
        .D(j202_soc_core_qspi_wb_addr[18]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_15_ ( 
        .D(j202_soc_core_qspi_wb_addr[17]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_14_ ( 
        .D(j202_soc_core_qspi_wb_addr[16]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_12_ ( 
        .D(j202_soc_core_qspi_wb_addr[14]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_11_ ( 
        .D(j202_soc_core_qspi_wb_addr[13]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_8_ ( 
        .D(j202_soc_core_qspi_wb_addr[10]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_7_ ( 
        .D(j202_soc_core_qspi_wb_addr[9]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_5_ ( 
        .D(j202_soc_core_qspi_wb_addr[7]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_4_ ( 
        .D(j202_soc_core_qspi_wb_addr[6]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_3_ ( 
        .D(j202_soc_core_qspi_wb_addr[5]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_2_ ( 
        .D(j202_soc_core_qspi_wb_addr[4]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_1_ ( 
        .D(j202_soc_core_qspi_wb_addr[3]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_state_reg_4_ ( .D(
        j202_soc_core_wbqspiflash_00_N728), .DE(
        j202_soc_core_wbqspiflash_00_N723), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_state[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_spd_reg ( .D(
        j202_soc_core_wbqspiflash_00_N592), .DE(
        j202_soc_core_wbqspiflash_00_N746), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_spd) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_spd_reg ( 
        .D(j202_soc_core_wbqspiflash_00_spi_spd), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N423), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_mod_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N356), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N354), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N358), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_interrupt_reg ( .D(
        j202_soc_core_wbqspiflash_00_N741), .DE(
        j202_soc_core_wbqspiflash_00_N740), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_int) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N23), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[20])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N323), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N359), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N324), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N360), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N325), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N361), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N326), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N362), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N327), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N363), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N328), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N364), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N329), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N365), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N330), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_8_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N366), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_8_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N331), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_9_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N367), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_9_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N332), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_10_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N368), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_10_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N333), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_11_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N369), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_11_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N334), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_12_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N370), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_12_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N335), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_13_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N371), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_13_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N336), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_14_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N372), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_14_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N337), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_15_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N373), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_15_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N338), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_16_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N374), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_16_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N339), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_17_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N375), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_17_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N340), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_18_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N376), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_18_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N341), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_19_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N377), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_19_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N342), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_20_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N378), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_20_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N343), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_21_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N379), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_21_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N344), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_22_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N380), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_22_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N345), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_23_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N381), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_23_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N346), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_24_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N382), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_24_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N347), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_25_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N383), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_25_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N348), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_26_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N384), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_26_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N349), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_27_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N385), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_27_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N350), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_28_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N386), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_28_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N351), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_29_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N387), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_29_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N352), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_30_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N388), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_input_reg_30_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N353), .DE(n25528), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_input[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_word_reg_31_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N389), .DE(n25529), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_out[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_dir_reg ( .D(
        j202_soc_core_wbqspiflash_00_N594), .DE(
        j202_soc_core_wbqspiflash_00_N747), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_dir) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_dir_reg ( 
        .D(j202_soc_core_wbqspiflash_00_spi_dir), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N423), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_r_dir) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_mod_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N355), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N354), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_cmd_reg ( .D(
        j202_soc_core_wbqspiflash_00_N663), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_cmd) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_31_ ( 
        .D(j202_soc_core_qspi_wb_wdat[31]), .DE(n25493), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_29_ ( 
        .D(j202_soc_core_qspi_wb_wdat[29]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_26_ ( 
        .D(j202_soc_core_qspi_wb_wdat[26]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_23_ ( 
        .D(j202_soc_core_qspi_wb_wdat[23]), .DE(n25493), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_22_ ( 
        .D(j202_soc_core_qspi_wb_wdat[22]), .DE(n25493), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_21_ ( 
        .D(j202_soc_core_qspi_wb_wdat[21]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_N718), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_20_ ( 
        .D(j202_soc_core_qspi_wb_wdat[20]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_N717), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_18_ ( 
        .D(j202_soc_core_qspi_wb_wdat[18]), .DE(n25493), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_N715), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_15_ ( 
        .D(j202_soc_core_qspi_wb_wdat[15]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_N712), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_14_ ( 
        .D(j202_soc_core_qspi_wb_wdat[14]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_N711), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_13_ ( 
        .D(j202_soc_core_qspi_wb_wdat[13]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_12_ ( 
        .D(j202_soc_core_qspi_wb_wdat[12]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_10_ ( 
        .D(j202_soc_core_qspi_wb_wdat[10]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_8_ ( 
        .D(j202_soc_core_qspi_wb_wdat[8]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_7_ ( 
        .D(j202_soc_core_qspi_wb_wdat[7]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_6_ ( 
        .D(j202_soc_core_qspi_wb_wdat[6]), .DE(n25493), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_6_ ( .D(
        n10528), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_5_ ( 
        .D(j202_soc_core_qspi_wb_wdat[5]), .DE(n25493), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_4_ ( 
        .D(j202_soc_core_qspi_wb_wdat[4]), .DE(n25493), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_4_ ( .D(
        n10530), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_3_ ( 
        .D(j202_soc_core_qspi_wb_wdat[3]), .DE(n25493), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_2_ ( 
        .D(j202_soc_core_qspi_wb_wdat[2]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_2_ ( .D(
        n10532), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_0_ ( 
        .D(j202_soc_core_qspi_wb_wdat[0]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_0_ ( .D(
        j202_soc_core_wbqspiflash_00_N628), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_N611), .DE(
        j202_soc_core_wbqspiflash_00_N750), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_N612), .DE(
        j202_soc_core_wbqspiflash_00_N750), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_N605), .DE(
        j202_soc_core_wbqspiflash_00_N749), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_N607), .DE(
        j202_soc_core_wbqspiflash_00_N749), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_N608), .DE(
        j202_soc_core_wbqspiflash_00_N749), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_N609), .DE(
        j202_soc_core_wbqspiflash_00_N749), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_N613), .DE(
        j202_soc_core_wbqspiflash_00_N749), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_N667), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_3_ ( .D(
        n10531), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_29_ ( 
        .D(j202_soc_core_wbqspiflash_00_N696), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_31_ ( 
        .D(j202_soc_core_wbqspiflash_00_N698), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_15_ ( 
        .D(n25261), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_13_ ( 
        .D(j202_soc_core_qspi_wb_addr[15]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_15_ ( .D(
        n25261), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3365), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3329), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3290), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2698), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2735), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[50]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2772), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[82]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2809), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[114]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2846), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[146]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2883), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[178]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2920), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[210]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2957), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[242]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N2994), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[274]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3031), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[306]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3068), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[338]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3105), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[370]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3142), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[402]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3179), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[434]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3216), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[466]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__18_ ( .D(
        j202_soc_core_j22_cpu_rf_N3253), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[498]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_18_ ( .D(n25466), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_16_ ( .D(
        j202_soc_core_j22_cpu_ml_N319), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_16_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[16]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_16_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[16]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_16_ ( .D(
        j202_soc_core_j22_cpu_ml_N354), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_0_ ( .D(
        j202_soc_core_j22_cpu_ml_N412), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_16_ ( .D(
        j202_soc_core_j22_cpu_rf_N314), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__16_ ( 
        .D(n25346), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[16]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_16_ ( 
        .D(j202_soc_core_qspi_wb_wdat[16]), .CLK(wb_clk_i), .RESET_B(n25731), 
        .Q(j202_soc_core_bldc_core_00_wdata[16]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_0_ ( .D(n70), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_uart_div1[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_16_ ( 
        .D(j202_soc_core_qspi_wb_wdat[16]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_N713), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_8_ ( .D(
        j202_soc_core_j22_cpu_ml_N311), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_8_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[8]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_8_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[8]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__q_ ( .D(
        j202_soc_core_j22_cpu_rf_N2638), .DE(j202_soc_core_j22_cpu_rf_N2637), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__q_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_8_ ( .D(
        j202_soc_core_j22_cpu_ml_N420), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_8_ ( .D(
        j202_soc_core_j22_cpu_rf_N306), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__24_ ( 
        .D(n25354), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[24]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_0_ ( .D(n69), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_uart_div0[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_24_ ( 
        .D(j202_soc_core_qspi_wb_wdat[24]), .DE(n25493), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_8_ ( .D(
        n25378), .DE(n11200), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_addr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_6_ ( 
        .D(j202_soc_core_qspi_wb_addr[8]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_8_ ( .D(
        n10526), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_8_ ( .D(
        n25378), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2aqu_00_aquco_reg_CE__0_ ( .D(
        j202_soc_core_ahb2aqu_00_N97), .DE(j202_soc_core_ahb2aqu_00_N95), 
        .CLK(wb_clk_i), .Q(j202_soc_core_aquc_CE__0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_state_reg_1_ ( 
        .D(n25483), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_22_ ( 
        .D(n68), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_21_ ( 
        .D(n67), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_20_ ( 
        .D(n66), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_18_ ( 
        .D(n65), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_16_ ( 
        .D(n64), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_15_ ( 
        .D(n63), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_14_ ( 
        .D(n62), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_13_ ( 
        .D(n61), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_12_ ( 
        .D(n60), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_11_ ( 
        .D(n59), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_period[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_10_ ( 
        .D(n58), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_period[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_8_ ( 
        .D(n57), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_period[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_7_ ( 
        .D(n56), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_period[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_6_ ( 
        .D(n55), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_period[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_5_ ( 
        .D(n54), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_period[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_4_ ( 
        .D(n53), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_period[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_3_ ( 
        .D(n52), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_period[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_2_ ( 
        .D(n51), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_period[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_0_ ( 
        .D(n50), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_period[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_23_ ( 
        .D(n49), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bcr_00_reg_o_reg_0_ ( 
        .D(n48), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_en) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ccr_00_reg_o_reg_0_ ( 
        .D(n47), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_comm[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ccr_00_reg_o_reg_2_ ( 
        .D(n46), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_comm[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_00_reg_o_reg_0_ ( 
        .D(n45), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_wen_1_reg ( 
        .D(n25404), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_wen) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_00_reg_o_reg_0_ ( 
        .D(n44), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_reg_0_ ( 
        .D(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_nxt_latch_status_0_), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bldc_int_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_nxt_bldc_int), 
        .CLK(wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_bldc_int) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[19])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_14_ ( .D(
        j202_soc_core_j22_cpu_ml_N317), .DE(j202_soc_core_j22_cpu_ml_N323), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_ml_bufa[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_14_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[14]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_14_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[14]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_14_ ( .D(
        j202_soc_core_j22_cpu_ml_N426), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_14_ ( .D(
        j202_soc_core_j22_cpu_rf_N312), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__30_ ( 
        .D(n25361), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[30]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_6_ ( .D(n43), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_uart_div0[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_30_ ( 
        .D(j202_soc_core_qspi_wb_wdat[30]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3367), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3331), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3292), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2700), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2737), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[52]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2774), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[84]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2811), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[116]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2848), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[148]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2885), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[180]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2922), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[212]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2959), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[244]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N2996), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[276]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3033), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[308]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3070), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[340]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3107), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[372]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3144), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[404]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3181), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[436]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3218), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[468]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__20_ ( .D(
        j202_soc_core_j22_cpu_rf_N3255), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[500]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_20_ ( .D(n25465), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_12_ ( .D(
        j202_soc_core_j22_cpu_ml_N315), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_12_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[12]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_12_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[12]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_12_ ( .D(
        j202_soc_core_j22_cpu_ml_N424), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_12_ ( .D(
        j202_soc_core_j22_cpu_rf_N310), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__28_ ( 
        .D(n25358), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[28]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_4_ ( .D(n42), .CLK(
        wb_clk_i), .RESET_B(n25734), .Q(j202_soc_core_uart_div0[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_28_ ( 
        .D(j202_soc_core_qspi_wb_wdat[28]), .DE(n25493), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_02_state_reg_0_ ( .D(n25436), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2apb_02_state[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_02_state_reg_2_ ( .D(n25487), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2apb_02_state[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_02_state_reg_1_ ( .D(n25486), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2apb_02_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_2_ ( 
        .D(n25339), .DE(n10559), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_0_ ( .D(
        n25446), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_hsize_buf_reg_1_ ( .D(
        n25428), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_02_hsize_buf[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_hsize_buf_reg_0_ ( .D(
        n25445), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_02_hsize_buf[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_hwrite_buf_reg ( .D(
        n25444), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_pwrite[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_7_ ( .D(
        n25443), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_6_ ( .D(
        n25442), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_5_ ( .D(
        n25441), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_4_ ( .D(
        n25440), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_3_ ( .D(
        n25439), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_2_ ( .D(
        n25438), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_haddr_buf_reg_1_ ( .D(
        n25437), .DE(j202_soc_core_ahb2apb_02_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_reg_addr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_31_ ( 
        .D(n25389), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_30_ ( 
        .D(n25284), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_29_ ( 
        .D(n25296), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_28_ ( 
        .D(n25395), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_26_ ( 
        .D(n25282), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_24_ ( 
        .D(n25264), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_23_ ( 
        .D(n25292), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_22_ ( 
        .D(n25289), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_21_ ( 
        .D(n25283), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_20_ ( 
        .D(n25265), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_18_ ( 
        .D(n25285), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_16_ ( 
        .D(n25266), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_15_ ( 
        .D(n25262), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_12_ ( 
        .D(n25267), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_10_ ( 
        .D(n25263), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_8_ ( 
        .D(n25268), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_7_ ( 
        .D(n25297), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_6_ ( 
        .D(n25298), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_5_ ( 
        .D(n25294), .DE(n25532), .CLK(wb_clk_i), .Q(gpio_en_o[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_4_ ( 
        .D(n25269), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_2_ ( 
        .D(n25286), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_0_ ( 
        .D(n25270), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_31_ ( 
        .D(n25389), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_30_ ( 
        .D(n25284), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_29_ ( 
        .D(n25296), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_28_ ( 
        .D(n25395), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_26_ ( 
        .D(n25282), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_24_ ( 
        .D(n25264), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_23_ ( 
        .D(n25292), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_22_ ( 
        .D(n25289), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_21_ ( 
        .D(n25283), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_20_ ( 
        .D(n25265), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_18_ ( 
        .D(n25285), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_16_ ( 
        .D(n25266), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_15_ ( 
        .D(n25262), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_12_ ( 
        .D(n25267), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_10_ ( 
        .D(n25263), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_8_ ( 
        .D(n25268), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_7_ ( 
        .D(n25297), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_6_ ( 
        .D(n25298), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_5_ ( 
        .D(n25294), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_4_ ( 
        .D(n25269), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_2_ ( 
        .D(n25286), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_0_ ( 
        .D(n25270), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_31_ ( 
        .D(n25389), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_30_ ( 
        .D(n25284), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_29_ ( 
        .D(n25296), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_28_ ( 
        .D(n25395), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_26_ ( 
        .D(n25282), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_24_ ( 
        .D(n25264), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_23_ ( 
        .D(n25292), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_22_ ( 
        .D(n25289), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_21_ ( 
        .D(n25283), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_20_ ( 
        .D(n25265), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_18_ ( 
        .D(n25285), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_16_ ( 
        .D(n25266), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_15_ ( 
        .D(n25262), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_12_ ( 
        .D(n25267), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_10_ ( 
        .D(n25263), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_8_ ( 
        .D(n25268), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_7_ ( 
        .D(n25297), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_6_ ( 
        .D(n25298), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_5_ ( 
        .D(n25294), .DE(n25533), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_4_ ( 
        .D(n25269), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_2_ ( 
        .D(n25286), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_0_ ( 
        .D(n25270), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_10_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N50), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_15_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N55), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_31_ ( 
        .D(n25389), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_31_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N71), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_31_ ( .D(
        j202_soc_core_ahb2apb_02_N159), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[63]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_30_ ( 
        .D(n25284), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_30_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N70), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_30_ ( .D(
        j202_soc_core_ahb2apb_02_N158), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[62]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_29_ ( 
        .D(n25296), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_29_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N69), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_29_ ( .D(
        j202_soc_core_ahb2apb_02_N157), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[61]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_28_ ( 
        .D(n25395), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_28_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N68), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_28_ ( .D(
        j202_soc_core_ahb2apb_02_N156), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[60]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_26_ ( 
        .D(n25282), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_26_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N66), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_26_ ( .D(
        j202_soc_core_ahb2apb_02_N154), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[58]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_24_ ( 
        .D(n25264), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_24_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N64), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_24_ ( .D(
        j202_soc_core_ahb2apb_02_N152), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[56]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_23_ ( 
        .D(n25292), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_23_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N63), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_23_ ( .D(
        j202_soc_core_ahb2apb_02_N151), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[55]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_22_ ( 
        .D(n25289), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_22_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N62), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_22_ ( .D(
        j202_soc_core_ahb2apb_02_N150), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[54]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_21_ ( 
        .D(n25283), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_21_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N61), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_21_ ( .D(
        j202_soc_core_ahb2apb_02_N149), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[53]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_20_ ( 
        .D(n25265), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_20_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N60), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_20_ ( .D(
        j202_soc_core_ahb2apb_02_N148), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[52]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_18_ ( 
        .D(n25285), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_18_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N58), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_18_ ( .D(
        j202_soc_core_ahb2apb_02_N146), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[50]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_16_ ( 
        .D(n25266), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_16_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N56), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_16_ ( .D(
        j202_soc_core_ahb2apb_02_N144), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[48]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_12_ ( 
        .D(n25267), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_12_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N52), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_12_ ( .D(
        j202_soc_core_ahb2apb_02_N140), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[44]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_8_ ( 
        .D(n25268), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_8_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N48), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_8_ ( .D(
        j202_soc_core_ahb2apb_02_N136), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[40]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_7_ ( 
        .D(n25297), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_7_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N47), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_7_ ( .D(
        j202_soc_core_ahb2apb_02_N135), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[39]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_6_ ( 
        .D(n25298), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_6_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N46), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_6_ ( .D(
        j202_soc_core_ahb2apb_02_N134), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[38]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_5_ ( 
        .D(n25294), .DE(n25534), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_5_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N45), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_5_ ( .D(
        j202_soc_core_ahb2apb_02_N133), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[37]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_4_ ( 
        .D(n25269), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_4_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N44), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_4_ ( .D(
        j202_soc_core_ahb2apb_02_N132), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[36]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_2_ ( 
        .D(n25286), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_2_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N42), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_2_ ( .D(
        j202_soc_core_ahb2apb_02_N130), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[34]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_0_ ( 
        .D(n25270), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N40), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_02_N128), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[32]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel_reg_1_ ( 
        .D(n25340), .DE(n10559), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_01_state_reg_0_ ( .D(n25463), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2apb_01_state[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_01_state_reg_2_ ( .D(n25485), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2apb_01_state[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_ahb2apb_01_state_reg_1_ ( .D(n25484), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahb2apb_01_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_0_ ( .D(
        n25462), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_hsize_buf_reg_1_ ( .D(
        n25429), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_01_hsize_buf[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_hsize_buf_reg_0_ ( .D(
        n25461), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahb2apb_01_hsize_buf[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_hwrite_buf_reg ( .D(
        n25460), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_pwrite[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_10_ ( .D(
        n25459), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_9_ ( .D(
        n25458), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_8_ ( .D(
        n25457), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_7_ ( .D(
        n25456), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_6_ ( .D(
        n25455), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_5_ ( .D(
        n25454), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_4_ ( .D(
        n25453), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_3_ ( .D(
        n25452), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_2_ ( .D(
        n25451), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_1_ ( .D(
        n25450), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_6_ ( .D(
        n25322), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_2_ ( .D(
        n25320), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_12_ ( 
        .D(n25272), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_10_ ( 
        .D(j202_soc_core_qspi_wb_addr[12]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_12_ ( .D(
        n25272), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_4_ ( .D(
        n25327), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_11_ ( .D(
        j202_soc_core_j22_cpu_ml_N314), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_11_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[11]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_11_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[11]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_11_ ( .D(
        j202_soc_core_j22_cpu_ml_N423), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_11_ ( .D(
        j202_soc_core_j22_cpu_rf_N309), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__27_ ( 
        .D(n25357), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[27]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div0_reg_3_ ( .D(n41), .CLK(
        wb_clk_i), .RESET_B(n25734), .Q(j202_soc_core_uart_div0[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_clr_reg ( .D(
        j202_soc_core_uart_BRG_N21), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps_clr) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_0_ ( .D(
        j202_soc_core_uart_BRG_N12), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_1_ ( .D(
        j202_soc_core_uart_BRG_N13), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_2_ ( .D(
        j202_soc_core_uart_BRG_N14), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_3_ ( .D(
        j202_soc_core_uart_BRG_N15), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_4_ ( .D(
        j202_soc_core_uart_BRG_N16), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_5_ ( .D(
        j202_soc_core_uart_BRG_N17), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_6_ ( .D(
        j202_soc_core_uart_BRG_N18), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_ps_reg_7_ ( .D(
        j202_soc_core_uart_BRG_N19), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_ps[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_27_ ( 
        .D(j202_soc_core_qspi_wb_wdat[27]), .DE(n25493), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_27_ ( 
        .D(n25291), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_27_ ( 
        .D(n25291), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_27_ ( 
        .D(n25291), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_27_ ( 
        .D(n25291), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_27_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N67), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_27_ ( .D(
        j202_soc_core_ahb2apb_02_N155), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[59]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_haddr_buf_reg_11_ ( .D(
        n25449), .DE(j202_soc_core_ahb2apb_01_N22), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_bs_addr[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_15__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_15__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N18), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[15])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_14__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_14__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N17), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[14])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_13__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_13__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N16), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[13])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_12__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_12__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N15), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[12])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_11__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_11__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N14), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[11])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_10__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_10__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N13), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[10])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_9__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_9__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N12), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_8__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_8__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N11), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_7__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_7__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N10), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_6__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_6__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N9), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_5__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_5__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N8), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_4__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_4__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N7), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_3__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_3__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N6), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_2__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_2__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N5), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_1__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_1__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N4), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_sint_label_0__rg_sint_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_0__rg_sint_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_sint[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N3), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[64]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[66]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[67]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[68]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[69]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[70]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[71]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[72]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[74]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[76]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[77]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[78]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[79]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[80]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[82]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[84]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[85]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[86]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[87]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[88]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[90]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[91]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[92]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[93]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[94]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[95]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[96]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[98]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[99]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[100]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[101]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[102]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[103]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[104]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[106]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[108]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[109]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[110]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[111]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[112]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[114]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[116]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[117]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[118]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[119]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[120]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[122]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[123]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[124]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[125]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[126]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[127]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[32]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[34]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[35]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[36]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[37]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[38]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[39]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[40]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[42]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[44]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[45]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[46]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[47]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[48]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[50]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[52]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[53]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[54]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[55]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[56]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[58]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[59]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[60]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[61]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[62]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[63]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[2]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[4]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[6]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[64]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[96]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[33]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[65]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[97]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[66]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[35]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[67]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[99]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[68]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[37]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[69]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[101]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[70]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[102]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[39]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[71]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[103]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[27]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[29]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[24]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[26]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[28]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[30]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[31]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[88]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[120]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[57]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[89]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[121]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[90]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[59]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[91]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[123]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[92]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[61]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[93]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[125]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[94]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[126]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[63]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[95]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[127]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[10]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[12]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[15]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[72]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[104]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[41]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[73]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[105]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[74]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[43]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[75]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[107]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[76]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[45]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[77]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[109]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[78]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[110]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[47]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[79]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[111]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_4_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N7), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_12_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N15), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_20_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N23), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[21]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N3), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[18]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_16_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N19), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[20]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_24_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N27), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_28_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N31), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[23]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_2_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N5), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[80]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_3_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N6), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[112]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_5_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N8), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[49]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_6_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N9), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[81]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_7_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N10), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[113]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_10_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N13), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[82]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[51]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[83]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_15_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N18), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[115]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[84]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_21_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N24), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[53]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_22_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N25), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[85]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_23_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N26), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[117]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_26_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N29), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[86]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_27_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N30), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[118]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_29_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N32), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[55]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_30_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N33), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[87]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_31_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N34), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[119]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_2_ ( .D(
        j202_soc_core_ahb2apb_01_N130), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[66]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_4_ ( .D(
        j202_soc_core_ahb2apb_01_N132), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[68]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_5_ ( .D(
        j202_soc_core_ahb2apb_01_N133), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[69]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_6_ ( .D(
        j202_soc_core_ahb2apb_01_N134), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[70]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_7_ ( .D(
        j202_soc_core_ahb2apb_01_N135), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[71]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_15_ ( .D(
        j202_soc_core_ahb2apb_01_N143), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[79]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_20_ ( .D(
        j202_soc_core_ahb2apb_01_N148), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[84]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_21_ ( .D(
        j202_soc_core_ahb2apb_01_N149), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[85]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_22_ ( .D(
        j202_soc_core_ahb2apb_01_N150), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[86]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_23_ ( .D(
        j202_soc_core_ahb2apb_01_N151), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[87]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_01_N128), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[64]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_10_ ( .D(
        j202_soc_core_ahb2apb_01_N138), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[74]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_24_ ( .D(
        j202_soc_core_ahb2apb_01_N152), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[88]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_26_ ( .D(
        j202_soc_core_ahb2apb_01_N154), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[90]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_27_ ( .D(
        j202_soc_core_ahb2apb_01_N155), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[91]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_28_ ( .D(
        j202_soc_core_ahb2apb_01_N156), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[92]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_29_ ( .D(
        j202_soc_core_ahb2apb_01_N157), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[93]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_30_ ( .D(
        j202_soc_core_ahb2apb_01_N158), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[94]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_31_ ( .D(
        j202_soc_core_ahb2apb_01_N159), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[95]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_13_ ( .D(
        n25332), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[13])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_11_ ( .D(
        n25331), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[11])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_9_ ( .D(
        n25330), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_5_ ( .D(
        n25328), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_3_ ( .D(
        n25325), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_11_ ( 
        .D(n25374), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_9_ ( 
        .D(j202_soc_core_qspi_wb_addr[11]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_bootrom_00_address_w_reg_11_ ( .D(
        n25374), .DE(n25542), .CLK(wb_clk_i), .Q(
        j202_soc_core_bootrom_00_address_w[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_12_ ( .D(
        n25323), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[12])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_10_ ( .D(
        n25317), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[10])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_8_ ( .D(
        n25318), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufa_reg_17_ ( .D(
        j202_soc_core_j22_cpu_ml_N320), .DE(n25537), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufa[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_mach_reg_17_ ( .D(
        j202_soc_core_j22_cpu_ml_machj[17]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_mach[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_j22_cpu_ml_macl_reg_17_ ( .D(
        j202_soc_core_j22_cpu_ml_maclj[17]), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_macl[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_17_ ( .D(
        j202_soc_core_j22_cpu_ml_N355), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_17_ ( .D(
        j202_soc_core_j22_cpu_rf_N315), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_1_ ( .D(
        j202_soc_core_j22_cpu_ml_N413), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_1_ ( .D(
        j202_soc_core_j22_cpu_rf_N299), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_1_ ( .D(
        j202_soc_core_j22_cpu_rf_N3346), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__1_ ( .D(
        n25306), .DE(n25488), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_1_ ( 
        .D(j202_soc_core_qspi_wb_wdat[1]), .CLK(wb_clk_i), .RESET_B(n25732), 
        .Q(j202_soc_core_bldc_core_00_wdata[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ccr_00_reg_o_reg_1_ ( 
        .D(n40), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_comm[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bcr_00_reg_o_reg_1_ ( 
        .D(n39), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_adc_en) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_1_ ( 
        .D(n38), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_pwm_period[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_din_i_reg_1_ ( .D(n37), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_uart_din_i[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_0__1_ ( .D(
        j202_soc_core_uart_din_i[1]), .DE(j202_soc_core_uart_TOP_tx_fifo_N32), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_1__1_ ( .D(
        j202_soc_core_uart_din_i[1]), .DE(j202_soc_core_uart_TOP_tx_fifo_N31), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_2__1_ ( .D(
        j202_soc_core_uart_din_i[1]), .DE(j202_soc_core_uart_TOP_tx_fifo_N30), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_mem_reg_3__1_ ( .D(
        j202_soc_core_uart_din_i[1]), .DE(j202_soc_core_uart_TOP_tx_fifo_N29), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_fifo_mem[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_1_ ( 
        .D(j202_soc_core_qspi_wb_wdat[1]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_1_ ( 
        .D(n36), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_cmt_core_00_const1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_1_ ( 
        .D(n35), .CLK(wb_clk_i), .RESET_B(n25732), .Q(
        j202_soc_core_cmt_core_00_const0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1_reg_reg_o_reg_1_ ( 
        .D(n34), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_cmt_core_00_cks1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0_reg_reg_o_reg_1_ ( 
        .D(n33), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_cmt_core_00_cks0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[0]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[1]), .CLK(wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[2]), .CLK(wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[3]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[4]), .CLK(wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[5]), .CLK(wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[6]), .CLK(wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[7]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[8]), .CLK(wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[9]), .CLK(wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmstr_reg_reg_o_reg_1_ ( 
        .D(n32), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_cmt_core_00_str1) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[9]), .CLK(wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[0]), .CLK(wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[2]), .CLK(wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cnt1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[2]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[3]), .CLK(wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_cmt_core_00_cnt1[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[3]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[4]), .CLK(wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_cmt_core_00_cnt1[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[4]), .CLK(wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[5]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_cmt_core_00_cnt1[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[5]), .CLK(wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[6]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cnt1[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[6]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[7]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cnt1[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[7]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[1]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[2]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[3]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[4]), .CLK(wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[5]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[6]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[7]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[8]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[0]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[8]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cnt1[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[8]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[1]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cnt1[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[1]), .CLK(wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_1_ ( 
        .D(j202_soc_core_qspi_wb_wdat[1]), .DE(n25493), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_1_ ( .D(
        j202_soc_core_wbqspiflash_00_N629), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_quad_mode_enabled_reg ( 
        .D(j202_soc_core_wbqspiflash_00_N739), .DE(
        j202_soc_core_wbqspiflash_00_N738), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_27_ ( 
        .D(j202_soc_core_wbqspiflash_00_N694), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_last_status_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_N606), .DE(
        j202_soc_core_wbqspiflash_00_N749), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_last_status[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[56]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[48]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[40]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[32]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[97]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[65]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[33]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_dout_reg_1_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N4), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_eimk[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_01_N129), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[65]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_1_ ( 
        .D(n25288), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_1_ ( 
        .D(n25288), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_1_ ( 
        .D(n25288), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_1_ ( 
        .D(n25288), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_1_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N41), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_02_N129), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[33]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__17_ ( 
        .D(n25347), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[17]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_17_ ( 
        .D(j202_soc_core_qspi_wb_wdat[17]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_bldc_core_00_wdata[17]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_17_ ( 
        .D(n31), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_17_ ( 
        .D(j202_soc_core_qspi_wb_wdat[17]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_N714), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[60]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[52]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[44]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[36]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[113]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[81]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[49]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_17_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N20), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_17_ ( .D(
        j202_soc_core_ahb2apb_01_N145), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[81]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_17_ ( 
        .D(n25293), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_17_ ( 
        .D(n25293), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_17_ ( 
        .D(n25293), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_17_ ( 
        .D(n25293), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[17]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_17_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N57), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_17_ ( .D(
        j202_soc_core_ahb2apb_02_N145), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[49]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_9_ ( .D(
        j202_soc_core_j22_cpu_rf_N307), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__25_ ( 
        .D(n25355), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_25_ ( 
        .D(j202_soc_core_qspi_wb_wdat[25]), .DE(n25493), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[62]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[54]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[46]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[38]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[121]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[89]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[57]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_25_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N28), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_25_ ( .D(
        j202_soc_core_ahb2apb_01_N153), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[89]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_25_ ( 
        .D(n25290), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_25_ ( 
        .D(n25290), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_25_ ( 
        .D(n25290), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_25_ ( 
        .D(n25290), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[25]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_25_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N65), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_25_ ( .D(
        j202_soc_core_ahb2apb_02_N153), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[57]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__9_ ( .D(
        n25368), .DE(n25488), .CLK(wb_clk_i), .Q(j202_soc_core_qspi_wb_wdat[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_9_ ( 
        .D(j202_soc_core_qspi_wb_wdat[9]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_bldc_core_00_wdata[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_9_ ( 
        .D(n30), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_pwm_period[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_apb_00_pwdata_1_reg_9_ ( 
        .D(j202_soc_core_qspi_wb_wdat[9]), .CLK(wb_clk_i), .RESET_B(n25733), 
        .Q(j202_soc_core_cmt_core_00_wdata_cnt0[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor1_reg_reg_o_reg_9_ ( 
        .D(n29), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_cmt_core_00_const1[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcor0_reg_reg_o_reg_9_ ( 
        .D(n28), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_cmt_core_00_const0[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[9]), .CLK(wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cnt0[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_9_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[9]), .CLK(wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[9]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmf0_o_reg ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt0_to1), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_cmt_core_00_cmf0) );
  sky130_fd_sc_hd__dfstp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[0]), .CLK(wb_clk_i), .SET_B(n25734), .Q(j202_soc_core_cmt_core_00_cnt0[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[0]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[0]), .CLK(wb_clk_i), 
        .RESET_B(n25730), .Q(j202_soc_core_prdata[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_0_ ( .D(
        j202_soc_core_ahb2apb_00_N128), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[96]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[1]), .CLK(wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_cmt_core_00_cnt0[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[1]), .CLK(wb_clk_i), .RESET_B(n25734), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[1]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_1_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[1]), .CLK(wb_clk_i), 
        .RESET_B(n25732), .Q(j202_soc_core_prdata[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_1_ ( .D(
        j202_soc_core_ahb2apb_00_N129), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[97]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[2]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cnt0[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[2]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_2_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[2]), .CLK(wb_clk_i), 
        .RESET_B(n25732), .Q(j202_soc_core_prdata[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_2_ ( .D(
        j202_soc_core_ahb2apb_00_N130), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[98]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[3]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cnt0[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[3]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[3]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_3_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[3]), .CLK(wb_clk_i), 
        .RESET_B(n25732), .Q(j202_soc_core_prdata[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_3_ ( .D(
        j202_soc_core_ahb2apb_00_N131), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[99]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[4]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cnt0[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[4]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[4]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_4_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[4]), .CLK(wb_clk_i), 
        .RESET_B(n25732), .Q(j202_soc_core_prdata[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_4_ ( .D(
        j202_soc_core_ahb2apb_00_N132), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[100])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[5]), .CLK(wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cnt0[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[5]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[5]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_5_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[5]), .CLK(wb_clk_i), 
        .RESET_B(n25732), .Q(j202_soc_core_prdata[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_5_ ( .D(
        j202_soc_core_ahb2apb_00_N133), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[101])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[6]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cnt0[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[6]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[6]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_6_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[6]), .CLK(wb_clk_i), 
        .RESET_B(n25732), .Q(j202_soc_core_prdata[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_6_ ( .D(
        j202_soc_core_ahb2apb_00_N134), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[102])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[7]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cnt0[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[7]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[8]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cnt0[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[8]), .CLK(wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[8]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_8_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[8]), .CLK(wb_clk_i), 
        .RESET_B(n25730), .Q(j202_soc_core_prdata[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_8_ ( .D(
        j202_soc_core_ahb2apb_00_N136), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[104])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[10]), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cnt0[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[10]), .CLK(wb_clk_i), .RESET_B(
        n25733), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[11]), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_cmt_core_00_cnt0[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[11]), .CLK(wb_clk_i), .RESET_B(
        n25730), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[11]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_11_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[11]), .CLK(wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_prdata[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_11_ ( .D(
        j202_soc_core_ahb2apb_00_N139), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[107])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[12]), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_cmt_core_00_cnt0[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[12]), .CLK(wb_clk_i), .RESET_B(
        n25730), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[13]), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cnt0[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[13]), .CLK(wb_clk_i), .RESET_B(
        n25733), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[14]), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cnt0[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[14]), .CLK(wb_clk_i), .RESET_B(
        n25733), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt0_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[15]), .CLK(
        wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_cmt_core_00_cnt0[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cnt0[15]), .CLK(wb_clk_i), .RESET_B(
        n25733), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_9_ ( 
        .D(j202_soc_core_qspi_wb_wdat[9]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_9_ ( .D(
        n10525), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[58]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[50]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[42]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[34]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[105]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[73]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[41]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_9_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N12), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_9_ ( .D(
        j202_soc_core_ahb2apb_01_N137), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[73]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_9_ ( 
        .D(n25275), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_9_ ( 
        .D(n25275), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_9_ ( 
        .D(n25275), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_9_ ( 
        .D(n25275), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[9]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_9_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N49), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_9_ ( .D(
        j202_soc_core_ahb2apb_02_N137), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[41]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pr_reg_21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3368), .DE(j202_soc_core_j22_cpu_rf_N3371), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_pr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_vbr_reg_21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3333), .DE(n25433), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_rf_vbr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gbr_reg_21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3294), .DE(j202_soc_core_j22_cpu_rf_N3301), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gbr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_0__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2702), .DE(j202_soc_core_j22_cpu_rf_N2709), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_1__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2739), .DE(j202_soc_core_j22_cpu_rf_N2746), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[53]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_2__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2776), .DE(j202_soc_core_j22_cpu_rf_N2783), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[85]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_3__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2813), .DE(j202_soc_core_j22_cpu_rf_N2820), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[117]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_4__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2850), .DE(j202_soc_core_j22_cpu_rf_N2857), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[149]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_5__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2887), .DE(j202_soc_core_j22_cpu_rf_N2894), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[181]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_6__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2924), .DE(j202_soc_core_j22_cpu_rf_N2931), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[213]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_7__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2961), .DE(j202_soc_core_j22_cpu_rf_N2968), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[245]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_8__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N2998), .DE(j202_soc_core_j22_cpu_rf_N3005), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[277]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_9__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3035), .DE(j202_soc_core_j22_cpu_rf_N3042), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[309]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_10__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3072), .DE(j202_soc_core_j22_cpu_rf_N3079), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[341]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_11__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3109), .DE(j202_soc_core_j22_cpu_rf_N3116), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[373]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_12__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3146), .DE(j202_soc_core_j22_cpu_rf_N3153), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[405]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_13__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3183), .DE(j202_soc_core_j22_cpu_rf_N3190), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[437]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_14__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3220), .DE(j202_soc_core_j22_cpu_rf_N3227), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[469]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_gpr_reg_15__21_ ( .D(
        j202_soc_core_j22_cpu_rf_N3257), .DE(j202_soc_core_j22_cpu_rf_N3264), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_gpr[501]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_tmp_reg_21_ ( .D(n25464), 
        .DE(n25489), .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rf_tmp[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_3_ ( .D(
        j202_soc_core_ahb2apb_01_N131), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[67]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_3_ ( 
        .D(n25287), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_3_ ( 
        .D(n25287), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_3_ ( 
        .D(n25287), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_3_ ( 
        .D(n25287), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_3_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N43), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_3_ ( .D(
        j202_soc_core_ahb2apb_02_N131), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[35]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ma_ahbc_reg_HWDATA__19_ ( 
        .D(n25349), .DE(n25488), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_wdat[19]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_wb_slave_00_reg_wdata_o_reg_19_ ( 
        .D(j202_soc_core_qspi_wb_wdat[19]), .CLK(wb_clk_i), .RESET_B(n25731), 
        .Q(j202_soc_core_bldc_core_00_wdata[19]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_ppr_00_reg_o_reg_19_ ( 
        .D(n27), .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_bldc_core_00_pwm_duty[7]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld_reg ( 
        .D(n26), .CLK(wb_clk_i), .RESET_B(n25730), .Q(
        j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_div1_reg_3_ ( .D(n25), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_uart_div1[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_19_ ( 
        .D(j202_soc_core_qspi_wb_wdat[19]), .DE(n25493), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_erased_sector_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_N716), .DE(
        j202_soc_core_wbqspiflash_00_N710), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_erased_sector[5]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[124]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[116]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[108]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[100]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[115]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[83]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[51]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_19_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N22), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_19_ ( .D(
        j202_soc_core_ahb2apb_01_N147), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[83]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_19_ ( 
        .D(n25295), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_19_ ( 
        .D(n25295), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_19_ ( 
        .D(n25295), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_19_ ( 
        .D(n25295), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[19]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_19_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N59), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_19_ ( .D(
        j202_soc_core_ahb2apb_02_N147), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[51]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_29_ ( .D(
        j202_soc_core_j22_cpu_ml_N368), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_13_ ( .D(
        j202_soc_core_j22_cpu_ml_N425), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_25_ ( 
        .D(j202_soc_core_wbqspiflash_00_N692), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_24_ ( 
        .D(j202_soc_core_wbqspiflash_00_N691), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_23_ ( 
        .D(j202_soc_core_wbqspiflash_00_N690), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_22_ ( 
        .D(j202_soc_core_wbqspiflash_00_N689), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_21_ ( 
        .D(j202_soc_core_wbqspiflash_00_N688), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_20_ ( 
        .D(j202_soc_core_wbqspiflash_00_N687), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_19_ ( 
        .D(j202_soc_core_wbqspiflash_00_N686), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_18_ ( 
        .D(j202_soc_core_wbqspiflash_00_N685), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_17_ ( 
        .D(j202_soc_core_wbqspiflash_00_N684), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_16_ ( 
        .D(j202_soc_core_wbqspiflash_00_N683), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_15_ ( 
        .D(j202_soc_core_wbqspiflash_00_N682), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_14_ ( 
        .D(j202_soc_core_wbqspiflash_00_N681), .DE(n25536), .CLK(wb_clk_i), 
        .Q(j202_soc_core_ahblite_interconnect_s_hrdata[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_13_ ( 
        .D(j202_soc_core_wbqspiflash_00_N680), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_12_ ( 
        .D(j202_soc_core_wbqspiflash_00_N679), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_11_ ( 
        .D(j202_soc_core_wbqspiflash_00_N678), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_10_ ( 
        .D(j202_soc_core_wbqspiflash_00_N677), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_9_ ( 
        .D(j202_soc_core_wbqspiflash_00_N676), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_8_ ( 
        .D(j202_soc_core_wbqspiflash_00_N675), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_N674), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_N673), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_id_opn_reg_inst__6_ ( .D(
        n25276), .DE(n25434), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_id_opn_inst__6_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_N672), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_N671), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_N670), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_N669), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_o_wb_data_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_N668), .DE(
        j202_soc_core_wbqspiflash_00_N755), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_24_ ( .D(
        n10510), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_25_ ( .D(
        n10509), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_26_ ( .D(
        n10508), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_6_ ( .D(
        j202_soc_core_j22_cpu_ml_N418), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_22_ ( 
        .D(n25277), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_20_ ( 
        .D(j202_soc_core_qspi_wb_addr[22]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[8]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_8_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N11), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_8_ ( .D(
        j202_soc_core_ahb2apb_01_N136), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[72]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_31_ ( .D(
        j202_soc_core_j22_cpu_ml_N370), .DE(n25481), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_15_ ( .D(
        j202_soc_core_j22_cpu_ml_N427), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_ml_bufb_reg_32_ ( .D(
        j202_soc_core_j22_cpu_ml_N429), .DE(n25491), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_ml_bufb[32]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_13_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N16), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_13_ ( .D(
        j202_soc_core_ahb2apb_01_N141), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[77]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_13_ ( 
        .D(n25278), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_13_ ( 
        .D(n25278), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_13_ ( 
        .D(n25278), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_13_ ( 
        .D(n25278), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[13]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_13_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N53), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_13_ ( .D(
        j202_soc_core_ahb2apb_02_N141), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[45]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__4_ ( .D(
        j202_soc_core_uart_TOP_rxr[6]), .DE(j202_soc_core_uart_TOP_rx_fifo_N32), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__3_ ( .D(
        j202_soc_core_uart_TOP_rxr[5]), .DE(j202_soc_core_uart_TOP_rx_fifo_N32), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__2_ ( .D(
        j202_soc_core_uart_TOP_rxr[4]), .DE(j202_soc_core_uart_TOP_rx_fifo_N32), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_rx_fifo_mem_reg_0__1_ ( .D(
        j202_soc_core_uart_TOP_rxr[3]), .DE(j202_soc_core_uart_TOP_rx_fifo_N32), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_rx_fifo_mem[25]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_dpll_state_reg_1_ ( .D(n24), 
        .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_uart_TOP_dpll_state[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_cnt_reg_0_ ( .D(
        j202_soc_core_uart_BRG_N56), .DE(j202_soc_core_uart_BRG_N55), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_BRG_cnt[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_cnt_reg_1_ ( .D(
        j202_soc_core_uart_BRG_N57), .DE(j202_soc_core_uart_BRG_N55), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_BRG_cnt[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_r_reg ( .D(n25399), 
        .CLK(wb_clk_i), .Q(j202_soc_core_uart_BRG_sio_ce_r) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_BRG_sio_ce_reg ( .D(
        j202_soc_core_uart_BRG_N59), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_sio_ce) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_txf_empty_r_reg ( .D(
        j202_soc_core_uart_TOP_N16), .DE(n10676), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_txf_empty_r) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_load_reg ( .D(
        j202_soc_core_uart_TOP_N137), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_load) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_bit_cnt_reg_1_ ( .D(
        j202_soc_core_uart_TOP_N59), .DE(j202_soc_core_uart_TOP_N57), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_bit_cnt[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_bit_cnt_reg_3_ ( .D(
        j202_soc_core_uart_TOP_N61), .DE(j202_soc_core_uart_TOP_N57), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_bit_cnt[3]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_uart_TOP_shift_en_reg ( .D(
        j202_soc_core_uart_TOP_N123), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_shift_en) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_shift_en_r_reg ( .D(n25401), 
        .DE(n10676), .CLK(wb_clk_i), .Q(j202_soc_core_uart_TOP_shift_en_r) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_bit_cnt_reg_0_ ( .D(
        j202_soc_core_uart_TOP_N58), .DE(j202_soc_core_uart_TOP_N57), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_bit_cnt[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_bit_cnt_reg_2_ ( .D(
        j202_soc_core_uart_TOP_N60), .DE(j202_soc_core_uart_TOP_N57), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_tx_bit_cnt[2]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_tx_fifo_rp_reg_0_ ( .D(n23), 
        .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_uart_TOP_tx_fifo_rp[0]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_uart_TOP_tx_fifo_rp_reg_1_ ( .D(n22), 
        .CLK(wb_clk_i), .RESET_B(n25733), .Q(
        j202_soc_core_uart_TOP_tx_fifo_rp[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_tx_fifo_gb_reg ( .D(
        j202_soc_core_uart_TOP_tx_fifo_N42), .DE(
        j202_soc_core_uart_TOP_tx_fifo_N41), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_TOP_tx_fifo_gb) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_8_ ( .D(
        j202_soc_core_uart_TOP_N33), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_7_ ( .D(
        j202_soc_core_uart_TOP_N32), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_6_ ( .D(
        j202_soc_core_uart_TOP_N31), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_5_ ( .D(
        j202_soc_core_uart_TOP_N30), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_4_ ( .D(
        j202_soc_core_uart_TOP_N29), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_3_ ( .D(
        j202_soc_core_uart_TOP_N28), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_2_ ( .D(
        j202_soc_core_uart_TOP_N27), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_1_ ( .D(
        j202_soc_core_uart_TOP_N26), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_hold_reg_reg_0_ ( .D(
        j202_soc_core_uart_TOP_N25), .DE(j202_soc_core_uart_TOP_N24), .CLK(
        wb_clk_i), .Q(j202_soc_core_uart_TOP_hold_reg[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_TOP_txd_o_reg ( .D(
        j202_soc_core_uart_TOP_N43), .DE(n10676), .CLK(wb_clk_i), .Q(io_out[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_0_ ( .D(
        j202_soc_core_uart_BRG_N35), .DE(n10675), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_7_ ( .D(
        j202_soc_core_uart_BRG_N42), .DE(n10675), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_6_ ( .D(
        j202_soc_core_uart_BRG_N41), .DE(n10675), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_5_ ( .D(
        j202_soc_core_uart_BRG_N40), .DE(n10675), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_4_ ( .D(
        j202_soc_core_uart_BRG_N39), .DE(n10675), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_3_ ( .D(
        j202_soc_core_uart_BRG_N38), .DE(n10675), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_2_ ( .D(
        j202_soc_core_uart_BRG_N37), .DE(n10675), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_uart_BRG_br_cnt_reg_1_ ( .D(
        j202_soc_core_uart_BRG_N36), .DE(n10675), .CLK(wb_clk_i), .Q(
        j202_soc_core_uart_BRG_br_cnt[1]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_14_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N17), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_14_ ( .D(
        j202_soc_core_ahb2apb_01_N142), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[78]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_14_ ( 
        .D(n25279), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_14_ ( 
        .D(n25279), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_14_ ( 
        .D(n25279), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_14_ ( 
        .D(n25279), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[14]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_14_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N54), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_14_ ( .D(
        j202_soc_core_ahb2apb_02_N142), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[46]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_rfuo_reg_sr__i__3_ ( .D(
        j202_soc_core_j22_cpu_rf_N3392), .DE(j202_soc_core_j22_cpu_rf_N3391), 
        .CLK(wb_clk_i), .Q(j202_soc_core_j22_cpu_rfuo_sr__i__3_) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_7_ ( .D(
        j202_soc_core_j22_cpu_rf_N305), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_23_ ( 
        .D(n25280), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_21_ ( 
        .D(j202_soc_core_qspi_wb_addr[23]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[10]), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cnt1[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[10]), .CLK(wb_clk_i), .RESET_B(
        n25731), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[10]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_10_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[10]), .CLK(wb_clk_i), .RESET_B(n25734), .Q(j202_soc_core_prdata[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_10_ ( .D(
        j202_soc_core_ahb2apb_00_N138), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[106])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[12]), .CLK(
        wb_clk_i), .RESET_B(n25732), .Q(j202_soc_core_cmt_core_00_cnt1[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[12]), .CLK(wb_clk_i), .RESET_B(
        n25734), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[12]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_12_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[12]), .CLK(wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_prdata[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_12_ ( .D(
        j202_soc_core_ahb2apb_00_N140), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[108])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[13]), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cnt1[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[13]), .CLK(wb_clk_i), .RESET_B(
        n25730), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[13]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_13_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[13]), .CLK(wb_clk_i), .RESET_B(n25733), .Q(j202_soc_core_prdata[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_13_ ( .D(
        j202_soc_core_ahb2apb_00_N141), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[109])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[14]), .CLK(
        wb_clk_i), .RESET_B(n25730), .Q(j202_soc_core_cmt_core_00_cnt1[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[14]), .CLK(wb_clk_i), .RESET_B(
        n25731), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[14]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_14_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[14]), .CLK(wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_prdata[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_14_ ( .D(
        j202_soc_core_ahb2apb_00_N142), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[110])
         );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[15]), .CLK(
        wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_cmt_core_00_cnt1[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cnt1[15]), .CLK(wb_clk_i), .RESET_B(
        n25731), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[15]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_15_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[15]), .CLK(wb_clk_i), .RESET_B(n25731), .Q(j202_soc_core_prdata[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_15_ ( .D(
        j202_soc_core_ahb2apb_00_N143), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[111])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_data_reg_11_ ( 
        .D(j202_soc_core_qspi_wb_wdat[11]), .DE(n25492), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_data[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[122]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[114]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[106]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_itgt[98]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[107]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[75]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[43]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ipr[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_irqc[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_rg_ie[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_11_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N14), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_11_ ( .D(
        j202_soc_core_ahb2apb_01_N139), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[75]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_odr_reg_reg_o_reg_11_ ( 
        .D(n25402), .DE(n10673), .CLK(wb_clk_i), .Q(la_data_out[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dr_reg_reg_o_reg_11_ ( 
        .D(n25402), .DE(n10672), .CLK(wb_clk_i), .Q(gpio_en_o[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_ier_reg_reg_o_reg_11_ ( 
        .D(n25402), .DE(n10671), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_dtr_reg_reg_o_reg_11_ ( 
        .D(n25402), .DE(n10670), .CLK(wb_clk_i), .Q(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_latch_status_reg_11_ ( 
        .D(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N51), .CLK(wb_clk_i), .Q(j202_soc_core_gpio_core_00_gpio_regs_00_isr[11]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N21), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[18])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_dout_reg_18_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N21), .CLK(wb_clk_i), .Q(j202_soc_core_intc_core_00_in_intreq[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_18_ ( .D(
        j202_soc_core_ahb2apb_01_N146), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[82]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_02_prdata_buf_reg_11_ ( .D(
        j202_soc_core_ahb2apb_02_N139), .DE(n25530), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[43]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_j22_cpu_rf_pc_reg_18_ ( .D(
        j202_soc_core_j22_cpu_rf_N316), .DE(n25490), .CLK(wb_clk_i), .Q(
        j202_soc_core_j22_cpu_pc[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2wbqspi_00_addr_temp_reg_21_ ( 
        .D(n25281), .DE(n11200), .CLK(wb_clk_i), .Q(
        j202_soc_core_qspi_wb_addr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spif_addr_reg_19_ ( 
        .D(j202_soc_core_qspi_wb_addr[21]), .DE(n25494), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_29_ ( .D(
        n10505), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[29]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_nxt_latch_status_0_), 
        .CLK(wb_clk_i), .RESET_B(n25731), .Q(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_0_) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_cmt_core_00_cmt_regs_00_rdata_reg_7_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[7]), .CLK(wb_clk_i), 
        .RESET_B(n25733), .Q(j202_soc_core_prdata[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_00_prdata_buf_reg_7_ ( .D(
        j202_soc_core_ahb2apb_00_N135), .DE(j202_soc_core_ahb2apb_00_N127), 
        .CLK(wb_clk_i), .Q(j202_soc_core_ahblite_interconnect_s_hrdata[103])
         );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N425), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N426), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N427), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N430), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_spi_len_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N428), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N424), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N391), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N392), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N393), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N394), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_4_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N395), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[4]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_10_ ( .D(
        n10524), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_11_ ( .D(
        n10523), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_22_ ( .D(
        n10512), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_23_ ( .D(
        n10511), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_28_ ( .D(
        n10506), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_5_ ( .D(
        n10529), .DE(n25535), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_5_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N396), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[5]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_6_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N397), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[6]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_7_ ( .D(
        n10527), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_7_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N398), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[7]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_8_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N399), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[8]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_9_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N400), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[9]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_10_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N401), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[10]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_11_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N402), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[11]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_12_ ( .D(
        n10522), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_12_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N403), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[12]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_13_ ( .D(
        n10521), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_13_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N404), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[13]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_14_ ( .D(
        n10520), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_14_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N405), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[14]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_15_ ( .D(
        n10519), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_15_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N406), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[15]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_16_ ( .D(
        n10518), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_16_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N407), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[16]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_17_ ( .D(
        n10517), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_17_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N408), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[17]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_18_ ( .D(
        n10516), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_18_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N409), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[18]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_19_ ( .D(
        n10515), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_19_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N410), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[19]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_20_ ( .D(
        n10514), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_20_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N411), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[20]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_21_ ( .D(
        n10513), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_21_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N412), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[21]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_22_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N413), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[22]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_23_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N414), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[23]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_24_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N415), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[24]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_25_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N416), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[25]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_26_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N417), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[26]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_27_ ( .D(
        n10507), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_27_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N418), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[27]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_28_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N419), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[28]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_29_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N420), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[29]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_dat_reg_1_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N317), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N315), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[1]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_spi_in_reg_30_ ( .D(
        n10504), .DE(j202_soc_core_wbqspiflash_00_N752), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_in[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_30_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N421), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[30]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_r_word_reg_31_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N422), .DE(n25527), .CLK(
        wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_lldriver_r_word[31]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_dat_reg_0_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N316), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N315), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[0]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_dat_reg_3_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N319), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N315), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[3]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_dat_reg_2_ ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N318), .DE(
        j202_soc_core_wbqspiflash_00_lldriver_N315), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[2]) );
  sky130_fd_sc_hd__edfxtp_1 j202_soc_core_ahb2apb_01_prdata_buf_reg_12_ ( .D(
        j202_soc_core_ahb2apb_01_N140), .DE(n25531), .CLK(wb_clk_i), .Q(
        j202_soc_core_ahblite_interconnect_s_hrdata[76]) );
  sky130_fd_sc_hd__fa_1 DP_OP_1501J1_126_8405_U6 ( .A(n25435), .B(n25482), 
        .CIN(DP_OP_1501J1_126_8405_n4), .COUT(DP_OP_1501J1_126_8405_n3), .SUM(
        U7_RSOP_1488_C3_DATA3_2) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_busy_reg ( 
        .D(j202_soc_core_wbqspiflash_00_lldriver_N321), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spi_busy) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_wbqspiflash_00_lldriver_o_valid_reg ( 
        .D(n25392), .CLK(wb_clk_i), .Q(j202_soc_core_wbqspiflash_00_spi_valid)
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_dout_reg_0_ ( 
        .D(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N3), .CLK(wb_clk_i), .Q(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_15_ ( .D(
        n25329), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[15])
         );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_7_ ( .D(
        n25326), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[7]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_memory0_ram_dout0_sel_reg_14_ ( .D(
        n25319), .CLK(wb_clk_i), .Q(j202_soc_core_memory0_ram_dout0_sel[14])
         );
  sky130_fd_sc_hd__dfstp_2 j202_soc_core_cmt_core_00_cmt_2ch_00_cmpcnt1_reg_0_ ( 
        .D(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[0]), .CLK(wb_clk_i), .SET_B(n25733), .Q(j202_soc_core_cmt_core_00_cnt1[0]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_02_pstrb_o_reg_2_ ( .GATE(
        j202_soc_core_ahb2apb_02_N123), .D(n10903), .RESET_B(
        j202_soc_core_pwrite[2]), .Q(j202_soc_core_pstrb[2]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_02_pstrb_o_reg_0_ ( .GATE(
        j202_soc_core_ahb2apb_02_N123), .D(n10901), .RESET_B(
        j202_soc_core_pwrite[2]), .Q(j202_soc_core_pstrb[0]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_01_pstrb_o_reg_1_ ( .GATE(
        j202_soc_core_ahb2apb_01_N123), .D(n10743), .RESET_B(
        j202_soc_core_pwrite[1]), .Q(j202_soc_core_pstrb[5]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_01_pstrb_o_reg_3_ ( .GATE(
        j202_soc_core_ahb2apb_01_N123), .D(n10745), .RESET_B(
        j202_soc_core_pwrite[1]), .Q(j202_soc_core_pstrb[7]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_02_pstrb_o_reg_1_ ( .GATE(
        j202_soc_core_ahb2apb_02_N123), .D(n10902), .RESET_B(
        j202_soc_core_pwrite[2]), .Q(j202_soc_core_pstrb[1]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_01_pstrb_o_reg_2_ ( .GATE(
        j202_soc_core_ahb2apb_01_N123), .D(n10744), .RESET_B(
        j202_soc_core_pwrite[1]), .Q(j202_soc_core_pstrb[6]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_02_pstrb_o_reg_3_ ( .GATE(
        j202_soc_core_ahb2apb_02_N123), .D(n10904), .RESET_B(
        j202_soc_core_pwrite[2]), .Q(j202_soc_core_pstrb[3]) );
  sky130_fd_sc_hd__dlrtp_1 j202_soc_core_ahb2apb_01_pstrb_o_reg_0_ ( .GATE(
        j202_soc_core_ahb2apb_01_N123), .D(n10742), .RESET_B(
        j202_soc_core_pwrite[1]), .Q(j202_soc_core_pstrb[4]) );
  sky130_fd_sc_hd__dfxtp_1 ready_reg ( .D(n25307), .CLK(wb_clk_i), .Q(
        wbs_ack_o) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_nega_o_reg ( 
        .D(n25397), .CLK(wb_clk_i), .RESET_B(n25733), .Q(io_out[17]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_posc_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posc), .CLK(wb_clk_i), .RESET_B(n25733), .Q(io_out[20]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_negb_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_negb), .CLK(wb_clk_i), .RESET_B(n25731), .Q(io_out[19]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_negc_o_reg ( 
        .D(n25398), .CLK(wb_clk_i), .RESET_B(n25733), .Q(io_out[21]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_posb_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posb), .CLK(wb_clk_i), .RESET_B(n25733), .Q(io_out[18]) );
  sky130_fd_sc_hd__dfrtp_1 j202_soc_core_bldc_core_00_bldc_pwm_00_pwm_posa_o_reg ( 
        .D(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posa), .CLK(wb_clk_i), .RESET_B(n25731), .Q(io_out[16]) );
  sky130_fd_sc_hd__dfxtp_1 j202_soc_core_wbqspiflash_00_spif_override_reg ( 
        .D(j202_soc_core_wbqspiflash_00_N742), .CLK(wb_clk_i), .Q(
        j202_soc_core_wbqspiflash_00_spif_override) );
  sky130_fd_sc_hd__dfxtp_4 j202_soc_core_rst_reg ( .D(j202_soc_core_rst1), 
        .CLK(wb_clk_i), .Q(j202_soc_core_rst) );
  sky130_fd_sc_hd__inv_4 U13287 ( .A(n10994), .Y(n10967) );
  sky130_fd_sc_hd__inv_4 U13288 ( .A(n25719), .Y(n10957) );
  sky130_fd_sc_hd__inv_4 U13289 ( .A(n10984), .Y(n10917) );
  sky130_fd_sc_hd__inv_4 U13290 ( .A(n10989), .Y(n10919) );
  sky130_fd_sc_hd__inv_4 U13291 ( .A(n10985), .Y(n10937) );
  sky130_fd_sc_hd__inv_4 U13292 ( .A(n10990), .Y(n10939) );
  sky130_fd_sc_hd__buf_2 U13312 ( .A(n10971), .X(n11178) );
  sky130_fd_sc_hd__clkbuf_1 U13315 ( .A(n20317), .X(n11179) );
  sky130_fd_sc_hd__clkbuf_1 U13316 ( .A(n21264), .X(n11172) );
  sky130_fd_sc_hd__clkbuf_1 U13317 ( .A(n21257), .X(n11171) );
  sky130_fd_sc_hd__clkbuf_1 U13318 ( .A(n20491), .X(n11180) );
  sky130_fd_sc_hd__clkbuf_1 U13319 ( .A(n21261), .X(n11173) );
  sky130_fd_sc_hd__clkbuf_1 U13320 ( .A(n21323), .X(n11174) );
  sky130_fd_sc_hd__clkbuf_1 U13321 ( .A(n21259), .X(n11176) );
  sky130_fd_sc_hd__clkbuf_1 U13322 ( .A(n21258), .X(n11175) );
  sky130_fd_sc_hd__inv_12 U13323 ( .A(n10970), .Y(n10971) );
  sky130_fd_sc_hd__nor2_1 U13324 ( .A(n21915), .B(n11036), .Y(n21262) );
  sky130_fd_sc_hd__nor2_1 U13325 ( .A(n22818), .B(n11036), .Y(n21260) );
  sky130_fd_sc_hd__nor2_1 U13326 ( .A(n21254), .B(n11036), .Y(n21255) );
  sky130_fd_sc_hd__inv_2 U13327 ( .A(n21243), .Y(n11177) );
  sky130_fd_sc_hd__nor2_1 U13328 ( .A(n21263), .B(n11036), .Y(n21264) );
  sky130_fd_sc_hd__nor2_1 U13329 ( .A(n21322), .B(n11036), .Y(n21323) );
  sky130_fd_sc_hd__nor2_1 U13330 ( .A(n22819), .B(n11036), .Y(n21261) );
  sky130_fd_sc_hd__nor2_1 U13331 ( .A(n22820), .B(n11036), .Y(n20491) );
  sky130_fd_sc_hd__nor2_1 U13332 ( .A(n22822), .B(n11036), .Y(n21259) );
  sky130_fd_sc_hd__nor2_1 U13333 ( .A(n22823), .B(n11036), .Y(n21258) );
  sky130_fd_sc_hd__nor2_1 U13334 ( .A(n22825), .B(n11036), .Y(n21257) );
  sky130_fd_sc_hd__nor2_1 U13335 ( .A(n21239), .B(n21242), .Y(n21240) );
  sky130_fd_sc_hd__nor2_2 U13339 ( .A(n11513), .B(n11531), .Y(n20301) );
  sky130_fd_sc_hd__inv_16 U13340 ( .A(n10917), .Y(n10918) );
  sky130_fd_sc_hd__inv_1 U13341 ( .A(n10981), .Y(n10984) );
  sky130_fd_sc_hd__inv_16 U13342 ( .A(n10919), .Y(n10920) );
  sky130_fd_sc_hd__inv_1 U13343 ( .A(n10986), .Y(n10989) );
  sky130_fd_sc_hd__inv_1 U13346 ( .A(n10996), .Y(n10999) );
  sky130_fd_sc_hd__inv_1 U13348 ( .A(n11001), .Y(n11004) );
  sky130_fd_sc_hd__inv_1 U13350 ( .A(n11006), .Y(n11009) );
  sky130_fd_sc_hd__inv_1 U13352 ( .A(n11011), .Y(n11014) );
  sky130_fd_sc_hd__inv_1 U13354 ( .A(n11016), .Y(n11019) );
  sky130_fd_sc_hd__inv_1 U13356 ( .A(n11021), .Y(n11024) );
  sky130_fd_sc_hd__inv_1 U13358 ( .A(n11026), .Y(n11029) );
  sky130_fd_sc_hd__inv_1 U13360 ( .A(n11031), .Y(n11034) );
  sky130_fd_sc_hd__inv_16 U13361 ( .A(n10937), .Y(n10938) );
  sky130_fd_sc_hd__inv_1 U13362 ( .A(n10981), .Y(n10985) );
  sky130_fd_sc_hd__inv_16 U13363 ( .A(n10939), .Y(n10940) );
  sky130_fd_sc_hd__inv_1 U13364 ( .A(n10986), .Y(n10990) );
  sky130_fd_sc_hd__inv_4 U13381 ( .A(n10957), .Y(n10958) );
  sky130_fd_sc_hd__inv_6 U13382 ( .A(n10957), .Y(n10959) );
  sky130_fd_sc_hd__inv_6 U13383 ( .A(n10957), .Y(n10960) );
  sky130_fd_sc_hd__inv_6 U13388 ( .A(n11178), .Y(n10964) );
  sky130_fd_sc_hd__inv_6 U13390 ( .A(n10964), .Y(n10966) );
  sky130_fd_sc_hd__inv_12 U13391 ( .A(n10967), .Y(n10968) );
  sky130_fd_sc_hd__inv_12 U13392 ( .A(n10967), .Y(n10969) );
  sky130_fd_sc_hd__inv_4 U13393 ( .A(n21240), .Y(n10970) );
  sky130_fd_sc_hd__inv_16 U13395 ( .A(n10972), .Y(n10974) );
  sky130_fd_sc_hd__inv_12 U13396 ( .A(n10972), .Y(n10976) );
  sky130_fd_sc_hd__buf_6 U13397 ( .A(n11178), .X(n10978) );
  sky130_fd_sc_hd__buf_12 U13398 ( .A(n11178), .X(n10979) );
  sky130_fd_sc_hd__clkinv_1 U13431 ( .A(j202_soc_core_j22_cpu_ml_bufa[20]), 
        .Y(n15783) );
  sky130_fd_sc_hd__clkinv_1 U13432 ( .A(n11169), .Y(n11170) );
  sky130_fd_sc_hd__inv_2 U13433 ( .A(j202_soc_core_memory0_ram_dout0_sel[13]), 
        .Y(n11303) );
  sky130_fd_sc_hd__clkinv_1 U13434 ( .A(n21147), .Y(n21108) );
  sky130_fd_sc_hd__clkinv_1 U13435 ( .A(j202_soc_core_memory0_ram_dout0_sel[9]), .Y(n11298) );
  sky130_fd_sc_hd__clkinv_1 U13438 ( .A(j202_soc_core_j22_cpu_ml_bufb[0]), .Y(
        n15962) );
  sky130_fd_sc_hd__clkinv_1 U13440 ( .A(n20257), .Y(n14060) );
  sky130_fd_sc_hd__clkinv_1 U13443 ( .A(n20986), .Y(n21574) );
  sky130_fd_sc_hd__clkinv_1 U13444 ( .A(n20260), .Y(n14047) );
  sky130_fd_sc_hd__clkinv_1 U13445 ( .A(n21624), .Y(n13094) );
  sky130_fd_sc_hd__clkinv_1 U13446 ( .A(io_in[15]), .Y(n14801) );
  sky130_fd_sc_hd__clkinv_1 U13447 ( .A(n22141), .Y(n20805) );
  sky130_fd_sc_hd__clkinv_1 U13448 ( .A(n21170), .Y(n21091) );
  sky130_fd_sc_hd__clkinv_1 U13451 ( .A(n19959), .Y(n20036) );
  sky130_fd_sc_hd__inv_1 U13452 ( .A(n22185), .Y(n21627) );
  sky130_fd_sc_hd__inv_1 U13453 ( .A(n22708), .Y(n22611) );
  sky130_fd_sc_hd__inv_1 U13454 ( .A(n20277), .Y(n20278) );
  sky130_fd_sc_hd__clkinv_1 U13455 ( .A(n22735), .Y(n22742) );
  sky130_fd_sc_hd__inv_1 U13456 ( .A(n22705), .Y(n22646) );
  sky130_fd_sc_hd__inv_1 U13457 ( .A(n22176), .Y(n22037) );
  sky130_fd_sc_hd__clkinv_1 U13458 ( .A(n21635), .Y(n22407) );
  sky130_fd_sc_hd__clkinv_1 U13459 ( .A(n24873), .Y(n21418) );
  sky130_fd_sc_hd__inv_2 U13461 ( .A(j202_soc_core_j22_cpu_ma_M_area[0]), .Y(
        n11288) );
  sky130_fd_sc_hd__clkinv_1 U13462 ( .A(n25377), .Y(n22333) );
  sky130_fd_sc_hd__clkinv_1 U13464 ( .A(n22662), .Y(n22757) );
  sky130_fd_sc_hd__clkinv_1 U13465 ( .A(n23300), .Y(n22368) );
  sky130_fd_sc_hd__nor2_1 U13466 ( .A(n22509), .B(n22687), .Y(n21137) );
  sky130_fd_sc_hd__clkinv_1 U13469 ( .A(n20983), .Y(n22734) );
  sky130_fd_sc_hd__clkinv_1 U13470 ( .A(n21480), .Y(n21403) );
  sky130_fd_sc_hd__inv_1 U13473 ( .A(n22283), .Y(n21483) );
  sky130_fd_sc_hd__clkinv_1 U13475 ( .A(n23343), .Y(n23297) );
  sky130_fd_sc_hd__clkinv_1 U13476 ( .A(n24444), .Y(n20114) );
  sky130_fd_sc_hd__clkinv_1 U13479 ( .A(n21019), .Y(n22487) );
  sky130_fd_sc_hd__nand2_1 U13480 ( .A(n21009), .B(n20880), .Y(n23321) );
  sky130_fd_sc_hd__clkinv_1 U13481 ( .A(n23239), .Y(n24894) );
  sky130_fd_sc_hd__inv_2 U13482 ( .A(j202_soc_core_j22_cpu_memop_MEM__2_), .Y(
        n23243) );
  sky130_fd_sc_hd__or2b_2 U13483 ( .A(n25339), .B_N(n25734), .X(
        j202_soc_core_ahb2apb_02_N22) );
  sky130_fd_sc_hd__inv_2 U13492 ( .A(n10978), .Y(n11167) );
  sky130_fd_sc_hd__nor2_1 U13493 ( .A(n18510), .B(n21904), .Y(n21249) );
  sky130_fd_sc_hd__clkinv_1 U13494 ( .A(n22221), .Y(n22224) );
  sky130_fd_sc_hd__clkinv_1 U13495 ( .A(n22785), .Y(n21393) );
  sky130_fd_sc_hd__clkinv_1 U13496 ( .A(n21365), .Y(n21385) );
  sky130_fd_sc_hd__or2_0 U13497 ( .A(n20994), .B(n21598), .X(n21496) );
  sky130_fd_sc_hd__clkinv_1 U13498 ( .A(n25375), .Y(n21263) );
  sky130_fd_sc_hd__clkinv_1 U13499 ( .A(n25373), .Y(n20316) );
  sky130_fd_sc_hd__or2_0 U13500 ( .A(n20330), .B(n21418), .X(n20340) );
  sky130_fd_sc_hd__or2_0 U13501 ( .A(n20639), .B(n20355), .X(n22270) );
  sky130_fd_sc_hd__or2_0 U13502 ( .A(n21046), .B(n20355), .X(n21890) );
  sky130_fd_sc_hd__or2_0 U13503 ( .A(n20856), .B(n20355), .X(n21971) );
  sky130_fd_sc_hd__or2_0 U13504 ( .A(n20356), .B(n20355), .X(n22081) );
  sky130_fd_sc_hd__or2_0 U13505 ( .A(n20382), .B(n20355), .X(n21981) );
  sky130_fd_sc_hd__clkinv_1 U13506 ( .A(n25381), .Y(n22328) );
  sky130_fd_sc_hd__clkinv_1 U13507 ( .A(n25387), .Y(n22309) );
  sky130_fd_sc_hd__or2_0 U13508 ( .A(n16507), .B(n16508), .X(n18997) );
  sky130_fd_sc_hd__or2_0 U13509 ( .A(n16026), .B(n16027), .X(n19223) );
  sky130_fd_sc_hd__or2_0 U13510 ( .A(n16028), .B(n16029), .X(n19226) );
  sky130_fd_sc_hd__or2_0 U13511 ( .A(n16013), .B(n16014), .X(n18866) );
  sky130_fd_sc_hd__or2_0 U13512 ( .A(n16015), .B(n16016), .X(n17045) );
  sky130_fd_sc_hd__or2_0 U13513 ( .A(n16517), .B(n16518), .X(n18853) );
  sky130_fd_sc_hd__or2_0 U13514 ( .A(n16519), .B(n16520), .X(n18856) );
  sky130_fd_sc_hd__or2_0 U13515 ( .A(n12717), .B(n12718), .X(n11181) );
  sky130_fd_sc_hd__or2_0 U13516 ( .A(n15978), .B(n15979), .X(n16633) );
  sky130_fd_sc_hd__or2_0 U13517 ( .A(n12683), .B(n12684), .X(n11186) );
  sky130_fd_sc_hd__or2_0 U13518 ( .A(n14037), .B(n14038), .X(n11185) );
  sky130_fd_sc_hd__or2_0 U13519 ( .A(n13997), .B(n13998), .X(n11189) );
  sky130_fd_sc_hd__or2_0 U13520 ( .A(n12843), .B(n12844), .X(n11190) );
  sky130_fd_sc_hd__or2_0 U13521 ( .A(n16572), .B(n16573), .X(n19094) );
  sky130_fd_sc_hd__or2_0 U13522 ( .A(n12785), .B(n12786), .X(n11188) );
  sky130_fd_sc_hd__or2_0 U13523 ( .A(n12751), .B(n12752), .X(n11192) );
  sky130_fd_sc_hd__or2_0 U13524 ( .A(j202_soc_core_rst), .B(n24491), .X(n24744) );
  sky130_fd_sc_hd__or2_0 U13525 ( .A(n16586), .B(n16587), .X(n19350) );
  sky130_fd_sc_hd__or2_0 U13526 ( .A(n15973), .B(n15974), .X(n19141) );
  sky130_fd_sc_hd__or2_0 U13527 ( .A(n14090), .B(n14091), .X(n11194) );
  sky130_fd_sc_hd__or2_0 U13528 ( .A(n19596), .B(n19354), .X(n19922) );
  sky130_fd_sc_hd__or2_0 U13529 ( .A(n15952), .B(n15953), .X(n16840) );
  sky130_fd_sc_hd__or2_0 U13530 ( .A(n12649), .B(n12650), .X(n11195) );
  sky130_fd_sc_hd__or2_0 U13531 ( .A(n20095), .B(n24495), .X(n24493) );
  sky130_fd_sc_hd__or2_0 U13532 ( .A(n16580), .B(n21728), .X(n15933) );
  sky130_fd_sc_hd__or2_0 U13533 ( .A(n19329), .B(n19596), .X(n19552) );
  sky130_fd_sc_hd__or2_0 U13534 ( .A(n19368), .B(n19596), .X(n19390) );
  sky130_fd_sc_hd__or2_0 U13535 ( .A(n19364), .B(n19596), .X(n20027) );
  sky130_fd_sc_hd__or2_0 U13536 ( .A(n19556), .B(n19596), .X(n19937) );
  sky130_fd_sc_hd__or2_0 U13537 ( .A(n20496), .B(n20495), .X(n25189) );
  sky130_fd_sc_hd__or2_0 U13538 ( .A(n13611), .B(n18100), .X(n18130) );
  sky130_fd_sc_hd__or2_0 U13539 ( .A(n14694), .B(n14693), .X(n14712) );
  sky130_fd_sc_hd__or2_0 U13540 ( .A(n18767), .B(n18512), .X(n18526) );
  sky130_fd_sc_hd__or2_0 U13541 ( .A(n13256), .B(n17969), .X(n13585) );
  sky130_fd_sc_hd__or2_0 U13542 ( .A(n18775), .B(n18512), .X(n16931) );
  sky130_fd_sc_hd__or2_0 U13543 ( .A(n24898), .B(j202_soc_core_rst), .X(
        j202_soc_core_wbqspiflash_00_N720) );
  sky130_fd_sc_hd__or2_0 U13544 ( .A(j202_soc_core_j22_cpu_ml_bufa[2]), .B(
        n15944), .X(n15946) );
  sky130_fd_sc_hd__or2_0 U13545 ( .A(n20839), .B(n20931), .X(n21141) );
  sky130_fd_sc_hd__or2_0 U13546 ( .A(n14598), .B(n14597), .X(n14599) );
  sky130_fd_sc_hd__nor3_2 U13547 ( .A(j202_soc_core_memory0_ram_dout0_sel[9]), 
        .B(n11291), .C(n11297), .Y(n18062) );
  sky130_fd_sc_hd__clkinv_1 U13548 ( .A(n12111), .Y(n11512) );
  sky130_fd_sc_hd__or2_0 U13549 ( .A(n13214), .B(n13213), .X(n18032) );
  sky130_fd_sc_hd__and2_0 U13550 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]), .B(n25734), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N10) );
  sky130_fd_sc_hd__and2_0 U13551 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[19]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N22) );
  sky130_fd_sc_hd__and2_0 U13552 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[18]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N21) );
  sky130_fd_sc_hd__and2_0 U13553 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N17) );
  sky130_fd_sc_hd__and2_0 U13554 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[10]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N13) );
  sky130_fd_sc_hd__and2_0 U13555 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N18) );
  sky130_fd_sc_hd__and2_0 U13556 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]), .B(n25734), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N4) );
  sky130_fd_sc_hd__and2_0 U13557 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]), .B(n25734), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N8) );
  sky130_fd_sc_hd__or2_0 U13558 ( .A(j202_soc_core_j22_cpu_ml_bufb[3]), .B(
        j202_soc_core_j22_cpu_ml_bufb[2]), .X(n11196) );
  sky130_fd_sc_hd__or2_0 U13559 ( .A(j202_soc_core_j22_cpu_ml_bufb[1]), .B(
        j202_soc_core_j22_cpu_ml_bufb[0]), .X(n15229) );
  sky130_fd_sc_hd__or2_0 U13560 ( .A(j202_soc_core_j22_cpu_ml_bufb[1]), .B(
        j202_soc_core_j22_cpu_ml_bufb[2]), .X(n11198) );
  sky130_fd_sc_hd__and2_0 U13561 ( .A(n25340), .B(n25334), .X(n25452) );
  sky130_fd_sc_hd__and2_0 U13562 ( .A(n25340), .B(n25333), .X(n25451) );
  sky130_fd_sc_hd__and2_0 U13563 ( .A(n25340), .B(n25391), .X(n25450) );
  sky130_fd_sc_hd__and2_1 U13565 ( .A(n25340), .B(n25375), .X(n25458) );
  sky130_fd_sc_hd__nand2b_2 U13567 ( .A_N(n25340), .B(n25730), .Y(
        j202_soc_core_ahb2apb_01_N22) );
  sky130_fd_sc_hd__and2_0 U13568 ( .A(n25340), .B(n25335), .X(n25453) );
  sky130_fd_sc_hd__and2_1 U13569 ( .A(n25340), .B(n25373), .X(n25459) );
  sky130_fd_sc_hd__and2_1 U13571 ( .A(n25340), .B(n25338), .X(n25456) );
  sky130_fd_sc_hd__and2_1 U13572 ( .A(n25340), .B(n25337), .X(n25455) );
  sky130_fd_sc_hd__and2_1 U13573 ( .A(n25340), .B(n25488), .X(n25460) );
  sky130_fd_sc_hd__and2_1 U13574 ( .A(n25340), .B(n21906), .X(n25429) );
  sky130_fd_sc_hd__and2_0 U13575 ( .A(n25340), .B(n25374), .X(n25449) );
  sky130_fd_sc_hd__and2_1 U13576 ( .A(n25340), .B(n25378), .X(n25457) );
  sky130_fd_sc_hd__and2_1 U13577 ( .A(n25340), .B(n22100), .X(n25461) );
  sky130_fd_sc_hd__clkinv_1 U13578 ( .A(n25325), .Y(n10543) );
  sky130_fd_sc_hd__clkinv_1 U13579 ( .A(n25326), .Y(n10547) );
  sky130_fd_sc_hd__clkinv_1 U13580 ( .A(n25319), .Y(n10554) );
  sky130_fd_sc_hd__clkinv_1 U13581 ( .A(n25328), .Y(n10545) );
  sky130_fd_sc_hd__clkinv_1 U13582 ( .A(n25330), .Y(n10549) );
  sky130_fd_sc_hd__clkinv_1 U13583 ( .A(n25323), .Y(n10552) );
  sky130_fd_sc_hd__clkinv_1 U13584 ( .A(n25317), .Y(n10550) );
  sky130_fd_sc_hd__clkinv_1 U13585 ( .A(n25322), .Y(n10546) );
  sky130_fd_sc_hd__clkinv_1 U13586 ( .A(n25329), .Y(n10555) );
  sky130_fd_sc_hd__clkinv_1 U13587 ( .A(n22824), .Y(n25541) );
  sky130_fd_sc_hd__clkinv_1 U13588 ( .A(n25321), .Y(n10540) );
  sky130_fd_sc_hd__clkinv_1 U13589 ( .A(n25324), .Y(n10541) );
  sky130_fd_sc_hd__clkinv_1 U13590 ( .A(n25331), .Y(n10551) );
  sky130_fd_sc_hd__clkinv_1 U13591 ( .A(n25318), .Y(n10548) );
  sky130_fd_sc_hd__clkinv_1 U13592 ( .A(n25320), .Y(n10542) );
  sky130_fd_sc_hd__clkinv_1 U13593 ( .A(n25332), .Y(n10553) );
  sky130_fd_sc_hd__clkinv_1 U13594 ( .A(n25327), .Y(n10544) );
  sky130_fd_sc_hd__clkinv_1 U13595 ( .A(n25362), .Y(n21307) );
  sky130_fd_sc_hd__clkinv_1 U13597 ( .A(n25361), .Y(n21305) );
  sky130_fd_sc_hd__and2_0 U13599 ( .A(n21980), .B(n21996), .X(n25477) );
  sky130_fd_sc_hd__clkinv_1 U13600 ( .A(n25359), .Y(n21301) );
  sky130_fd_sc_hd__nor2_1 U13613 ( .A(n20316), .B(n21253), .Y(n20317) );
  sky130_fd_sc_hd__clkinv_1 U13617 ( .A(n22403), .Y(n22829) );
  sky130_fd_sc_hd__clkinv_1 U13618 ( .A(n25358), .Y(n21299) );
  sky130_fd_sc_hd__clkinv_1 U13619 ( .A(n25345), .Y(n21273) );
  sky130_fd_sc_hd__and2_0 U13626 ( .A(n22079), .B(n21996), .X(n25432) );
  sky130_fd_sc_hd__clkinv_1 U13629 ( .A(n25357), .Y(n21297) );
  sky130_fd_sc_hd__clkinv_1 U13636 ( .A(n25343), .Y(n21269) );
  sky130_fd_sc_hd__clkinv_1 U13639 ( .A(n14956), .Y(n14958) );
  sky130_fd_sc_hd__clkinv_1 U13640 ( .A(n25356), .Y(n21295) );
  sky130_fd_sc_hd__clkinv_1 U13641 ( .A(n25353), .Y(n21289) );
  sky130_fd_sc_hd__clkinv_1 U13642 ( .A(n22194), .Y(n22197) );
  sky130_fd_sc_hd__clkinv_1 U13643 ( .A(n25366), .Y(n21315) );
  sky130_fd_sc_hd__clkinv_1 U13644 ( .A(n25342), .Y(n21267) );
  sky130_fd_sc_hd__clkinv_1 U13645 ( .A(n25355), .Y(n21293) );
  sky130_fd_sc_hd__clkinv_1 U13646 ( .A(n25301), .Y(n20312) );
  sky130_fd_sc_hd__clkinv_1 U13647 ( .A(n25344), .Y(n21271) );
  sky130_fd_sc_hd__clkinv_1 U13648 ( .A(n21884), .Y(n21886) );
  sky130_fd_sc_hd__clkinv_1 U13649 ( .A(n25368), .Y(n21319) );
  sky130_fd_sc_hd__clkinv_1 U13650 ( .A(n25365), .Y(n21313) );
  sky130_fd_sc_hd__clkinv_1 U13651 ( .A(n25300), .Y(n20310) );
  sky130_fd_sc_hd__clkinv_1 U13652 ( .A(n25367), .Y(n21317) );
  sky130_fd_sc_hd__clkinv_1 U13653 ( .A(n25351), .Y(n21285) );
  sky130_fd_sc_hd__clkinv_1 U13654 ( .A(n25352), .Y(n21287) );
  sky130_fd_sc_hd__clkinv_1 U13655 ( .A(n21742), .Y(n21744) );
  sky130_fd_sc_hd__clkinv_1 U13656 ( .A(n25354), .Y(n21291) );
  sky130_fd_sc_hd__clkinv_1 U13657 ( .A(n22086), .Y(n22088) );
  sky130_fd_sc_hd__clkinv_1 U13658 ( .A(n22506), .Y(n22508) );
  sky130_fd_sc_hd__clkinv_1 U13659 ( .A(n25363), .Y(n21309) );
  sky130_fd_sc_hd__clkinv_1 U13660 ( .A(n25349), .Y(n21281) );
  sky130_fd_sc_hd__clkinv_1 U13661 ( .A(n25348), .Y(n21279) );
  sky130_fd_sc_hd__clkinv_1 U13662 ( .A(n21793), .Y(n21794) );
  sky130_fd_sc_hd__clkinv_1 U13663 ( .A(n25360), .Y(n21303) );
  sky130_fd_sc_hd__clkinv_1 U13664 ( .A(n21813), .Y(n21814) );
  sky130_fd_sc_hd__clkinv_1 U13665 ( .A(n25306), .Y(n20489) );
  sky130_fd_sc_hd__clkinv_1 U13666 ( .A(n25347), .Y(n21277) );
  sky130_fd_sc_hd__clkinv_1 U13667 ( .A(n25346), .Y(n21275) );
  sky130_fd_sc_hd__clkinv_1 U13668 ( .A(n18472), .Y(n21075) );
  sky130_fd_sc_hd__clkinv_1 U13669 ( .A(n25341), .Y(n21265) );
  sky130_fd_sc_hd__clkinv_1 U13670 ( .A(n25302), .Y(n20314) );
  sky130_fd_sc_hd__clkinv_1 U13671 ( .A(n21892), .Y(n21896) );
  sky130_fd_sc_hd__clkinv_1 U13672 ( .A(n25364), .Y(n21311) );
  sky130_fd_sc_hd__clkinv_1 U13673 ( .A(n22208), .Y(n22209) );
  sky130_fd_sc_hd__clkinv_1 U13674 ( .A(n21692), .Y(n21719) );
  sky130_fd_sc_hd__clkinv_1 U13675 ( .A(n21918), .Y(n21919) );
  sky130_fd_sc_hd__clkinv_1 U13676 ( .A(n25350), .Y(n21283) );
  sky130_fd_sc_hd__clkinv_1 U13678 ( .A(n14961), .Y(n14964) );
  sky130_fd_sc_hd__and2_1 U13679 ( .A(n22017), .B(n21996), .X(n25465) );
  sky130_fd_sc_hd__clkinv_1 U13680 ( .A(n22027), .Y(n22028) );
  sky130_fd_sc_hd__a21o_1 U13681 ( .A1(n14396), .A2(n11194), .B1(n14092), .X(
        n14093) );
  sky130_fd_sc_hd__clkinv_1 U13682 ( .A(n21694), .Y(n21714) );
  sky130_fd_sc_hd__clkinv_1 U13683 ( .A(n18506), .Y(n14962) );
  sky130_fd_sc_hd__clkinv_1 U13684 ( .A(n21952), .Y(n21956) );
  sky130_fd_sc_hd__clkinv_1 U13685 ( .A(n19499), .Y(n19502) );
  sky130_fd_sc_hd__clkinv_1 U13686 ( .A(n22210), .Y(n22211) );
  sky130_fd_sc_hd__clkinv_1 U13687 ( .A(n19291), .Y(n16785) );
  sky130_fd_sc_hd__clkinv_1 U13688 ( .A(n25257), .Y(n14948) );
  sky130_fd_sc_hd__clkinv_1 U13689 ( .A(n22252), .Y(n22256) );
  sky130_fd_sc_hd__clkinv_1 U13690 ( .A(n21945), .Y(n21946) );
  sky130_fd_sc_hd__clkinv_1 U13691 ( .A(n21541), .Y(n21521) );
  sky130_fd_sc_hd__clkinv_1 U13692 ( .A(n25305), .Y(n20350) );
  sky130_fd_sc_hd__clkinv_1 U13693 ( .A(n22220), .Y(n22222) );
  sky130_fd_sc_hd__clkinv_1 U13694 ( .A(n22212), .Y(n22214) );
  sky130_fd_sc_hd__clkinv_1 U13695 ( .A(n21765), .Y(n21769) );
  sky130_fd_sc_hd__clkinv_1 U13696 ( .A(n21940), .Y(n21941) );
  sky130_fd_sc_hd__clkinv_1 U13697 ( .A(n21773), .Y(n21774) );
  sky130_fd_sc_hd__clkinv_1 U13698 ( .A(n18998), .Y(n19129) );
  sky130_fd_sc_hd__clkinv_1 U13699 ( .A(n21704), .Y(n21705) );
  sky130_fd_sc_hd__clkinv_1 U13700 ( .A(n21703), .Y(n21706) );
  sky130_fd_sc_hd__clkinv_1 U13701 ( .A(n21593), .Y(n21595) );
  sky130_fd_sc_hd__clkinv_1 U13702 ( .A(n21839), .Y(n21844) );
  sky130_fd_sc_hd__clkinv_1 U13704 ( .A(n24861), .Y(n21600) );
  sky130_fd_sc_hd__clkinv_1 U13705 ( .A(n21739), .Y(n21740) );
  sky130_fd_sc_hd__clkinv_1 U13706 ( .A(n21823), .Y(n21827) );
  sky130_fd_sc_hd__clkinv_1 U13707 ( .A(n21504), .Y(n21512) );
  sky130_fd_sc_hd__clkinv_1 U13709 ( .A(n17079), .Y(n18876) );
  sky130_fd_sc_hd__clkinv_1 U13710 ( .A(n21877), .Y(n21882) );
  sky130_fd_sc_hd__clkinv_1 U13711 ( .A(n24843), .Y(n23225) );
  sky130_fd_sc_hd__clkinv_1 U13712 ( .A(n18859), .Y(n18975) );
  sky130_fd_sc_hd__clkinv_1 U13713 ( .A(n21473), .Y(n21482) );
  sky130_fd_sc_hd__clkinv_1 U13714 ( .A(n21974), .Y(n21978) );
  sky130_fd_sc_hd__clkinv_1 U13715 ( .A(n19361), .Y(n19216) );
  sky130_fd_sc_hd__clkinv_1 U13716 ( .A(n21406), .Y(n22797) );
  sky130_fd_sc_hd__clkinv_1 U13717 ( .A(n22327), .Y(n21990) );
  sky130_fd_sc_hd__clkinv_1 U13718 ( .A(n21643), .Y(n21645) );
  sky130_fd_sc_hd__clkinv_1 U13719 ( .A(n22020), .Y(n22024) );
  sky130_fd_sc_hd__clkinv_1 U13720 ( .A(n21756), .Y(n21760) );
  sky130_fd_sc_hd__clkinv_1 U13721 ( .A(n16625), .Y(n19299) );
  sky130_fd_sc_hd__clkinv_1 U13722 ( .A(n21913), .Y(n21247) );
  sky130_fd_sc_hd__clkinv_1 U13723 ( .A(n22107), .Y(n22332) );
  sky130_fd_sc_hd__clkinv_1 U13724 ( .A(n25254), .Y(n18502) );
  sky130_fd_sc_hd__clkinv_1 U13725 ( .A(n24849), .Y(n21327) );
  sky130_fd_sc_hd__clkinv_1 U13726 ( .A(n20743), .Y(n20744) );
  sky130_fd_sc_hd__clkinv_1 U13727 ( .A(n20332), .Y(n20988) );
  sky130_fd_sc_hd__clkinv_1 U13728 ( .A(n21786), .Y(n21791) );
  sky130_fd_sc_hd__clkinv_1 U13729 ( .A(n21564), .Y(n22387) );
  sky130_fd_sc_hd__clkinv_1 U13730 ( .A(n24871), .Y(n20992) );
  sky130_fd_sc_hd__clkinv_1 U13731 ( .A(n17082), .Y(n19007) );
  sky130_fd_sc_hd__clkinv_1 U13732 ( .A(n22115), .Y(n22120) );
  sky130_fd_sc_hd__clkinv_1 U13733 ( .A(n21510), .Y(n21632) );
  sky130_fd_sc_hd__clkinv_1 U13734 ( .A(n19801), .Y(n19835) );
  sky130_fd_sc_hd__clkinv_1 U13735 ( .A(n22329), .Y(n22108) );
  sky130_fd_sc_hd__clkinv_1 U13736 ( .A(n22307), .Y(n22280) );
  sky130_fd_sc_hd__clkinv_1 U13737 ( .A(n21412), .Y(n21456) );
  sky130_fd_sc_hd__clkinv_1 U13738 ( .A(n19834), .Y(n19796) );
  sky130_fd_sc_hd__clkinv_1 U13739 ( .A(n22282), .Y(n21430) );
  sky130_fd_sc_hd__clkinv_1 U13740 ( .A(n21536), .Y(n21461) );
  sky130_fd_sc_hd__clkinv_1 U13741 ( .A(n16832), .Y(n19859) );
  sky130_fd_sc_hd__clkinv_1 U13742 ( .A(n25273), .Y(n21245) );
  sky130_fd_sc_hd__clkinv_1 U13743 ( .A(n21457), .Y(n20995) );
  sky130_fd_sc_hd__clkinv_1 U13744 ( .A(n24853), .Y(n21631) );
  sky130_fd_sc_hd__clkinv_1 U13745 ( .A(n16605), .Y(n19224) );
  sky130_fd_sc_hd__clkinv_1 U13746 ( .A(n21244), .Y(n19836) );
  sky130_fd_sc_hd__clkinv_1 U13747 ( .A(n21435), .Y(n20742) );
  sky130_fd_sc_hd__clkinv_1 U13748 ( .A(n22373), .Y(n22380) );
  sky130_fd_sc_hd__clkinv_1 U13749 ( .A(n21907), .Y(n21238) );
  sky130_fd_sc_hd__clkinv_1 U13750 ( .A(n22419), .Y(n20768) );
  sky130_fd_sc_hd__a21oi_1 U13751 ( .A1(n18494), .A2(n11181), .B1(n12719), .Y(
        n13545) );
  sky130_fd_sc_hd__clkinv_1 U13752 ( .A(n20975), .Y(n21548) );
  sky130_fd_sc_hd__clkinv_1 U13753 ( .A(n20331), .Y(n21569) );
  sky130_fd_sc_hd__clkinv_1 U13754 ( .A(n21474), .Y(n21634) );
  sky130_fd_sc_hd__clkinv_1 U13755 ( .A(n21506), .Y(n20772) );
  sky130_fd_sc_hd__clkinv_1 U13756 ( .A(n14959), .Y(n14945) );
  sky130_fd_sc_hd__clkinv_1 U13757 ( .A(n25378), .Y(n21915) );
  sky130_fd_sc_hd__clkinv_1 U13758 ( .A(n23321), .Y(n21820) );
  sky130_fd_sc_hd__clkinv_1 U13759 ( .A(n22733), .Y(n21572) );
  sky130_fd_sc_hd__clkinv_1 U13760 ( .A(n20759), .Y(n21331) );
  sky130_fd_sc_hd__clkinv_1 U13761 ( .A(n22273), .Y(n22279) );
  sky130_fd_sc_hd__clkinv_1 U13762 ( .A(n20396), .Y(n20383) );
  sky130_fd_sc_hd__clkinv_1 U13763 ( .A(n21422), .Y(n21409) );
  sky130_fd_sc_hd__clkinv_1 U13764 ( .A(n21336), .Y(n21534) );
  sky130_fd_sc_hd__clkinv_1 U13765 ( .A(n23547), .Y(n23549) );
  sky130_fd_sc_hd__clkinv_1 U13766 ( .A(n25272), .Y(n19798) );
  sky130_fd_sc_hd__clkinv_1 U13767 ( .A(n25374), .Y(n19832) );
  sky130_fd_sc_hd__clkinv_1 U13768 ( .A(n18989), .Y(n19111) );
  sky130_fd_sc_hd__clkinv_1 U13769 ( .A(n22816), .Y(n25391) );
  sky130_fd_sc_hd__clkinv_1 U13770 ( .A(n22390), .Y(n21563) );
  sky130_fd_sc_hd__clkinv_1 U13771 ( .A(n17042), .Y(n18867) );
  sky130_fd_sc_hd__and2_0 U13773 ( .A(n25379), .B(n21908), .X(n21239) );
  sky130_fd_sc_hd__clkinv_1 U13774 ( .A(n21332), .Y(n21486) );
  sky130_fd_sc_hd__clkinv_1 U13775 ( .A(n23241), .Y(
        j202_soc_core_j22_cpu_ifetch) );
  sky130_fd_sc_hd__clkinv_1 U13776 ( .A(n20993), .Y(n20342) );
  sky130_fd_sc_hd__clkinv_1 U13777 ( .A(n21171), .Y(n21140) );
  sky130_fd_sc_hd__clkinv_1 U13778 ( .A(n20760), .Y(n21547) );
  sky130_fd_sc_hd__clkinv_1 U13779 ( .A(n20673), .Y(n20679) );
  sky130_fd_sc_hd__clkinv_1 U13780 ( .A(n21122), .Y(n21106) );
  sky130_fd_sc_hd__clkinv_1 U13781 ( .A(n21861), .Y(n21866) );
  sky130_fd_sc_hd__clkinv_1 U13782 ( .A(n22389), .Y(n21424) );
  sky130_fd_sc_hd__clkinv_1 U13783 ( .A(n16805), .Y(n19957) );
  sky130_fd_sc_hd__clkinv_1 U13784 ( .A(n21801), .Y(n22306) );
  sky130_fd_sc_hd__clkinv_1 U13785 ( .A(n21413), .Y(n21492) );
  sky130_fd_sc_hd__clkinv_1 U13786 ( .A(n19438), .Y(n19439) );
  sky130_fd_sc_hd__clkinv_1 U13787 ( .A(n19437), .Y(n19440) );
  sky130_fd_sc_hd__clkinv_1 U13788 ( .A(n21381), .Y(n21353) );
  sky130_fd_sc_hd__clkinv_1 U13789 ( .A(n21533), .Y(n20343) );
  sky130_fd_sc_hd__clkinv_1 U13790 ( .A(n20752), .Y(n21487) );
  sky130_fd_sc_hd__clkinv_1 U13791 ( .A(n20737), .Y(n21455) );
  sky130_fd_sc_hd__clkinv_1 U13792 ( .A(n20985), .Y(n21575) );
  sky130_fd_sc_hd__clkinv_1 U13793 ( .A(n21734), .Y(n20978) );
  sky130_fd_sc_hd__clkinv_1 U13794 ( .A(n22516), .Y(n20902) );
  sky130_fd_sc_hd__a21oi_1 U13795 ( .A1(n18829), .A2(n11195), .B1(n12651), .Y(
        n18809) );
  sky130_fd_sc_hd__clkinv_1 U13796 ( .A(n21361), .Y(n21377) );
  sky130_fd_sc_hd__clkinv_1 U13797 ( .A(n21366), .Y(n21367) );
  sky130_fd_sc_hd__clkinv_1 U13798 ( .A(n20335), .Y(n19322) );
  sky130_fd_sc_hd__clkinv_1 U13799 ( .A(n21573), .Y(n20741) );
  sky130_fd_sc_hd__clkinv_1 U13800 ( .A(n19736), .Y(n19520) );
  sky130_fd_sc_hd__clkinv_1 U13801 ( .A(n21735), .Y(n20341) );
  sky130_fd_sc_hd__clkinv_1 U13802 ( .A(n16615), .Y(n16616) );
  sky130_fd_sc_hd__clkinv_1 U13803 ( .A(n16614), .Y(n16617) );
  sky130_fd_sc_hd__clkinv_1 U13804 ( .A(n21530), .Y(n21004) );
  sky130_fd_sc_hd__clkinv_1 U13805 ( .A(n16787), .Y(n16790) );
  sky130_fd_sc_hd__clkinv_1 U13806 ( .A(n18973), .Y(n18974) );
  sky130_fd_sc_hd__clkinv_1 U13807 ( .A(n24857), .Y(n22337) );
  sky130_fd_sc_hd__clkinv_1 U13808 ( .A(n21623), .Y(n21622) );
  sky130_fd_sc_hd__clkinv_1 U13809 ( .A(n18972), .Y(n18976) );
  sky130_fd_sc_hd__clkinv_1 U13810 ( .A(n16621), .Y(n16622) );
  sky130_fd_sc_hd__clkinv_1 U13811 ( .A(n25386), .Y(n24827) );
  sky130_fd_sc_hd__clkinv_1 U13812 ( .A(n16620), .Y(n16623) );
  sky130_fd_sc_hd__clkinv_1 U13813 ( .A(n16788), .Y(n16789) );
  sky130_fd_sc_hd__clkinv_1 U13814 ( .A(n22047), .Y(n19532) );
  sky130_fd_sc_hd__clkinv_1 U13815 ( .A(n24835), .Y(n24845) );
  sky130_fd_sc_hd__clkinv_1 U13816 ( .A(n19664), .Y(n19667) );
  sky130_fd_sc_hd__clkinv_1 U13817 ( .A(n19665), .Y(n19666) );
  sky130_fd_sc_hd__clkinv_1 U13818 ( .A(n21559), .Y(n21560) );
  sky130_fd_sc_hd__clkinv_1 U13819 ( .A(n21994), .Y(n21995) );
  sky130_fd_sc_hd__clkinv_1 U13820 ( .A(n25304), .Y(n19479) );
  sky130_fd_sc_hd__o21ai_2 U13821 ( .A1(n20323), .A2(n20324), .B1(n21134), .Y(
        j202_soc_core_j22_cpu_rf_N3190) );
  sky130_fd_sc_hd__clkinv_1 U13822 ( .A(n19300), .Y(n16626) );
  sky130_fd_sc_hd__clkinv_1 U13823 ( .A(n24874), .Y(n21501) );
  sky130_fd_sc_hd__clkinv_1 U13824 ( .A(n19213), .Y(n19214) );
  sky130_fd_sc_hd__o21ai_2 U13825 ( .A1(n20319), .A2(n20320), .B1(n21068), .Y(
        j202_soc_core_j22_cpu_rf_N3116) );
  sky130_fd_sc_hd__clkinv_1 U13826 ( .A(n24885), .Y(n24886) );
  sky130_fd_sc_hd__clkinv_1 U13827 ( .A(n18873), .Y(n18875) );
  sky130_fd_sc_hd__clkinv_1 U13828 ( .A(n19217), .Y(n19219) );
  sky130_fd_sc_hd__clkinv_1 U13829 ( .A(n16600), .Y(n19215) );
  sky130_fd_sc_hd__clkinv_1 U13830 ( .A(n17034), .Y(n17036) );
  sky130_fd_sc_hd__clkinv_1 U13831 ( .A(n16822), .Y(n16824) );
  sky130_fd_sc_hd__clkinv_1 U13832 ( .A(n17032), .Y(n18861) );
  sky130_fd_sc_hd__o21ai_2 U13833 ( .A1(n20319), .A2(n20325), .B1(n21205), .Y(
        j202_soc_core_j22_cpu_rf_N3079) );
  sky130_fd_sc_hd__clkinv_1 U13834 ( .A(n21583), .Y(n20776) );
  sky130_fd_sc_hd__o21ai_2 U13835 ( .A1(n20322), .A2(n20325), .B1(n21192), .Y(
        j202_soc_core_j22_cpu_rf_N2783) );
  sky130_fd_sc_hd__clkinv_1 U13836 ( .A(n19131), .Y(n19133) );
  sky130_fd_sc_hd__clkinv_1 U13837 ( .A(n19002), .Y(n19004) );
  sky130_fd_sc_hd__clkinv_1 U13838 ( .A(n18948), .Y(n19080) );
  sky130_fd_sc_hd__clkinv_1 U13839 ( .A(n19850), .Y(n19852) );
  sky130_fd_sc_hd__clkinv_1 U13840 ( .A(n21607), .Y(n21040) );
  sky130_fd_sc_hd__clkinv_1 U13841 ( .A(n18979), .Y(n18981) );
  sky130_fd_sc_hd__o21ai_2 U13842 ( .A1(n20279), .A2(n20481), .B1(n22369), .Y(
        j202_soc_core_j22_cpu_rf_N3371) );
  sky130_fd_sc_hd__clkinv_1 U13843 ( .A(n19100), .Y(n18978) );
  sky130_fd_sc_hd__clkinv_1 U13844 ( .A(n18860), .Y(n17033) );
  sky130_fd_sc_hd__o21ai_2 U13845 ( .A1(n20268), .A2(n20324), .B1(n21195), .Y(
        j202_soc_core_j22_cpu_rf_N3153) );
  sky130_fd_sc_hd__clkinv_1 U13846 ( .A(n16791), .Y(n19950) );
  sky130_fd_sc_hd__clkinv_1 U13847 ( .A(n22521), .Y(n20800) );
  sky130_fd_sc_hd__clkinv_1 U13848 ( .A(n21196), .Y(n21216) );
  sky130_fd_sc_hd__clkinv_1 U13849 ( .A(n25385), .Y(n20761) );
  sky130_fd_sc_hd__clkinv_1 U13850 ( .A(n25315), .Y(n19480) );
  sky130_fd_sc_hd__clkinv_1 U13851 ( .A(n22416), .Y(n21605) );
  sky130_fd_sc_hd__clkinv_1 U13852 ( .A(n24880), .Y(n24890) );
  sky130_fd_sc_hd__clkinv_1 U13853 ( .A(n18977), .Y(n19101) );
  sky130_fd_sc_hd__clkinv_1 U13854 ( .A(n19949), .Y(n16792) );
  sky130_fd_sc_hd__clkinv_1 U13855 ( .A(n24844), .Y(n24888) );
  sky130_fd_sc_hd__clkinv_1 U13856 ( .A(n19295), .Y(n19297) );
  sky130_fd_sc_hd__clkinv_1 U13857 ( .A(n16793), .Y(n16795) );
  sky130_fd_sc_hd__clkinv_1 U13858 ( .A(n17083), .Y(n18879) );
  sky130_fd_sc_hd__clkinv_1 U13859 ( .A(n25393), .Y(n22904) );
  sky130_fd_sc_hd__clkinv_1 U13860 ( .A(n19855), .Y(n19857) );
  sky130_fd_sc_hd__clkinv_1 U13861 ( .A(n18964), .Y(n18965) );
  sky130_fd_sc_hd__clkinv_1 U13862 ( .A(n22531), .Y(n20879) );
  sky130_fd_sc_hd__clkinv_1 U13863 ( .A(n18996), .Y(n16509) );
  sky130_fd_sc_hd__clkinv_1 U13864 ( .A(n16604), .Y(n19222) );
  sky130_fd_sc_hd__clkinv_1 U13865 ( .A(n18963), .Y(n18966) );
  sky130_fd_sc_hd__clkinv_1 U13866 ( .A(n19107), .Y(n19109) );
  sky130_fd_sc_hd__clkinv_1 U13867 ( .A(n19127), .Y(n16510) );
  sky130_fd_sc_hd__clkinv_1 U13868 ( .A(n22000), .Y(n20035) );
  sky130_fd_sc_hd__clkinv_1 U13869 ( .A(n18999), .Y(n19128) );
  sky130_fd_sc_hd__clkinv_1 U13870 ( .A(j202_soc_core_j22_cpu_rf_N2627), .Y(
        n22729) );
  sky130_fd_sc_hd__clkinv_1 U13871 ( .A(n18878), .Y(n17084) );
  sky130_fd_sc_hd__clkinv_1 U13872 ( .A(n19225), .Y(n16030) );
  sky130_fd_sc_hd__clkinv_1 U13873 ( .A(n17076), .Y(n17078) );
  sky130_fd_sc_hd__clkinv_1 U13874 ( .A(n10562), .Y(n20499) );
  sky130_fd_sc_hd__clkinv_1 U13875 ( .A(n16829), .Y(n16831) );
  sky130_fd_sc_hd__clkinv_1 U13876 ( .A(n18986), .Y(n18988) );
  sky130_fd_sc_hd__clkinv_1 U13877 ( .A(n17085), .Y(n17087) );
  sky130_fd_sc_hd__clkinv_1 U13878 ( .A(n22906), .Y(n22898) );
  sky130_fd_sc_hd__clkinv_1 U13879 ( .A(n16802), .Y(n16804) );
  sky130_fd_sc_hd__clkinv_1 U13880 ( .A(n19941), .Y(n19943) );
  sky130_fd_sc_hd__clkinv_1 U13881 ( .A(n19292), .Y(n16613) );
  sky130_fd_sc_hd__o21ai_2 U13882 ( .A1(n23236), .A2(n20481), .B1(n22366), .Y(
        j202_soc_core_j22_cpu_rf_N3301) );
  sky130_fd_sc_hd__clkinv_1 U13883 ( .A(n19954), .Y(n19956) );
  sky130_fd_sc_hd__clkinv_1 U13884 ( .A(n18855), .Y(n16521) );
  sky130_fd_sc_hd__clkinv_1 U13885 ( .A(n20546), .Y(n22527) );
  sky130_fd_sc_hd__clkinv_1 U13886 ( .A(n19287), .Y(n19289) );
  sky130_fd_sc_hd__clkinv_1 U13887 ( .A(n22538), .Y(n22539) );
  sky130_fd_sc_hd__clkinv_1 U13888 ( .A(n20778), .Y(n22522) );
  sky130_fd_sc_hd__clkinv_1 U13889 ( .A(n22528), .Y(n20617) );
  sky130_fd_sc_hd__clkinv_1 U13890 ( .A(n17330), .Y(n17333) );
  sky130_fd_sc_hd__clkinv_1 U13891 ( .A(n16782), .Y(n18852) );
  sky130_fd_sc_hd__clkinv_1 U13892 ( .A(n22523), .Y(n20928) );
  sky130_fd_sc_hd__clkinv_1 U13893 ( .A(n17320), .Y(n17323) );
  sky130_fd_sc_hd__clkinv_1 U13894 ( .A(n21398), .Y(n20666) );
  sky130_fd_sc_hd__clkinv_1 U13895 ( .A(n22721), .Y(n22124) );
  sky130_fd_sc_hd__clkinv_1 U13896 ( .A(n22728), .Y(n22718) );
  sky130_fd_sc_hd__clkinv_1 U13897 ( .A(n23224), .Y(n23227) );
  sky130_fd_sc_hd__clkinv_1 U13898 ( .A(n17044), .Y(n16017) );
  sky130_fd_sc_hd__clkinv_1 U13899 ( .A(n18865), .Y(n17043) );
  sky130_fd_sc_hd__clkinv_1 U13900 ( .A(n22541), .Y(n19890) );
  sky130_fd_sc_hd__clkinv_1 U13901 ( .A(n19097), .Y(n17028) );
  sky130_fd_sc_hd__clkinv_1 U13902 ( .A(n21045), .Y(n22517) );
  sky130_fd_sc_hd__clkinv_1 U13903 ( .A(n20196), .Y(n20202) );
  sky130_fd_sc_hd__clkinv_1 U13904 ( .A(n19095), .Y(n16575) );
  sky130_fd_sc_hd__clkinv_1 U13905 ( .A(n19093), .Y(n16574) );
  sky130_fd_sc_hd__clkinv_1 U13906 ( .A(n22525), .Y(n18465) );
  sky130_fd_sc_hd__clkinv_1 U13907 ( .A(n19012), .Y(n19014) );
  sky130_fd_sc_hd__clkinv_1 U13908 ( .A(n16632), .Y(n15980) );
  sky130_fd_sc_hd__clkinv_1 U13909 ( .A(n19307), .Y(n19309) );
  sky130_fd_sc_hd__clkinv_1 U13910 ( .A(n17228), .Y(n17221) );
  sky130_fd_sc_hd__clkinv_1 U13911 ( .A(n18967), .Y(n18969) );
  sky130_fd_sc_hd__clkinv_1 U13912 ( .A(n21155), .Y(n20809) );
  sky130_fd_sc_hd__clkinv_1 U13913 ( .A(n20825), .Y(n20826) );
  sky130_fd_sc_hd__clkinv_1 U13914 ( .A(n19668), .Y(n19670) );
  sky130_fd_sc_hd__clkinv_1 U13915 ( .A(n19140), .Y(n15975) );
  sky130_fd_sc_hd__inv_1 U13916 ( .A(n13537), .Y(n13538) );
  sky130_fd_sc_hd__clkinv_1 U13917 ( .A(n19348), .Y(n19349) );
  sky130_fd_sc_hd__clkinv_1 U13918 ( .A(n19875), .Y(n19157) );
  sky130_fd_sc_hd__clkinv_1 U13919 ( .A(n21163), .Y(n21118) );
  sky130_fd_sc_hd__clkinv_1 U13920 ( .A(n18883), .Y(n18885) );
  sky130_fd_sc_hd__clkinv_1 U13921 ( .A(n21154), .Y(n21029) );
  sky130_fd_sc_hd__clkinv_1 U13922 ( .A(n17094), .Y(n17096) );
  sky130_fd_sc_hd__clkinv_1 U13923 ( .A(n21166), .Y(n21049) );
  sky130_fd_sc_hd__clkinv_1 U13924 ( .A(n21387), .Y(n21390) );
  sky130_fd_sc_hd__clkinv_1 U13925 ( .A(n19864), .Y(n19866) );
  sky130_fd_sc_hd__clkinv_1 U13926 ( .A(n21382), .Y(n21350) );
  sky130_fd_sc_hd__clkinv_1 U13927 ( .A(n21167), .Y(n21053) );
  sky130_fd_sc_hd__clkinv_1 U13928 ( .A(n21116), .Y(n21153) );
  sky130_fd_sc_hd__clkinv_1 U13929 ( .A(n21156), .Y(n21157) );
  sky130_fd_sc_hd__clkinv_1 U13930 ( .A(n20651), .Y(n20714) );
  sky130_fd_sc_hd__clkinv_1 U13931 ( .A(n16839), .Y(n15954) );
  sky130_fd_sc_hd__clkinv_1 U13932 ( .A(n21375), .Y(n21359) );
  sky130_fd_sc_hd__clkinv_1 U13933 ( .A(n21379), .Y(n21347) );
  sky130_fd_sc_hd__clkinv_1 U13934 ( .A(n19921), .Y(n19355) );
  sky130_fd_sc_hd__clkinv_1 U13935 ( .A(n22883), .Y(n22877) );
  sky130_fd_sc_hd__clkinv_1 U13936 ( .A(n22298), .Y(n22304) );
  sky130_fd_sc_hd__clkinv_1 U13937 ( .A(n21085), .Y(n21144) );
  sky130_fd_sc_hd__clkinv_1 U13938 ( .A(n19880), .Y(n16668) );
  sky130_fd_sc_hd__clkinv_1 U13939 ( .A(n22592), .Y(n19153) );
  sky130_fd_sc_hd__clkinv_1 U13940 ( .A(n23298), .Y(n22375) );
  sky130_fd_sc_hd__clkinv_1 U13941 ( .A(n22070), .Y(n22068) );
  sky130_fd_sc_hd__clkinv_1 U13942 ( .A(n22183), .Y(n22754) );
  sky130_fd_sc_hd__clkinv_1 U13943 ( .A(n16298), .Y(n16269) );
  sky130_fd_sc_hd__clkinv_1 U13944 ( .A(n23313), .Y(n22599) );
  sky130_fd_sc_hd__clkinv_1 U13945 ( .A(n16346), .Y(n16336) );
  sky130_fd_sc_hd__clkinv_1 U13946 ( .A(n16270), .Y(n16236) );
  sky130_fd_sc_hd__clkinv_1 U13947 ( .A(n23301), .Y(n22116) );
  sky130_fd_sc_hd__clkinv_1 U13948 ( .A(n16543), .Y(n16562) );
  sky130_fd_sc_hd__clkinv_1 U13949 ( .A(n23344), .Y(n22607) );
  sky130_fd_sc_hd__clkinv_1 U13950 ( .A(n22441), .Y(n22651) );
  sky130_fd_sc_hd__clkinv_1 U13951 ( .A(n22874), .Y(n22878) );
  sky130_fd_sc_hd__clkinv_1 U13952 ( .A(n23316), .Y(n21878) );
  sky130_fd_sc_hd__clkinv_1 U13953 ( .A(n18629), .Y(n18759) );
  sky130_fd_sc_hd__clkinv_1 U13954 ( .A(n23322), .Y(n21840) );
  sky130_fd_sc_hd__clkinv_1 U13955 ( .A(n24292), .Y(n20083) );
  sky130_fd_sc_hd__clkinv_1 U13956 ( .A(n22351), .Y(n22164) );
  sky130_fd_sc_hd__clkinv_1 U13957 ( .A(n22064), .Y(n22161) );
  sky130_fd_sc_hd__clkinv_1 U13958 ( .A(n22314), .Y(n22169) );
  sky130_fd_sc_hd__clkinv_1 U13959 ( .A(n18282), .Y(n18284) );
  sky130_fd_sc_hd__clkinv_1 U13960 ( .A(n22300), .Y(n22159) );
  sky130_fd_sc_hd__clkinv_1 U13961 ( .A(n21985), .Y(n23336) );
  sky130_fd_sc_hd__clkinv_1 U13962 ( .A(n18146), .Y(n18148) );
  sky130_fd_sc_hd__clkinv_1 U13963 ( .A(n14715), .Y(n14409) );
  sky130_fd_sc_hd__clkinv_1 U13964 ( .A(n22349), .Y(n22355) );
  sky130_fd_sc_hd__clkinv_1 U13965 ( .A(n22074), .Y(n23333) );
  sky130_fd_sc_hd__clkinv_1 U13966 ( .A(n20481), .Y(n20236) );
  sky130_fd_sc_hd__clkinv_1 U13967 ( .A(n22711), .Y(n22179) );
  sky130_fd_sc_hd__clkinv_1 U13968 ( .A(n23614), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N393) );
  sky130_fd_sc_hd__clkinv_1 U13969 ( .A(n18099), .Y(n18003) );
  sky130_fd_sc_hd__clkinv_1 U13970 ( .A(n23613), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N392) );
  sky130_fd_sc_hd__clkinv_1 U13971 ( .A(n22602), .Y(n23327) );
  sky130_fd_sc_hd__clkinv_1 U13972 ( .A(n21807), .Y(n22166) );
  sky130_fd_sc_hd__clkinv_1 U13973 ( .A(n19936), .Y(n19557) );
  sky130_fd_sc_hd__clkinv_1 U13974 ( .A(n19591), .Y(n19560) );
  sky130_fd_sc_hd__clkinv_1 U13975 ( .A(n19625), .Y(n19626) );
  sky130_fd_sc_hd__clkinv_1 U13976 ( .A(n18029), .Y(n13218) );
  sky130_fd_sc_hd__clkinv_1 U13977 ( .A(n19803), .Y(n19594) );
  sky130_fd_sc_hd__clkinv_1 U13978 ( .A(n19769), .Y(n19771) );
  sky130_fd_sc_hd__clkinv_1 U13979 ( .A(n20026), .Y(n19365) );
  sky130_fd_sc_hd__clkinv_1 U13980 ( .A(n19419), .Y(n19421) );
  sky130_fd_sc_hd__clkinv_1 U13981 ( .A(n18663), .Y(n11349) );
  sky130_fd_sc_hd__clkinv_1 U13982 ( .A(n19441), .Y(n19443) );
  sky130_fd_sc_hd__clkinv_1 U13983 ( .A(n10559), .Y(n22808) );
  sky130_fd_sc_hd__clkinv_1 U13984 ( .A(n19550), .Y(n19551) );
  sky130_fd_sc_hd__clkinv_1 U13985 ( .A(n19694), .Y(n19696) );
  sky130_fd_sc_hd__clkinv_1 U13986 ( .A(n19389), .Y(n19369) );
  sky130_fd_sc_hd__clkinv_1 U13987 ( .A(n19523), .Y(n19525) );
  sky130_fd_sc_hd__clkinv_1 U13988 ( .A(n17536), .Y(n17802) );
  sky130_fd_sc_hd__clkinv_1 U13989 ( .A(n14355), .Y(n14356) );
  sky130_fd_sc_hd__clkinv_1 U13990 ( .A(n18433), .Y(n17590) );
  sky130_fd_sc_hd__clkinv_1 U13991 ( .A(n21806), .Y(n21811) );
  sky130_fd_sc_hd__clkinv_1 U13992 ( .A(n17917), .Y(n17658) );
  sky130_fd_sc_hd__clkinv_1 U13994 ( .A(n14736), .Y(n14741) );
  sky130_fd_sc_hd__clkinv_1 U13995 ( .A(n21018), .Y(n20365) );
  sky130_fd_sc_hd__clkinv_1 U13996 ( .A(n20151), .Y(n20187) );
  sky130_fd_sc_hd__clkinv_1 U13997 ( .A(n16659), .Y(n22581) );
  sky130_fd_sc_hd__clkinv_1 U13998 ( .A(n17872), .Y(n18352) );
  sky130_fd_sc_hd__clkinv_1 U13999 ( .A(n17947), .Y(n18404) );
  sky130_fd_sc_hd__clkinv_1 U14000 ( .A(n24893), .Y(n23238) );
  sky130_fd_sc_hd__clkinv_1 U14001 ( .A(n19743), .Y(n19745) );
  sky130_fd_sc_hd__clkinv_1 U14002 ( .A(n17511), .Y(n17500) );
  sky130_fd_sc_hd__clkinv_1 U14003 ( .A(n22579), .Y(n22604) );
  sky130_fd_sc_hd__clkinv_1 U14004 ( .A(n14423), .Y(n14444) );
  sky130_fd_sc_hd__clkinv_1 U14005 ( .A(n11381), .Y(n11373) );
  sky130_fd_sc_hd__clkinv_1 U14006 ( .A(n11375), .Y(n15191) );
  sky130_fd_sc_hd__clkinv_1 U14007 ( .A(n14156), .Y(n14160) );
  sky130_fd_sc_hd__clkinv_1 U14008 ( .A(n23250), .Y(n25543) );
  sky130_fd_sc_hd__clkinv_1 U14009 ( .A(n17961), .Y(n18085) );
  sky130_fd_sc_hd__clkinv_1 U14010 ( .A(n17525), .Y(n17556) );
  sky130_fd_sc_hd__clkinv_1 U14011 ( .A(n14731), .Y(n14732) );
  sky130_fd_sc_hd__clkinv_1 U14012 ( .A(n16595), .Y(n21728) );
  sky130_fd_sc_hd__clkinv_1 U14013 ( .A(n17378), .Y(n17381) );
  sky130_fd_sc_hd__clkinv_1 U14014 ( .A(n18030), .Y(n17965) );
  sky130_fd_sc_hd__clkinv_1 U14015 ( .A(n22584), .Y(n22146) );
  sky130_fd_sc_hd__clkinv_1 U14016 ( .A(n22631), .Y(n20955) );
  sky130_fd_sc_hd__clkinv_1 U14017 ( .A(n11266), .Y(n13308) );
  sky130_fd_sc_hd__clkinv_1 U14018 ( .A(n20496), .Y(n20430) );
  sky130_fd_sc_hd__clkinv_1 U14019 ( .A(n22313), .Y(n22318) );
  sky130_fd_sc_hd__clkinv_1 U14020 ( .A(n22591), .Y(n22608) );
  sky130_fd_sc_hd__clkinv_1 U14021 ( .A(n21616), .Y(n21620) );
  sky130_fd_sc_hd__clkinv_1 U14022 ( .A(n18774), .Y(n18516) );
  sky130_fd_sc_hd__clkinv_1 U14023 ( .A(n21657), .Y(n21672) );
  sky130_fd_sc_hd__clkinv_1 U14024 ( .A(n17258), .Y(n17261) );
  sky130_fd_sc_hd__clkinv_1 U14025 ( .A(n15151), .Y(n18255) );
  sky130_fd_sc_hd__clkinv_1 U14026 ( .A(n16988), .Y(n17001) );
  sky130_fd_sc_hd__clkinv_1 U14027 ( .A(n13240), .Y(n18044) );
  sky130_fd_sc_hd__clkinv_1 U14028 ( .A(n18134), .Y(n13208) );
  sky130_fd_sc_hd__clkinv_1 U14029 ( .A(n17300), .Y(n17303) );
  sky130_fd_sc_hd__clkinv_1 U14030 ( .A(n20154), .Y(n20143) );
  sky130_fd_sc_hd__clkinv_1 U14031 ( .A(n18112), .Y(n18143) );
  sky130_fd_sc_hd__clkinv_1 U14032 ( .A(n17940), .Y(n17869) );
  sky130_fd_sc_hd__clkinv_1 U14033 ( .A(n17257), .Y(n17253) );
  sky130_fd_sc_hd__clkinv_1 U14034 ( .A(n21174), .Y(n20845) );
  sky130_fd_sc_hd__clkinv_1 U14035 ( .A(n17971), .Y(n18039) );
  sky130_fd_sc_hd__clkinv_1 U14036 ( .A(n21010), .Y(n19167) );
  sky130_fd_sc_hd__clkinv_1 U14037 ( .A(n18659), .Y(n18679) );
  sky130_fd_sc_hd__clkinv_1 U14038 ( .A(n18136), .Y(n18043) );
  sky130_fd_sc_hd__clkinv_1 U14039 ( .A(n18263), .Y(n18265) );
  sky130_fd_sc_hd__clkinv_1 U14040 ( .A(n17748), .Y(n17937) );
  sky130_fd_sc_hd__clkinv_1 U14041 ( .A(n14217), .Y(n14334) );
  sky130_fd_sc_hd__clkinv_1 U14042 ( .A(n14833), .Y(n14451) );
  sky130_fd_sc_hd__clkinv_1 U14043 ( .A(n17293), .Y(n17296) );
  sky130_fd_sc_hd__clkinv_1 U14044 ( .A(n17902), .Y(n16766) );
  sky130_fd_sc_hd__clkinv_1 U14045 ( .A(n13432), .Y(n13438) );
  sky130_fd_sc_hd__clkinv_1 U14046 ( .A(n14849), .Y(n14855) );
  sky130_fd_sc_hd__clkinv_1 U14047 ( .A(n21926), .Y(n21933) );
  sky130_fd_sc_hd__clkinv_1 U14048 ( .A(n17670), .Y(n17876) );
  sky130_fd_sc_hd__clkinv_1 U14049 ( .A(n17773), .Y(n17615) );
  sky130_fd_sc_hd__clkinv_1 U14050 ( .A(n17865), .Y(n17845) );
  sky130_fd_sc_hd__clkinv_1 U14051 ( .A(n17928), .Y(n17502) );
  sky130_fd_sc_hd__clkinv_1 U14052 ( .A(n15036), .Y(n15011) );
  sky130_fd_sc_hd__clkinv_1 U14053 ( .A(n18641), .Y(n18782) );
  sky130_fd_sc_hd__clkinv_1 U14054 ( .A(n17739), .Y(n17537) );
  sky130_fd_sc_hd__clkinv_1 U14055 ( .A(n18266), .Y(n16908) );
  sky130_fd_sc_hd__clkinv_1 U14056 ( .A(n16759), .Y(n17843) );
  sky130_fd_sc_hd__clkinv_1 U14057 ( .A(j202_soc_core_ahbcs_6__HREADY_), .Y(
        n20488) );
  sky130_fd_sc_hd__clkinv_1 U14058 ( .A(n17805), .Y(n17801) );
  sky130_fd_sc_hd__clkinv_1 U14059 ( .A(n18670), .Y(n18677) );
  sky130_fd_sc_hd__clkinv_1 U14060 ( .A(n17551), .Y(n17747) );
  sky130_fd_sc_hd__clkinv_1 U14061 ( .A(n21796), .Y(n17099) );
  sky130_fd_sc_hd__clkinv_1 U14062 ( .A(n22866), .Y(n21235) );
  sky130_fd_sc_hd__clkinv_1 U14063 ( .A(n13584), .Y(n18035) );
  sky130_fd_sc_hd__clkinv_1 U14064 ( .A(n17942), .Y(n17656) );
  sky130_fd_sc_hd__clkinv_1 U14065 ( .A(n17516), .Y(n17613) );
  sky130_fd_sc_hd__clkinv_1 U14066 ( .A(n25370), .Y(n21344) );
  sky130_fd_sc_hd__clkinv_1 U14067 ( .A(n20905), .Y(n20641) );
  sky130_fd_sc_hd__clkinv_1 U14068 ( .A(n21027), .Y(n21028) );
  sky130_fd_sc_hd__clkinv_1 U14069 ( .A(n18444), .Y(n18401) );
  sky130_fd_sc_hd__and2_0 U14070 ( .A(n21139), .B(n17107), .X(n20904) );
  sky130_fd_sc_hd__clkinv_1 U14071 ( .A(n16977), .Y(n18709) );
  sky130_fd_sc_hd__clkinv_1 U14072 ( .A(n14618), .Y(n14622) );
  sky130_fd_sc_hd__clkinv_1 U14073 ( .A(n16907), .Y(n18688) );
  sky130_fd_sc_hd__clkinv_1 U14074 ( .A(n17495), .Y(n18430) );
  sky130_fd_sc_hd__clkinv_1 U14075 ( .A(n18554), .Y(n18527) );
  sky130_fd_sc_hd__clkinv_1 U14076 ( .A(n17557), .Y(n17744) );
  sky130_fd_sc_hd__clkinv_1 U14077 ( .A(n17943), .Y(n17620) );
  sky130_fd_sc_hd__clkinv_1 U14078 ( .A(n17554), .Y(n17600) );
  sky130_fd_sc_hd__clkinv_1 U14079 ( .A(n19317), .Y(n20020) );
  sky130_fd_sc_hd__clkinv_1 U14080 ( .A(n17863), .Y(n17941) );
  sky130_fd_sc_hd__clkinv_1 U14081 ( .A(n17591), .Y(n17592) );
  sky130_fd_sc_hd__clkinv_1 U14082 ( .A(n18379), .Y(n18245) );
  sky130_fd_sc_hd__clkinv_1 U14083 ( .A(n16997), .Y(n16998) );
  sky130_fd_sc_hd__clkinv_1 U14084 ( .A(n19953), .Y(n20038) );
  sky130_fd_sc_hd__clkinv_1 U14085 ( .A(n18144), .Y(n18114) );
  sky130_fd_sc_hd__clkinv_1 U14086 ( .A(n14323), .Y(n14324) );
  sky130_fd_sc_hd__clkinv_1 U14087 ( .A(n22863), .Y(n22864) );
  sky130_fd_sc_hd__clkinv_1 U14088 ( .A(n17972), .Y(n13554) );
  sky130_fd_sc_hd__clkinv_1 U14089 ( .A(n18135), .Y(n13220) );
  sky130_fd_sc_hd__clkinv_1 U14090 ( .A(n13254), .Y(n13242) );
  sky130_fd_sc_hd__clkinv_1 U14091 ( .A(n13234), .Y(n17969) );
  sky130_fd_sc_hd__clkinv_1 U14092 ( .A(n13215), .Y(n18102) );
  sky130_fd_sc_hd__clkinv_1 U14093 ( .A(n13586), .Y(n17958) );
  sky130_fd_sc_hd__clkinv_1 U14094 ( .A(n18037), .Y(n13247) );
  sky130_fd_sc_hd__clkinv_1 U14095 ( .A(n13257), .Y(n18123) );
  sky130_fd_sc_hd__clkinv_1 U14096 ( .A(n14195), .Y(n14345) );
  sky130_fd_sc_hd__clkinv_1 U14097 ( .A(n18343), .Y(n18416) );
  sky130_fd_sc_hd__clkinv_1 U14098 ( .A(n11357), .Y(n18595) );
  sky130_fd_sc_hd__clkinv_1 U14099 ( .A(n15118), .Y(n18533) );
  sky130_fd_sc_hd__clkinv_1 U14100 ( .A(n18790), .Y(n18589) );
  sky130_fd_sc_hd__clkinv_1 U14101 ( .A(n18700), .Y(n18768) );
  sky130_fd_sc_hd__clkinv_1 U14102 ( .A(n13600), .Y(n18015) );
  sky130_fd_sc_hd__clkinv_1 U14103 ( .A(n18537), .Y(n16978) );
  sky130_fd_sc_hd__clkinv_1 U14104 ( .A(n14695), .Y(n14778) );
  sky130_fd_sc_hd__clkinv_1 U14105 ( .A(n14885), .Y(n14768) );
  sky130_fd_sc_hd__clkinv_1 U14106 ( .A(n22289), .Y(n22294) );
  sky130_fd_sc_hd__clkinv_1 U14107 ( .A(n17725), .Y(n17654) );
  sky130_fd_sc_hd__clkinv_1 U14108 ( .A(n14692), .Y(n14457) );
  sky130_fd_sc_hd__clkinv_1 U14109 ( .A(n15065), .Y(n11256) );
  sky130_fd_sc_hd__clkinv_1 U14110 ( .A(n13111), .Y(n13300) );
  sky130_fd_sc_hd__clkinv_1 U14111 ( .A(n13502), .Y(n11258) );
  sky130_fd_sc_hd__clkinv_1 U14112 ( .A(n13172), .Y(n13485) );
  sky130_fd_sc_hd__clkinv_1 U14113 ( .A(n13457), .Y(n11277) );
  sky130_fd_sc_hd__clkinv_1 U14114 ( .A(n11278), .Y(n13126) );
  sky130_fd_sc_hd__clkinv_1 U14115 ( .A(n14446), .Y(n14401) );
  sky130_fd_sc_hd__clkinv_1 U14116 ( .A(n25065), .Y(n25047) );
  sky130_fd_sc_hd__clkinv_1 U14117 ( .A(n11511), .Y(n11445) );
  sky130_fd_sc_hd__clkinv_1 U14118 ( .A(n14766), .Y(n14877) );
  sky130_fd_sc_hd__clkinv_1 U14119 ( .A(n14486), .Y(n14462) );
  sky130_fd_sc_hd__clkinv_1 U14120 ( .A(n16916), .Y(n18564) );
  sky130_fd_sc_hd__clkinv_1 U14121 ( .A(n17984), .Y(n18115) );
  sky130_fd_sc_hd__clkinv_1 U14122 ( .A(n13307), .Y(n13453) );
  sky130_fd_sc_hd__clkinv_1 U14123 ( .A(n11264), .Y(n13112) );
  sky130_fd_sc_hd__clkinv_1 U14124 ( .A(n14597), .Y(n13037) );
  sky130_fd_sc_hd__clkinv_1 U14125 ( .A(n18680), .Y(n18643) );
  sky130_fd_sc_hd__clkinv_1 U14126 ( .A(n18522), .Y(n16987) );
  sky130_fd_sc_hd__clkinv_1 U14127 ( .A(n16901), .Y(n18644) );
  sky130_fd_sc_hd__clkinv_1 U14128 ( .A(n13487), .Y(n13411) );
  sky130_fd_sc_hd__clkinv_1 U14129 ( .A(n15527), .Y(n15621) );
  sky130_fd_sc_hd__clkinv_1 U14130 ( .A(n15182), .Y(n18592) );
  sky130_fd_sc_hd__clkinv_1 U14131 ( .A(n13608), .Y(n18086) );
  sky130_fd_sc_hd__clkinv_1 U14132 ( .A(n14454), .Y(n14772) );
  sky130_fd_sc_hd__clkinv_1 U14133 ( .A(n13237), .Y(n18034) );
  sky130_fd_sc_hd__clkinv_1 U14134 ( .A(n17875), .Y(n17746) );
  sky130_fd_sc_hd__clkinv_1 U14135 ( .A(n17997), .Y(n18118) );
  sky130_fd_sc_hd__clkinv_1 U14136 ( .A(n13589), .Y(n11224) );
  sky130_fd_sc_hd__clkinv_1 U14137 ( .A(n18675), .Y(n15153) );
  sky130_fd_sc_hd__clkinv_1 U14138 ( .A(n18514), .Y(n18687) );
  sky130_fd_sc_hd__clkinv_1 U14139 ( .A(n13493), .Y(n13435) );
  sky130_fd_sc_hd__clkinv_1 U14140 ( .A(n18710), .Y(n18698) );
  sky130_fd_sc_hd__clkinv_1 U14141 ( .A(n18584), .Y(n18569) );
  sky130_fd_sc_hd__clkinv_1 U14142 ( .A(n16925), .Y(n18770) );
  sky130_fd_sc_hd__clkinv_1 U14143 ( .A(n13312), .Y(n13330) );
  sky130_fd_sc_hd__clkinv_1 U14144 ( .A(n17866), .Y(n18347) );
  sky130_fd_sc_hd__clkinv_1 U14145 ( .A(n18702), .Y(n18639) );
  sky130_fd_sc_hd__clkinv_1 U14146 ( .A(n18005), .Y(n18119) );
  sky130_fd_sc_hd__clkinv_1 U14147 ( .A(n11280), .Y(n11263) );
  sky130_fd_sc_hd__clkinv_1 U14148 ( .A(n13167), .Y(n11234) );
  sky130_fd_sc_hd__clkinv_1 U14149 ( .A(n15121), .Y(n18660) );
  sky130_fd_sc_hd__clkinv_1 U14150 ( .A(n13042), .Y(n13043) );
  sky130_fd_sc_hd__clkinv_1 U14151 ( .A(n18524), .Y(n18681) );
  sky130_fd_sc_hd__clkinv_1 U14152 ( .A(n13422), .Y(n13380) );
  sky130_fd_sc_hd__clkinv_1 U14153 ( .A(n15122), .Y(n16924) );
  sky130_fd_sc_hd__clkinv_1 U14154 ( .A(n13607), .Y(n13555) );
  sky130_fd_sc_hd__clkinv_1 U14155 ( .A(n16996), .Y(n18642) );
  sky130_fd_sc_hd__clkinv_1 U14156 ( .A(n17963), .Y(n18179) );
  sky130_fd_sc_hd__clkinv_1 U14157 ( .A(n18512), .Y(n18521) );
  sky130_fd_sc_hd__clkinv_1 U14158 ( .A(n11227), .Y(n13170) );
  sky130_fd_sc_hd__clkinv_1 U14159 ( .A(n18673), .Y(n18713) );
  sky130_fd_sc_hd__clkinv_1 U14160 ( .A(n18341), .Y(n17611) );
  sky130_fd_sc_hd__clkinv_1 U14161 ( .A(n13236), .Y(n13255) );
  sky130_fd_sc_hd__clkinv_1 U14162 ( .A(n15194), .Y(n18784) );
  sky130_fd_sc_hd__clkinv_1 U14163 ( .A(n14567), .Y(n14579) );
  sky130_fd_sc_hd__clkinv_1 U14164 ( .A(n14162), .Y(n14811) );
  sky130_fd_sc_hd__clkinv_1 U14165 ( .A(n14146), .Y(n14417) );
  sky130_fd_sc_hd__clkinv_1 U14166 ( .A(n18397), .Y(n17617) );
  sky130_fd_sc_hd__clkinv_1 U14167 ( .A(n16195), .Y(n15454) );
  sky130_fd_sc_hd__clkinv_1 U14168 ( .A(n14448), .Y(n14416) );
  sky130_fd_sc_hd__clkinv_1 U14169 ( .A(n17618), .Y(n18436) );
  sky130_fd_sc_hd__clkinv_1 U14170 ( .A(n14808), .Y(n14814) );
  sky130_fd_sc_hd__clkinv_1 U14171 ( .A(n18392), .Y(n17757) );
  sky130_fd_sc_hd__clkinv_1 U14172 ( .A(n13235), .Y(n18101) );
  sky130_fd_sc_hd__clkinv_1 U14173 ( .A(n20161), .Y(n20167) );
  sky130_fd_sc_hd__clkinv_1 U14174 ( .A(n14474), .Y(n14458) );
  sky130_fd_sc_hd__clkinv_1 U14175 ( .A(n17478), .Y(n18418) );
  sky130_fd_sc_hd__clkinv_1 U14176 ( .A(n13041), .Y(n13007) );
  sky130_fd_sc_hd__clkinv_1 U14177 ( .A(n17916), .Y(n17868) );
  sky130_fd_sc_hd__clkinv_1 U14178 ( .A(n17784), .Y(n17534) );
  sky130_fd_sc_hd__clkinv_1 U14179 ( .A(n17945), .Y(n17653) );
  sky130_fd_sc_hd__clkinv_1 U14180 ( .A(n14157), .Y(n14494) );
  sky130_fd_sc_hd__clkinv_1 U14181 ( .A(n13324), .Y(n13369) );
  sky130_fd_sc_hd__clkinv_1 U14182 ( .A(n17509), .Y(n16764) );
  sky130_fd_sc_hd__clkinv_1 U14183 ( .A(n14881), .Y(n14782) );
  sky130_fd_sc_hd__clkinv_1 U14184 ( .A(n17774), .Y(n17596) );
  sky130_fd_sc_hd__clkinv_1 U14185 ( .A(n17910), .Y(n17779) );
  sky130_fd_sc_hd__clkinv_1 U14186 ( .A(n18446), .Y(n17944) );
  sky130_fd_sc_hd__clkinv_1 U14187 ( .A(n18346), .Y(n17752) );
  sky130_fd_sc_hd__clkinv_1 U14188 ( .A(n14337), .Y(n14338) );
  sky130_fd_sc_hd__clkinv_1 U14189 ( .A(n14625), .Y(n14277) );
  sky130_fd_sc_hd__clkinv_1 U14190 ( .A(n23462), .Y(n23464) );
  sky130_fd_sc_hd__clkinv_1 U14191 ( .A(n18703), .Y(n18558) );
  sky130_fd_sc_hd__clkinv_1 U14192 ( .A(n17717), .Y(n15069) );
  sky130_fd_sc_hd__clkinv_1 U14193 ( .A(n17662), .Y(n17678) );
  sky130_fd_sc_hd__clkinv_1 U14194 ( .A(n15368), .Y(n15523) );
  sky130_fd_sc_hd__clkinv_1 U14195 ( .A(n18031), .Y(n13224) );
  sky130_fd_sc_hd__clkinv_1 U14196 ( .A(n23589), .Y(n23751) );
  sky130_fd_sc_hd__clkinv_1 U14197 ( .A(n18543), .Y(n15199) );
  sky130_fd_sc_hd__clkinv_1 U14198 ( .A(n14880), .Y(n14481) );
  sky130_fd_sc_hd__clkinv_1 U14199 ( .A(n18168), .Y(n18026) );
  sky130_fd_sc_hd__clkinv_1 U14200 ( .A(n14553), .Y(n14592) );
  sky130_fd_sc_hd__clkinv_1 U14201 ( .A(n18045), .Y(n13587) );
  sky130_fd_sc_hd__clkinv_1 U14202 ( .A(n18289), .Y(n18312) );
  sky130_fd_sc_hd__clkinv_1 U14203 ( .A(n17675), .Y(n17795) );
  sky130_fd_sc_hd__clkinv_1 U14204 ( .A(n16184), .Y(n16436) );
  sky130_fd_sc_hd__clkinv_1 U14205 ( .A(n21651), .Y(n21656) );
  sky130_fd_sc_hd__clkinv_1 U14206 ( .A(n16983), .Y(n16984) );
  sky130_fd_sc_hd__clkinv_1 U14207 ( .A(n18557), .Y(n16974) );
  sky130_fd_sc_hd__clkinv_1 U14208 ( .A(n14860), .Y(n14433) );
  sky130_fd_sc_hd__clkinv_1 U14209 ( .A(n23528), .Y(n25064) );
  sky130_fd_sc_hd__clkinv_1 U14210 ( .A(n21011), .Y(n22707) );
  sky130_fd_sc_hd__clkinv_1 U14211 ( .A(n17799), .Y(n18248) );
  sky130_fd_sc_hd__clkinv_1 U14212 ( .A(n22034), .Y(n22041) );
  sky130_fd_sc_hd__clkinv_1 U14213 ( .A(n21237), .Y(n16690) );
  sky130_fd_sc_hd__clkinv_1 U14214 ( .A(n18435), .Y(n17771) );
  sky130_fd_sc_hd__clkinv_1 U14215 ( .A(n17737), .Y(n16737) );
  sky130_fd_sc_hd__clkinv_1 U14216 ( .A(n16898), .Y(n18290) );
  sky130_fd_sc_hd__clkinv_1 U14217 ( .A(n14477), .Y(n14872) );
  sky130_fd_sc_hd__clkinv_1 U14218 ( .A(n17768), .Y(n17593) );
  sky130_fd_sc_hd__clkinv_1 U14219 ( .A(n14876), .Y(n14490) );
  sky130_fd_sc_hd__clkinv_1 U14220 ( .A(n14419), .Y(n14422) );
  sky130_fd_sc_hd__clkinv_1 U14221 ( .A(n17624), .Y(n18345) );
  sky130_fd_sc_hd__clkinv_1 U14222 ( .A(n18674), .Y(n18559) );
  sky130_fd_sc_hd__clkinv_1 U14223 ( .A(n16968), .Y(n15189) );
  sky130_fd_sc_hd__clkinv_1 U14224 ( .A(n17911), .Y(n17727) );
  sky130_fd_sc_hd__clkinv_1 U14225 ( .A(n14142), .Y(n14679) );
  sky130_fd_sc_hd__clkinv_1 U14226 ( .A(n17923), .Y(n17860) );
  sky130_fd_sc_hd__clkinv_1 U14227 ( .A(n23600), .Y(n23601) );
  sky130_fd_sc_hd__clkinv_1 U14228 ( .A(n15318), .Y(n15434) );
  sky130_fd_sc_hd__clkinv_1 U14229 ( .A(n18253), .Y(n18291) );
  sky130_fd_sc_hd__clkinv_1 U14230 ( .A(n23602), .Y(n23603) );
  sky130_fd_sc_hd__clkinv_1 U14231 ( .A(n17672), .Y(n17935) );
  sky130_fd_sc_hd__clkinv_1 U14232 ( .A(n14414), .Y(n14784) );
  sky130_fd_sc_hd__clkinv_1 U14233 ( .A(n14777), .Y(n13547) );
  sky130_fd_sc_hd__clkinv_1 U14234 ( .A(n18588), .Y(n18766) );
  sky130_fd_sc_hd__clkinv_1 U14235 ( .A(n14154), .Y(n14476) );
  sky130_fd_sc_hd__clkinv_1 U14236 ( .A(n19239), .Y(n19891) );
  sky130_fd_sc_hd__clkinv_1 U14237 ( .A(n18399), .Y(n17619) );
  sky130_fd_sc_hd__clkinv_1 U14239 ( .A(n14822), .Y(n14781) );
  sky130_fd_sc_hd__clkinv_1 U14240 ( .A(n11389), .Y(n18361) );
  sky130_fd_sc_hd__clkinv_1 U14241 ( .A(n14447), .Y(n14828) );
  sky130_fd_sc_hd__clkinv_1 U14242 ( .A(n17548), .Y(n17621) );
  sky130_fd_sc_hd__clkinv_1 U14243 ( .A(n14854), .Y(n14861) );
  sky130_fd_sc_hd__clkinv_1 U14244 ( .A(n19232), .Y(n19233) );
  sky130_fd_sc_hd__clkinv_1 U14245 ( .A(n17912), .Y(n17498) );
  sky130_fd_sc_hd__clkinv_1 U14246 ( .A(n14570), .Y(n14581) );
  sky130_fd_sc_hd__clkinv_1 U14247 ( .A(n14459), .Y(n14460) );
  sky130_fd_sc_hd__clkinv_1 U14248 ( .A(n17791), .Y(n17847) );
  sky130_fd_sc_hd__clkinv_1 U14249 ( .A(n14991), .Y(n17785) );
  sky130_fd_sc_hd__clkinv_1 U14250 ( .A(n21212), .Y(n19379) );
  sky130_fd_sc_hd__clkinv_1 U14251 ( .A(n18638), .Y(n15184) );
  sky130_fd_sc_hd__clkinv_1 U14252 ( .A(n18585), .Y(n18662) );
  sky130_fd_sc_hd__clkinv_1 U14253 ( .A(n13919), .Y(n11814) );
  sky130_fd_sc_hd__clkinv_1 U14254 ( .A(n13920), .Y(n11817) );
  sky130_fd_sc_hd__clkinv_1 U14255 ( .A(n18007), .Y(n18041) );
  sky130_fd_sc_hd__clkinv_1 U14256 ( .A(n18173), .Y(n18040) );
  sky130_fd_sc_hd__clkinv_1 U14257 ( .A(n11265), .Y(n13311) );
  sky130_fd_sc_hd__clkinv_1 U14258 ( .A(n13567), .Y(n13241) );
  sky130_fd_sc_hd__clkinv_1 U14259 ( .A(n13333), .Y(n13480) );
  sky130_fd_sc_hd__clkinv_1 U14260 ( .A(n13581), .Y(n13553) );
  sky130_fd_sc_hd__clkinv_1 U14261 ( .A(n13454), .Y(n13314) );
  sky130_fd_sc_hd__clkinv_1 U14262 ( .A(n13212), .Y(n13595) );
  sky130_fd_sc_hd__clkinv_1 U14263 ( .A(n13001), .Y(n14300) );
  sky130_fd_sc_hd__clkinv_1 U14264 ( .A(n21250), .Y(n21252) );
  sky130_fd_sc_hd__clkinv_1 U14265 ( .A(n14284), .Y(n14330) );
  sky130_fd_sc_hd__clkinv_1 U14266 ( .A(n14344), .Y(n14554) );
  sky130_fd_sc_hd__clkinv_1 U14267 ( .A(n13334), .Y(n13134) );
  sky130_fd_sc_hd__clkinv_1 U14268 ( .A(n14550), .Y(n14358) );
  sky130_fd_sc_hd__clkinv_1 U14269 ( .A(n12116), .Y(n12121) );
  sky130_fd_sc_hd__clkinv_1 U14270 ( .A(n13040), .Y(n14538) );
  sky130_fd_sc_hd__clkinv_1 U14271 ( .A(n13223), .Y(n17991) );
  sky130_fd_sc_hd__clkinv_1 U14272 ( .A(n18100), .Y(n18133) );
  sky130_fd_sc_hd__clkinv_1 U14273 ( .A(n23345), .Y(n23296) );
  sky130_fd_sc_hd__clkinv_1 U14274 ( .A(n13123), .Y(n11259) );
  sky130_fd_sc_hd__clkinv_1 U14275 ( .A(n13434), .Y(n13492) );
  sky130_fd_sc_hd__clkinv_1 U14276 ( .A(n23756), .Y(n23762) );
  sky130_fd_sc_hd__clkinv_1 U14277 ( .A(n14188), .Y(n14189) );
  sky130_fd_sc_hd__clkinv_1 U14278 ( .A(n18125), .Y(n13551) );
  sky130_fd_sc_hd__clkinv_1 U14279 ( .A(n13440), .Y(n13494) );
  sky130_fd_sc_hd__clkinv_1 U14280 ( .A(n14155), .Y(n14683) );
  sky130_fd_sc_hd__clkinv_1 U14281 ( .A(n13136), .Y(n13329) );
  sky130_fd_sc_hd__clkinv_1 U14282 ( .A(n18092), .Y(n13253) );
  sky130_fd_sc_hd__clkinv_1 U14283 ( .A(n17988), .Y(n14680) );
  sky130_fd_sc_hd__clkinv_1 U14284 ( .A(n18091), .Y(n18081) );
  sky130_fd_sc_hd__clkinv_1 U14285 ( .A(n13165), .Y(n13433) );
  sky130_fd_sc_hd__clkinv_1 U14286 ( .A(n14022), .Y(n14068) );
  sky130_fd_sc_hd__clkinv_1 U14287 ( .A(n22147), .Y(n12948) );
  sky130_fd_sc_hd__clkinv_1 U14288 ( .A(n14113), .Y(n14119) );
  sky130_fd_sc_hd__clkinv_1 U14289 ( .A(n21676), .Y(n12951) );
  sky130_fd_sc_hd__clkinv_1 U14290 ( .A(n23450), .Y(n23366) );
  sky130_fd_sc_hd__clkinv_1 U14291 ( .A(n22692), .Y(n22668) );
  sky130_fd_sc_hd__clkinv_1 U14292 ( .A(n20248), .Y(n12915) );
  sky130_fd_sc_hd__clkinv_1 U14293 ( .A(n17711), .Y(n17712) );
  sky130_fd_sc_hd__clkinv_1 U14294 ( .A(n14404), .Y(n14103) );
  sky130_fd_sc_hd__clkinv_1 U14295 ( .A(n17469), .Y(n14412) );
  sky130_fd_sc_hd__clkinv_1 U14296 ( .A(n14314), .Y(n14110) );
  sky130_fd_sc_hd__clkinv_1 U14297 ( .A(n15272), .Y(n15347) );
  sky130_fd_sc_hd__clkinv_1 U14298 ( .A(n24073), .Y(n20130) );
  sky130_fd_sc_hd__clkinv_1 U14299 ( .A(n11347), .Y(n13412) );
  sky130_fd_sc_hd__clkinv_1 U14300 ( .A(n14296), .Y(n14104) );
  sky130_fd_sc_hd__clkinv_1 U14301 ( .A(n12539), .Y(n12425) );
  sky130_fd_sc_hd__clkinv_1 U14302 ( .A(n14293), .Y(n14571) );
  sky130_fd_sc_hd__clkinv_1 U14303 ( .A(n11363), .Y(n11209) );
  sky130_fd_sc_hd__clkinv_1 U14304 ( .A(n13032), .Y(n14161) );
  sky130_fd_sc_hd__clkinv_1 U14305 ( .A(n21339), .Y(n20347) );
  sky130_fd_sc_hd__clkinv_1 U14306 ( .A(n13328), .Y(n13124) );
  sky130_fd_sc_hd__clkinv_1 U14307 ( .A(n14837), .Y(n14117) );
  sky130_fd_sc_hd__clkinv_1 U14308 ( .A(n15334), .Y(n15423) );
  sky130_fd_sc_hd__clkinv_1 U14309 ( .A(n15335), .Y(n15416) );
  sky130_fd_sc_hd__clkinv_1 U14310 ( .A(n17413), .Y(n17415) );
  sky130_fd_sc_hd__clkinv_1 U14311 ( .A(n22058), .Y(n22055) );
  sky130_fd_sc_hd__clkinv_1 U14312 ( .A(n20098), .Y(n12949) );
  sky130_fd_sc_hd__clkinv_1 U14313 ( .A(n15357), .Y(n15319) );
  sky130_fd_sc_hd__clkinv_1 U14314 ( .A(n18268), .Y(n18518) );
  sky130_fd_sc_hd__clkinv_1 U14315 ( .A(n16594), .Y(n16597) );
  sky130_fd_sc_hd__clkinv_1 U14316 ( .A(n21723), .Y(n15244) );
  sky130_fd_sc_hd__clkinv_1 U14317 ( .A(n16740), .Y(n14997) );
  sky130_fd_sc_hd__clkinv_1 U14318 ( .A(n14576), .Y(n13028) );
  sky130_fd_sc_hd__clkinv_1 U14319 ( .A(n22374), .Y(n22756) );
  sky130_fd_sc_hd__clkinv_1 U14320 ( .A(n13008), .Y(n13031) );
  sky130_fd_sc_hd__clkinv_1 U14321 ( .A(n13065), .Y(n14578) );
  sky130_fd_sc_hd__clkinv_1 U14322 ( .A(n23356), .Y(n23789) );
  sky130_fd_sc_hd__clkinv_1 U14323 ( .A(n13016), .Y(n14235) );
  sky130_fd_sc_hd__clkinv_1 U14324 ( .A(n14988), .Y(n13598) );
  sky130_fd_sc_hd__clkinv_1 U14325 ( .A(n21222), .Y(n19764) );
  sky130_fd_sc_hd__clkinv_1 U14326 ( .A(n13596), .Y(n13597) );
  sky130_fd_sc_hd__clkinv_1 U14327 ( .A(n25018), .Y(n23479) );
  sky130_fd_sc_hd__clkinv_1 U14328 ( .A(n14120), .Y(n13196) );
  sky130_fd_sc_hd__clkinv_1 U14329 ( .A(n20829), .Y(n20831) );
  sky130_fd_sc_hd__clkinv_1 U14330 ( .A(n21681), .Y(n20100) );
  sky130_fd_sc_hd__clkinv_1 U14331 ( .A(n14184), .Y(n14283) );
  sky130_fd_sc_hd__clkinv_1 U14332 ( .A(n13373), .Y(n13375) );
  sky130_fd_sc_hd__clkinv_1 U14333 ( .A(n15140), .Y(n15142) );
  sky130_fd_sc_hd__clkinv_1 U14334 ( .A(n13195), .Y(n13213) );
  sky130_fd_sc_hd__clkinv_1 U14335 ( .A(n17533), .Y(n15010) );
  sky130_fd_sc_hd__clkinv_1 U14336 ( .A(n14723), .Y(n14309) );
  sky130_fd_sc_hd__clkinv_1 U14337 ( .A(n15009), .Y(n17931) );
  sky130_fd_sc_hd__clkinv_1 U14338 ( .A(n17441), .Y(n17930) );
  sky130_fd_sc_hd__clkinv_1 U14339 ( .A(n20839), .Y(n20840) );
  sky130_fd_sc_hd__clkinv_1 U14340 ( .A(n19565), .Y(n19963) );
  sky130_fd_sc_hd__clkinv_1 U14341 ( .A(n16744), .Y(n14979) );
  sky130_fd_sc_hd__clkinv_1 U14342 ( .A(n19981), .Y(n19843) );
  sky130_fd_sc_hd__clkinv_1 U14343 ( .A(n13017), .Y(n14572) );
  sky130_fd_sc_hd__clkinv_1 U14344 ( .A(n20085), .Y(n20101) );
  sky130_fd_sc_hd__clkinv_1 U14345 ( .A(n18161), .Y(n18183) );
  sky130_fd_sc_hd__clkinv_1 U14346 ( .A(n14943), .Y(n14944) );
  sky130_fd_sc_hd__clkinv_1 U14347 ( .A(n13246), .Y(n13193) );
  sky130_fd_sc_hd__clkinv_1 U14348 ( .A(n25290), .Y(n24393) );
  sky130_fd_sc_hd__clkinv_1 U14349 ( .A(n14348), .Y(n14631) );
  sky130_fd_sc_hd__clkinv_1 U14350 ( .A(n24069), .Y(n20125) );
  sky130_fd_sc_hd__clkinv_1 U14351 ( .A(n16741), .Y(n11225) );
  sky130_fd_sc_hd__clkinv_1 U14352 ( .A(n14102), .Y(n14575) );
  sky130_fd_sc_hd__clkinv_1 U14353 ( .A(n15093), .Y(n15149) );
  sky130_fd_sc_hd__clkinv_1 U14354 ( .A(n24473), .Y(n25270) );
  sky130_fd_sc_hd__clkinv_1 U14355 ( .A(n14310), .Y(n14549) );
  sky130_fd_sc_hd__clkinv_1 U14356 ( .A(n17108), .Y(n16665) );
  sky130_fd_sc_hd__clkinv_1 U14357 ( .A(n24430), .Y(n25279) );
  sky130_fd_sc_hd__clkinv_1 U14358 ( .A(n24432), .Y(n25262) );
  sky130_fd_sc_hd__clkinv_1 U14359 ( .A(n13006), .Y(n13413) );
  sky130_fd_sc_hd__clkinv_1 U14360 ( .A(n24481), .Y(n25269) );
  sky130_fd_sc_hd__clkinv_1 U14361 ( .A(n18155), .Y(n18172) );
  sky130_fd_sc_hd__clkinv_1 U14362 ( .A(n12991), .Y(n11233) );
  sky130_fd_sc_hd__clkinv_1 U14363 ( .A(n14399), .Y(n14413) );
  sky130_fd_sc_hd__clkinv_1 U14364 ( .A(n11356), .Y(n13374) );
  sky130_fd_sc_hd__clkinv_1 U14365 ( .A(n24424), .Y(n25402) );
  sky130_fd_sc_hd__clkinv_1 U14366 ( .A(n23535), .Y(n23433) );
  sky130_fd_sc_hd__clkinv_1 U14367 ( .A(n11348), .Y(n11337) );
  sky130_fd_sc_hd__clkinv_1 U14368 ( .A(n15241), .Y(n16596) );
  sky130_fd_sc_hd__clkinv_1 U14369 ( .A(n24443), .Y(n25265) );
  sky130_fd_sc_hd__clkinv_1 U14370 ( .A(n20249), .Y(n12973) );
  sky130_fd_sc_hd__clkinv_1 U14371 ( .A(n23292), .Y(n25109) );
  sky130_fd_sc_hd__clkinv_1 U14372 ( .A(n23412), .Y(n22856) );
  sky130_fd_sc_hd__clkinv_1 U14373 ( .A(n24392), .Y(n25264) );
  sky130_fd_sc_hd__clkinv_1 U14374 ( .A(n20479), .Y(n20226) );
  sky130_fd_sc_hd__clkinv_1 U14375 ( .A(n23398), .Y(n25001) );
  sky130_fd_sc_hd__clkinv_1 U14376 ( .A(n11471), .Y(n11470) );
  sky130_fd_sc_hd__clkinv_1 U14377 ( .A(n14339), .Y(n14645) );
  sky130_fd_sc_hd__clkinv_1 U14378 ( .A(n14292), .Y(n14294) );
  sky130_fd_sc_hd__clkinv_1 U14379 ( .A(n12280), .Y(n12426) );
  sky130_fd_sc_hd__clkinv_1 U14380 ( .A(n13652), .Y(n13653) );
  sky130_fd_sc_hd__clkinv_1 U14381 ( .A(n15063), .Y(n25245) );
  sky130_fd_sc_hd__clkinv_1 U14382 ( .A(n24418), .Y(n25268) );
  sky130_fd_sc_hd__clkinv_1 U14383 ( .A(n14099), .Y(n13192) );
  sky130_fd_sc_hd__clkinv_1 U14384 ( .A(n24426), .Y(n25267) );
  sky130_fd_sc_hd__clkinv_1 U14385 ( .A(n11338), .Y(n11334) );
  sky130_fd_sc_hd__clkinv_1 U14386 ( .A(n24452), .Y(n24327) );
  sky130_fd_sc_hd__clkinv_1 U14387 ( .A(n14615), .Y(n14244) );
  sky130_fd_sc_hd__clkinv_1 U14388 ( .A(n24434), .Y(n25266) );
  sky130_fd_sc_hd__clkinv_1 U14389 ( .A(n20234), .Y(n12938) );
  sky130_fd_sc_hd__clkinv_1 U14390 ( .A(n14980), .Y(n11339) );
  sky130_fd_sc_hd__clkinv_1 U14391 ( .A(n24422), .Y(n25263) );
  sky130_fd_sc_hd__clkinv_1 U14392 ( .A(n20231), .Y(n20232) );
  sky130_fd_sc_hd__clkinv_1 U14394 ( .A(n25282), .Y(n24395) );
  sky130_fd_sc_hd__clkinv_1 U14395 ( .A(n19172), .Y(n21017) );
  sky130_fd_sc_hd__clkinv_1 U14396 ( .A(n12904), .Y(n11438) );
  sky130_fd_sc_hd__clkinv_1 U14397 ( .A(n14201), .Y(n12987) );
  sky130_fd_sc_hd__clkinv_1 U14398 ( .A(n11542), .Y(n11534) );
  sky130_fd_sc_hd__clkinv_1 U14399 ( .A(n23236), .Y(n20485) );
  sky130_fd_sc_hd__clkinv_1 U14400 ( .A(n13018), .Y(n13012) );
  sky130_fd_sc_hd__clkinv_1 U14401 ( .A(n25284), .Y(n24402) );
  sky130_fd_sc_hd__clkinv_1 U14402 ( .A(n14841), .Y(n14884) );
  sky130_fd_sc_hd__clkinv_1 U14403 ( .A(n15390), .Y(n15275) );
  sky130_fd_sc_hd__clkinv_1 U14404 ( .A(n15394), .Y(n15274) );
  sky130_fd_sc_hd__clkinv_1 U14405 ( .A(n13005), .Y(n14295) );
  sky130_fd_sc_hd__clkinv_1 U14406 ( .A(n15016), .Y(n15019) );
  sky130_fd_sc_hd__clkinv_1 U14407 ( .A(n20155), .Y(n20142) );
  sky130_fd_sc_hd__clkinv_1 U14408 ( .A(n20274), .Y(n20279) );
  sky130_fd_sc_hd__clkinv_1 U14409 ( .A(n25291), .Y(n24397) );
  sky130_fd_sc_hd__clkinv_1 U14410 ( .A(n17532), .Y(n15008) );
  sky130_fd_sc_hd__clkinv_1 U14411 ( .A(n14989), .Y(n14473) );
  sky130_fd_sc_hd__clkinv_1 U14412 ( .A(n14990), .Y(n17731) );
  sky130_fd_sc_hd__clkinv_1 U14413 ( .A(n25289), .Y(n24389) );
  sky130_fd_sc_hd__clkinv_1 U14414 ( .A(n13093), .Y(n11439) );
  sky130_fd_sc_hd__clkinv_1 U14415 ( .A(n14111), .Y(n13198) );
  sky130_fd_sc_hd__clkinv_1 U14416 ( .A(n13015), .Y(n13027) );
  sky130_fd_sc_hd__clkinv_1 U14417 ( .A(n15417), .Y(n15419) );
  sky130_fd_sc_hd__clkinv_1 U14418 ( .A(n22803), .Y(n19325) );
  sky130_fd_sc_hd__clkinv_1 U14419 ( .A(n17177), .Y(n17196) );
  sky130_fd_sc_hd__clkinv_1 U14420 ( .A(n15414), .Y(n15415) );
  sky130_fd_sc_hd__clkinv_1 U14421 ( .A(n25202), .Y(n18244) );
  sky130_fd_sc_hd__clkinv_1 U14422 ( .A(n11213), .Y(n14096) );
  sky130_fd_sc_hd__clkinv_1 U14423 ( .A(n14978), .Y(n14982) );
  sky130_fd_sc_hd__clkinv_1 U14424 ( .A(n24420), .Y(n25275) );
  sky130_fd_sc_hd__clkinv_1 U14425 ( .A(n14108), .Y(n14986) );
  sky130_fd_sc_hd__clkinv_1 U14426 ( .A(n11535), .Y(n11531) );
  sky130_fd_sc_hd__clkinv_1 U14427 ( .A(n20836), .Y(n16663) );
  sky130_fd_sc_hd__clkinv_1 U14428 ( .A(n24399), .Y(n25395) );
  sky130_fd_sc_hd__clkinv_1 U14429 ( .A(n11537), .Y(n11533) );
  sky130_fd_sc_hd__clkinv_1 U14430 ( .A(n14977), .Y(n14981) );
  sky130_fd_sc_hd__clkinv_1 U14431 ( .A(n25292), .Y(n24390) );
  sky130_fd_sc_hd__clkinv_1 U14432 ( .A(n25283), .Y(n24387) );
  sky130_fd_sc_hd__clkinv_1 U14433 ( .A(n14866), .Y(n14882) );
  sky130_fd_sc_hd__clkinv_1 U14434 ( .A(n14236), .Y(n14604) );
  sky130_fd_sc_hd__clkinv_1 U14435 ( .A(n14101), .Y(n14472) );
  sky130_fd_sc_hd__clkinv_1 U14436 ( .A(n13464), .Y(n13496) );
  sky130_fd_sc_hd__clkinv_1 U14437 ( .A(n11566), .Y(n11567) );
  sky130_fd_sc_hd__clkinv_1 U14438 ( .A(n15387), .Y(n15389) );
  sky130_fd_sc_hd__clkinv_1 U14439 ( .A(n15370), .Y(n15246) );
  sky130_fd_sc_hd__clkinv_1 U14440 ( .A(n14639), .Y(n14613) );
  sky130_fd_sc_hd__clkinv_1 U14441 ( .A(n18189), .Y(n18047) );
  sky130_fd_sc_hd__clkinv_1 U14442 ( .A(n15284), .Y(n15393) );
  sky130_fd_sc_hd__clkinv_1 U14443 ( .A(n15391), .Y(n15392) );
  sky130_fd_sc_hd__clkinv_1 U14444 ( .A(n15361), .Y(n15363) );
  sky130_fd_sc_hd__clkinv_1 U14445 ( .A(n14352), .Y(n14619) );
  sky130_fd_sc_hd__clkinv_1 U14446 ( .A(n14815), .Y(n14888) );
  sky130_fd_sc_hd__clkinv_1 U14447 ( .A(n15297), .Y(n15299) );
  sky130_fd_sc_hd__clkinv_1 U14448 ( .A(n13449), .Y(n14098) );
  sky130_fd_sc_hd__clkinv_1 U14449 ( .A(n14313), .Y(n12995) );
  sky130_fd_sc_hd__clkinv_1 U14450 ( .A(n12916), .Y(n11557) );
  sky130_fd_sc_hd__clkinv_1 U14451 ( .A(n14605), .Y(n12989) );
  sky130_fd_sc_hd__clkinv_1 U14452 ( .A(n15435), .Y(n15340) );
  sky130_fd_sc_hd__clkinv_1 U14453 ( .A(n20097), .Y(n12953) );
  sky130_fd_sc_hd__clkinv_1 U14454 ( .A(n25005), .Y(n23451) );
  sky130_fd_sc_hd__clkinv_1 U14455 ( .A(n11336), .Y(n14095) );
  sky130_fd_sc_hd__clkinv_1 U14456 ( .A(n15430), .Y(n15432) );
  sky130_fd_sc_hd__inv_1 U14457 ( .A(n20245), .Y(n20268) );
  sky130_fd_sc_hd__clkinv_1 U14458 ( .A(n15411), .Y(n15413) );
  sky130_fd_sc_hd__clkinv_1 U14459 ( .A(n15310), .Y(n15283) );
  sky130_fd_sc_hd__clkinv_1 U14460 ( .A(n15309), .Y(n15333) );
  sky130_fd_sc_hd__clkinv_1 U14461 ( .A(n15332), .Y(n15287) );
  sky130_fd_sc_hd__clkinv_1 U14462 ( .A(n14562), .Y(n14563) );
  sky130_fd_sc_hd__clkinv_1 U14463 ( .A(n17368), .Y(n17369) );
  sky130_fd_sc_hd__clkinv_1 U14464 ( .A(n12019), .Y(n12942) );
  sky130_fd_sc_hd__clkinv_1 U14465 ( .A(n15214), .Y(n15220) );
  sky130_fd_sc_hd__clkinv_1 U14466 ( .A(n11555), .Y(n12020) );
  sky130_fd_sc_hd__clkinv_1 U14467 ( .A(n14308), .Y(n14617) );
  sky130_fd_sc_hd__clkinv_1 U14468 ( .A(n21905), .Y(n21903) );
  sky130_fd_sc_hd__clkinv_1 U14469 ( .A(n21328), .Y(n22336) );
  sky130_fd_sc_hd__clkinv_1 U14470 ( .A(n16658), .Y(n16657) );
  sky130_fd_sc_hd__clkinv_1 U14471 ( .A(n20198), .Y(n20205) );
  sky130_fd_sc_hd__clkinv_1 U14472 ( .A(n15420), .Y(n15380) );
  sky130_fd_sc_hd__clkinv_1 U14473 ( .A(n24469), .Y(n24379) );
  sky130_fd_sc_hd__clkinv_1 U14474 ( .A(n22509), .Y(n17107) );
  sky130_fd_sc_hd__clkinv_1 U14475 ( .A(n15348), .Y(n15350) );
  sky130_fd_sc_hd__clkinv_1 U14476 ( .A(n15344), .Y(n15345) );
  sky130_fd_sc_hd__clkinv_1 U14477 ( .A(n15268), .Y(n15346) );
  sky130_fd_sc_hd__clkinv_1 U14478 ( .A(n21678), .Y(n12950) );
  sky130_fd_sc_hd__clkinv_1 U14479 ( .A(n21724), .Y(n16591) );
  sky130_fd_sc_hd__clkinv_1 U14480 ( .A(n21654), .Y(n21679) );
  sky130_fd_sc_hd__clkinv_1 U14481 ( .A(n18147), .Y(n18178) );
  sky130_fd_sc_hd__clkinv_1 U14482 ( .A(n14972), .Y(n14951) );
  sky130_fd_sc_hd__clkinv_1 U14483 ( .A(j202_soc_core_j22_cpu_rf_gpr[27]), .Y(
        n13823) );
  sky130_fd_sc_hd__clkinv_1 U14484 ( .A(j202_soc_core_j22_cpu_ml_macl[3]), .Y(
        n18888) );
  sky130_fd_sc_hd__clkinv_1 U14485 ( .A(j202_soc_core_intc_core_00_rg_ipr[74]), 
        .Y(n24606) );
  sky130_fd_sc_hd__clkinv_1 U14486 ( .A(j202_soc_core_j22_cpu_ml_macl[19]), 
        .Y(n20037) );
  sky130_fd_sc_hd__clkinv_1 U14487 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .Y(n14094) );
  sky130_fd_sc_hd__clkinv_1 U14488 ( .A(j202_soc_core_j22_cpu_ml_mach[0]), .Y(
        n15704) );
  sky130_fd_sc_hd__clkinv_1 U14489 ( .A(j202_soc_core_j22_cpu_rf_gpr[5]), .Y(
        n12259) );
  sky130_fd_sc_hd__clkinv_1 U14490 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[3]), 
        .Y(n16664) );
  sky130_fd_sc_hd__clkinv_1 U14491 ( .A(j202_soc_core_j22_cpu_ml_mach[5]), .Y(
        n19136) );
  sky130_fd_sc_hd__clkinv_1 U14492 ( .A(j202_soc_core_intr_vec__3_), .Y(n22905) );
  sky130_fd_sc_hd__clkinv_1 U14493 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .Y(n14985) );
  sky130_fd_sc_hd__clkinv_1 U14494 ( .A(j202_soc_core_j22_cpu_regop_imm__5_), 
        .Y(n12168) );
  sky130_fd_sc_hd__clkinv_1 U14495 ( .A(j202_soc_core_j22_cpu_ml_mach[21]), 
        .Y(n19367) );
  sky130_fd_sc_hd__clkinv_1 U14496 ( .A(j202_soc_core_j22_cpu_rf_gpr[16]), .Y(
        n11734) );
  sky130_fd_sc_hd__clkinv_1 U14497 ( .A(j202_soc_core_j22_cpu_ml_macl[23]), 
        .Y(n15875) );
  sky130_fd_sc_hd__clkinv_1 U14498 ( .A(j202_soc_core_j22_cpu_rf_gpr[26]), .Y(
        n13956) );
  sky130_fd_sc_hd__clkinv_1 U14499 ( .A(j202_soc_core_j22_cpu_rf_pr[4]), .Y(
        n17063) );
  sky130_fd_sc_hd__clkinv_1 U14500 ( .A(j202_soc_core_j22_cpu_ml_macl[7]), .Y(
        n16636) );
  sky130_fd_sc_hd__clkinv_1 U14501 ( .A(j202_soc_core_j22_cpu_ml_bufa[12]), 
        .Y(n22098) );
  sky130_fd_sc_hd__clkinv_1 U14502 ( .A(j202_soc_core_j22_cpu_pc[15]), .Y(
        n12675) );
  sky130_fd_sc_hd__clkinv_1 U14503 ( .A(j202_soc_core_intc_core_00_rg_ipr[34]), 
        .Y(n24353) );
  sky130_fd_sc_hd__clkinv_1 U14504 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__0_), 
        .Y(n17064) );
  sky130_fd_sc_hd__clkinv_1 U14505 ( .A(j202_soc_core_j22_cpu_ml_bufa[14]), 
        .Y(n21900) );
  sky130_fd_sc_hd__clkinv_1 U14506 ( .A(j202_soc_core_j22_cpu_rf_pr[15]), .Y(
        n15218) );
  sky130_fd_sc_hd__clkinv_1 U14507 ( .A(j202_soc_core_j22_cpu_rf_gbr[4]), .Y(
        n17065) );
  sky130_fd_sc_hd__clkinv_1 U14508 ( .A(j202_soc_core_intc_core_00_rg_ipr[3]), 
        .Y(n24530) );
  sky130_fd_sc_hd__clkinv_1 U14509 ( .A(j202_soc_core_intc_core_00_rg_ipr[72]), 
        .Y(n24589) );
  sky130_fd_sc_hd__clkinv_1 U14510 ( .A(j202_soc_core_j22_cpu_ml_mach[23]), 
        .Y(n19327) );
  sky130_fd_sc_hd__clkinv_1 U14511 ( .A(j202_soc_core_j22_cpu_ml_macl[0]), .Y(
        n19235) );
  sky130_fd_sc_hd__clkinv_1 U14512 ( .A(j202_soc_core_intc_core_00_rg_ipr[71]), 
        .Y(n24330) );
  sky130_fd_sc_hd__clkinv_1 U14513 ( .A(j202_soc_core_intc_core_00_rg_ipr[18]), 
        .Y(n24385) );
  sky130_fd_sc_hd__clkinv_1 U14514 ( .A(j202_soc_core_intc_core_00_rg_ipr[23]), 
        .Y(n24391) );
  sky130_fd_sc_hd__clkinv_1 U14515 ( .A(j202_soc_core_intc_core_00_rg_ipr[67]), 
        .Y(n24531) );
  sky130_fd_sc_hd__clkinv_1 U14516 ( .A(j202_soc_core_intc_core_00_bs_addr[2]), 
        .Y(n24293) );
  sky130_fd_sc_hd__clkinv_1 U14517 ( .A(j202_soc_core_intc_core_00_rg_ipr[17]), 
        .Y(n24666) );
  sky130_fd_sc_hd__clkinv_1 U14518 ( .A(j202_soc_core_j22_cpu_ml_bufa[23]), 
        .Y(n19377) );
  sky130_fd_sc_hd__clkinv_1 U14519 ( .A(j202_soc_core_j22_cpu_ml_macl[21]), 
        .Y(n15925) );
  sky130_fd_sc_hd__clkinv_1 U14520 ( .A(j202_soc_core_intc_core_00_rg_ipr[21]), 
        .Y(n24388) );
  sky130_fd_sc_hd__clkinv_1 U14521 ( .A(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .Y(n15235) );
  sky130_fd_sc_hd__clkinv_1 U14522 ( .A(j202_soc_core_intc_core_00_rg_ipr[70]), 
        .Y(n24562) );
  sky130_fd_sc_hd__clkinv_1 U14523 ( .A(j202_soc_core_intc_core_00_rg_ipr[19]), 
        .Y(n24680) );
  sky130_fd_sc_hd__clkinv_1 U14524 ( .A(j202_soc_core_j22_cpu_rf_gpr[13]), .Y(
        n12642) );
  sky130_fd_sc_hd__clkinv_1 U14525 ( .A(j202_soc_core_j22_cpu_rf_gbr[5]), .Y(
        n19181) );
  sky130_fd_sc_hd__clkinv_1 U14526 ( .A(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .Y(n15236) );
  sky130_fd_sc_hd__clkinv_1 U14527 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__1_), 
        .Y(n19180) );
  sky130_fd_sc_hd__clkinv_1 U14528 ( .A(j202_soc_core_intc_core_00_rg_ipr[22]), 
        .Y(n24706) );
  sky130_fd_sc_hd__clkinv_1 U14529 ( .A(j202_soc_core_intc_core_00_rg_ipr[77]), 
        .Y(n24633) );
  sky130_fd_sc_hd__clkinv_1 U14530 ( .A(j202_soc_core_j22_cpu_rf_pr[5]), .Y(
        n19179) );
  sky130_fd_sc_hd__clkinv_1 U14531 ( .A(j202_soc_core_j22_cpu_ml_macl[5]), .Y(
        n19144) );
  sky130_fd_sc_hd__clkinv_1 U14532 ( .A(j202_soc_core_intc_core_00_rg_ipr[73]), 
        .Y(n24597) );
  sky130_fd_sc_hd__clkinv_1 U14533 ( .A(j202_soc_core_j22_cpu_rf_gpr[15]), .Y(
        n12676) );
  sky130_fd_sc_hd__clkinv_1 U14534 ( .A(j202_soc_core_j22_cpu_ml_mach[20]), 
        .Y(n19427) );
  sky130_fd_sc_hd__clkinv_1 U14535 ( .A(j202_soc_core_j22_cpu_ml_bufa[5]), .Y(
        n22031) );
  sky130_fd_sc_hd__clkinv_1 U14536 ( .A(j202_soc_core_intc_core_00_rg_ipr[69]), 
        .Y(n24329) );
  sky130_fd_sc_hd__clkinv_1 U14537 ( .A(j202_soc_core_intc_core_00_rg_ipr[14]), 
        .Y(n24641) );
  sky130_fd_sc_hd__clkinv_1 U14538 ( .A(j202_soc_core_j22_cpu_rf_gpr[4]), .Y(
        n12343) );
  sky130_fd_sc_hd__clkinv_1 U14539 ( .A(j202_soc_core_intc_core_00_rg_ipr[13]), 
        .Y(n24632) );
  sky130_fd_sc_hd__clkinv_1 U14540 ( .A(j202_soc_core_j22_cpu_ml_mach[19]), 
        .Y(n19363) );
  sky130_fd_sc_hd__clkinv_1 U14541 ( .A(j202_soc_core_intc_core_00_rg_ipr[12]), 
        .Y(n24623) );
  sky130_fd_sc_hd__clkinv_1 U14542 ( .A(j202_soc_core_intc_core_00_rg_ipr[65]), 
        .Y(n24511) );
  sky130_fd_sc_hd__clkinv_1 U14543 ( .A(j202_soc_core_j22_cpu_ml_mach[6]), .Y(
        n15617) );
  sky130_fd_sc_hd__clkinv_1 U14544 ( .A(j202_soc_core_intr_vec__2_), .Y(n22903) );
  sky130_fd_sc_hd__clkinv_1 U14545 ( .A(j202_soc_core_intc_core_00_rg_ipr[10]), 
        .Y(n24609) );
  sky130_fd_sc_hd__clkinv_1 U14546 ( .A(j202_soc_core_j22_cpu_regop_imm__4_), 
        .Y(n12223) );
  sky130_fd_sc_hd__clkinv_1 U14547 ( .A(j202_soc_core_j22_cpu_ml_macl[16]), 
        .Y(n15942) );
  sky130_fd_sc_hd__clkinv_1 U14548 ( .A(j202_soc_core_intc_core_00_rg_ipr[15]), 
        .Y(n24653) );
  sky130_fd_sc_hd__clkinv_1 U14549 ( .A(j202_soc_core_intc_core_00_rg_ipr[31]), 
        .Y(n24407) );
  sky130_fd_sc_hd__clkinv_1 U14550 ( .A(j202_soc_core_intc_core_00_rg_ipr[20]), 
        .Y(n24386) );
  sky130_fd_sc_hd__clkinv_1 U14551 ( .A(j202_soc_core_intc_core_00_rg_ipr[9]), 
        .Y(n24600) );
  sky130_fd_sc_hd__clkinv_1 U14552 ( .A(j202_soc_core_j22_cpu_rf_gpr[31]), .Y(
        n13696) );
  sky130_fd_sc_hd__clkinv_1 U14553 ( .A(j202_soc_core_j22_cpu_ml_mach[15]), 
        .Y(n16582) );
  sky130_fd_sc_hd__clkinv_1 U14554 ( .A(j202_soc_core_intc_core_00_rg_ipr[78]), 
        .Y(n24642) );
  sky130_fd_sc_hd__clkinv_1 U14555 ( .A(j202_soc_core_intc_core_00_rg_ipr[1]), 
        .Y(n24510) );
  sky130_fd_sc_hd__clkinv_1 U14556 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[4]), .Y(n25174) );
  sky130_fd_sc_hd__clkinv_1 U14557 ( .A(j202_soc_core_intc_core_00_rg_ipr[28]), 
        .Y(n24747) );
  sky130_fd_sc_hd__clkinv_1 U14558 ( .A(j202_soc_core_j22_cpu_ml_macl[15]), 
        .Y(n16608) );
  sky130_fd_sc_hd__clkinv_1 U14559 ( .A(j202_soc_core_intc_core_00_rg_ipr[5]), 
        .Y(n24381) );
  sky130_fd_sc_hd__clkinv_1 U14560 ( .A(j202_soc_core_intc_core_00_rg_ipr[75]), 
        .Y(n24616) );
  sky130_fd_sc_hd__clkinv_1 U14561 ( .A(j202_soc_core_intc_core_00_rg_ipr[6]), 
        .Y(n24561) );
  sky130_fd_sc_hd__clkinv_1 U14562 ( .A(j202_soc_core_intc_core_00_rg_ipr[30]), 
        .Y(n24403) );
  sky130_fd_sc_hd__clkinv_1 U14563 ( .A(j202_soc_core_j22_cpu_ml_macl[22]), 
        .Y(n19533) );
  sky130_fd_sc_hd__clkinv_1 U14564 ( .A(j202_soc_core_intc_core_00_rg_ipr[7]), 
        .Y(n24382) );
  sky130_fd_sc_hd__clkinv_1 U14565 ( .A(j202_soc_core_intc_core_00_rg_ipr[26]), 
        .Y(n24396) );
  sky130_fd_sc_hd__clkinv_1 U14566 ( .A(j202_soc_core_j22_cpu_ml_mach[24]), 
        .Y(n19549) );
  sky130_fd_sc_hd__clkinv_1 U14567 ( .A(j202_soc_core_intc_core_00_rg_ipr[29]), 
        .Y(n24401) );
  sky130_fd_sc_hd__clkinv_1 U14568 ( .A(j202_soc_core_j22_cpu_ml_bufa[13]), 
        .Y(n22232) );
  sky130_fd_sc_hd__clkinv_1 U14569 ( .A(j202_soc_core_j22_cpu_ml_macl[6]), .Y(
        n19017) );
  sky130_fd_sc_hd__clkinv_1 U14570 ( .A(j202_soc_core_intc_core_00_rg_ipr[0]), 
        .Y(n24500) );
  sky130_fd_sc_hd__clkinv_1 U14571 ( .A(j202_soc_core_intc_core_00_rg_ipr[8]), 
        .Y(n24588) );
  sky130_fd_sc_hd__clkinv_1 U14572 ( .A(j202_soc_core_intc_core_00_rg_ipr[2]), 
        .Y(n24520) );
  sky130_fd_sc_hd__clkinv_1 U14573 ( .A(j202_soc_core_intc_core_00_rg_ipr[64]), 
        .Y(n24501) );
  sky130_fd_sc_hd__clkinv_1 U14574 ( .A(j202_soc_core_j22_cpu_regop_imm__3_), 
        .Y(n12279) );
  sky130_fd_sc_hd__clkinv_1 U14575 ( .A(j202_soc_core_intr_vec__1_), .Y(n22899) );
  sky130_fd_sc_hd__clkinv_1 U14576 ( .A(j202_soc_core_j22_cpu_ml_mach[18]), 
        .Y(n19331) );
  sky130_fd_sc_hd__clkinv_1 U14577 ( .A(j202_soc_core_j22_cpu_rf_gbr[6]), .Y(
        n19053) );
  sky130_fd_sc_hd__clkinv_1 U14578 ( .A(j202_soc_core_j22_cpu_ml_mach[22]), 
        .Y(n19330) );
  sky130_fd_sc_hd__clkinv_1 U14579 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__2_), 
        .Y(n19052) );
  sky130_fd_sc_hd__clkinv_1 U14580 ( .A(j202_soc_core_j22_cpu_rf_pr[6]), .Y(
        n19051) );
  sky130_fd_sc_hd__clkinv_1 U14581 ( .A(j202_soc_core_j22_cpu_rf_tmp[12]), .Y(
        n17057) );
  sky130_fd_sc_hd__clkinv_1 U14582 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__1_), 
        .Y(n20318) );
  sky130_fd_sc_hd__clkinv_1 U14583 ( .A(j202_soc_core_j22_cpu_rf_gpr[21]), .Y(
        n11497) );
  sky130_fd_sc_hd__clkinv_1 U14584 ( .A(j202_soc_core_j22_cpu_pc[12]), .Y(
        n17053) );
  sky130_fd_sc_hd__clkinv_1 U14585 ( .A(j202_soc_core_j22_cpu_rf_pr[12]), .Y(
        n17052) );
  sky130_fd_sc_hd__clkinv_1 U14586 ( .A(j202_soc_core_j22_cpu_rf_gbr[12]), .Y(
        n17056) );
  sky130_fd_sc_hd__clkinv_1 U14587 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__3_), 
        .Y(n20263) );
  sky130_fd_sc_hd__clkinv_1 U14588 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[15]), .Y(n24987) );
  sky130_fd_sc_hd__clkinv_1 U14589 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]), .Y(n24944) );
  sky130_fd_sc_hd__clkinv_1 U14590 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__2_), 
        .Y(n20255) );
  sky130_fd_sc_hd__clkinv_1 U14591 ( .A(j202_soc_core_j22_cpu_ml_mach[16]), 
        .Y(n19339) );
  sky130_fd_sc_hd__clkinv_1 U14592 ( .A(j202_soc_core_j22_cpu_ml_macl[13]), 
        .Y(n19112) );
  sky130_fd_sc_hd__clkinv_1 U14593 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[10]), .Y(n24922) );
  sky130_fd_sc_hd__clkinv_1 U14594 ( .A(j202_soc_core_intc_core_00_rg_ipr[59]), 
        .Y(n24372) );
  sky130_fd_sc_hd__clkinv_1 U14595 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[11]), .Y(n24925) );
  sky130_fd_sc_hd__clkinv_1 U14596 ( .A(j202_soc_core_intc_core_00_rg_ipr[50]), 
        .Y(n24365) );
  sky130_fd_sc_hd__clkinv_1 U14597 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[6]), .Y(n24909) );
  sky130_fd_sc_hd__clkinv_1 U14598 ( .A(j202_soc_core_j22_cpu_ml_macl[29]), 
        .Y(n15796) );
  sky130_fd_sc_hd__clkinv_1 U14599 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[4]), .Y(n24905) );
  sky130_fd_sc_hd__clkinv_1 U14600 ( .A(j202_soc_core_intc_core_00_rg_ipr[56]), 
        .Y(n24719) );
  sky130_fd_sc_hd__clkinv_1 U14601 ( .A(j202_soc_core_j22_cpu_ml_mach[27]), 
        .Y(n19592) );
  sky130_fd_sc_hd__clkinv_1 U14602 ( .A(j202_soc_core_intc_core_00_bs_addr[7]), 
        .Y(n24573) );
  sky130_fd_sc_hd__clkinv_1 U14603 ( .A(j202_soc_core_intc_core_00_rg_ipr[57]), 
        .Y(n24370) );
  sky130_fd_sc_hd__clkinv_1 U14604 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[8]), .Y(n24940) );
  sky130_fd_sc_hd__clkinv_1 U14605 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .Y(n23567) );
  sky130_fd_sc_hd__clkinv_1 U14606 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]), .Y(n25019) );
  sky130_fd_sc_hd__clkinv_1 U14607 ( .A(j202_soc_core_intc_core_00_rg_ipr[63]), 
        .Y(n24377) );
  sky130_fd_sc_hd__clkinv_1 U14608 ( .A(j202_soc_core_qspi_wb_addr[23]), .Y(
        n25088) );
  sky130_fd_sc_hd__clkinv_1 U14609 ( .A(j202_soc_core_intc_core_00_rg_ipr[58]), 
        .Y(n24371) );
  sky130_fd_sc_hd__clkinv_1 U14610 ( .A(j202_soc_core_j22_cpu_rf_gpr[8]), .Y(
        n12487) );
  sky130_fd_sc_hd__clkinv_1 U14611 ( .A(j202_soc_core_j22_cpu_rf_gpr[22]), .Y(
        n11469) );
  sky130_fd_sc_hd__clkinv_1 U14612 ( .A(j202_soc_core_pwrite[2]), .Y(n24067)
         );
  sky130_fd_sc_hd__clkinv_1 U14613 ( .A(j202_soc_core_ahb2apb_02_state[2]), 
        .Y(n21218) );
  sky130_fd_sc_hd__clkinv_1 U14614 ( .A(j202_soc_core_intc_core_00_rg_ipr[60]), 
        .Y(n24743) );
  sky130_fd_sc_hd__clkinv_1 U14615 ( .A(j202_soc_core_j22_cpu_rf_gpr[11]), .Y(
        n12406) );
  sky130_fd_sc_hd__clkinv_1 U14616 ( .A(j202_soc_core_j22_cpu_rf_pr[9]), .Y(
        n19972) );
  sky130_fd_sc_hd__clkinv_1 U14617 ( .A(j202_soc_core_j22_cpu_ml_mach[29]), 
        .Y(n19586) );
  sky130_fd_sc_hd__clkinv_1 U14618 ( .A(j202_soc_core_j22_cpu_ml_mach[8]), .Y(
        n19303) );
  sky130_fd_sc_hd__clkinv_1 U14619 ( .A(j202_soc_core_j22_cpu_rf_gpr[19]), .Y(
        n11580) );
  sky130_fd_sc_hd__clkinv_1 U14620 ( .A(j202_soc_core_j22_cpu_regop_imm__10_), 
        .Y(n12362) );
  sky130_fd_sc_hd__clkinv_1 U14621 ( .A(j202_soc_core_j22_cpu_rf_gpr[10]), .Y(
        n12570) );
  sky130_fd_sc_hd__clkinv_1 U14622 ( .A(j202_soc_core_j22_cpu_ml_macl[11]), 
        .Y(n18869) );
  sky130_fd_sc_hd__clkinv_1 U14623 ( .A(j202_soc_core_j22_cpu_rf_gbr[11]), .Y(
        n18930) );
  sky130_fd_sc_hd__clkinv_1 U14624 ( .A(j202_soc_core_j22_cpu_rf_pr[11]), .Y(
        n18926) );
  sky130_fd_sc_hd__clkinv_1 U14625 ( .A(j202_soc_core_j22_cpu_pc[11]), .Y(
        n18927) );
  sky130_fd_sc_hd__clkinv_1 U14626 ( .A(j202_soc_core_j22_cpu_rf_tmp[11]), .Y(
        n18931) );
  sky130_fd_sc_hd__clkinv_1 U14627 ( .A(j202_soc_core_intc_core_00_bs_addr[8]), 
        .Y(n24448) );
  sky130_fd_sc_hd__clkinv_1 U14628 ( .A(j202_soc_core_j22_cpu_ml_macl[27]), 
        .Y(n15853) );
  sky130_fd_sc_hd__clkinv_1 U14629 ( .A(j202_soc_core_j22_cpu_regop_We__3_), 
        .Y(n20237) );
  sky130_fd_sc_hd__clkinv_1 U14630 ( .A(j202_soc_core_j22_cpu_ml_macl[30]), 
        .Y(n15709) );
  sky130_fd_sc_hd__clkinv_1 U14631 ( .A(j202_soc_core_j22_cpu_ml_macl[14]), 
        .Y(n18992) );
  sky130_fd_sc_hd__clkinv_1 U14632 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__2_), 
        .Y(n20230) );
  sky130_fd_sc_hd__clkinv_1 U14633 ( .A(j202_soc_core_j22_cpu_regop_imm__9_), 
        .Y(n12538) );
  sky130_fd_sc_hd__clkinv_1 U14634 ( .A(j202_soc_core_j22_cpu_ml_macl[12]), 
        .Y(n17048) );
  sky130_fd_sc_hd__clkinv_1 U14635 ( .A(j202_soc_core_j22_cpu_ml_mach[3]), .Y(
        n15602) );
  sky130_fd_sc_hd__clkinv_1 U14636 ( .A(j202_soc_core_j22_cpu_ml_mach[9]), .Y(
        n20006) );
  sky130_fd_sc_hd__clkinv_1 U14637 ( .A(j202_soc_core_j22_cpu_ml_mach[28]), 
        .Y(n19588) );
  sky130_fd_sc_hd__clkinv_1 U14638 ( .A(j202_soc_core_j22_cpu_rf_gpr[9]), .Y(
        n19984) );
  sky130_fd_sc_hd__clkinv_1 U14639 ( .A(j202_soc_core_j22_cpu_rf_gpr[20]), .Y(
        n11608) );
  sky130_fd_sc_hd__clkinv_1 U14640 ( .A(j202_soc_core_j22_cpu_rf_gpr[30]), .Y(
        n13671) );
  sky130_fd_sc_hd__clkinv_1 U14641 ( .A(j202_soc_core_j22_cpu_rf_gpr[18]), .Y(
        n11661) );
  sky130_fd_sc_hd__clkinv_1 U14642 ( .A(j202_soc_core_j22_cpu_macop_MAC_[3]), 
        .Y(n21669) );
  sky130_fd_sc_hd__clkinv_1 U14643 ( .A(j202_soc_core_wbqspiflash_00_spi_valid), .Y(n23363) );
  sky130_fd_sc_hd__clkinv_1 U14644 ( .A(j202_soc_core_j22_cpu_rf_gbr[10]), .Y(
        n16880) );
  sky130_fd_sc_hd__clkinv_1 U14645 ( .A(j202_soc_core_j22_cpu_ml_macl[10]), 
        .Y(n16808) );
  sky130_fd_sc_hd__clkinv_1 U14646 ( .A(j202_soc_core_j22_cpu_rf_pr[10]), .Y(
        n16876) );
  sky130_fd_sc_hd__clkinv_1 U14647 ( .A(j202_soc_core_j22_cpu_ml_macl[28]), 
        .Y(n15804) );
  sky130_fd_sc_hd__clkinv_1 U14648 ( .A(j202_soc_core_j22_cpu_ml_mach[17]), 
        .Y(n19328) );
  sky130_fd_sc_hd__clkinv_1 U14649 ( .A(j202_soc_core_j22_cpu_pc[10]), .Y(
        n16877) );
  sky130_fd_sc_hd__clkinv_1 U14650 ( .A(j202_soc_core_j22_cpu_ml_macl[26]), 
        .Y(n15841) );
  sky130_fd_sc_hd__clkinv_1 U14651 ( .A(j202_soc_core_j22_cpu_rf_tmp[10]), .Y(
        n16881) );
  sky130_fd_sc_hd__clkinv_1 U14652 ( .A(j202_soc_core_ahb2apb_02_state[0]), 
        .Y(n20123) );
  sky130_fd_sc_hd__clkinv_1 U14653 ( .A(j202_soc_core_j22_cpu_rf_pr[13]), .Y(
        n19117) );
  sky130_fd_sc_hd__clkinv_1 U14654 ( .A(j202_soc_core_j22_cpu_pc[13]), .Y(
        n19121) );
  sky130_fd_sc_hd__clkinv_1 U14655 ( .A(j202_soc_core_j22_cpu_rfuo_sr__q_), 
        .Y(n19201) );
  sky130_fd_sc_hd__clkinv_1 U14656 ( .A(j202_soc_core_intc_core_00_rg_ipr[41]), 
        .Y(n24359) );
  sky130_fd_sc_hd__clkinv_1 U14657 ( .A(j202_soc_core_j22_cpu_rf_gbr[8]), .Y(
        n19202) );
  sky130_fd_sc_hd__clkinv_1 U14658 ( .A(j202_soc_core_j22_cpu_rf_gbr[13]), .Y(
        n19116) );
  sky130_fd_sc_hd__clkinv_1 U14659 ( .A(j202_soc_core_intc_core_00_rg_ipr[42]), 
        .Y(n24360) );
  sky130_fd_sc_hd__clkinv_1 U14660 ( .A(j202_soc_core_j22_cpu_ml_mach[25]), 
        .Y(n19555) );
  sky130_fd_sc_hd__clkinv_1 U14661 ( .A(j202_soc_core_j22_cpu_rf_gpr[24]), .Y(
        n12856) );
  sky130_fd_sc_hd__clkinv_1 U14662 ( .A(j202_soc_core_intc_core_00_rg_ipr[43]), 
        .Y(n24615) );
  sky130_fd_sc_hd__clkinv_1 U14663 ( .A(j202_soc_core_intc_core_00_rg_ipr[40]), 
        .Y(n24358) );
  sky130_fd_sc_hd__clkinv_1 U14664 ( .A(j202_soc_core_pwrite[1]), .Y(n24447)
         );
  sky130_fd_sc_hd__clkinv_1 U14665 ( .A(j202_soc_core_j22_cpu_rf_gbr[29]), .Y(
        n14078) );
  sky130_fd_sc_hd__clkinv_1 U14666 ( .A(j202_soc_core_j22_cpu_rf_pr[29]), .Y(
        n14080) );
  sky130_fd_sc_hd__clkinv_1 U14667 ( .A(j202_soc_core_j22_cpu_pc[29]), .Y(
        n14074) );
  sky130_fd_sc_hd__clkinv_1 U14668 ( .A(j202_soc_core_j22_cpu_rf_gpr[29]), .Y(
        n14076) );
  sky130_fd_sc_hd__clkinv_1 U14669 ( .A(j202_soc_core_j22_cpu_rf_tmp[29]), .Y(
        n14070) );
  sky130_fd_sc_hd__clkinv_1 U14670 ( .A(j202_soc_core_wbqspiflash_00_spi_spd), 
        .Y(n23735) );
  sky130_fd_sc_hd__clkinv_1 U14671 ( .A(j202_soc_core_j22_cpu_regop_imm__6_), 
        .Y(n12143) );
  sky130_fd_sc_hd__clkinv_1 U14672 ( .A(j202_soc_core_intr_vec__4_), .Y(n22900) );
  sky130_fd_sc_hd__clkinv_1 U14673 ( .A(j202_soc_core_j22_cpu_rf_tmp[26]), .Y(
        n13954) );
  sky130_fd_sc_hd__clkinv_1 U14674 ( .A(j202_soc_core_j22_cpu_pc[26]), .Y(
        n13955) );
  sky130_fd_sc_hd__clkinv_1 U14675 ( .A(j202_soc_core_j22_cpu_rf_pr[26]), .Y(
        n13958) );
  sky130_fd_sc_hd__clkinv_1 U14676 ( .A(j202_soc_core_j22_cpu_rf_gbr[26]), .Y(
        n13957) );
  sky130_fd_sc_hd__clkinv_1 U14677 ( .A(j202_soc_core_intc_core_00_rg_ipr[39]), 
        .Y(n24357) );
  sky130_fd_sc_hd__clkinv_1 U14678 ( .A(j202_soc_core_j22_cpu_rf_gpr[6]), .Y(
        n12204) );
  sky130_fd_sc_hd__clkinv_1 U14679 ( .A(j202_soc_core_j22_cpu_ml_mach[4]), .Y(
        n17092) );
  sky130_fd_sc_hd__clkinv_1 U14680 ( .A(j202_soc_core_j22_cpu_rf_gpr[25]), .Y(
        n13879) );
  sky130_fd_sc_hd__clkinv_1 U14681 ( .A(j202_soc_core_j22_cpu_ml_mach[1]), .Y(
        n19860) );
  sky130_fd_sc_hd__clkinv_1 U14682 ( .A(j202_soc_core_j22_cpu_ml_macl[8]), .Y(
        n19312) );
  sky130_fd_sc_hd__clkinv_1 U14683 ( .A(j202_soc_core_intc_core_00_rg_ipr[36]), 
        .Y(n24355) );
  sky130_fd_sc_hd__clkinv_1 U14684 ( .A(j202_soc_core_j22_cpu_rf_pr[7]), .Y(
        n16691) );
  sky130_fd_sc_hd__clkinv_1 U14685 ( .A(j202_soc_core_j22_cpu_rf_gpr[12]), .Y(
        n11944) );
  sky130_fd_sc_hd__clkinv_1 U14686 ( .A(j202_soc_core_j22_cpu_ml_macl[24]), 
        .Y(n15880) );
  sky130_fd_sc_hd__clkinv_1 U14687 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__3_), 
        .Y(n16692) );
  sky130_fd_sc_hd__clkinv_1 U14688 ( .A(j202_soc_core_j22_cpu_ml_macl[20]), 
        .Y(n15609) );
  sky130_fd_sc_hd__clkinv_1 U14689 ( .A(j202_soc_core_j22_cpu_rf_gbr[7]), .Y(
        n16693) );
  sky130_fd_sc_hd__clkinv_1 U14690 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .Y(n18479) );
  sky130_fd_sc_hd__clkinv_1 U14691 ( .A(j202_soc_core_intc_core_00_rg_ipr[38]), 
        .Y(n24356) );
  sky130_fd_sc_hd__clkinv_1 U14692 ( .A(j202_soc_core_j22_cpu_rf_tmp[9]), .Y(
        n19982) );
  sky130_fd_sc_hd__clkinv_1 U14693 ( .A(j202_soc_core_j22_cpu_ml_bufa[8]), .Y(
        n21922) );
  sky130_fd_sc_hd__clkinv_1 U14694 ( .A(j202_soc_core_j22_cpu_pc[9]), .Y(
        n19978) );
  sky130_fd_sc_hd__clkinv_1 U14695 ( .A(j202_soc_core_intc_core_00_rg_ipr[61]), 
        .Y(n24373) );
  sky130_fd_sc_hd__clkinv_1 U14696 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .Y(n24903) );
  sky130_fd_sc_hd__clkinv_1 U14697 ( .A(j202_soc_core_j22_cpu_rfuo_sr__m_), 
        .Y(n19974) );
  sky130_fd_sc_hd__clkinv_1 U14698 ( .A(j202_soc_core_j22_cpu_ml_macl[9]), .Y(
        n20013) );
  sky130_fd_sc_hd__clkinv_1 U14699 ( .A(j202_soc_core_j22_cpu_regop_imm__11_), 
        .Y(n11890) );
  sky130_fd_sc_hd__clkinv_1 U14700 ( .A(j202_soc_core_j22_cpu_ml_macl[25]), 
        .Y(n15894) );
  sky130_fd_sc_hd__clkinv_1 U14701 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[11]), .Y(n25184) );
  sky130_fd_sc_hd__clkinv_1 U14702 ( .A(j202_soc_core_intc_core_00_rg_ipr[62]), 
        .Y(n24374) );
  sky130_fd_sc_hd__clkinv_1 U14703 ( .A(j202_soc_core_qspi_wb_addr[10]), .Y(
        n20139) );
  sky130_fd_sc_hd__clkinv_1 U14704 ( .A(j202_soc_core_qspi_wb_addr[2]), .Y(
        n25053) );
  sky130_fd_sc_hd__clkinv_1 U14705 ( .A(j202_soc_core_intc_core_00_rg_ipr[54]), 
        .Y(n24702) );
  sky130_fd_sc_hd__clkinv_1 U14706 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[1]), .Y(n25156) );
  sky130_fd_sc_hd__clkinv_1 U14707 ( .A(j202_soc_core_j22_cpu_rf_gpr[17]), .Y(
        n11685) );
  sky130_fd_sc_hd__clkinv_1 U14708 ( .A(j202_soc_core_qspi_wb_addr[3]), .Y(
        n23409) );
  sky130_fd_sc_hd__clkinv_1 U14709 ( .A(j202_soc_core_j22_cpu_rf_gbr[15]), .Y(
        n15217) );
  sky130_fd_sc_hd__clkinv_1 U14710 ( .A(j202_soc_core_j22_cpu_ml_bufa[7]), .Y(
        n22235) );
  sky130_fd_sc_hd__clkinv_1 U14711 ( .A(j202_soc_core_j22_cpu_ml_bufa[9]), .Y(
        n21817) );
  sky130_fd_sc_hd__clkinv_1 U14712 ( .A(j202_soc_core_intc_core_00_rg_ipr[53]), 
        .Y(n24368) );
  sky130_fd_sc_hd__clkinv_1 U14713 ( .A(j202_soc_core_j22_cpu_ml_mach[26]), 
        .Y(n19558) );
  sky130_fd_sc_hd__clkinv_1 U14714 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]), .Y(n25069) );
  sky130_fd_sc_hd__clkinv_1 U14715 ( .A(j202_soc_core_j22_cpu_rf_gpr[23]), .Y(
        n12800) );
  sky130_fd_sc_hd__clkinv_1 U14716 ( .A(j202_soc_core_intc_core_00_rg_ipr[49]), 
        .Y(n24665) );
  sky130_fd_sc_hd__clkinv_1 U14717 ( .A(j202_soc_core_qspi_wb_addr[21]), .Y(
        n25067) );
  sky130_fd_sc_hd__clkinv_1 U14718 ( .A(j202_soc_core_intc_core_00_rg_ipr[51]), 
        .Y(n24366) );
  sky130_fd_sc_hd__clkinv_1 U14719 ( .A(j202_soc_core_j22_cpu_ml_mach[7]), .Y(
        n16628) );
  sky130_fd_sc_hd__clkinv_1 U14720 ( .A(j202_soc_core_intc_core_00_rg_ipr[48]), 
        .Y(n24364) );
  sky130_fd_sc_hd__clkinv_1 U14721 ( .A(j202_soc_core_j22_cpu_regop_imm__7_), 
        .Y(n12454) );
  sky130_fd_sc_hd__clkinv_1 U14722 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[8]), .Y(n25182) );
  sky130_fd_sc_hd__clkinv_1 U14723 ( .A(j202_soc_core_j22_cpu_rf_gpr[7]), .Y(
        n12517) );
  sky130_fd_sc_hd__clkinv_1 U14724 ( .A(j202_soc_core_j22_cpu_ml_mach[2]), .Y(
        n16835) );
  sky130_fd_sc_hd__clkinv_1 U14725 ( .A(j202_soc_core_intc_core_00_rg_ipr[32]), 
        .Y(n24351) );
  sky130_fd_sc_hd__clkinv_1 U14726 ( .A(j202_soc_core_j22_cpu_ml_mach[10]), 
        .Y(n16798) );
  sky130_fd_sc_hd__clkinv_1 U14727 ( .A(j202_soc_core_intc_core_00_rg_ipr[47]), 
        .Y(n24651) );
  sky130_fd_sc_hd__clkinv_1 U14728 ( .A(j202_soc_core_bldc_core_00_pwm_duty[3]), .Y(n25188) );
  sky130_fd_sc_hd__clkinv_1 U14729 ( .A(j202_soc_core_j22_cpu_rf_tmp[13]), .Y(
        n19120) );
  sky130_fd_sc_hd__clkinv_1 U14730 ( .A(j202_soc_core_j22_cpu_rf_pr[8]), .Y(
        n19200) );
  sky130_fd_sc_hd__clkinv_1 U14731 ( .A(j202_soc_core_intc_core_00_rg_ipr[46]), 
        .Y(n24363) );
  sky130_fd_sc_hd__clkinv_1 U14732 ( .A(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[4]), .Y(n12957) );
  sky130_fd_sc_hd__clkinv_1 U14733 ( .A(j202_soc_core_j22_cpu_ml_mach[14]), 
        .Y(n15467) );
  sky130_fd_sc_hd__clkinv_1 U14734 ( .A(j202_soc_core_j22_cpu_opst[3]), .Y(
        n20773) );
  sky130_fd_sc_hd__clkinv_1 U14735 ( .A(j202_soc_core_j22_cpu_regop_Ra__1_), 
        .Y(n12042) );
  sky130_fd_sc_hd__clkinv_1 U14736 ( .A(j202_soc_core_j22_cpu_opst[2]), .Y(
        n22417) );
  sky130_fd_sc_hd__clkinv_1 U14737 ( .A(j202_soc_core_intr_req_), .Y(n21399)
         );
  sky130_fd_sc_hd__clkinv_1 U14738 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[7]), .Y(n25180) );
  sky130_fd_sc_hd__clkinv_1 U14739 ( .A(j202_soc_core_j22_cpu_opst[1]), .Y(
        n21441) );
  sky130_fd_sc_hd__clkinv_1 U14740 ( .A(j202_soc_core_j22_cpu_ml_bufa[10]), 
        .Y(n21799) );
  sky130_fd_sc_hd__clkinv_1 U14741 ( .A(j202_soc_core_j22_cpu_regop_Rn__0_), 
        .Y(n11448) );
  sky130_fd_sc_hd__clkinv_1 U14742 ( .A(j202_soc_core_j22_cpu_macop_MAC_[1]), 
        .Y(n22923) );
  sky130_fd_sc_hd__clkinv_1 U14743 ( .A(j202_soc_core_j22_cpu_memop_MEM__1_), 
        .Y(n23242) );
  sky130_fd_sc_hd__clkinv_1 U14745 ( .A(j202_soc_core_j22_cpu_regop_Rn__2_), 
        .Y(n11447) );
  sky130_fd_sc_hd__clkinv_1 U14746 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[0]), 
        .Y(n22790) );
  sky130_fd_sc_hd__clkinv_1 U14747 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[2]), .Y(n12947) );
  sky130_fd_sc_hd__clkinv_1 U14748 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .Y(n20102) );
  sky130_fd_sc_hd__clkinv_1 U14749 ( .A(
        j202_soc_core_wbqspiflash_00_w_qspi_sck), .Y(n23587) );
  sky130_fd_sc_hd__clkinv_1 U14750 ( .A(j202_soc_core_j22_cpu_rf_pr[1]), .Y(
        n19837) );
  sky130_fd_sc_hd__clkinv_1 U14751 ( .A(j202_soc_core_j22_cpu_regop_Rn__1_), 
        .Y(n11446) );
  sky130_fd_sc_hd__clkinv_1 U14752 ( .A(j202_soc_core_j22_cpu_ml_mach[12]), 
        .Y(n17039) );
  sky130_fd_sc_hd__clkinv_1 U14753 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[6]), .Y(n11241) );
  sky130_fd_sc_hd__clkinv_1 U14754 ( .A(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]), .Y(n15239) );
  sky130_fd_sc_hd__clkinv_1 U14756 ( .A(j202_soc_core_j22_cpu_rf_tmp[3]), .Y(
        n18917) );
  sky130_fd_sc_hd__clkinv_1 U14757 ( .A(j202_soc_core_j22_cpu_rf_pr[3]), .Y(
        n18914) );
  sky130_fd_sc_hd__clkinv_1 U14758 ( .A(j202_soc_core_j22_cpu_pc[3]), .Y(
        n18918) );
  sky130_fd_sc_hd__clkinv_1 U14759 ( .A(j202_soc_core_j22_cpu_rf_gpr[3]), .Y(
        n12313) );
  sky130_fd_sc_hd__clkinv_1 U14760 ( .A(j202_soc_core_j22_cpu_rf_gbr[3]), .Y(
        n18913) );
  sky130_fd_sc_hd__clkinv_1 U14761 ( .A(j202_soc_core_j22_cpu_rfuo_sr__s_), 
        .Y(n21653) );
  sky130_fd_sc_hd__clkinv_1 U14762 ( .A(j202_soc_core_j22_cpu_ml_macl[17]), 
        .Y(n15941) );
  sky130_fd_sc_hd__clkinv_1 U14763 ( .A(j202_soc_core_j22_cpu_rf_gbr[1]), .Y(
        n19838) );
  sky130_fd_sc_hd__clkinv_1 U14764 ( .A(j202_soc_core_j22_cpu_regop_Rn__3_), 
        .Y(n11449) );
  sky130_fd_sc_hd__clkinv_1 U14765 ( .A(j202_soc_core_j22_cpu_rf_gbr[28]), .Y(
        n13861) );
  sky130_fd_sc_hd__clkinv_1 U14766 ( .A(j202_soc_core_j22_cpu_rf_pr[28]), .Y(
        n13862) );
  sky130_fd_sc_hd__clkinv_1 U14767 ( .A(j202_soc_core_j22_cpu_regop_Ra__0_), 
        .Y(n12971) );
  sky130_fd_sc_hd__clkinv_1 U14768 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[0]), .Y(n25172) );
  sky130_fd_sc_hd__clkinv_1 U14769 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__0_), 
        .Y(n20269) );
  sky130_fd_sc_hd__clkinv_1 U14770 ( .A(j202_soc_core_j22_cpu_memop_Ma__0_), 
        .Y(n13096) );
  sky130_fd_sc_hd__clkinv_1 U14771 ( .A(j202_soc_core_j22_cpu_pc[28]), .Y(
        n13859) );
  sky130_fd_sc_hd__clkinv_1 U14772 ( .A(j202_soc_core_j22_cpu_regop_Rb__0_), 
        .Y(n12930) );
  sky130_fd_sc_hd__clkinv_1 U14773 ( .A(j202_soc_core_j22_cpu_regop_Rs__0_), 
        .Y(n12931) );
  sky130_fd_sc_hd__clkinv_1 U14774 ( .A(j202_soc_core_j22_cpu_rf_tmp[28]), .Y(
        n13858) );
  sky130_fd_sc_hd__clkinv_1 U14775 ( .A(j202_soc_core_j22_cpu_rf_gpr[1]), .Y(
        n12022) );
  sky130_fd_sc_hd__clkinv_1 U14776 ( .A(j202_soc_core_j22_cpu_regop_We__2_), 
        .Y(n20478) );
  sky130_fd_sc_hd__clkinv_1 U14777 ( .A(j202_soc_core_j22_cpu_regop_imm__1_), 
        .Y(n11951) );
  sky130_fd_sc_hd__clkinv_1 U14778 ( .A(j202_soc_core_j22_cpu_regop_Rm__3_), 
        .Y(n11538) );
  sky130_fd_sc_hd__clkinv_1 U14779 ( .A(j202_soc_core_j22_cpu_ml_mach[13]), 
        .Y(n19104) );
  sky130_fd_sc_hd__clkinv_1 U14780 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[5]), 
        .Y(n22670) );
  sky130_fd_sc_hd__clkinv_1 U14781 ( .A(j202_soc_core_ahb2wbqspi_00_stb_o), 
        .Y(n20103) );
  sky130_fd_sc_hd__clkinv_1 U14782 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .Y(n16652) );
  sky130_fd_sc_hd__clkinv_1 U14784 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[3]), .Y(n18283) );
  sky130_fd_sc_hd__clkinv_1 U14785 ( .A(j202_soc_core_j22_cpu_regop_Rm__1_), 
        .Y(n11529) );
  sky130_fd_sc_hd__clkinv_1 U14786 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[4]), .Y(n11428) );
  sky130_fd_sc_hd__clkinv_1 U14787 ( .A(j202_soc_core_ahb2apb_00_state[0]), 
        .Y(n22764) );
  sky130_fd_sc_hd__clkinv_1 U14788 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[1]), .Y(n11430) );
  sky130_fd_sc_hd__clkinv_1 U14789 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[1]), 
        .Y(n22715) );
  sky130_fd_sc_hd__clkinv_1 U14790 ( .A(j202_soc_core_j22_cpu_macop_MAC_[4]), 
        .Y(n23247) );
  sky130_fd_sc_hd__clkinv_1 U14791 ( .A(j202_soc_core_j22_cpu_rf_gpr[28]), .Y(
        n13860) );
  sky130_fd_sc_hd__clkinv_1 U14792 ( .A(j202_soc_core_j22_cpu_ml_bufa[2]), .Y(
        n22238) );
  sky130_fd_sc_hd__clkinv_1 U14793 ( .A(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[0]), .Y(n21659) );
  sky130_fd_sc_hd__clkinv_1 U14794 ( .A(j202_soc_core_j22_cpu_regop_imm__0_), 
        .Y(n11987) );
  sky130_fd_sc_hd__clkinv_1 U14795 ( .A(j202_soc_core_j22_cpu_ml_bufa[11]), 
        .Y(n21960) );
  sky130_fd_sc_hd__clkinv_1 U14796 ( .A(j202_soc_core_j22_cpu_ma_M_address[1]), 
        .Y(n16650) );
  sky130_fd_sc_hd__clkinv_1 U14797 ( .A(j202_soc_core_j22_cpu_rf_gpr[0]), .Y(
        n19278) );
  sky130_fd_sc_hd__clkinv_1 U14798 ( .A(j202_soc_core_j22_cpu_regop_imm__12_), 
        .Y(n11472) );
  sky130_fd_sc_hd__clkinv_1 U14799 ( .A(j202_soc_core_aquc_ADR__2_), .Y(n15064) );
  sky130_fd_sc_hd__clkinv_1 U14801 ( .A(j202_soc_core_aquc_WE_), .Y(n11247) );
  sky130_fd_sc_hd__clkinv_1 U14802 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__1_), 
        .Y(n20235) );
  sky130_fd_sc_hd__clkinv_1 U14803 ( .A(j202_soc_core_j22_cpu_ml_macl[2]), .Y(
        n16843) );
  sky130_fd_sc_hd__inv_1 U14804 ( .A(j202_soc_core_memory0_ram_dout0_sel[3]), 
        .Y(n11312) );
  sky130_fd_sc_hd__clkinv_1 U14805 ( .A(j202_soc_core_j22_cpu_rf_tmp[0]), .Y(
        n19277) );
  sky130_fd_sc_hd__clkinv_1 U14806 ( .A(j202_soc_core_aquc_ADR__4_), .Y(n11255) );
  sky130_fd_sc_hd__clkinv_1 U14807 ( .A(j202_soc_core_j22_cpu_ml_macl[1]), .Y(
        n19869) );
  sky130_fd_sc_hd__clkinv_1 U14808 ( .A(j202_soc_core_memory0_ram_dout0_sel[5]), .Y(n11293) );
  sky130_fd_sc_hd__clkinv_1 U14809 ( .A(j202_soc_core_j22_cpu_regop_other__0_), 
        .Y(n11556) );
  sky130_fd_sc_hd__clkinv_1 U14810 ( .A(j202_soc_core_j22_cpu_ifetchl), .Y(
        n22807) );
  sky130_fd_sc_hd__clkinv_1 U14811 ( .A(j202_soc_core_j22_cpu_pc[0]), .Y(
        n21630) );
  sky130_fd_sc_hd__clkinv_1 U14812 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__3_), 
        .Y(n20487) );
  sky130_fd_sc_hd__clkinv_1 U14813 ( .A(j202_soc_core_j22_cpu_istall), .Y(
        n12914) );
  sky130_fd_sc_hd__clkinv_1 U14814 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[0]), 
        .Y(n25206) );
  sky130_fd_sc_hd__clkinv_1 U14815 ( .A(j202_soc_core_j22_cpu_regop_other__1_), 
        .Y(n12941) );
  sky130_fd_sc_hd__clkinv_1 U14816 ( .A(j202_soc_core_j22_cpu_pc[1]), .Y(
        n21647) );
  sky130_fd_sc_hd__clkinv_1 U14817 ( .A(
        j202_soc_core_memory0_ram_dout0_sel[12]), .Y(n11289) );
  sky130_fd_sc_hd__clkinv_1 U14818 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[3]), .Y(n22128) );
  sky130_fd_sc_hd__clkinv_1 U14819 ( .A(j202_soc_core_j22_cpu_rf_gbr[0]), .Y(
        n19274) );
  sky130_fd_sc_hd__clkinv_1 U14820 ( .A(j202_soc_core_j22_cpu_rf_gpr[2]), .Y(
        n12041) );
  sky130_fd_sc_hd__clkinv_1 U14821 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[1]), 
        .Y(n25203) );
  sky130_fd_sc_hd__clkinv_1 U14822 ( .A(j202_soc_core_memory0_ram_dout0_sel[8]), .Y(n11291) );
  sky130_fd_sc_hd__clkinv_1 U14823 ( .A(
        j202_soc_core_memory0_ram_dout0_sel[10]), .Y(n11290) );
  sky130_fd_sc_hd__clkinv_1 U14824 ( .A(j202_soc_core_memory0_ram_dout0_sel[2]), .Y(n11309) );
  sky130_fd_sc_hd__clkinv_1 U14825 ( .A(j202_soc_core_j22_cpu_ml_mach[11]), 
        .Y(n15262) );
  sky130_fd_sc_hd__clkinv_1 U14826 ( .A(j202_soc_core_j22_cpu_ml_macl[18]), 
        .Y(n15951) );
  sky130_fd_sc_hd__clkinv_1 U14827 ( .A(j202_soc_core_j22_cpu_rf_pr[0]), .Y(
        n19273) );
  sky130_fd_sc_hd__nor2_2 U14951 ( .A(n11512), .B(n11511), .Y(n14089) );
  sky130_fd_sc_hd__nand2_1 U14953 ( .A(n11520), .B(
        j202_soc_core_j22_cpu_regop_Rm__0_), .Y(n11539) );
  sky130_fd_sc_hd__nor2_2 U14954 ( .A(n11540), .B(n11539), .Y(n20296) );
  sky130_fd_sc_hd__nor2_2 U14955 ( .A(n11534), .B(n11533), .Y(n11193) );
  sky130_fd_sc_hd__inv_6 U14956 ( .A(n11167), .Y(n11168) );
  sky130_fd_sc_hd__clkinv_1 U14957 ( .A(n13395), .Y(n12787) );
  sky130_fd_sc_hd__clkinv_1 U14958 ( .A(n14273), .Y(n13999) );
  sky130_fd_sc_hd__clkinv_1 U14959 ( .A(n18828), .Y(n12651) );
  sky130_fd_sc_hd__clkinv_1 U14960 ( .A(n18493), .Y(n12719) );
  sky130_fd_sc_hd__clkinv_1 U14961 ( .A(n19096), .Y(n19920) );
  sky130_fd_sc_hd__clkinv_1 U14962 ( .A(n14180), .Y(n14039) );
  sky130_fd_sc_hd__a21boi_0 U14963 ( .A1(n22531), .A2(n16647), .B1_N(n16646), 
        .Y(n16648) );
  sky130_fd_sc_hd__clkinv_1 U14964 ( .A(n13102), .Y(n12845) );
  sky130_fd_sc_hd__clkinv_1 U14965 ( .A(n19653), .Y(n12685) );
  sky130_fd_sc_hd__nand3_1 U14966 ( .A(n12982), .B(n12981), .C(n12980), .Y(
        n13537) );
  sky130_fd_sc_hd__nor2_1 U14967 ( .A(n12969), .B(n22801), .Y(n12981) );
  sky130_fd_sc_hd__clkinv_1 U14968 ( .A(n13188), .Y(n12753) );
  sky130_fd_sc_hd__nand2_1 U14969 ( .A(j202_soc_core_ahbcs_6__HREADY_), .B(
        n12909), .Y(n21657) );
  sky130_fd_sc_hd__clkinv_1 U14970 ( .A(j202_soc_core_j22_cpu_ml_bufa[19]), 
        .Y(n20042) );
  sky130_fd_sc_hd__clkinv_1 U14971 ( .A(n22112), .Y(n23303) );
  sky130_fd_sc_hd__nand3_1 U14972 ( .A(n17106), .B(n17105), .C(n17104), .Y(
        n22484) );
  sky130_fd_sc_hd__clkinv_1 U14973 ( .A(n22378), .Y(n22759) );
  sky130_fd_sc_hd__maj3_1 U14974 ( .A(n17320), .B(n17321), .C(n17219), .X(
        n17220) );
  sky130_fd_sc_hd__nor2_1 U14975 ( .A(n16190), .B(n16595), .Y(n16581) );
  sky130_fd_sc_hd__clkinv_1 U14976 ( .A(n16581), .Y(n16546) );
  sky130_fd_sc_hd__nand2_1 U14977 ( .A(n21796), .B(n15244), .Y(n16595) );
  sky130_fd_sc_hd__nand2_1 U14978 ( .A(n15232), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .Y(n16191) );
  sky130_fd_sc_hd__clkinv_1 U14979 ( .A(n21683), .Y(n22565) );
  sky130_fd_sc_hd__clkinv_1 U14980 ( .A(n14042), .Y(n13681) );
  sky130_fd_sc_hd__nor2_1 U14981 ( .A(j202_soc_core_j22_cpu_regop_Rm__0_), .B(
        n11529), .Y(n11537) );
  sky130_fd_sc_hd__clkinv_1 U14982 ( .A(n19247), .Y(n12124) );
  sky130_fd_sc_hd__a21oi_1 U14983 ( .A1(n19920), .A2(n19667), .B1(n19666), .Y(
        n19672) );
  sky130_fd_sc_hd__nand2_1 U14984 ( .A(n16593), .B(n20007), .Y(n19953) );
  sky130_fd_sc_hd__nand2_1 U14985 ( .A(n16592), .B(n16191), .Y(n19959) );
  sky130_fd_sc_hd__clkinv_1 U14986 ( .A(n22136), .Y(n22556) );
  sky130_fd_sc_hd__and2_0 U14987 ( .A(n15944), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15945) );
  sky130_fd_sc_hd__nand3_1 U14988 ( .A(n16590), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .C(n21659), .Y(n20007) );
  sky130_fd_sc_hd__a2bb2oi_1 U14989 ( .B1(n21722), .B2(n21721), .A1_N(n21720), 
        .A2_N(n21721), .Y(n21729) );
  sky130_fd_sc_hd__nor2_1 U14990 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[4]), .B(n15239), .Y(n15241) );
  sky130_fd_sc_hd__a21boi_0 U14991 ( .A1(n17165), .A2(n17223), .B1_N(n17222), 
        .Y(n21382) );
  sky130_fd_sc_hd__nand2_1 U14992 ( .A(n20488), .B(n12967), .Y(n23235) );
  sky130_fd_sc_hd__a21boi_0 U14993 ( .A1(n17254), .A2(n17311), .B1_N(n17310), 
        .Y(n21375) );
  sky130_fd_sc_hd__clkinv_1 U14994 ( .A(n25380), .Y(n21420) );
  sky130_fd_sc_hd__clkinv_1 U14995 ( .A(n23304), .Y(n21787) );
  sky130_fd_sc_hd__nand3_1 U14996 ( .A(n12027), .B(n12026), .C(n12025), .Y(
        n22183) );
  sky130_fd_sc_hd__clkinv_1 U14997 ( .A(n25260), .Y(n21248) );
  sky130_fd_sc_hd__nand2_1 U14998 ( .A(n21249), .B(n21246), .Y(n19799) );
  sky130_fd_sc_hd__clkinv_1 U14999 ( .A(n22156), .Y(n21862) );
  sky130_fd_sc_hd__clkinv_1 U15000 ( .A(n22154), .Y(n22275) );
  sky130_fd_sc_hd__clkinv_1 U15001 ( .A(n21731), .Y(n22190) );
  sky130_fd_sc_hd__clkinv_1 U15002 ( .A(j202_soc_core_j22_cpu_ml_bufa[22]), 
        .Y(n19536) );
  sky130_fd_sc_hd__clkinv_1 U15003 ( .A(n22131), .Y(n22084) );
  sky130_fd_sc_hd__clkinv_1 U15004 ( .A(n22270), .Y(n22274) );
  sky130_fd_sc_hd__clkinv_1 U15005 ( .A(n22269), .Y(n20671) );
  sky130_fd_sc_hd__and2_0 U15006 ( .A(n25388), .B(n22530), .X(n20639) );
  sky130_fd_sc_hd__nand2_1 U15007 ( .A(n21009), .B(n20903), .Y(n23300) );
  sky130_fd_sc_hd__a21oi_1 U15008 ( .A1(n20926), .A2(n21137), .B1(n20925), .Y(
        n22371) );
  sky130_fd_sc_hd__clkinv_1 U15009 ( .A(n21803), .Y(n22168) );
  sky130_fd_sc_hd__nand3_1 U15010 ( .A(n20543), .B(n20542), .C(n20541), .Y(
        n21924) );
  sky130_fd_sc_hd__and2_0 U15011 ( .A(n22524), .B(n22530), .X(n21104) );
  sky130_fd_sc_hd__clkinv_1 U15012 ( .A(n21834), .Y(n21838) );
  sky130_fd_sc_hd__clkinv_1 U15013 ( .A(n13293), .Y(n13295) );
  sky130_fd_sc_hd__and2_0 U15014 ( .A(n21135), .B(n22530), .X(n21136) );
  sky130_fd_sc_hd__clkinv_1 U15015 ( .A(n21874), .Y(n21204) );
  sky130_fd_sc_hd__clkinv_1 U15016 ( .A(n22514), .Y(n22158) );
  sky130_fd_sc_hd__a21boi_0 U15017 ( .A1(n20587), .A2(n21152), .B1_N(n20586), 
        .Y(n20589) );
  sky130_fd_sc_hd__clkinv_1 U15018 ( .A(n22515), .Y(n22350) );
  sky130_fd_sc_hd__and2_0 U15019 ( .A(n21009), .B(n20953), .X(n21949) );
  sky130_fd_sc_hd__nand3_1 U15020 ( .A(n20798), .B(n20797), .C(n20796), .Y(
        n21752) );
  sky130_fd_sc_hd__and2_0 U15021 ( .A(n21009), .B(n20801), .X(n22112) );
  sky130_fd_sc_hd__nand2_1 U15022 ( .A(n22216), .B(n22218), .Y(n22221) );
  sky130_fd_sc_hd__nand2_1 U15023 ( .A(n21729), .B(n21728), .Y(n22218) );
  sky130_fd_sc_hd__clkinv_1 U15024 ( .A(n22216), .Y(n22213) );
  sky130_fd_sc_hd__clkinv_1 U15025 ( .A(n22198), .Y(n22219) );
  sky130_fd_sc_hd__a21boi_1 U15026 ( .A1(n25274), .A2(n19895), .B1_N(n19894), 
        .Y(n22662) );
  sky130_fd_sc_hd__clkinv_1 U15027 ( .A(n23324), .Y(n22605) );
  sky130_fd_sc_hd__and2_0 U15028 ( .A(n22541), .B(n22530), .X(n21078) );
  sky130_fd_sc_hd__clkinv_1 U15029 ( .A(n21761), .Y(n21764) );
  sky130_fd_sc_hd__clkinv_1 U15030 ( .A(n23319), .Y(n22613) );
  sky130_fd_sc_hd__nand3_1 U15031 ( .A(n12110), .B(n12109), .C(n12108), .Y(
        n22185) );
  sky130_fd_sc_hd__clkinv_1 U15032 ( .A(n14802), .Y(n14804) );
  sky130_fd_sc_hd__nand2_1 U15033 ( .A(n23239), .B(n20243), .Y(n21188) );
  sky130_fd_sc_hd__and2_0 U15034 ( .A(n21009), .B(n20827), .X(n22512) );
  sky130_fd_sc_hd__nand3_1 U15035 ( .A(n16864), .B(n16863), .C(n16862), .Y(
        n22547) );
  sky130_fd_sc_hd__clkinv_1 U15036 ( .A(n22372), .Y(n22345) );
  sky130_fd_sc_hd__nand3_1 U15037 ( .A(n19271), .B(n19270), .C(n19269), .Y(
        n21613) );
  sky130_fd_sc_hd__a21boi_0 U15038 ( .A1(n22725), .A2(n19266), .B1_N(n19265), 
        .Y(n19270) );
  sky130_fd_sc_hd__clkinv_1 U15039 ( .A(n22081), .Y(n23335) );
  sky130_fd_sc_hd__clkinv_1 U15040 ( .A(n21850), .Y(n20515) );
  sky130_fd_sc_hd__clkinv_1 U15041 ( .A(n22555), .Y(n22492) );
  sky130_fd_sc_hd__clkinv_1 U15042 ( .A(n22033), .Y(n20514) );
  sky130_fd_sc_hd__clkinv_1 U15043 ( .A(n22554), .Y(n22299) );
  sky130_fd_sc_hd__clkinv_1 U15044 ( .A(n25369), .Y(n22342) );
  sky130_fd_sc_hd__nand4_1 U15045 ( .A(n20221), .B(
        j202_soc_core_ahbcs_6__HREADY_), .C(n21599), .D(n12914), .Y(n12983) );
  sky130_fd_sc_hd__and2_0 U15046 ( .A(n20981), .B(n25385), .X(n24826) );
  sky130_fd_sc_hd__nand3_1 U15047 ( .A(n18894), .B(n18893), .C(n18892), .Y(
        n22013) );
  sky130_fd_sc_hd__a21oi_1 U15048 ( .A1(n19115), .A2(n14086), .B1(n12647), .Y(
        n22300) );
  sky130_fd_sc_hd__clkinv_1 U15049 ( .A(n21981), .Y(n23338) );
  sky130_fd_sc_hd__clkinv_1 U15050 ( .A(n14531), .Y(n14533) );
  sky130_fd_sc_hd__clkinv_1 U15051 ( .A(n22512), .Y(n23329) );
  sky130_fd_sc_hd__clkinv_1 U15052 ( .A(n13967), .Y(n12901) );
  sky130_fd_sc_hd__nand3_1 U15053 ( .A(n17133), .B(n17132), .C(n17131), .Y(
        n22057) );
  sky130_fd_sc_hd__nand2_1 U15054 ( .A(n21009), .B(n21008), .Y(n23348) );
  sky130_fd_sc_hd__nor2_1 U15055 ( .A(n21624), .B(n21623), .Y(n22360) );
  sky130_fd_sc_hd__clkinv_1 U15056 ( .A(n22484), .Y(n22536) );
  sky130_fd_sc_hd__and2_0 U15057 ( .A(n19470), .B(n19192), .X(n19619) );
  sky130_fd_sc_hd__nand3_1 U15058 ( .A(n19023), .B(n19022), .C(n19021), .Y(
        n22045) );
  sky130_fd_sc_hd__and2_0 U15059 ( .A(n19547), .B(n19064), .X(n19767) );
  sky130_fd_sc_hd__clkinv_1 U15060 ( .A(n22495), .Y(n22290) );
  sky130_fd_sc_hd__and2_0 U15061 ( .A(n20065), .B(n18924), .X(n19830) );
  sky130_fd_sc_hd__nand2_1 U15062 ( .A(n21009), .B(n20779), .Y(n23309) );
  sky130_fd_sc_hd__clkinv_1 U15063 ( .A(n23307), .Y(n22642) );
  sky130_fd_sc_hd__clkinv_1 U15064 ( .A(n13541), .Y(n13543) );
  sky130_fd_sc_hd__fa_1 U15065 ( .A(n14677), .B(n14676), .CIN(n14093), .COUT(
        n20674), .SUM(n21892) );
  sky130_fd_sc_hd__clkinv_1 U15066 ( .A(n21890), .Y(n23342) );
  sky130_fd_sc_hd__a21boi_0 U15067 ( .A1(n24869), .A2(n20768), .B1_N(n22741), 
        .Y(n21580) );
  sky130_fd_sc_hd__a21oi_1 U15068 ( .A1(n18912), .A2(n14086), .B1(n12318), .Y(
        n22711) );
  sky130_fd_sc_hd__clkinv_1 U15069 ( .A(n25372), .Y(n22330) );
  sky130_fd_sc_hd__clkinv_1 U15071 ( .A(n22360), .Y(n22752) );
  sky130_fd_sc_hd__and2_0 U15072 ( .A(n22540), .B(n22530), .X(n20406) );
  sky130_fd_sc_hd__clkinv_1 U15073 ( .A(n23310), .Y(n22640) );
  sky130_fd_sc_hd__clkinv_1 U15074 ( .A(n13403), .Y(n13405) );
  sky130_fd_sc_hd__clkinv_1 U15075 ( .A(n22181), .Y(n22264) );
  sky130_fd_sc_hd__clkinv_1 U15076 ( .A(n21644), .Y(n24863) );
  sky130_fd_sc_hd__nand2_1 U15077 ( .A(n23239), .B(n25731), .Y(n21592) );
  sky130_fd_sc_hd__nor2_1 U15078 ( .A(n19324), .B(n21592), .Y(n24879) );
  sky130_fd_sc_hd__and2_0 U15080 ( .A(n25339), .B(n25391), .X(n25437) );
  sky130_fd_sc_hd__and2_0 U15081 ( .A(n25339), .B(n25333), .X(n25438) );
  sky130_fd_sc_hd__and2_0 U15082 ( .A(n25339), .B(n25334), .X(n25439) );
  sky130_fd_sc_hd__and2_0 U15083 ( .A(n25339), .B(n25335), .X(n25440) );
  sky130_fd_sc_hd__and2_0 U15084 ( .A(n25339), .B(n25336), .X(n25441) );
  sky130_fd_sc_hd__and2_0 U15085 ( .A(n25339), .B(n25337), .X(n25442) );
  sky130_fd_sc_hd__and2_0 U15086 ( .A(n25339), .B(n25338), .X(n25443) );
  sky130_fd_sc_hd__and2_0 U15087 ( .A(n25339), .B(n22100), .X(n25445) );
  sky130_fd_sc_hd__and2_0 U15088 ( .A(n25339), .B(n21906), .X(n25428) );
  sky130_fd_sc_hd__and2_0 U15089 ( .A(n25339), .B(n25379), .X(n25446) );
  sky130_fd_sc_hd__nand3_1 U15090 ( .A(n18222), .B(n18221), .C(n18220), .Y(
        n25381) );
  sky130_fd_sc_hd__nand2_1 U15091 ( .A(n18219), .B(n18218), .Y(n25377) );
  sky130_fd_sc_hd__clkinv_1 U15092 ( .A(j202_soc_core_j22_cpu_ml_macl[31]), 
        .Y(n16190) );
  sky130_fd_sc_hd__clkinv_1 U15093 ( .A(n16399), .Y(n16384) );
  sky130_fd_sc_hd__clkinv_1 U15094 ( .A(n19345), .Y(n19341) );
  sky130_fd_sc_hd__nand4bb_1 U15095 ( .A_N(n14728), .B_N(n14727), .C(n14726), 
        .D(n14725), .Y(n14729) );
  sky130_fd_sc_hd__nand4bb_1 U15096 ( .A_N(n14719), .B_N(n14738), .C(n14718), 
        .D(n14717), .Y(n14722) );
  sky130_fd_sc_hd__and2_0 U15097 ( .A(n15016), .B(
        j202_soc_core_bootrom_00_address_w[3]), .X(n14851) );
  sky130_fd_sc_hd__and2_0 U15098 ( .A(n14456), .B(
        j202_soc_core_bootrom_00_address_w[9]), .X(n13199) );
  sky130_fd_sc_hd__clkinv_1 U15099 ( .A(n22839), .Y(n20174) );
  sky130_fd_sc_hd__clkinv_1 U15100 ( .A(n19629), .Y(n19596) );
  sky130_fd_sc_hd__inv_2 U15101 ( .A(n12920), .Y(n11477) );
  sky130_fd_sc_hd__clkinv_1 U15102 ( .A(n19253), .Y(n19255) );
  sky130_fd_sc_hd__clkinv_1 U15103 ( .A(n21145), .Y(n20385) );
  sky130_fd_sc_hd__and2_0 U15104 ( .A(n22691), .B(n22589), .X(n20370) );
  sky130_fd_sc_hd__nand4bb_1 U15105 ( .A_N(n22469), .B_N(n22468), .C(n22467), 
        .D(n22466), .Y(n22675) );
  sky130_fd_sc_hd__clkinv_1 U15106 ( .A(n22435), .Y(n22443) );
  sky130_fd_sc_hd__and2_0 U15107 ( .A(n14456), .B(
        j202_soc_core_bootrom_00_address_w[10]), .X(n14850) );
  sky130_fd_sc_hd__and2_0 U15108 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .B(j202_soc_core_bootrom_00_address_w[11]), .X(n14724) );
  sky130_fd_sc_hd__and2_0 U15109 ( .A(n14774), .B(n14773), .X(n14775) );
  sky130_fd_sc_hd__and2_0 U15110 ( .A(n13589), .B(
        j202_soc_core_bootrom_00_address_w[9]), .X(n17975) );
  sky130_fd_sc_hd__and2_0 U15111 ( .A(n14279), .B(n13054), .X(n14583) );
  sky130_fd_sc_hd__and2_0 U15112 ( .A(n14188), .B(n13014), .X(n14565) );
  sky130_fd_sc_hd__a21boi_0 U15113 ( .A1(n14313), .A2(n14314), .B1_N(n13013), 
        .Y(n14542) );
  sky130_fd_sc_hd__and2_0 U15114 ( .A(n14399), .B(n13014), .X(n13056) );
  sky130_fd_sc_hd__and2_0 U15115 ( .A(n13440), .B(n13014), .X(n13114) );
  sky130_fd_sc_hd__and2_0 U15116 ( .A(n13440), .B(
        j202_soc_core_bootrom_00_address_w[2]), .X(n13463) );
  sky130_fd_sc_hd__clkinv_1 U15117 ( .A(j202_soc_core_intr_level__1_), .Y(
        n14927) );
  sky130_fd_sc_hd__clkinv_1 U15118 ( .A(n21963), .Y(n22643) );
  sky130_fd_sc_hd__clkinv_1 U15119 ( .A(n22577), .Y(n22641) );
  sky130_fd_sc_hd__clkinv_1 U15120 ( .A(n21775), .Y(n22566) );
  sky130_fd_sc_hd__and2_0 U15121 ( .A(n20206), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]), .X(n20207) );
  sky130_fd_sc_hd__clkinv_1 U15122 ( .A(n16580), .Y(n19623) );
  sky130_fd_sc_hd__clkinv_1 U15123 ( .A(j202_soc_core_j22_cpu_ml_mach[30]), 
        .Y(n19621) );
  sky130_fd_sc_hd__clkinv_1 U15124 ( .A(n22133), .Y(n22563) );
  sky130_fd_sc_hd__clkinv_1 U15125 ( .A(n21935), .Y(n22568) );
  sky130_fd_sc_hd__clkinv_1 U15126 ( .A(n21867), .Y(n22567) );
  sky130_fd_sc_hd__clkinv_1 U15127 ( .A(n22576), .Y(n22610) );
  sky130_fd_sc_hd__clkinv_1 U15128 ( .A(n14071), .Y(n14020) );
  sky130_fd_sc_hd__clkinv_1 U15129 ( .A(n14079), .Y(n14027) );
  sky130_fd_sc_hd__clkinv_1 U15130 ( .A(n14075), .Y(n14026) );
  sky130_fd_sc_hd__clkinv_1 U15131 ( .A(n14073), .Y(n14025) );
  sky130_fd_sc_hd__clkinv_1 U15132 ( .A(n15933), .Y(n16189) );
  sky130_fd_sc_hd__nor2_1 U15133 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]), .B(n12957), .Y(n15232) );
  sky130_fd_sc_hd__clkinv_1 U15134 ( .A(n22706), .Y(n22594) );
  sky130_fd_sc_hd__clkinv_1 U15135 ( .A(n22574), .Y(n22606) );
  sky130_fd_sc_hd__clkinv_1 U15136 ( .A(n21828), .Y(n22614) );
  sky130_fd_sc_hd__nor2_1 U15137 ( .A(n11477), .B(n20258), .Y(n13904) );
  sky130_fd_sc_hd__nor2_1 U15138 ( .A(n11477), .B(n20302), .Y(n13921) );
  sky130_fd_sc_hd__nor2_1 U15139 ( .A(n11477), .B(n20241), .Y(n13923) );
  sky130_fd_sc_hd__nor2_1 U15140 ( .A(n11477), .B(n20266), .Y(n13912) );
  sky130_fd_sc_hd__nor2_1 U15141 ( .A(n11477), .B(n20272), .Y(n13896) );
  sky130_fd_sc_hd__nor2_1 U15142 ( .A(n11477), .B(n20280), .Y(n13922) );
  sky130_fd_sc_hd__nor2_1 U15143 ( .A(n11477), .B(n20291), .Y(n13894) );
  sky130_fd_sc_hd__and2_0 U15144 ( .A(n11470), .B(n12971), .X(n11184) );
  sky130_fd_sc_hd__nor2_1 U15145 ( .A(n11477), .B(n20289), .Y(n13903) );
  sky130_fd_sc_hd__nor2_1 U15146 ( .A(n11477), .B(n20294), .Y(n13895) );
  sky130_fd_sc_hd__nor2_1 U15147 ( .A(n11477), .B(n20305), .Y(n13902) );
  sky130_fd_sc_hd__nor2_1 U15148 ( .A(n11477), .B(n20283), .Y(n13911) );
  sky130_fd_sc_hd__and2_0 U15149 ( .A(j202_soc_core_j22_cpu_regop_Rn__1_), .B(
        j202_soc_core_j22_cpu_regop_Rn__0_), .X(n11473) );
  sky130_fd_sc_hd__inv_2 U15150 ( .A(n20270), .Y(n14059) );
  sky130_fd_sc_hd__inv_2 U15151 ( .A(n20265), .Y(n14058) );
  sky130_fd_sc_hd__clkinv_1 U15152 ( .A(n21063), .Y(n21143) );
  sky130_fd_sc_hd__nand2_1 U15153 ( .A(n21139), .B(n16870), .Y(n20905) );
  sky130_fd_sc_hd__clkinv_1 U15154 ( .A(n22573), .Y(n22601) );
  sky130_fd_sc_hd__nor2_1 U15155 ( .A(n19153), .B(n16662), .Y(n21164) );
  sky130_fd_sc_hd__clkinv_1 U15156 ( .A(n22578), .Y(n22600) );
  sky130_fd_sc_hd__and2_0 U15157 ( .A(n13166), .B(n13311), .X(n13456) );
  sky130_fd_sc_hd__nand2_1 U15158 ( .A(n11468), .B(
        j202_soc_core_j22_cpu_regop_Ra__0_), .Y(n13919) );
  sky130_fd_sc_hd__clkinv_1 U15159 ( .A(n21150), .Y(n21089) );
  sky130_fd_sc_hd__nor2_1 U15160 ( .A(n16653), .B(n20931), .Y(n21170) );
  sky130_fd_sc_hd__clkinv_1 U15161 ( .A(n20904), .Y(n20908) );
  sky130_fd_sc_hd__and2_0 U15162 ( .A(j202_soc_core_j22_cpu_regop_Rn__2_), .B(
        j202_soc_core_j22_cpu_regop_Rn__3_), .X(n11476) );
  sky130_fd_sc_hd__clkinv_1 U15163 ( .A(n14077), .Y(n14028) );
  sky130_fd_sc_hd__nand2_1 U15164 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[0]), .Y(n22509) );
  sky130_fd_sc_hd__and2_0 U15165 ( .A(n14403), .B(n14451), .X(n14145) );
  sky130_fd_sc_hd__clkinv_1 U15166 ( .A(n14720), .Y(n14871) );
  sky130_fd_sc_hd__clkinv_1 U15167 ( .A(n13121), .Y(n13500) );
  sky130_fd_sc_hd__clkinv_1 U15168 ( .A(n13489), .Y(n17468) );
  sky130_fd_sc_hd__clkinv_1 U15169 ( .A(n13483), .Y(n17730) );
  sky130_fd_sc_hd__clkinv_1 U15170 ( .A(j202_soc_core_memory0_ram_dout0_sel[6]), .Y(n11301) );
  sky130_fd_sc_hd__clkinv_1 U15171 ( .A(j202_soc_core_bootrom_00_address_w[3]), 
        .Y(n14100) );
  sky130_fd_sc_hd__clkinv_1 U15172 ( .A(n16990), .Y(n18645) );
  sky130_fd_sc_hd__and2_0 U15173 ( .A(n11302), .B(
        j202_soc_core_memory0_ram_dout0_sel[12]), .X(n18745) );
  sky130_fd_sc_hd__and2_0 U15174 ( .A(n17639), .B(
        j202_soc_core_memory0_ram_dout0_sel[7]), .X(n18744) );
  sky130_fd_sc_hd__and2_0 U15175 ( .A(n11299), .B(
        j202_soc_core_memory0_ram_dout0_sel[10]), .X(n18740) );
  sky130_fd_sc_hd__clkinv_1 U15176 ( .A(j202_soc_core_bootrom_00_address_w[10]), .Y(n14983) );
  sky130_fd_sc_hd__nor2_1 U15177 ( .A(n11292), .B(n11297), .Y(n17639) );
  sky130_fd_sc_hd__clkinv_1 U15178 ( .A(j202_soc_core_bootrom_00_address_w[11]), .Y(n15017) );
  sky130_fd_sc_hd__clkinv_1 U15179 ( .A(j202_soc_core_intr_level__3_), .Y(
        n14926) );
  sky130_fd_sc_hd__clkinv_1 U15180 ( .A(j202_soc_core_intr_level__2_), .Y(
        n14925) );
  sky130_fd_sc_hd__clkinv_1 U15181 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .Y(n14998) );
  sky130_fd_sc_hd__clkinv_1 U15182 ( .A(j202_soc_core_bootrom_00_address_w[7]), 
        .Y(n14999) );
  sky130_fd_sc_hd__clkinv_1 U15183 ( .A(n16736), .Y(n18354) );
  sky130_fd_sc_hd__clkinv_1 U15184 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[1]), 
        .Y(n16643) );
  sky130_fd_sc_hd__clkinv_1 U15185 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[0]), 
        .Y(n20352) );
  sky130_fd_sc_hd__clkinv_1 U15186 ( .A(n18276), .Y(n18281) );
  sky130_fd_sc_hd__clkinv_1 U15187 ( .A(j202_soc_core_j22_cpu_rf_gpr[489]), 
        .Y(n19987) );
  sky130_fd_sc_hd__clkinv_1 U15188 ( .A(j202_soc_core_j22_cpu_rf_gbr[9]), .Y(
        n19976) );
  sky130_fd_sc_hd__clkinv_1 U15189 ( .A(j202_soc_core_j22_cpu_rf_vbr[17]), .Y(
        n19909) );
  sky130_fd_sc_hd__clkinv_1 U15190 ( .A(j202_soc_core_j22_cpu_rf_gpr[481]), 
        .Y(n19841) );
  sky130_fd_sc_hd__clkinv_1 U15191 ( .A(n24776), .Y(n24705) );
  sky130_fd_sc_hd__clkinv_1 U15192 ( .A(
        j202_soc_core_intc_core_00_in_intreq[7]), .Y(n24572) );
  sky130_fd_sc_hd__clkinv_1 U15193 ( .A(j202_soc_core_intc_core_00_bs_addr[6]), 
        .Y(n24468) );
  sky130_fd_sc_hd__clkinv_1 U15194 ( .A(j202_soc_core_intc_core_00_bs_addr[3]), 
        .Y(n24453) );
  sky130_fd_sc_hd__and2_0 U15195 ( .A(j202_soc_core_intc_core_00_bs_addr[6]), 
        .B(j202_soc_core_intc_core_00_bs_addr[4]), .X(n24457) );
  sky130_fd_sc_hd__clkinv_1 U15196 ( .A(n22789), .Y(n21215) );
  sky130_fd_sc_hd__clkinv_1 U15197 ( .A(n25261), .Y(n21246) );
  sky130_fd_sc_hd__clkinv_1 U15198 ( .A(j202_soc_core_j22_cpu_rf_vbr[30]), .Y(
        n19756) );
  sky130_fd_sc_hd__clkinv_1 U15199 ( .A(j202_soc_core_j22_cpu_rf_vbr[24]), .Y(
        n19709) );
  sky130_fd_sc_hd__nand2_1 U15200 ( .A(n11445), .B(n11568), .Y(n13706) );
  sky130_fd_sc_hd__clkinv_1 U15201 ( .A(j202_soc_core_j22_cpu_rf_vbr[31]), .Y(
        n19641) );
  sky130_fd_sc_hd__clkinv_1 U15202 ( .A(j202_soc_core_j22_cpu_ml_mach[31]), 
        .Y(n19622) );
  sky130_fd_sc_hd__clkinv_1 U15203 ( .A(j202_soc_core_j22_cpu_ml_bufa[27]), 
        .Y(n19811) );
  sky130_fd_sc_hd__clkinv_1 U15204 ( .A(n19507), .Y(n19508) );
  sky130_fd_sc_hd__clkinv_1 U15205 ( .A(n21795), .Y(n20040) );
  sky130_fd_sc_hd__clkinv_1 U15206 ( .A(j202_soc_core_j22_cpu_rf_gpr[480]), 
        .Y(n19279) );
  sky130_fd_sc_hd__nor2_1 U15207 ( .A(n19959), .B(n19953), .Y(n21796) );
  sky130_fd_sc_hd__clkinv_1 U15208 ( .A(n20005), .Y(n20032) );
  sky130_fd_sc_hd__clkinv_1 U15209 ( .A(n16191), .Y(n20025) );
  sky130_fd_sc_hd__nor2_1 U15210 ( .A(n16598), .B(n16607), .Y(n20005) );
  sky130_fd_sc_hd__clkinv_1 U15211 ( .A(n22695), .Y(n22510) );
  sky130_fd_sc_hd__and2_0 U15212 ( .A(n11541), .B(n11536), .X(n20250) );
  sky130_fd_sc_hd__nor2_1 U15213 ( .A(n12929), .B(n20479), .Y(n20256) );
  sky130_fd_sc_hd__nand2_1 U15214 ( .A(n20277), .B(
        j202_soc_core_j22_cpu_regop_We__2_), .Y(n20248) );
  sky130_fd_sc_hd__clkinv_1 U15215 ( .A(j202_soc_core_j22_cpu_regop_We__1_), 
        .Y(n20275) );
  sky130_fd_sc_hd__clkinv_1 U15216 ( .A(n20616), .Y(n20707) );
  sky130_fd_sc_hd__nand2_1 U15217 ( .A(n16643), .B(
        j202_soc_core_j22_cpu_ma_M_MEM[0]), .Y(n22551) );
  sky130_fd_sc_hd__nor2_1 U15218 ( .A(j202_soc_core_j22_cpu_regop_We__3_), .B(
        n20506), .Y(n20277) );
  sky130_fd_sc_hd__clkinv_1 U15219 ( .A(j202_soc_core_j22_cpu_rf_gpr[486]), 
        .Y(n19057) );
  sky130_fd_sc_hd__clkinv_1 U15220 ( .A(j202_soc_core_j22_cpu_pc[6]), .Y(
        n19054) );
  sky130_fd_sc_hd__clkinv_1 U15221 ( .A(j202_soc_core_j22_cpu_rf_pr[2]), .Y(
        n16814) );
  sky130_fd_sc_hd__clkinv_1 U15222 ( .A(j202_soc_core_j22_cpu_rf_gbr[2]), .Y(
        n16813) );
  sky130_fd_sc_hd__clkinv_1 U15223 ( .A(j202_soc_core_j22_cpu_rf_gpr[482]), 
        .Y(n16815) );
  sky130_fd_sc_hd__clkinv_1 U15224 ( .A(j202_soc_core_j22_cpu_rf_vbr[20]), .Y(
        n19411) );
  sky130_fd_sc_hd__clkinv_1 U15225 ( .A(j202_soc_core_j22_cpu_rf_gpr[484]), 
        .Y(n17069) );
  sky130_fd_sc_hd__clkinv_1 U15226 ( .A(j202_soc_core_j22_cpu_pc[4]), .Y(
        n17066) );
  sky130_fd_sc_hd__clkinv_1 U15227 ( .A(j202_soc_core_j22_cpu_rf_gpr[485]), 
        .Y(n19185) );
  sky130_fd_sc_hd__clkinv_1 U15228 ( .A(j202_soc_core_j22_cpu_pc[5]), .Y(
        n19182) );
  sky130_fd_sc_hd__clkinv_1 U15229 ( .A(j202_soc_core_j22_cpu_rf_gpr[487]), 
        .Y(n16697) );
  sky130_fd_sc_hd__clkinv_1 U15230 ( .A(j202_soc_core_j22_cpu_pc[7]), .Y(
        n16694) );
  sky130_fd_sc_hd__clkinv_1 U15231 ( .A(j202_soc_core_j22_cpu_rf_gpr[483]), 
        .Y(n18916) );
  sky130_fd_sc_hd__clkinv_1 U15232 ( .A(n21137), .Y(n20638) );
  sky130_fd_sc_hd__clkinv_1 U15233 ( .A(j202_soc_core_j22_cpu_rf_gpr[488]), 
        .Y(n19206) );
  sky130_fd_sc_hd__clkinv_1 U15234 ( .A(j202_soc_core_j22_cpu_pc[8]), .Y(
        n19203) );
  sky130_fd_sc_hd__clkinv_1 U15235 ( .A(n20483), .Y(n20505) );
  sky130_fd_sc_hd__clkinv_1 U15236 ( .A(n17833), .Y(n17124) );
  sky130_fd_sc_hd__clkinv_1 U15237 ( .A(j202_soc_core_j22_cpu_rf_gpr[493]), 
        .Y(n19119) );
  sky130_fd_sc_hd__and2_0 U15238 ( .A(j202_soc_core_aquc_WE_), .B(
        j202_soc_core_aquc_CE__1_), .X(n22104) );
  sky130_fd_sc_hd__and2_0 U15239 ( .A(n17639), .B(n18360), .X(n18752) );
  sky130_fd_sc_hd__clkinv_1 U15240 ( .A(n16682), .Y(n21178) );
  sky130_fd_sc_hd__clkinv_1 U15241 ( .A(j202_soc_core_j22_cpu_rf_pr[14]), .Y(
        n18952) );
  sky130_fd_sc_hd__clkinv_1 U15242 ( .A(j202_soc_core_j22_cpu_pc[14]), .Y(
        n18953) );
  sky130_fd_sc_hd__and2_0 U15243 ( .A(n11537), .B(n11519), .X(n11183) );
  sky130_fd_sc_hd__nor2_1 U15244 ( .A(n20275), .B(n20248), .Y(n20309) );
  sky130_fd_sc_hd__clkinv_1 U15245 ( .A(n20256), .Y(n20306) );
  sky130_fd_sc_hd__a21oi_1 U15246 ( .A1(n20271), .A2(n20306), .B1(n24894), .Y(
        n20307) );
  sky130_fd_sc_hd__nand2_1 U15247 ( .A(n15219), .B(n12020), .Y(n14071) );
  sky130_fd_sc_hd__clkinv_1 U15248 ( .A(n18939), .Y(n19509) );
  sky130_fd_sc_hd__clkinv_1 U15249 ( .A(n18941), .Y(n18942) );
  sky130_fd_sc_hd__clkinv_1 U15250 ( .A(n18940), .Y(n18943) );
  sky130_fd_sc_hd__clkinv_1 U15251 ( .A(j202_soc_core_j22_cpu_rf_gpr[491]), 
        .Y(n18929) );
  sky130_fd_sc_hd__clkinv_1 U15252 ( .A(n20355), .Y(n21007) );
  sky130_fd_sc_hd__clkinv_1 U15253 ( .A(n22687), .Y(n22690) );
  sky130_fd_sc_hd__clkinv_1 U15254 ( .A(n22693), .Y(n22689) );
  sky130_fd_sc_hd__nand2_1 U15255 ( .A(n16858), .B(n16857), .Y(n19895) );
  sky130_fd_sc_hd__clkinv_1 U15256 ( .A(n20706), .Y(n16858) );
  sky130_fd_sc_hd__and2_0 U15257 ( .A(j202_soc_core_j22_cpu_ma_M_address[1]), 
        .B(n16860), .X(n19889) );
  sky130_fd_sc_hd__clkinv_1 U15258 ( .A(n21208), .Y(n19833) );
  sky130_fd_sc_hd__and2_0 U15259 ( .A(n18267), .B(n16977), .X(n18560) );
  sky130_fd_sc_hd__and2_0 U15260 ( .A(n14961), .B(n14394), .X(n14530) );
  sky130_fd_sc_hd__clkinv_1 U15261 ( .A(n21234), .Y(n21324) );
  sky130_fd_sc_hd__clkinv_1 U15262 ( .A(n25000), .Y(n23491) );
  sky130_fd_sc_hd__and2_0 U15263 ( .A(n20119), .B(n20111), .X(n23525) );
  sky130_fd_sc_hd__clkinv_1 U15264 ( .A(n23529), .Y(n23788) );
  sky130_fd_sc_hd__and2_0 U15265 ( .A(n23403), .B(n23564), .X(n22775) );
  sky130_fd_sc_hd__and2_0 U15266 ( .A(n20217), .B(j202_soc_core_qspi_wb_we), 
        .X(n23404) );
  sky130_fd_sc_hd__clkinv_1 U15267 ( .A(j202_soc_core_wbqspiflash_00_state[2]), 
        .Y(n24899) );
  sky130_fd_sc_hd__clkinv_1 U15268 ( .A(j202_soc_core_wbqspiflash_00_state[4]), 
        .Y(n23513) );
  sky130_fd_sc_hd__clkinv_1 U15269 ( .A(n23754), .Y(n25099) );
  sky130_fd_sc_hd__clkinv_1 U15270 ( .A(n14395), .Y(n14092) );
  sky130_fd_sc_hd__clkinv_1 U15271 ( .A(n22575), .Y(n21048) );
  sky130_fd_sc_hd__and2_0 U15272 ( .A(n14185), .B(n14184), .X(n14187) );
  sky130_fd_sc_hd__clkinv_1 U15273 ( .A(n18761), .Y(n14906) );
  sky130_fd_sc_hd__clkinv_1 U15274 ( .A(n17123), .Y(n17834) );
  sky130_fd_sc_hd__clkinv_1 U15275 ( .A(n17122), .Y(n19045) );
  sky130_fd_sc_hd__nand2_1 U15276 ( .A(n11558), .B(n12940), .Y(n14079) );
  sky130_fd_sc_hd__nand2_1 U15277 ( .A(n11558), .B(n15212), .Y(n14073) );
  sky130_fd_sc_hd__nand2_1 U15278 ( .A(n11558), .B(n11557), .Y(n14075) );
  sky130_fd_sc_hd__clkinv_1 U15279 ( .A(j202_soc_core_j22_cpu_regop_Rb__1_), 
        .Y(n14086) );
  sky130_fd_sc_hd__clkinv_1 U15280 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[2]), .Y(n18277) );
  sky130_fd_sc_hd__and2_0 U15281 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .B(j202_soc_core_bootrom_00_address_w[7]), .X(n17606) );
  sky130_fd_sc_hd__and2_0 U15282 ( .A(n11315), .B(
        j202_soc_core_memory0_ram_dout0_sel[5]), .X(n18735) );
  sky130_fd_sc_hd__and2_0 U15283 ( .A(n17481), .B(n17846), .X(n17674) );
  sky130_fd_sc_hd__clkinv_1 U15284 ( .A(n18513), .Y(n18783) );
  sky130_fd_sc_hd__nand3_1 U15285 ( .A(n11206), .B(n11242), .C(n11205), .Y(
        n18212) );
  sky130_fd_sc_hd__and2_0 U15286 ( .A(n11204), .B(n11203), .X(n11205) );
  sky130_fd_sc_hd__clkinv_1 U15287 ( .A(n18792), .Y(n18651) );
  sky130_fd_sc_hd__clkinv_1 U15288 ( .A(n18212), .Y(n14668) );
  sky130_fd_sc_hd__clkinv_1 U15289 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .Y(n13210) );
  sky130_fd_sc_hd__clkinv_1 U15290 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .Y(n13231) );
  sky130_fd_sc_hd__clkinv_1 U15291 ( .A(n17639), .Y(n18736) );
  sky130_fd_sc_hd__and2_0 U15292 ( .A(n18446), .B(n15020), .X(n15022) );
  sky130_fd_sc_hd__and2_0 U15293 ( .A(n17470), .B(n17768), .X(n17528) );
  sky130_fd_sc_hd__clkinv_1 U15294 ( .A(n17812), .Y(n18445) );
  sky130_fd_sc_hd__clkinv_1 U15295 ( .A(n17606), .Y(n18423) );
  sky130_fd_sc_hd__and2_0 U15296 ( .A(n25159), .B(n17711), .X(n17427) );
  sky130_fd_sc_hd__clkinv_1 U15297 ( .A(n17543), .Y(n18437) );
  sky130_fd_sc_hd__clkinv_1 U15298 ( .A(j202_soc_core_j22_cpu_rf_gpr[492]), 
        .Y(n17055) );
  sky130_fd_sc_hd__clkinv_1 U15299 ( .A(n22551), .Y(n22530) );
  sky130_fd_sc_hd__clkinv_1 U15300 ( .A(n20774), .Y(n21443) );
  sky130_fd_sc_hd__clkinv_1 U15301 ( .A(j202_soc_core_j22_cpu_rf_gpr[490]), 
        .Y(n16879) );
  sky130_fd_sc_hd__clkinv_1 U15302 ( .A(n16679), .Y(n19725) );
  sky130_fd_sc_hd__clkinv_1 U15304 ( .A(n24074), .Y(n24079) );
  sky130_fd_sc_hd__clkinv_1 U15305 ( .A(n19931), .Y(n20043) );
  sky130_fd_sc_hd__clkinv_1 U15306 ( .A(j202_soc_core_j22_cpu_rf_gpr[495]), 
        .Y(n15222) );
  sky130_fd_sc_hd__clkinv_1 U15307 ( .A(n19983), .Y(n19842) );
  sky130_fd_sc_hd__clkinv_1 U15308 ( .A(j202_soc_core_j22_cpu_regop_Rs__1_), 
        .Y(n19969) );
  sky130_fd_sc_hd__clkinv_1 U15309 ( .A(n15076), .Y(n17828) );
  sky130_fd_sc_hd__nor2_1 U15310 ( .A(n12908), .B(n12986), .Y(n21624) );
  sky130_fd_sc_hd__nand3_1 U15311 ( .A(n19078), .B(n13092), .C(n13096), .Y(
        n13095) );
  sky130_fd_sc_hd__and2_0 U15312 ( .A(j202_soc_core_j22_cpu_ifetchl), .B(
        n21647), .X(n11182) );
  sky130_fd_sc_hd__clkinv_1 U15313 ( .A(n24471), .Y(n24446) );
  sky130_fd_sc_hd__clkinv_1 U15314 ( .A(n23590), .Y(n23593) );
  sky130_fd_sc_hd__clkinv_1 U15315 ( .A(n23734), .Y(n23740) );
  sky130_fd_sc_hd__clkinv_1 U15316 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[13]), .Y(n24975) );
  sky130_fd_sc_hd__clkinv_1 U15317 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[12]), .Y(n24967) );
  sky130_fd_sc_hd__clkinv_1 U15318 ( .A(j202_soc_core_qspi_wb_addr[15]), .Y(
        n24986) );
  sky130_fd_sc_hd__clkinv_1 U15319 ( .A(n25055), .Y(n25081) );
  sky130_fd_sc_hd__clkinv_1 U15320 ( .A(n23612), .Y(n23747) );
  sky130_fd_sc_hd__and2_0 U15321 ( .A(n23747), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[2]), .X(n25435) );
  sky130_fd_sc_hd__clkinv_1 U15322 ( .A(n23742), .Y(n23694) );
  sky130_fd_sc_hd__and2_0 U15323 ( .A(n23199), .B(n23202), .X(n23206) );
  sky130_fd_sc_hd__clkinv_1 U15324 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[0]), 
        .Y(n25123) );
  sky130_fd_sc_hd__clkinv_1 U15325 ( .A(j202_soc_core_intc_core_00_rg_ipr[83]), 
        .Y(n24682) );
  sky130_fd_sc_hd__clkinv_1 U15326 ( .A(n25295), .Y(n24440) );
  sky130_fd_sc_hd__clkinv_1 U15327 ( .A(j202_soc_core_bldc_core_00_pwm_duty[7]), .Y(n25126) );
  sky130_fd_sc_hd__clkinv_1 U15328 ( .A(n21970), .Y(n20878) );
  sky130_fd_sc_hd__and2_0 U15329 ( .A(j202_soc_core_cmt_core_00_cnt0[4]), .B(
        n23058), .X(n23060) );
  sky130_fd_sc_hd__clkinv_1 U15330 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[9]), .Y(n25153) );
  sky130_fd_sc_hd__clkinv_1 U15331 ( .A(n25293), .Y(n24436) );
  sky130_fd_sc_hd__clkinv_1 U15332 ( .A(j202_soc_core_bldc_core_00_pwm_duty[5]), .Y(n25135) );
  sky130_fd_sc_hd__clkinv_1 U15333 ( .A(n25288), .Y(n24475) );
  sky130_fd_sc_hd__clkinv_1 U15334 ( .A(n17824), .Y(n17826) );
  sky130_fd_sc_hd__clkinv_1 U15335 ( .A(n24746), .Y(n24766) );
  sky130_fd_sc_hd__clkinv_1 U15336 ( .A(n24681), .Y(n24771) );
  sky130_fd_sc_hd__clkinv_1 U15337 ( .A(n24744), .Y(n24770) );
  sky130_fd_sc_hd__clkinv_1 U15338 ( .A(n24498), .Y(n20084) );
  sky130_fd_sc_hd__clkinv_1 U15339 ( .A(n24289), .Y(n20497) );
  sky130_fd_sc_hd__clkinv_1 U15340 ( .A(n24492), .Y(n20092) );
  sky130_fd_sc_hd__clkinv_1 U15341 ( .A(n24291), .Y(n20115) );
  sky130_fd_sc_hd__clkinv_1 U15342 ( .A(n24548), .Y(n20082) );
  sky130_fd_sc_hd__clkinv_1 U15343 ( .A(j202_soc_core_intc_core_00_rg_ipr[37]), 
        .Y(n24559) );
  sky130_fd_sc_hd__clkinv_1 U15344 ( .A(n24491), .Y(n24350) );
  sky130_fd_sc_hd__clkinv_1 U15345 ( .A(n24497), .Y(n24294) );
  sky130_fd_sc_hd__clkinv_1 U15346 ( .A(j202_soc_core_intc_core_00_rg_ipr[76]), 
        .Y(n24626) );
  sky130_fd_sc_hd__clkinv_1 U15347 ( .A(j202_soc_core_intc_core_00_rg_ipr[66]), 
        .Y(n24521) );
  sky130_fd_sc_hd__clkinv_1 U15348 ( .A(j202_soc_core_intc_core_00_rg_ipr[24]), 
        .Y(n24718) );
  sky130_fd_sc_hd__clkinv_1 U15349 ( .A(n25296), .Y(n24400) );
  sky130_fd_sc_hd__clkinv_1 U15350 ( .A(n25285), .Y(n24438) );
  sky130_fd_sc_hd__clkinv_1 U15351 ( .A(n24495), .Y(n24408) );
  sky130_fd_sc_hd__clkinv_1 U15352 ( .A(n25297), .Y(n24488) );
  sky130_fd_sc_hd__clkinv_1 U15353 ( .A(n25298), .Y(n24485) );
  sky130_fd_sc_hd__clkinv_1 U15354 ( .A(n25294), .Y(n24483) );
  sky130_fd_sc_hd__clkinv_1 U15355 ( .A(n25287), .Y(n24479) );
  sky130_fd_sc_hd__clkinv_1 U15356 ( .A(n25286), .Y(n24477) );
  sky130_fd_sc_hd__clkinv_1 U15357 ( .A(j202_soc_core_uart_div0[3]), .Y(n24807) );
  sky130_fd_sc_hd__clkinv_1 U15358 ( .A(j202_soc_core_uart_div0[4]), .Y(n24804) );
  sky130_fd_sc_hd__clkinv_1 U15359 ( .A(j202_soc_core_uart_div0[7]), .Y(n24805) );
  sky130_fd_sc_hd__clkinv_1 U15360 ( .A(j202_soc_core_uart_div0[2]), .Y(n24815) );
  sky130_fd_sc_hd__clkinv_1 U15361 ( .A(n18837), .Y(n18839) );
  sky130_fd_sc_hd__clkinv_1 U15362 ( .A(n20689), .Y(n22564) );
  sky130_fd_sc_hd__clkinv_1 U15363 ( .A(j202_soc_core_ahb2apb_01_state[2]), 
        .Y(n21224) );
  sky130_fd_sc_hd__clkinv_1 U15364 ( .A(n23872), .Y(n24061) );
  sky130_fd_sc_hd__clkinv_1 U15365 ( .A(j202_soc_core_j22_cpu_rf_vbr[28]), .Y(
        n19786) );
  sky130_fd_sc_hd__clkinv_1 U15366 ( .A(n18817), .Y(n18819) );
  sky130_fd_sc_hd__a21boi_0 U15367 ( .A1(n21700), .A2(n20030), .B1_N(n17041), 
        .Y(n22095) );
  sky130_fd_sc_hd__clkinv_1 U15368 ( .A(n20720), .Y(n22560) );
  sky130_fd_sc_hd__nand3_1 U15369 ( .A(n20428), .B(n20427), .C(n20426), .Y(
        n22017) );
  sky130_fd_sc_hd__clkinv_1 U15370 ( .A(n21152), .Y(n22562) );
  sky130_fd_sc_hd__or3b_2 U15371 ( .A(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[0]), .B(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[2]), .C_N(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[1]), .X(n20495) );
  sky130_fd_sc_hd__clkinv_1 U15372 ( .A(j202_soc_core_bldc_core_00_pwm_duty[0]), .Y(n25128) );
  sky130_fd_sc_hd__clkinv_1 U15373 ( .A(j202_soc_core_bldc_core_00_pwm_duty[6]), .Y(n25136) );
  sky130_fd_sc_hd__clkinv_1 U15374 ( .A(j202_soc_core_bldc_core_00_pwm_duty[9]), .Y(n25139) );
  sky130_fd_sc_hd__clkinv_1 U15375 ( .A(n25189), .Y(n25193) );
  sky130_fd_sc_hd__and2_0 U15376 ( .A(j202_soc_core_aquc_STB_), .B(
        j202_soc_core_aquc_CE__0_), .X(n21228) );
  sky130_fd_sc_hd__clkinv_1 U15377 ( .A(j202_soc_core_qspi_wb_addr[8]), .Y(
        n24939) );
  sky130_fd_sc_hd__clkinv_1 U15378 ( .A(n22171), .Y(n21929) );
  sky130_fd_sc_hd__clkinv_1 U15379 ( .A(n19721), .Y(n19723) );
  sky130_fd_sc_hd__clkinv_1 U15380 ( .A(n20721), .Y(n22558) );
  sky130_fd_sc_hd__clkinv_1 U15381 ( .A(n19917), .Y(n20064) );
  sky130_fd_sc_hd__clkinv_1 U15382 ( .A(n21782), .Y(n20952) );
  sky130_fd_sc_hd__clkinv_1 U15383 ( .A(n23757), .Y(n23760) );
  sky130_fd_sc_hd__clkinv_1 U15384 ( .A(n25108), .Y(n23787) );
  sky130_fd_sc_hd__clkinv_1 U15385 ( .A(n23509), .Y(n20120) );
  sky130_fd_sc_hd__clkinv_1 U15386 ( .A(n24954), .Y(n24960) );
  sky130_fd_sc_hd__clkinv_1 U15387 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .Y(n24901) );
  sky130_fd_sc_hd__clkinv_1 U15388 ( .A(n25009), .Y(n25041) );
  sky130_fd_sc_hd__clkinv_1 U15389 ( .A(j202_soc_core_qspi_wb_we), .Y(n23494)
         );
  sky130_fd_sc_hd__clkinv_1 U15390 ( .A(n23738), .Y(n23689) );
  sky130_fd_sc_hd__clkinv_1 U15391 ( .A(n23435), .Y(n23384) );
  sky130_fd_sc_hd__clkinv_1 U15392 ( .A(j202_soc_core_j22_cpu_rf_vbr[29]), .Y(
        n19611) );
  sky130_fd_sc_hd__clkinv_1 U15393 ( .A(j202_soc_core_j22_cpu_rf_vbr[26]), .Y(
        n19576) );
  sky130_fd_sc_hd__a21boi_0 U15394 ( .A1(n19376), .A2(n20040), .B1_N(n19375), 
        .Y(n21833) );
  sky130_fd_sc_hd__clkinv_1 U15395 ( .A(j202_soc_core_j22_cpu_rf_vbr[22]), .Y(
        n19538) );
  sky130_fd_sc_hd__a21boi_0 U15396 ( .A1(n19451), .A2(n20040), .B1_N(n19450), 
        .Y(n21780) );
  sky130_fd_sc_hd__clkinv_1 U15397 ( .A(n22246), .Y(n22225) );
  sky130_fd_sc_hd__o31ai_1 U15398 ( .A1(n22556), .A2(n22145), .A3(n22150), 
        .B1(n21682), .Y(n22131) );
  sky130_fd_sc_hd__a31o_1 U15399 ( .A1(n22143), .A2(n21678), .A3(n21677), .B1(
        n22126), .X(n22132) );
  sky130_fd_sc_hd__clkinv_1 U15400 ( .A(n21675), .Y(n21677) );
  sky130_fd_sc_hd__clkinv_1 U15401 ( .A(j202_soc_core_j22_cpu_ml_bufa[15]), 
        .Y(n22229) );
  sky130_fd_sc_hd__clkinv_1 U15402 ( .A(n22195), .Y(n22206) );
  sky130_fd_sc_hd__nand3_1 U15403 ( .A(n20663), .B(n20662), .C(n20661), .Y(
        n22269) );
  sky130_fd_sc_hd__clkinv_1 U15404 ( .A(n19511), .Y(n19513) );
  sky130_fd_sc_hd__clkinv_1 U15405 ( .A(n20935), .Y(n22557) );
  sky130_fd_sc_hd__clkinv_1 U15406 ( .A(n21925), .Y(n22173) );
  sky130_fd_sc_hd__a21boi_0 U15407 ( .A1(n22147), .A2(n20088), .B1_N(n23347), 
        .Y(n23345) );
  sky130_fd_sc_hd__clkinv_1 U15408 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]), .Y(n20086) );
  sky130_fd_sc_hd__clkinv_1 U15409 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .Y(n20087) );
  sky130_fd_sc_hd__clkinv_1 U15410 ( .A(n23318), .Y(n22513) );
  sky130_fd_sc_hd__nand3_1 U15411 ( .A(n21181), .B(n21180), .C(n21179), .Y(
        n21874) );
  sky130_fd_sc_hd__clkinv_1 U15412 ( .A(n21858), .Y(n20591) );
  sky130_fd_sc_hd__o21a_1 U15413 ( .A1(n20638), .A2(n20637), .B1(n20636), .X(
        n22072) );
  sky130_fd_sc_hd__clkinv_1 U15414 ( .A(n22346), .Y(n20615) );
  sky130_fd_sc_hd__clkinv_1 U15415 ( .A(n23330), .Y(n22609) );
  sky130_fd_sc_hd__clkinv_1 U15416 ( .A(n21947), .Y(n21951) );
  sky130_fd_sc_hd__clkinv_1 U15417 ( .A(n21752), .Y(n20799) );
  sky130_fd_sc_hd__clkinv_1 U15418 ( .A(n22111), .Y(n20824) );
  sky130_fd_sc_hd__clkinv_1 U15419 ( .A(n22149), .Y(n22186) );
  sky130_fd_sc_hd__clkinv_1 U15420 ( .A(n22187), .Y(n22153) );
  sky130_fd_sc_hd__nor2_1 U15421 ( .A(n22148), .B(n22274), .Y(n23343) );
  sky130_fd_sc_hd__nand2_1 U15422 ( .A(n23297), .B(n23296), .Y(n23339) );
  sky130_fd_sc_hd__a21boi_0 U15423 ( .A1(n21696), .A2(n20030), .B1_N(n19106), 
        .Y(n22207) );
  sky130_fd_sc_hd__clkinv_1 U15424 ( .A(n20648), .Y(n22561) );
  sky130_fd_sc_hd__clkinv_1 U15425 ( .A(n20699), .Y(n22559) );
  sky130_fd_sc_hd__clkinv_1 U15426 ( .A(n19173), .Y(n22580) );
  sky130_fd_sc_hd__clkinv_1 U15427 ( .A(j202_soc_core_j22_cpu_ml_bufa[3]), .Y(
        n22002) );
  sky130_fd_sc_hd__clkinv_1 U15428 ( .A(n22583), .Y(n22488) );
  sky130_fd_sc_hd__clkinv_1 U15429 ( .A(j202_soc_core_j22_cpu_ml_bufa[0]), .Y(
        n22247) );
  sky130_fd_sc_hd__and2_0 U15430 ( .A(n22135), .B(n20100), .X(n22143) );
  sky130_fd_sc_hd__nand2_1 U15431 ( .A(n16591), .B(n16590), .Y(n22246) );
  sky130_fd_sc_hd__clkinv_1 U15432 ( .A(j202_soc_core_j22_cpu_ml_bufa[6]), .Y(
        n22049) );
  sky130_fd_sc_hd__nand2_1 U15433 ( .A(n22221), .B(n22190), .Y(n22245) );
  sky130_fd_sc_hd__clkinv_1 U15434 ( .A(n20007), .Y(n22204) );
  sky130_fd_sc_hd__clkinv_1 U15435 ( .A(j202_soc_core_j22_cpu_macop_MAC_[2]), 
        .Y(n21680) );
  sky130_fd_sc_hd__clkinv_1 U15436 ( .A(j202_soc_core_j22_cpu_macop_MAC_[0]), 
        .Y(n22125) );
  sky130_fd_sc_hd__nand3_1 U15437 ( .A(n19904), .B(n19903), .C(n19902), .Y(
        n22122) );
  sky130_fd_sc_hd__clkinv_1 U15438 ( .A(n22122), .Y(n20757) );
  sky130_fd_sc_hd__a21oi_1 U15439 ( .A1(n20704), .A2(n21137), .B1(n20703), .Y(
        n22319) );
  sky130_fd_sc_hd__clkinv_1 U15440 ( .A(n21819), .Y(n20927) );
  sky130_fd_sc_hd__nand2_1 U15441 ( .A(n19083), .B(n18948), .Y(n19736) );
  sky130_fd_sc_hd__clkinv_1 U15442 ( .A(n19731), .Y(n19657) );
  sky130_fd_sc_hd__clkinv_1 U15443 ( .A(n19243), .Y(n19245) );
  sky130_fd_sc_hd__and2_0 U15444 ( .A(j202_soc_core_uart_WRTXD1), .B(n23254), 
        .X(n25201) );
  sky130_fd_sc_hd__clkinv_1 U15445 ( .A(n25379), .Y(n22817) );
  sky130_fd_sc_hd__clkinv_1 U15446 ( .A(n22259), .Y(n22267) );
  sky130_fd_sc_hd__clkinv_1 U15447 ( .A(n21199), .Y(n21102) );
  sky130_fd_sc_hd__clkinv_1 U15448 ( .A(n21198), .Y(n21199) );
  sky130_fd_sc_hd__nand2_1 U15449 ( .A(n23239), .B(n20253), .Y(n21190) );
  sky130_fd_sc_hd__clkinv_1 U15450 ( .A(n21190), .Y(n21191) );
  sky130_fd_sc_hd__and2_0 U15451 ( .A(n20546), .B(n22530), .X(n20382) );
  sky130_fd_sc_hd__nor2_1 U15452 ( .A(n20278), .B(n20483), .Y(n22367) );
  sky130_fd_sc_hd__nor2_1 U15453 ( .A(n22345), .B(n22367), .Y(n22369) );
  sky130_fd_sc_hd__nand3_1 U15454 ( .A(n18911), .B(n18910), .C(n18909), .Y(
        n22006) );
  sky130_fd_sc_hd__inv_2 U15455 ( .A(n23348), .Y(n22358) );
  sky130_fd_sc_hd__clkinv_1 U15456 ( .A(n22366), .Y(n22344) );
  sky130_fd_sc_hd__clkinv_1 U15457 ( .A(j202_soc_core_j22_cpu_regop_We__0_), 
        .Y(n20506) );
  sky130_fd_sc_hd__nand3_1 U15458 ( .A(n16874), .B(n16873), .C(n16872), .Y(
        n22258) );
  sky130_fd_sc_hd__clkinv_1 U15459 ( .A(n22248), .Y(n22251) );
  sky130_fd_sc_hd__clkinv_1 U15460 ( .A(n22547), .Y(n22486) );
  sky130_fd_sc_hd__clkinv_1 U15461 ( .A(n22258), .Y(n20520) );
  sky130_fd_sc_hd__clkinv_1 U15462 ( .A(n22013), .Y(n22519) );
  sky130_fd_sc_hd__clkinv_1 U15463 ( .A(n22006), .Y(n20519) );
  sky130_fd_sc_hd__clkinv_1 U15464 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__0_), 
        .Y(n20484) );
  sky130_fd_sc_hd__nand3_1 U15465 ( .A(n20505), .B(
        j202_soc_core_j22_cpu_regop_We__3_), .C(n20506), .Y(n21196) );
  sky130_fd_sc_hd__nand2_1 U15466 ( .A(n21196), .B(n21217), .Y(n21197) );
  sky130_fd_sc_hd__clkinv_1 U15467 ( .A(j202_soc_core_j22_cpu_opst[0]), .Y(
        n22418) );
  sky130_fd_sc_hd__clkinv_1 U15468 ( .A(n19500), .Y(n19907) );
  sky130_fd_sc_hd__clkinv_1 U15469 ( .A(j202_soc_core_j22_cpu_ml_bufa[18]), 
        .Y(n19452) );
  sky130_fd_sc_hd__clkinv_1 U15470 ( .A(j202_soc_core_j22_cpu_rf_vbr[18]), .Y(
        n19454) );
  sky130_fd_sc_hd__clkinv_1 U15471 ( .A(j202_soc_core_j22_cpu_ml_bufa[21]), 
        .Y(n19400) );
  sky130_fd_sc_hd__clkinv_1 U15472 ( .A(j202_soc_core_j22_cpu_rf_vbr[21]), .Y(
        n19402) );
  sky130_fd_sc_hd__clkinv_1 U15473 ( .A(j202_soc_core_j22_cpu_rf_vbr[23]), .Y(
        n19380) );
  sky130_fd_sc_hd__clkinv_1 U15474 ( .A(n23234), .Y(n23237) );
  sky130_fd_sc_hd__clkinv_1 U15475 ( .A(j202_soc_core_j22_cpu_memop_MEM__0_), 
        .Y(n23240) );
  sky130_fd_sc_hd__clkinv_1 U15476 ( .A(j202_soc_core_j22_cpu_memop_MEM__3_), 
        .Y(n23245) );
  sky130_fd_sc_hd__clkinv_1 U15477 ( .A(n22792), .Y(n22793) );
  sky130_fd_sc_hd__clkinv_1 U15478 ( .A(n25213), .Y(n25212) );
  sky130_fd_sc_hd__clkinv_1 U15479 ( .A(n22010), .Y(n22011) );
  sky130_fd_sc_hd__nand3_1 U15480 ( .A(n20405), .B(n20404), .C(n20403), .Y(
        n21980) );
  sky130_fd_sc_hd__nand3_1 U15481 ( .A(n20381), .B(n20380), .C(n20379), .Y(
        n22079) );
  sky130_fd_sc_hd__clkinv_1 U15482 ( .A(n21236), .Y(n21996) );
  sky130_fd_sc_hd__and2_0 U15483 ( .A(n19691), .B(n19286), .X(n19719) );
  sky130_fd_sc_hd__nand3_1 U15484 ( .A(n20505), .B(
        j202_soc_core_j22_cpu_regop_We__0_), .C(
        j202_soc_core_j22_cpu_regop_We__3_), .Y(n21236) );
  sky130_fd_sc_hd__clkinv_1 U15485 ( .A(n22483), .Y(n22647) );
  sky130_fd_sc_hd__clkinv_1 U15486 ( .A(n25228), .Y(n25227) );
  sky130_fd_sc_hd__clkinv_1 U15487 ( .A(n25230), .Y(n25229) );
  sky130_fd_sc_hd__clkinv_1 U15488 ( .A(n25335), .Y(n22822) );
  sky130_fd_sc_hd__clkinv_1 U15489 ( .A(n17125), .Y(n17127) );
  sky130_fd_sc_hd__nand3_1 U15490 ( .A(n19178), .B(n19177), .C(n19176), .Y(
        n22033) );
  sky130_fd_sc_hd__nand3_1 U15491 ( .A(n19151), .B(n19150), .C(n19149), .Y(
        n22555) );
  sky130_fd_sc_hd__clkinv_1 U15492 ( .A(j202_soc_core_uart_div1[4]), .Y(n24793) );
  sky130_fd_sc_hd__clkinv_1 U15493 ( .A(j202_soc_core_uart_div1[3]), .Y(n24790) );
  sky130_fd_sc_hd__clkinv_1 U15494 ( .A(j202_soc_core_uart_div1[0]), .Y(n24787) );
  sky130_fd_sc_hd__clkinv_1 U15495 ( .A(j202_soc_core_uart_div1[2]), .Y(n24797) );
  sky130_fd_sc_hd__and2_0 U15496 ( .A(n21467), .B(n21466), .X(n22402) );
  sky130_fd_sc_hd__clkinv_1 U15497 ( .A(n19072), .Y(n19074) );
  sky130_fd_sc_hd__clkinv_1 U15498 ( .A(n25336), .Y(n22820) );
  sky130_fd_sc_hd__clkinv_1 U15499 ( .A(n19040), .Y(n19042) );
  sky130_fd_sc_hd__clkinv_1 U15500 ( .A(n20530), .Y(n22612) );
  sky130_fd_sc_hd__clkinv_1 U15501 ( .A(n25337), .Y(n22818) );
  sky130_fd_sc_hd__nand3_1 U15502 ( .A(n19050), .B(n19049), .C(n19048), .Y(
        n21850) );
  sky130_fd_sc_hd__a21boi_0 U15503 ( .A1(n19039), .A2(n20530), .B1_N(n19038), 
        .Y(n19049) );
  sky130_fd_sc_hd__clkinv_1 U15504 ( .A(n22286), .Y(n20545) );
  sky130_fd_sc_hd__and2_0 U15505 ( .A(n22974), .B(n22973), .X(n23023) );
  sky130_fd_sc_hd__clkinv_1 U15506 ( .A(n23209), .Y(n23217) );
  sky130_fd_sc_hd__clkinv_1 U15507 ( .A(n23202), .Y(n23192) );
  sky130_fd_sc_hd__clkinv_1 U15508 ( .A(n23198), .Y(n23196) );
  sky130_fd_sc_hd__clkinv_1 U15509 ( .A(n22725), .Y(n22723) );
  sky130_fd_sc_hd__clkinv_1 U15510 ( .A(n21613), .Y(n22720) );
  sky130_fd_sc_hd__clkinv_1 U15511 ( .A(n18805), .Y(n18807) );
  sky130_fd_sc_hd__clkinv_1 U15512 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]), .Y(n25052) );
  sky130_fd_sc_hd__clkinv_1 U15513 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .Y(n23571) );
  sky130_fd_sc_hd__clkinv_1 U15514 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .Y(n23569) );
  sky130_fd_sc_hd__clkinv_1 U15515 ( .A(n25492), .Y(n20219) );
  sky130_fd_sc_hd__nand3_1 U15516 ( .A(n19078), .B(
        j202_soc_core_j22_cpu_memop_Ma__1_), .C(
        j202_soc_core_j22_cpu_memop_Ma__0_), .Y(n14919) );
  sky130_fd_sc_hd__clkinv_1 U15517 ( .A(n19734), .Y(n19517) );
  sky130_fd_sc_hd__clkinv_1 U15518 ( .A(n18481), .Y(n18483) );
  sky130_fd_sc_hd__clkinv_1 U15519 ( .A(n19078), .Y(n19732) );
  sky130_fd_sc_hd__clkinv_1 U15520 ( .A(j202_soc_core_ahb2apb_01_state[0]), 
        .Y(n20076) );
  sky130_fd_sc_hd__clkinv_1 U15521 ( .A(n25240), .Y(n25239) );
  sky130_fd_sc_hd__clkinv_1 U15522 ( .A(j202_soc_core_ahb2apb_00_state[2]), 
        .Y(n22768) );
  sky130_fd_sc_hd__clkinv_1 U15523 ( .A(j202_soc_core_ahb2apb_00_state[1]), 
        .Y(n22767) );
  sky130_fd_sc_hd__nand3_1 U15524 ( .A(n21249), .B(n21248), .C(n21247), .Y(
        n22824) );
  sky130_fd_sc_hd__clkinv_1 U15525 ( .A(n23610), .Y(n20116) );
  sky130_fd_sc_hd__and2_0 U15526 ( .A(n21234), .B(n23731), .X(n22886) );
  sky130_fd_sc_hd__and2_0 U15527 ( .A(n23591), .B(n23612), .X(n23598) );
  sky130_fd_sc_hd__nand3_1 U15528 ( .A(j202_soc_core_wbqspiflash_00_w_qspi_sck), .B(n23592), .C(n25731), .Y(n23731) );
  sky130_fd_sc_hd__clkinv_1 U15529 ( .A(n22862), .Y(n22880) );
  sky130_fd_sc_hd__clkinv_1 U15530 ( .A(j202_soc_core_wbqspiflash_00_state[1]), 
        .Y(n22847) );
  sky130_fd_sc_hd__and2_0 U15531 ( .A(n25024), .B(
        j202_soc_core_ahb2wbqspi_00_stb_o), .X(n23461) );
  sky130_fd_sc_hd__clkinv_1 U15532 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]), .Y(n25089) );
  sky130_fd_sc_hd__clkinv_1 U15533 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[0]), .Y(n23697) );
  sky130_fd_sc_hd__clkinv_1 U15534 ( .A(n23500), .Y(n25027) );
  sky130_fd_sc_hd__clkinv_1 U15535 ( .A(j202_soc_core_wbqspiflash_00_spi_wr), 
        .Y(n23396) );
  sky130_fd_sc_hd__and2_0 U15536 ( .A(n23289), .B(n23396), .X(n23290) );
  sky130_fd_sc_hd__clkinv_1 U15537 ( .A(n25042), .Y(n25046) );
  sky130_fd_sc_hd__clkinv_1 U15538 ( .A(j202_soc_core_wbqspiflash_00_state[3]), 
        .Y(n23395) );
  sky130_fd_sc_hd__clkinv_1 U15539 ( .A(n23364), .Y(n23523) );
  sky130_fd_sc_hd__clkinv_1 U15540 ( .A(j202_soc_core_qspi_wb_cyc), .Y(n25111)
         );
  sky130_fd_sc_hd__clkinv_1 U15541 ( .A(io_in[14]), .Y(n14971) );
  sky130_fd_sc_hd__clkinv_1 U15542 ( .A(n23340), .Y(n22603) );
  sky130_fd_sc_hd__nor4_1 U15543 ( .A(n14173), .B(n14172), .C(n14171), .D(
        n14170), .Y(n22542) );
  sky130_fd_sc_hd__nor2_1 U15544 ( .A(n11333), .B(j202_soc_core_j22_cpu_pc[1]), 
        .Y(n19089) );
  sky130_fd_sc_hd__and3_1 U15545 ( .A(n11420), .B(j202_soc_core_j22_cpu_pc[1]), 
        .C(n11419), .X(n19087) );
  sky130_fd_sc_hd__clkinv_1 U15546 ( .A(n25334), .Y(n22823) );
  sky130_fd_sc_hd__nor2_1 U15547 ( .A(n12913), .B(n21329), .Y(n23229) );
  sky130_fd_sc_hd__clkinv_1 U15548 ( .A(n18664), .Y(n18771) );
  sky130_fd_sc_hd__clkinv_1 U15549 ( .A(n18655), .Y(n18779) );
  sky130_fd_sc_hd__nor2_1 U15550 ( .A(n11246), .B(n11410), .Y(n18727) );
  sky130_fd_sc_hd__nor2_1 U15551 ( .A(n18288), .B(n18306), .Y(n18725) );
  sky130_fd_sc_hd__nand2_1 U15552 ( .A(n11288), .B(n11287), .Y(n18761) );
  sky130_fd_sc_hd__clkinv_1 U15553 ( .A(n18722), .Y(n18605) );
  sky130_fd_sc_hd__nor2_1 U15554 ( .A(n11268), .B(n18212), .Y(n18798) );
  sky130_fd_sc_hd__nand3_1 U15555 ( .A(n14668), .B(n13210), .C(n13231), .Y(
        n18722) );
  sky130_fd_sc_hd__nor2_1 U15556 ( .A(n18282), .B(n17717), .Y(n18629) );
  sky130_fd_sc_hd__clkinv_1 U15558 ( .A(n17609), .Y(n18720) );
  sky130_fd_sc_hd__clkinv_1 U15559 ( .A(n18798), .Y(n18552) );
  sky130_fd_sc_hd__clkinv_1 U15560 ( .A(n18610), .Y(n18666) );
  sky130_fd_sc_hd__clkinv_1 U15561 ( .A(n21368), .Y(n21371) );
  sky130_fd_sc_hd__clkinv_1 U15562 ( .A(n24493), .Y(n20096) );
  sky130_fd_sc_hd__nand2_1 U15563 ( .A(n16612), .B(
        j202_soc_core_j22_cpu_memop_MEM__1_), .Y(n20067) );
  sky130_fd_sc_hd__nand2_1 U15564 ( .A(n21622), .B(n21621), .Y(n22753) );
  sky130_fd_sc_hd__clkinv_1 U15565 ( .A(n25258), .Y(n22762) );
  sky130_fd_sc_hd__clkinv_1 U15566 ( .A(n24879), .Y(n22401) );
  sky130_fd_sc_hd__clkinv_1 U15567 ( .A(n19726), .Y(n16680) );
  sky130_fd_sc_hd__clkinv_1 U15568 ( .A(n22496), .Y(n22645) );
  sky130_fd_sc_hd__clkinv_1 U15569 ( .A(n25338), .Y(n22819) );
  sky130_fd_sc_hd__a21oi_1 U15570 ( .A1(n21041), .A2(n21040), .B1(n24863), .Y(
        n22283) );
  sky130_fd_sc_hd__clkinv_1 U15571 ( .A(n20067), .Y(n20019) );
  sky130_fd_sc_hd__and2_0 U15572 ( .A(n19464), .B(n16704), .X(n19651) );
  sky130_fd_sc_hd__clkinv_1 U15573 ( .A(n15073), .Y(n15075) );
  sky130_fd_sc_hd__clkinv_1 U15574 ( .A(n14919), .Y(n19737) );
  sky130_fd_sc_hd__clkinv_1 U15576 ( .A(n25333), .Y(n22825) );
  sky130_fd_sc_hd__nor2_1 U15577 ( .A(n21209), .B(n22099), .Y(n21210) );
  sky130_fd_sc_hd__a21boi_0 U15578 ( .A1(n21634), .A2(n21330), .B1_N(n24884), 
        .Y(n21537) );
  sky130_fd_sc_hd__clkinv_1 U15579 ( .A(n23229), .Y(n21599) );
  sky130_fd_sc_hd__and2_0 U15580 ( .A(n20348), .B(n22418), .X(n24878) );
  sky130_fd_sc_hd__clkinv_1 U15581 ( .A(n25316), .Y(n24872) );
  sky130_fd_sc_hd__nand3_1 U15582 ( .A(n14958), .B(n14957), .C(n21074), .Y(
        n22403) );
  sky130_fd_sc_hd__and2_0 U15583 ( .A(n25251), .B(n14959), .X(n14957) );
  sky130_fd_sc_hd__clkinv_1 U15584 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[5]), .Y(n18288) );
  sky130_fd_sc_hd__nand3_1 U15585 ( .A(n14976), .B(n14975), .C(n14974), .Y(
        n21207) );
  sky130_fd_sc_hd__clkinv_1 U15586 ( .A(n21076), .Y(n14976) );
  sky130_fd_sc_hd__clkinv_1 U15587 ( .A(n25149), .Y(n22963) );
  sky130_fd_sc_hd__clkinv_1 U15588 ( .A(gpio_en_o[1]), .Y(io_oeb[1]) );
  sky130_fd_sc_hd__clkinv_1 U15589 ( .A(gpio_en_o[2]), .Y(io_oeb[2]) );
  sky130_fd_sc_hd__clkinv_1 U15590 ( .A(gpio_en_o[3]), .Y(io_oeb[3]) );
  sky130_fd_sc_hd__clkinv_1 U15591 ( .A(gpio_en_o[5]), .Y(io_oeb[7]) );
  sky130_fd_sc_hd__clkinv_1 U15592 ( .A(gpio_en_o[6]), .Y(io_oeb[26]) );
  sky130_fd_sc_hd__clkinv_1 U15593 ( .A(gpio_en_o[7]), .Y(io_oeb[27]) );
  sky130_fd_sc_hd__clkinv_1 U15594 ( .A(gpio_en_o[9]), .Y(io_oeb[29]) );
  sky130_fd_sc_hd__clkinv_1 U15595 ( .A(gpio_en_o[10]), .Y(io_oeb[30]) );
  sky130_fd_sc_hd__clkinv_1 U15596 ( .A(gpio_en_o[11]), .Y(io_oeb[31]) );
  sky130_fd_sc_hd__clkinv_1 U15597 ( .A(gpio_en_o[12]), .Y(io_oeb[32]) );
  sky130_fd_sc_hd__clkinv_1 U15598 ( .A(gpio_en_o[13]), .Y(io_oeb[33]) );
  sky130_fd_sc_hd__clkinv_1 U15599 ( .A(gpio_en_o[14]), .Y(io_oeb[34]) );
  sky130_fd_sc_hd__clkinv_1 U15600 ( .A(gpio_en_o[15]), .Y(io_oeb[35]) );
  sky130_fd_sc_hd__clkinv_1 U15601 ( .A(gpio_en_o[17]), .Y(io_oeb[37]) );
  sky130_fd_sc_hd__clkinv_1 U15602 ( .A(n23534), .Y(io_out[8]) );
  sky130_fd_sc_hd__clkbuf_1 U15603 ( .A(n20498), .X(n25307) );
  sky130_fd_sc_hd__clkinv_1 U15604 ( .A(j202_soc_core_intr_vec__0_), .Y(n22901) );
  sky130_fd_sc_hd__clkinv_1 U15605 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]), .Y(n24935) );
  sky130_fd_sc_hd__clkinv_1 U15606 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[7]), .Y(n24914) );
  sky130_fd_sc_hd__clkinv_1 U15607 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[5]), .Y(n24907) );
  sky130_fd_sc_hd__and2_0 U15608 ( .A(j202_soc_core_wbqspiflash_00_spi_in[0]), 
        .B(n23690), .X(j202_soc_core_wbqspiflash_00_lldriver_N391) );
  sky130_fd_sc_hd__clkinv_1 U15609 ( .A(n24261), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N21) );
  sky130_fd_sc_hd__clkinv_1 U15610 ( .A(j202_soc_core_intc_core_00_rg_ipr[11]), 
        .Y(n24383) );
  sky130_fd_sc_hd__o2bb2ai_1 U15611 ( .B1(n24424), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[114]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o2bb2ai_1 U15612 ( .B1(n20477), .B2(n24424), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[122]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__and2_0 U15613 ( .A(n21970), .B(n21996), .X(n25464) );
  sky130_fd_sc_hd__clkinv_1 U15614 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[9]), .Y(n24919) );
  sky130_fd_sc_hd__clkinv_1 U15615 ( .A(j202_soc_core_intc_core_00_rg_ipr[25]), 
        .Y(n24394) );
  sky130_fd_sc_hd__o2bb2ai_1 U15616 ( .B1(n24393), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[54]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__clkinv_1 U15617 ( .A(j202_soc_core_intc_core_00_rg_ipr[81]), 
        .Y(n24333) );
  sky130_fd_sc_hd__and2_0 U15618 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[17]), .B(n25734), .X(
        j202_soc_core_wbqspiflash_00_N714) );
  sky130_fd_sc_hd__clkinv_1 U15619 ( .A(j202_soc_core_intc_core_00_rg_ipr[33]), 
        .Y(n24352) );
  sky130_fd_sc_hd__clkinv_1 U15620 ( .A(n22750), .Y(n22751) );
  sky130_fd_sc_hd__clkinv_1 U15621 ( .A(j202_soc_core_intc_core_00_rg_ipr[55]), 
        .Y(n24369) );
  sky130_fd_sc_hd__clkinv_1 U15622 ( .A(j202_soc_core_intc_core_00_rg_ipr[52]), 
        .Y(n24367) );
  sky130_fd_sc_hd__clkinv_1 U15623 ( .A(j202_soc_core_intc_core_00_rg_ipr[45]), 
        .Y(n24362) );
  sky130_fd_sc_hd__clkinv_1 U15624 ( .A(j202_soc_core_intc_core_00_rg_ipr[44]), 
        .Y(n24361) );
  sky130_fd_sc_hd__clkinv_1 U15625 ( .A(j202_soc_core_intc_core_00_rg_ipr[35]), 
        .Y(n24354) );
  sky130_fd_sc_hd__clkinv_1 U15626 ( .A(j202_soc_core_intc_core_00_rg_ipr[82]), 
        .Y(n24334) );
  sky130_fd_sc_hd__clkinv_1 U15627 ( .A(j202_soc_core_intc_core_00_rg_ipr[79]), 
        .Y(n24331) );
  sky130_fd_sc_hd__clkinv_1 U15628 ( .A(j202_soc_core_intc_core_00_rg_ipr[68]), 
        .Y(n24328) );
  sky130_fd_sc_hd__clkinv_1 U15629 ( .A(j202_soc_core_intc_core_00_rg_ipr[27]), 
        .Y(n24398) );
  sky130_fd_sc_hd__clkinv_1 U15630 ( .A(j202_soc_core_intc_core_00_rg_ipr[16]), 
        .Y(n24384) );
  sky130_fd_sc_hd__clkinv_1 U15631 ( .A(j202_soc_core_intc_core_00_rg_ipr[4]), 
        .Y(n24380) );
  sky130_fd_sc_hd__clkinv_1 U15632 ( .A(j202_soc_core_ahb2apb_01_state[1]), 
        .Y(n21229) );
  sky130_fd_sc_hd__nor2_1 U15634 ( .A(n19797), .B(n19799), .Y(n25339) );
  sky130_fd_sc_hd__clkinv_1 U15635 ( .A(j202_soc_core_ahb2apb_02_state[1]), 
        .Y(n21231) );
  sky130_fd_sc_hd__o2bb2ai_1 U15636 ( .B1(n21189), .B2(n23312), .A1_N(n21189), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N3255) );
  sky130_fd_sc_hd__o2bb2ai_1 U15637 ( .B1(n21187), .B2(n23312), .A1_N(n21187), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N3218) );
  sky130_fd_sc_hd__o2bb2ai_1 U15638 ( .B1(n21186), .B2(n23312), .A1_N(n21186), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N3181) );
  sky130_fd_sc_hd__o2bb2ai_1 U15639 ( .B1(n21071), .B2(n23312), .A1_N(n21071), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N3144) );
  sky130_fd_sc_hd__o2bb2ai_1 U15640 ( .B1(n21184), .B2(n23312), .A1_N(n21184), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N3107) );
  sky130_fd_sc_hd__o2bb2ai_1 U15641 ( .B1(n21206), .B2(n23312), .A1_N(n21206), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N3070) );
  sky130_fd_sc_hd__o2bb2ai_1 U15642 ( .B1(n21199), .B2(n23312), .A1_N(n21199), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N3033) );
  sky130_fd_sc_hd__o2bb2ai_1 U15643 ( .B1(n21069), .B2(n23312), .A1_N(n21069), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N2996) );
  sky130_fd_sc_hd__o2bb2ai_1 U15644 ( .B1(n21183), .B2(n23312), .A1_N(n21183), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N2959) );
  sky130_fd_sc_hd__o2bb2ai_1 U15645 ( .B1(n21185), .B2(n23312), .A1_N(n21185), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N2922) );
  sky130_fd_sc_hd__o2bb2ai_1 U15646 ( .B1(n21201), .B2(n23312), .A1_N(n21201), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N2885) );
  sky130_fd_sc_hd__o2bb2ai_1 U15647 ( .B1(n21070), .B2(n23312), .A1_N(n21070), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N2848) );
  sky130_fd_sc_hd__o2bb2ai_1 U15648 ( .B1(n21182), .B2(n23312), .A1_N(n21182), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N2811) );
  sky130_fd_sc_hd__o2bb2ai_1 U15649 ( .B1(n21103), .B2(n23312), .A1_N(n21103), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N2774) );
  sky130_fd_sc_hd__o2bb2ai_1 U15650 ( .B1(n21203), .B2(n23312), .A1_N(n21203), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N2737) );
  sky130_fd_sc_hd__clkinv_1 U15651 ( .A(j202_soc_core_bldc_core_00_pwm_duty[8]), .Y(n25191) );
  sky130_fd_sc_hd__and2_0 U15652 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[16]), .B(n25734), .X(
        j202_soc_core_wbqspiflash_00_N713) );
  sky130_fd_sc_hd__and2_0 U15653 ( .A(n21782), .B(n21996), .X(n25466) );
  sky130_fd_sc_hd__clkinv_1 U15654 ( .A(n23306), .Y(n21783) );
  sky130_fd_sc_hd__and2_0 U15655 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[15]), .B(n25734), .X(
        j202_soc_core_wbqspiflash_00_N712) );
  sky130_fd_sc_hd__and2_0 U15656 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[20]), .B(n25734), .X(
        j202_soc_core_wbqspiflash_00_N717) );
  sky130_fd_sc_hd__clkinv_1 U15657 ( .A(n23585), .Y(
        j202_soc_core_wbqspiflash_00_N710) );
  sky130_fd_sc_hd__and2_0 U15658 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[21]), .B(n25734), .X(
        j202_soc_core_wbqspiflash_00_N718) );
  sky130_fd_sc_hd__clkinv_1 U15659 ( .A(j202_soc_core_j22_cpu_ml_bufa[31]), 
        .Y(n22191) );
  sky130_fd_sc_hd__and2_0 U15660 ( .A(n22269), .B(n21996), .X(n25467) );
  sky130_fd_sc_hd__and2_0 U15661 ( .A(n21924), .B(n21996), .X(n25468) );
  sky130_fd_sc_hd__and2_0 U15662 ( .A(n21834), .B(n21996), .X(n25469) );
  sky130_fd_sc_hd__clkinv_1 U15663 ( .A(n21937), .Y(n21836) );
  sky130_fd_sc_hd__and2_0 U15664 ( .A(n21874), .B(n21996), .X(n25470) );
  sky130_fd_sc_hd__and2_0 U15665 ( .A(n21858), .B(n21996), .X(n25471) );
  sky130_fd_sc_hd__and2_0 U15666 ( .A(n22346), .B(n21996), .X(n25472) );
  sky130_fd_sc_hd__and2_0 U15667 ( .A(n21947), .B(n21996), .X(n25447) );
  sky130_fd_sc_hd__and2_0 U15668 ( .A(n21752), .B(n21996), .X(n25473) );
  sky130_fd_sc_hd__clkinv_1 U15669 ( .A(n23309), .Y(n21753) );
  sky130_fd_sc_hd__and2_0 U15670 ( .A(n22111), .B(n21996), .X(n25430) );
  sky130_fd_sc_hd__and2_0 U15671 ( .A(n25491), .B(n22153), .X(n25481) );
  sky130_fd_sc_hd__clkinv_1 U15672 ( .A(n21668), .Y(n21670) );
  sky130_fd_sc_hd__and2_0 U15673 ( .A(n22122), .B(n21996), .X(n25474) );
  sky130_fd_sc_hd__and2_0 U15674 ( .A(n21761), .B(n21996), .X(n25427) );
  sky130_fd_sc_hd__clkinv_1 U15675 ( .A(n23326), .Y(n21079) );
  sky130_fd_sc_hd__and2_0 U15676 ( .A(n21819), .B(n21996), .X(n25475) );
  sky130_fd_sc_hd__clkinv_1 U15677 ( .A(n21625), .Y(n21626) );
  sky130_fd_sc_hd__clkinv_1 U15678 ( .A(n21397), .Y(n21400) );
  sky130_fd_sc_hd__clkinv_1 U15679 ( .A(n21851), .Y(n21848) );
  sky130_fd_sc_hd__clkinv_1 U15680 ( .A(n22262), .Y(n22263) );
  sky130_fd_sc_hd__and2_0 U15681 ( .A(n21613), .B(n21996), .X(n25478) );
  sky130_fd_sc_hd__and2_0 U15682 ( .A(n22286), .B(n21996), .X(n25431) );
  sky130_fd_sc_hd__and2_0 U15683 ( .A(n21850), .B(n21996), .X(n25476) );
  sky130_fd_sc_hd__and2_0 U15684 ( .A(n22033), .B(n21996), .X(n25479) );
  sky130_fd_sc_hd__and2_0 U15685 ( .A(n22258), .B(n21996), .X(n25480) );
  sky130_fd_sc_hd__and2_0 U15686 ( .A(n24826), .B(n24825), .X(n24834) );
  sky130_fd_sc_hd__clkinv_1 U15687 ( .A(j202_soc_core_j22_cpu_intack), .Y(
        n19326) );
  sky130_fd_sc_hd__clkinv_1 U15688 ( .A(n22009), .Y(n22015) );
  sky130_fd_sc_hd__and2_0 U15689 ( .A(n22248), .B(n21996), .X(n25448) );
  sky130_fd_sc_hd__nand4bb_1 U15690 ( .A_N(n21464), .B_N(n24867), .C(n21463), 
        .D(n21462), .Y(n21469) );
  sky130_fd_sc_hd__and2_0 U15691 ( .A(n18631), .B(n18630), .X(n18632) );
  sky130_fd_sc_hd__and2_1 U15692 ( .A(n21249), .B(n25260), .X(n25376) );
  sky130_fd_sc_hd__nand2_1 U15693 ( .A(n22824), .B(n25731), .Y(
        j202_soc_core_ahb2apb_00_N22) );
  sky130_fd_sc_hd__nor2_1 U15694 ( .A(n18477), .B(n21904), .Y(n25249) );
  sky130_fd_sc_hd__nand3_1 U15695 ( .A(n18225), .B(n18224), .C(n18223), .Y(
        n25380) );
  sky130_fd_sc_hd__and2_1 U15696 ( .A(n25299), .B(
        j202_soc_core_ahbcs_6__HREADY_), .X(j202_soc_core_j22_cpu_id_N7) );
  sky130_fd_sc_hd__and2_0 U15697 ( .A(n22789), .B(n21647), .X(n17822) );
  sky130_fd_sc_hd__or4_1 U15698 ( .A(n17494), .B(n17493), .C(n17492), .D(
        n17491), .X(n25274) );
  sky130_fd_sc_hd__clkinv_1 U15699 ( .A(n21343), .Y(n25544) );
  sky130_fd_sc_hd__clkinv_1 U15700 ( .A(n21617), .Y(n20228) );
  sky130_fd_sc_hd__clkinv_1 U15701 ( .A(n22821), .Y(n25488) );
  sky130_fd_sc_hd__nand3_1 U15702 ( .A(n20351), .B(n20350), .C(n20349), .Y(
        n10582) );
  sky130_fd_sc_hd__and2_0 U15703 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[31]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N34) );
  sky130_fd_sc_hd__and2_0 U15704 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[30]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N33) );
  sky130_fd_sc_hd__and2_0 U15705 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[29]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N32) );
  sky130_fd_sc_hd__and2_0 U15706 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[27]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N30) );
  sky130_fd_sc_hd__and2_0 U15707 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[26]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N29) );
  sky130_fd_sc_hd__and2_0 U15708 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[25]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N28) );
  sky130_fd_sc_hd__and2_0 U15709 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[24]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N27) );
  sky130_fd_sc_hd__and2_0 U15710 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[23]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N26) );
  sky130_fd_sc_hd__and2_0 U15711 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[22]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N25) );
  sky130_fd_sc_hd__and2_0 U15712 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[21]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N24) );
  sky130_fd_sc_hd__and2_0 U15713 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[17]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N20) );
  sky130_fd_sc_hd__and2_0 U15714 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N19) );
  sky130_fd_sc_hd__and2_0 U15715 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N16) );
  sky130_fd_sc_hd__and2_0 U15716 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[12]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N15) );
  sky130_fd_sc_hd__and2_0 U15717 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[11]), .B(n25734), 
        .X(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N14) );
  sky130_fd_sc_hd__and2_0 U15718 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[9]), .B(n25734), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N12) );
  sky130_fd_sc_hd__and2_0 U15719 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]), .B(n25734), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N11) );
  sky130_fd_sc_hd__and2_0 U15720 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]), .B(n25734), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N9) );
  sky130_fd_sc_hd__and2_0 U15721 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[4]), .B(n25734), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N7) );
  sky130_fd_sc_hd__and2_0 U15722 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]), .B(n25734), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N6) );
  sky130_fd_sc_hd__and2_0 U15723 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[0]), .B(n25734), .X(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N3) );
  sky130_fd_sc_hd__nor2b_1 U15724 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[28]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N31) );
  sky130_fd_sc_hd__nor2b_1 U15725 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[26]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N29) );
  sky130_fd_sc_hd__nor2b_1 U15726 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[24]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N27) );
  sky130_fd_sc_hd__nor2b_1 U15727 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[22]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N25) );
  sky130_fd_sc_hd__and2_0 U15728 ( .A(n25307), .B(wbs_dat_i[0]), .X(n5) );
  sky130_fd_sc_hd__and2_0 U15729 ( .A(n25307), .B(wbs_dat_i[1]), .X(n6) );
  sky130_fd_sc_hd__and2_0 U15730 ( .A(n25307), .B(wbs_dat_i[2]), .X(n7) );
  sky130_fd_sc_hd__and2_0 U15731 ( .A(n25307), .B(wbs_dat_i[3]), .X(n8) );
  sky130_fd_sc_hd__and2_0 U15732 ( .A(n25307), .B(wbs_dat_i[4]), .X(n9) );
  sky130_fd_sc_hd__and2_0 U15733 ( .A(n25307), .B(wbs_dat_i[5]), .X(n10) );
  sky130_fd_sc_hd__and2_0 U15734 ( .A(n25307), .B(wbs_dat_i[6]), .X(n11) );
  sky130_fd_sc_hd__a31o_1 U15735 ( .A1(n25307), .A2(wbs_we_i), .A3(
        wbs_sel_i[0]), .B1(wb_rst_i), .X(n4) );
  sky130_fd_sc_hd__and2_0 U15736 ( .A(n25307), .B(wbs_dat_i[7]), .X(n12) );
  sky130_fd_sc_hd__and2_0 U15737 ( .A(n20498), .B(wbs_dat_i[8]), .X(n14) );
  sky130_fd_sc_hd__and2_0 U15738 ( .A(n20498), .B(wbs_dat_i[9]), .X(n15) );
  sky130_fd_sc_hd__and2_0 U15739 ( .A(n20498), .B(wbs_dat_i[10]), .X(n16) );
  sky130_fd_sc_hd__and2_0 U15740 ( .A(n20498), .B(wbs_dat_i[11]), .X(n17) );
  sky130_fd_sc_hd__and2_0 U15741 ( .A(n20498), .B(wbs_dat_i[12]), .X(n18) );
  sky130_fd_sc_hd__and2_0 U15742 ( .A(n20498), .B(wbs_dat_i[13]), .X(n19) );
  sky130_fd_sc_hd__and2_0 U15743 ( .A(n20498), .B(wbs_dat_i[14]), .X(n20) );
  sky130_fd_sc_hd__a31o_1 U15744 ( .A1(n25307), .A2(wbs_we_i), .A3(
        wbs_sel_i[1]), .B1(wb_rst_i), .X(n13) );
  sky130_fd_sc_hd__and2_0 U15745 ( .A(n20498), .B(wbs_dat_i[15]), .X(n21) );
  sky130_fd_sc_hd__and2_0 U15746 ( .A(n20498), .B(wbs_dat_i[16]), .X(n230) );
  sky130_fd_sc_hd__and2_0 U15747 ( .A(n20498), .B(wbs_dat_i[17]), .X(n240) );
  sky130_fd_sc_hd__and2_0 U15748 ( .A(n20498), .B(wbs_dat_i[18]), .X(n250) );
  sky130_fd_sc_hd__and2_0 U15749 ( .A(n20498), .B(wbs_dat_i[19]), .X(n260) );
  sky130_fd_sc_hd__and2_0 U15750 ( .A(n25307), .B(wbs_dat_i[20]), .X(n270) );
  sky130_fd_sc_hd__and2_0 U15751 ( .A(n25307), .B(wbs_dat_i[21]), .X(n280) );
  sky130_fd_sc_hd__and2_0 U15752 ( .A(n25307), .B(wbs_dat_i[22]), .X(n290) );
  sky130_fd_sc_hd__a31o_1 U15753 ( .A1(n25307), .A2(wbs_we_i), .A3(
        wbs_sel_i[2]), .B1(wb_rst_i), .X(n220) );
  sky130_fd_sc_hd__and2_0 U15754 ( .A(n25307), .B(wbs_dat_i[23]), .X(n300) );
  sky130_fd_sc_hd__and2_0 U15755 ( .A(n20498), .B(wbs_dat_i[24]), .X(n320) );
  sky130_fd_sc_hd__and2_0 U15756 ( .A(n25307), .B(wbs_dat_i[25]), .X(n330) );
  sky130_fd_sc_hd__and2_0 U15757 ( .A(n25307), .B(wbs_dat_i[26]), .X(n340) );
  sky130_fd_sc_hd__and2_0 U15758 ( .A(n25307), .B(wbs_dat_i[27]), .X(n350) );
  sky130_fd_sc_hd__and2_0 U15759 ( .A(n25307), .B(wbs_dat_i[28]), .X(n360) );
  sky130_fd_sc_hd__and2_0 U15760 ( .A(n25307), .B(wbs_dat_i[29]), .X(n370) );
  sky130_fd_sc_hd__and2_0 U15761 ( .A(n25307), .B(wbs_dat_i[30]), .X(n380) );
  sky130_fd_sc_hd__a31o_1 U15762 ( .A1(n25307), .A2(wbs_we_i), .A3(
        wbs_sel_i[3]), .B1(wb_rst_i), .X(n310) );
  sky130_fd_sc_hd__and2_0 U15763 ( .A(n25307), .B(wbs_dat_i[31]), .X(n390) );
  sky130_fd_sc_hd__buf_4 U15764 ( .A(n21320), .X(n25526) );
  sky130_fd_sc_hd__nor2_1 U15765 ( .A(n21319), .B(n11036), .Y(n21320) );
  sky130_fd_sc_hd__buf_4 U15766 ( .A(n21318), .X(n25525) );
  sky130_fd_sc_hd__nor2_1 U15767 ( .A(n21317), .B(n11036), .Y(n21318) );
  sky130_fd_sc_hd__buf_4 U15768 ( .A(n21316), .X(n25524) );
  sky130_fd_sc_hd__nor2_1 U15769 ( .A(n21315), .B(n11036), .Y(n21316) );
  sky130_fd_sc_hd__buf_4 U15770 ( .A(n21314), .X(n25522) );
  sky130_fd_sc_hd__nor2_1 U15771 ( .A(n21313), .B(n11036), .Y(n21314) );
  sky130_fd_sc_hd__buf_4 U15772 ( .A(n21312), .X(n25521) );
  sky130_fd_sc_hd__nor2_1 U15773 ( .A(n21311), .B(n11036), .Y(n21312) );
  sky130_fd_sc_hd__buf_4 U15774 ( .A(n21310), .X(n25520) );
  sky130_fd_sc_hd__nor2_1 U15775 ( .A(n21309), .B(n11036), .Y(n21310) );
  sky130_fd_sc_hd__buf_4 U15776 ( .A(n21308), .X(n25519) );
  sky130_fd_sc_hd__nor2_1 U15777 ( .A(n21307), .B(n11036), .Y(n21308) );
  sky130_fd_sc_hd__buf_4 U15778 ( .A(n21306), .X(n25518) );
  sky130_fd_sc_hd__nor2_1 U15779 ( .A(n21305), .B(n11036), .Y(n21306) );
  sky130_fd_sc_hd__buf_4 U15780 ( .A(n21304), .X(n25517) );
  sky130_fd_sc_hd__nor2_1 U15781 ( .A(n21303), .B(n11036), .Y(n21304) );
  sky130_fd_sc_hd__buf_4 U15782 ( .A(n21302), .X(n25516) );
  sky130_fd_sc_hd__nor2_1 U15783 ( .A(n21301), .B(n11036), .Y(n21302) );
  sky130_fd_sc_hd__nor2_1 U15784 ( .A(n21297), .B(n11036), .Y(n21298) );
  sky130_fd_sc_hd__nor2_1 U15786 ( .A(n21295), .B(n11036), .Y(n21296) );
  sky130_fd_sc_hd__buf_4 U15787 ( .A(n21294), .X(n25512) );
  sky130_fd_sc_hd__nor2_1 U15788 ( .A(n21293), .B(n11036), .Y(n21294) );
  sky130_fd_sc_hd__buf_4 U15789 ( .A(n21292), .X(n25511) );
  sky130_fd_sc_hd__nor2_1 U15790 ( .A(n21291), .B(n11036), .Y(n21292) );
  sky130_fd_sc_hd__buf_4 U15791 ( .A(n21290), .X(n25510) );
  sky130_fd_sc_hd__nor2_1 U15792 ( .A(n21289), .B(n11036), .Y(n21290) );
  sky130_fd_sc_hd__buf_4 U15793 ( .A(n21288), .X(n25509) );
  sky130_fd_sc_hd__nor2_1 U15794 ( .A(n21287), .B(n11036), .Y(n21288) );
  sky130_fd_sc_hd__buf_4 U15795 ( .A(n21286), .X(n25508) );
  sky130_fd_sc_hd__nor2_1 U15796 ( .A(n21285), .B(n11036), .Y(n21286) );
  sky130_fd_sc_hd__buf_4 U15797 ( .A(n21284), .X(n25507) );
  sky130_fd_sc_hd__nor2_1 U15798 ( .A(n21283), .B(n11036), .Y(n21284) );
  sky130_fd_sc_hd__buf_4 U15799 ( .A(n21282), .X(n25505) );
  sky130_fd_sc_hd__nor2_1 U15800 ( .A(n21281), .B(n11036), .Y(n21282) );
  sky130_fd_sc_hd__buf_4 U15801 ( .A(n21280), .X(n25504) );
  sky130_fd_sc_hd__nor2_1 U15802 ( .A(n21279), .B(n11036), .Y(n21280) );
  sky130_fd_sc_hd__buf_4 U15803 ( .A(n21278), .X(n25503) );
  sky130_fd_sc_hd__nor2_1 U15804 ( .A(n21277), .B(n11036), .Y(n21278) );
  sky130_fd_sc_hd__buf_4 U15805 ( .A(n21276), .X(n25502) );
  sky130_fd_sc_hd__nor2_1 U15806 ( .A(n21275), .B(n11036), .Y(n21276) );
  sky130_fd_sc_hd__buf_4 U15807 ( .A(n21274), .X(n25501) );
  sky130_fd_sc_hd__nor2_1 U15808 ( .A(n21273), .B(n11036), .Y(n21274) );
  sky130_fd_sc_hd__buf_4 U15809 ( .A(n21270), .X(n25497) );
  sky130_fd_sc_hd__nor2_1 U15810 ( .A(n21269), .B(n11036), .Y(n21270) );
  sky130_fd_sc_hd__buf_4 U15811 ( .A(n21268), .X(n25496) );
  sky130_fd_sc_hd__nor2_1 U15812 ( .A(n21267), .B(n11036), .Y(n21268) );
  sky130_fd_sc_hd__buf_4 U15813 ( .A(n21266), .X(n25495) );
  sky130_fd_sc_hd__nor2_1 U15814 ( .A(n21265), .B(n11036), .Y(n21266) );
  sky130_fd_sc_hd__clkinv_1 U15815 ( .A(j202_soc_core_j22_cpu_ml_bufb[32]), 
        .Y(n11169) );
  sky130_fd_sc_hd__nand3_1 U15816 ( .A(n14955), .B(n14954), .C(n14953), .Y(
        n21253) );
  sky130_fd_sc_hd__and2b_1 U15817 ( .B(n20475), .A_N(j202_soc_core_rst), .X(
        n20473) );
  sky130_fd_sc_hd__nor2_1 U15819 ( .A(n21104), .B(n20355), .Y(n21937) );
  sky130_fd_sc_hd__nor2_1 U15820 ( .A(n20406), .B(n20355), .Y(n23312) );
  sky130_fd_sc_hd__clkinv_1 U15821 ( .A(n23312), .Y(n20409) );
  sky130_fd_sc_hd__nor2_1 U15822 ( .A(n21078), .B(n20355), .Y(n23326) );
  sky130_fd_sc_hd__and4_1 U15825 ( .A(n12306), .B(n12305), .C(n12304), .D(
        n12303), .X(n11187) );
  sky130_fd_sc_hd__nor2_1 U15827 ( .A(n21136), .B(n20355), .Y(n23318) );
  sky130_fd_sc_hd__clkinv_1 U15828 ( .A(n21132), .Y(n21185) );
  sky130_fd_sc_hd__clkinv_1 U15829 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .Y(n13014) );
  sky130_fd_sc_hd__clkinv_1 U15830 ( .A(j202_soc_core_j22_cpu_regop_Rm__2_), 
        .Y(n11520) );
  sky130_fd_sc_hd__clkinv_1 U15831 ( .A(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .Y(n24784) );
  sky130_fd_sc_hd__nor2_1 U15832 ( .A(j202_soc_core_j22_cpu_pc_hold), .B(
        n21592), .Y(n24858) );
  sky130_fd_sc_hd__clkinv_1 U15833 ( .A(n24858), .Y(n24882) );
  sky130_fd_sc_hd__a21boi_1 U15834 ( .A1(n20735), .A2(n21137), .B1_N(n20734), 
        .Y(n21805) );
  sky130_fd_sc_hd__clkinv_1 U15835 ( .A(n21073), .Y(n21187) );
  sky130_fd_sc_hd__clkinv_1 U15836 ( .A(n21205), .Y(n21206) );
  sky130_fd_sc_hd__clkinv_1 U15837 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[2]), 
        .Y(n22697) );
  sky130_fd_sc_hd__clkinv_1 U15838 ( .A(n22322), .Y(n20705) );
  sky130_fd_sc_hd__nand2_1 U15839 ( .A(n20307), .B(n20273), .Y(n21192) );
  sky130_fd_sc_hd__clkinv_1 U15840 ( .A(n21192), .Y(n21103) );
  sky130_fd_sc_hd__clkinv_1 U15841 ( .A(n11522), .Y(n11519) );
  sky130_fd_sc_hd__nand2_1 U15842 ( .A(n20307), .B(n20262), .Y(n21195) );
  sky130_fd_sc_hd__clkinv_1 U15843 ( .A(n21195), .Y(n21071) );
  sky130_fd_sc_hd__nand2_1 U15844 ( .A(n20307), .B(n20259), .Y(n21193) );
  sky130_fd_sc_hd__clkinv_1 U15845 ( .A(n21193), .Y(n21069) );
  sky130_fd_sc_hd__nand2_1 U15846 ( .A(n20307), .B(n20267), .Y(n21194) );
  sky130_fd_sc_hd__clkinv_1 U15847 ( .A(n21194), .Y(n21070) );
  sky130_fd_sc_hd__clkinv_1 U15848 ( .A(n21133), .Y(n21183) );
  sky130_fd_sc_hd__clkinv_1 U15849 ( .A(n21068), .Y(n21184) );
  sky130_fd_sc_hd__clkinv_1 U15850 ( .A(n21072), .Y(n21182) );
  sky130_fd_sc_hd__clkinv_1 U15851 ( .A(n21134), .Y(n21186) );
  sky130_fd_sc_hd__and4_1 U15852 ( .A(n11961), .B(n11960), .C(n11959), .D(
        n11958), .X(n11197) );
  sky130_fd_sc_hd__clkinv_1 U15853 ( .A(n21202), .Y(n21203) );
  sky130_fd_sc_hd__clkinv_1 U15854 ( .A(j202_soc_core_j22_cpu_ml_bufa[1]), .Y(
        n15666) );
  sky130_fd_sc_hd__a21oi_1 U15855 ( .A1(n21892), .A2(n21178), .B1(n21067), .Y(
        n11199) );
  sky130_fd_sc_hd__and2_1 U15856 ( .A(n25249), .B(n18478), .X(n11200) );
  sky130_fd_sc_hd__clkinv_1 U15857 ( .A(j202_soc_core_j22_cpu_rfuo_sr__t_), 
        .Y(n11202) );
  sky130_fd_sc_hd__a21oi_1 U15858 ( .A1(n22426), .A2(n21178), .B1(n21038), .Y(
        n11201) );
  sky130_fd_sc_hd__clkinv_1 U15859 ( .A(n20219), .Y(n25493) );
  sky130_fd_sc_hd__clkinv_1 U15860 ( .A(n25382), .Y(n19483) );
  sky130_fd_sc_hd__nand2b_1 U15861 ( .A_N(n16157), .B(n16155), .Y(n19336) );
  sky130_fd_sc_hd__nand2_1 U15862 ( .A(n16599), .B(n21664), .Y(n16580) );
  sky130_fd_sc_hd__nor2_1 U15863 ( .A(n11477), .B(n20299), .Y(n13893) );
  sky130_fd_sc_hd__nor2_1 U15864 ( .A(n11477), .B(n20261), .Y(n13913) );
  sky130_fd_sc_hd__nor2_1 U15865 ( .A(n11477), .B(n20297), .Y(n13901) );
  sky130_fd_sc_hd__nor2_1 U15866 ( .A(n11477), .B(n20286), .Y(n13914) );
  sky130_fd_sc_hd__nor2_1 U15867 ( .A(n12127), .B(n12128), .Y(n15073) );
  sky130_fd_sc_hd__nor2_1 U15868 ( .A(j202_soc_core_j22_cpu_regop_Rn__1_), .B(
        n11448), .Y(n11461) );
  sky130_fd_sc_hd__nand2_1 U15869 ( .A(n21139), .B(n16665), .Y(n21174) );
  sky130_fd_sc_hd__nand3_1 U15870 ( .A(n16682), .B(n21011), .C(n20638), .Y(
        n20931) );
  sky130_fd_sc_hd__nand3_1 U15871 ( .A(n16642), .B(n16641), .C(n16640), .Y(
        n16682) );
  sky130_fd_sc_hd__nor2_1 U15872 ( .A(n11244), .B(n17717), .Y(n18379) );
  sky130_fd_sc_hd__nor2_1 U15873 ( .A(n20091), .B(n24292), .Y(n24579) );
  sky130_fd_sc_hd__nor2_1 U15874 ( .A(n24293), .B(n24378), .Y(n24349) );
  sky130_fd_sc_hd__a21oi_1 U15875 ( .A1(n17051), .A2(n14086), .B1(n11949), .Y(
        n22064) );
  sky130_fd_sc_hd__nand2_1 U15876 ( .A(n19670), .B(n19669), .Y(n19671) );
  sky130_fd_sc_hd__nor2_1 U15877 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[3]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[5]), .Y(n22687) );
  sky130_fd_sc_hd__nand2_1 U15878 ( .A(n20708), .B(n20354), .Y(n20355) );
  sky130_fd_sc_hd__clkinv_1 U15880 ( .A(n20931), .Y(n21139) );
  sky130_fd_sc_hd__nand2_1 U15881 ( .A(n20275), .B(
        j202_soc_core_j22_cpu_regop_We__3_), .Y(n20479) );
  sky130_fd_sc_hd__o21a_1 U15882 ( .A1(n16859), .A2(n20353), .B1(n16648), .X(
        n20708) );
  sky130_fd_sc_hd__clkinv_1 U15883 ( .A(n23457), .Y(n23442) );
  sky130_fd_sc_hd__nand2_1 U15884 ( .A(n12985), .B(n12984), .Y(n19078) );
  sky130_fd_sc_hd__clkinv_1 U15885 ( .A(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n18758) );
  sky130_fd_sc_hd__nor2_1 U15886 ( .A(n22125), .B(n21795), .Y(n20016) );
  sky130_fd_sc_hd__nand2_1 U15887 ( .A(n21619), .B(n21617), .Y(n21623) );
  sky130_fd_sc_hd__nand2_1 U15888 ( .A(n13653), .B(n16689), .Y(n21212) );
  sky130_fd_sc_hd__nor2_1 U15889 ( .A(j202_soc_core_intc_core_00_bs_addr[1]), 
        .B(j202_soc_core_intc_core_00_bs_addr[0]), .Y(n24471) );
  sky130_fd_sc_hd__nor2_1 U15890 ( .A(j202_soc_core_rst), .B(n24497), .Y(
        n24776) );
  sky130_fd_sc_hd__clkinv_1 U15891 ( .A(n13706), .Y(n20677) );
  sky130_fd_sc_hd__xor2_1 U15892 ( .A(n19672), .B(n19671), .X(n21731) );
  sky130_fd_sc_hd__nand2_1 U15893 ( .A(n21663), .B(n16599), .Y(n20030) );
  sky130_fd_sc_hd__nand2_1 U15894 ( .A(n21729), .B(n21725), .Y(n22216) );
  sky130_fd_sc_hd__o211ai_1 U15895 ( .A1(n20242), .A2(n20241), .B1(n20240), 
        .C1(n20239), .Y(n20243) );
  sky130_fd_sc_hd__nand2b_1 U15896 ( .A_N(n20355), .B(n22551), .Y(n21009) );
  sky130_fd_sc_hd__nand2_1 U15897 ( .A(n13654), .B(
        j202_soc_core_j22_cpu_memop_MEM__3_), .Y(n19917) );
  sky130_fd_sc_hd__nor2_1 U15898 ( .A(n23243), .B(n21241), .Y(n19905) );
  sky130_fd_sc_hd__nor2_1 U15899 ( .A(n24379), .B(n24378), .Y(n24576) );
  sky130_fd_sc_hd__nor3_1 U15900 ( .A(n22972), .B(n22969), .C(n22975), .Y(
        n23021) );
  sky130_fd_sc_hd__nand3_1 U15901 ( .A(n19242), .B(n19241), .C(n19240), .Y(
        n22725) );
  sky130_fd_sc_hd__nor2_1 U15902 ( .A(j202_soc_core_rst), .B(n24496), .Y(
        n24768) );
  sky130_fd_sc_hd__nor2_1 U15903 ( .A(n23417), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n25086) );
  sky130_fd_sc_hd__nand2_1 U15904 ( .A(n19734), .B(n19078), .Y(n19661) );
  sky130_fd_sc_hd__nand3_1 U15905 ( .A(n13182), .B(n13181), .C(n13180), .Y(
        n22531) );
  sky130_fd_sc_hd__nor2_1 U15906 ( .A(n18277), .B(n11410), .Y(n18726) );
  sky130_fd_sc_hd__nor2_1 U15907 ( .A(n11239), .B(n18212), .Y(n18610) );
  sky130_fd_sc_hd__o22ai_1 U15908 ( .A1(n21620), .A2(n21623), .B1(n21619), 
        .B2(n21618), .Y(n22378) );
  sky130_fd_sc_hd__nand2_1 U15909 ( .A(wbs_stb_i), .B(wbs_cyc_i), .Y(n20072)
         );
  sky130_fd_sc_hd__o21a_1 U15910 ( .A1(n21324), .A2(n22860), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd), .X(n23732) );
  sky130_fd_sc_hd__nor2b_1 U15911 ( .B_N(n25122), .A(n21325), .Y(n23853) );
  sky130_fd_sc_hd__clkinv_1 U15912 ( .A(n25392), .Y(n23699) );
  sky130_fd_sc_hd__clkinv_1 U15913 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .Y(n25070) );
  sky130_fd_sc_hd__nor2_1 U15914 ( .A(n21731), .B(n22216), .Y(n22198) );
  sky130_fd_sc_hd__clkinv_1 U15915 ( .A(n21924), .Y(n20544) );
  sky130_fd_sc_hd__clkinv_1 U15916 ( .A(n22093), .Y(n22163) );
  sky130_fd_sc_hd__clkinv_1 U15917 ( .A(n21949), .Y(n23332) );
  sky130_fd_sc_hd__nand2_1 U15918 ( .A(n21009), .B(n20929), .Y(n23306) );
  sky130_fd_sc_hd__clkinv_1 U15919 ( .A(n21971), .Y(n23315) );
  sky130_fd_sc_hd__clkinv_1 U15920 ( .A(n21188), .Y(n21189) );
  sky130_fd_sc_hd__o211ai_1 U15921 ( .A1(n20309), .A2(n20285), .B1(n20284), 
        .C1(n20307), .Y(n21198) );
  sky130_fd_sc_hd__clkinv_1 U15922 ( .A(n21200), .Y(n21201) );
  sky130_fd_sc_hd__nand3_1 U15923 ( .A(n23239), .B(n20277), .C(n20233), .Y(
        n22366) );
  sky130_fd_sc_hd__nand3_1 U15924 ( .A(n16685), .B(n16684), .C(n16683), .Y(
        n22286) );
  sky130_fd_sc_hd__clkinv_1 U15925 ( .A(n22045), .Y(n22520) );
  sky130_fd_sc_hd__o21a_1 U15927 ( .A1(n20638), .A2(n20568), .B1(n20567), .X(
        n22297) );
  sky130_fd_sc_hd__clkinv_1 U15928 ( .A(n22143), .Y(n22145) );
  sky130_fd_sc_hd__nand2_1 U15929 ( .A(n22104), .B(j202_soc_core_aquc_SEL__2_), 
        .Y(n22813) );
  sky130_fd_sc_hd__nand2_1 U15930 ( .A(n24576), .B(j202_soc_core_pwrite[1]), 
        .Y(n24404) );
  sky130_fd_sc_hd__nor2_1 U15931 ( .A(n24899), .B(n23491), .Y(n24898) );
  sky130_fd_sc_hd__nand2_1 U15932 ( .A(n24689), .B(
        j202_soc_core_intc_core_00_bs_addr[7]), .Y(n24777) );
  sky130_fd_sc_hd__clkinv_1 U15933 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .Y(n23690) );
  sky130_fd_sc_hd__a21oi_1 U15934 ( .A1(n25274), .A2(n19737), .B1(n17832), .Y(
        n22816) );
  sky130_fd_sc_hd__nor3_1 U15935 ( .A(wb_rst_i), .B(wbs_ack_o), .C(n20072), 
        .Y(n20498) );
  sky130_fd_sc_hd__nor2_1 U15936 ( .A(n21299), .B(n11036), .Y(n21300) );
  sky130_fd_sc_hd__nor2_1 U15937 ( .A(n21271), .B(n11036), .Y(n21272) );
  sky130_fd_sc_hd__nor2_1 U15938 ( .A(n23697), .B(n23731), .Y(n25392) );
  sky130_fd_sc_hd__o2bb2ai_1 U15939 ( .B1(n24424), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[98]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__clkinv_1 U15940 ( .A(n24428), .Y(n25278) );
  sky130_fd_sc_hd__o2bb2ai_1 U15941 ( .B1(n24440), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[116]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o2bb2ai_1 U15942 ( .B1(n24420), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[50]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o2bb2ai_1 U15943 ( .B1(n24393), .B2(n24442), .A1_N(
        j202_soc_core_intc_core_00_rg_ie[25]), .A2_N(n20114), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o2bb2ai_1 U15944 ( .B1(n24436), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[36]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o2bb2ai_1 U15945 ( .B1(n24475), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[32]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o2bb2ai_1 U15946 ( .B1(n20477), .B2(n24475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[56]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__nand2_1 U15947 ( .A(n18851), .B(n18850), .Y(n25374) );
  sky130_fd_sc_hd__o2bb2ai_1 U15948 ( .B1(n24405), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[119]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o2bb2ai_1 U15949 ( .B1(n24432), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[115]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o2bb2ai_1 U15950 ( .B1(n23940), .B2(n20473), .A1_N(n20475), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[19]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o2bb2ai_1 U15951 ( .B1(n24405), .B2(n20477), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[127]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o2bb2ai_1 U15952 ( .B1(n20477), .B2(n24397), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[126]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o2bb2ai_1 U15953 ( .B1(n20477), .B2(n24477), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[88]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o2bb2ai_1 U15954 ( .B1(n24389), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[69]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o2bb2ai_1 U15955 ( .B1(n23918), .B2(n20115), .A1_N(n24290), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[2]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o2bb2ai_1 U15956 ( .B1(n24405), .B2(n24442), .A1_N(
        j202_soc_core_intc_core_00_rg_ie[31]), .A2_N(n20114), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__clkinv_1 U15957 ( .A(n24279), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N14) );
  sky130_fd_sc_hd__clkbuf_1 U15958 ( .A(n10671), .X(n25533) );
  sky130_fd_sc_hd__nor2_1 U15959 ( .A(j202_soc_core_rst), .B(n23909), .Y(
        n25297) );
  sky130_fd_sc_hd__clkbuf_1 U15960 ( .A(n10672), .X(n25532) );
  sky130_fd_sc_hd__nor2_1 U15961 ( .A(n25378), .B(n22025), .Y(
        j202_soc_core_ahb2aqu_00_N97) );
  sky130_fd_sc_hd__a21oi_1 U15962 ( .A1(n20122), .A2(n23368), .B1(
        j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N755) );
  sky130_fd_sc_hd__clkbuf_1 U15963 ( .A(n20090), .X(n25491) );
  sky130_fd_sc_hd__nand3_1 U15964 ( .A(n19498), .B(n19497), .C(n19496), .Y(
        n25379) );
  sky130_fd_sc_hd__nor2_1 U15965 ( .A(n22817), .B(n22824), .Y(
        j202_soc_core_ahb2apb_00_N23) );
  sky130_fd_sc_hd__nand2_1 U15966 ( .A(n18836), .B(n18835), .Y(n25271) );
  sky130_fd_sc_hd__clkbuf_1 U15967 ( .A(j202_soc_core_j22_cpu_ml_N323), .X(
        n25537) );
  sky130_fd_sc_hd__nor2_1 U15968 ( .A(n22822), .B(n22824), .Y(
        j202_soc_core_ahb2apb_00_N27) );
  sky130_fd_sc_hd__nor2_1 U15969 ( .A(n25232), .B(n25231), .Y(
        j202_soc_core_uart_TOP_rx_fifo_N29) );
  sky130_fd_sc_hd__nor2_1 U15970 ( .A(n22820), .B(n22824), .Y(
        j202_soc_core_ahb2apb_00_N28) );
  sky130_fd_sc_hd__nor2_1 U15971 ( .A(n21915), .B(n22025), .Y(
        j202_soc_core_ahb2aqu_00_N98) );
  sky130_fd_sc_hd__nor3_1 U15972 ( .A(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[1]), .B(n20431), .C(n24781), 
        .Y(n25403) );
  sky130_fd_sc_hd__clkbuf_1 U15973 ( .A(j202_soc_core_wbqspiflash_00_N752), 
        .X(n25535) );
  sky130_fd_sc_hd__nand3_1 U15974 ( .A(n18340), .B(n18339), .C(n18338), .Y(
        n25387) );
  sky130_fd_sc_hd__nand3_1 U15975 ( .A(n22103), .B(n21912), .C(n21911), .Y(
        j202_soc_core_ahb2aqu_00_N164) );
  sky130_fd_sc_hd__and3_1 U15976 ( .A(n22802), .B(n17823), .C(n17822), .X(
        n25434) );
  sky130_fd_sc_hd__nand2_1 U15977 ( .A(n21618), .B(n20229), .Y(n25490) );
  sky130_fd_sc_hd__buf_4 U15979 ( .A(n21298), .X(n25514) );
  sky130_fd_sc_hd__buf_4 U15980 ( .A(n21272), .X(n25499) );
  sky130_fd_sc_hd__clkbuf_1 U15981 ( .A(io_oeb[12]), .X(io_oeb[13]) );
  sky130_fd_sc_hd__clkbuf_1 U15982 ( .A(la_data_out[1]), .X(io_out[1]) );
  sky130_fd_sc_hd__clkbuf_1 U15983 ( .A(la_data_out[10]), .X(io_out[30]) );
  sky130_fd_sc_hd__nand2_1 U15984 ( .A(n11202), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n12117) );
  sky130_fd_sc_hd__nand2_1 U15985 ( .A(n13210), .B(
        j202_soc_core_bootrom_00_address_w[8]), .Y(n11207) );
  sky130_fd_sc_hd__nor3b_1 U15986 ( .C_N(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[6]), .A(j202_soc_core_bootrom_00_address_w[17]), .B(
        j202_soc_core_bootrom_00_address_w[16]), .Y(n11206) );
  sky130_fd_sc_hd__nor2_1 U15987 ( .A(j202_soc_core_j22_cpu_ma_M_area[0]), .B(
        n11287), .Y(n11242) );
  sky130_fd_sc_hd__nor2_1 U15988 ( .A(j202_soc_core_bootrom_00_address_w[14]), 
        .B(j202_soc_core_bootrom_00_address_w[13]), .Y(n11204) );
  sky130_fd_sc_hd__nor2_1 U15989 ( .A(j202_soc_core_bootrom_00_address_w[15]), 
        .B(j202_soc_core_bootrom_00_address_w[12]), .Y(n11203) );
  sky130_fd_sc_hd__nor2_1 U15990 ( .A(n11207), .B(n18212), .Y(n17609) );
  sky130_fd_sc_hd__nand2_1 U15991 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .B(j202_soc_core_bootrom_00_address_w[5]), .Y(n14639) );
  sky130_fd_sc_hd__nor2_1 U15992 ( .A(j202_soc_core_bootrom_00_address_w[7]), 
        .B(n14983), .Y(n14399) );
  sky130_fd_sc_hd__nand2_1 U15993 ( .A(n14399), .B(n15017), .Y(n14120) );
  sky130_fd_sc_hd__nor2_1 U15994 ( .A(n14639), .B(n14120), .Y(n13334) );
  sky130_fd_sc_hd__nand2_1 U15995 ( .A(n13334), .B(n13014), .Y(n13487) );
  sky130_fd_sc_hd__nor2_1 U15996 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .B(n14985), .Y(n14348) );
  sky130_fd_sc_hd__nand2b_1 U15997 ( .A_N(n14120), .B(n14348), .Y(n13465) );
  sky130_fd_sc_hd__nor2_1 U15998 ( .A(n13014), .B(n13465), .Y(n13332) );
  sky130_fd_sc_hd__nor2_1 U15999 ( .A(n13411), .B(n13332), .Y(n11210) );
  sky130_fd_sc_hd__nor2_1 U16000 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .B(j202_soc_core_bootrom_00_address_w[4]), .Y(n14352) );
  sky130_fd_sc_hd__nand2_1 U16001 ( .A(n14352), .B(
        j202_soc_core_bootrom_00_address_w[11]), .Y(n11356) );
  sky130_fd_sc_hd__nand2_1 U16002 ( .A(n14983), .B(
        j202_soc_core_bootrom_00_address_w[7]), .Y(n11213) );
  sky130_fd_sc_hd__nand2_1 U16003 ( .A(n13374), .B(n14096), .Y(n11276) );
  sky130_fd_sc_hd__nor2_1 U16004 ( .A(n13014), .B(n11276), .Y(n11232) );
  sky130_fd_sc_hd__nand2_1 U16005 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .B(j202_soc_core_bootrom_00_address_w[2]), .Y(n14101) );
  sky130_fd_sc_hd__nor2_1 U16006 ( .A(n15017), .B(n14101), .Y(n14990) );
  sky130_fd_sc_hd__nand2_1 U16007 ( .A(n14990), .B(n14096), .Y(n18125) );
  sky130_fd_sc_hd__nor2_1 U16008 ( .A(n14094), .B(n18125), .Y(n11227) );
  sky130_fd_sc_hd__nand2_1 U16009 ( .A(n14983), .B(
        j202_soc_core_bootrom_00_address_w[5]), .Y(n11208) );
  sky130_fd_sc_hd__nor2_1 U16010 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .B(n13014), .Y(n15016) );
  sky130_fd_sc_hd__nand2_1 U16011 ( .A(n15016), .B(
        j202_soc_core_bootrom_00_address_w[11]), .Y(n15009) );
  sky130_fd_sc_hd__nor2_1 U16012 ( .A(n11208), .B(n15009), .Y(n18250) );
  sky130_fd_sc_hd__nand2_1 U16013 ( .A(n18250), .B(n14999), .Y(n13312) );
  sky130_fd_sc_hd__nor2_1 U16014 ( .A(n11227), .B(n13330), .Y(n13169) );
  sky130_fd_sc_hd__nand2_1 U16015 ( .A(n14985), .B(n13014), .Y(n14111) );
  sky130_fd_sc_hd__nand2_1 U16016 ( .A(n13198), .B(
        j202_soc_core_bootrom_00_address_w[11]), .Y(n17442) );
  sky130_fd_sc_hd__nor2_1 U16017 ( .A(n11213), .B(n17442), .Y(n13589) );
  sky130_fd_sc_hd__nand2_1 U16018 ( .A(n13589), .B(
        j202_soc_core_bootrom_00_address_w[5]), .Y(n13111) );
  sky130_fd_sc_hd__nand2_1 U16019 ( .A(n13169), .B(n13111), .Y(n13107) );
  sky130_fd_sc_hd__nand2_1 U16020 ( .A(n14348), .B(n15017), .Y(n11363) );
  sky130_fd_sc_hd__nand2_1 U16021 ( .A(j202_soc_core_bootrom_00_address_w[10]), 
        .B(j202_soc_core_bootrom_00_address_w[7]), .Y(n13449) );
  sky130_fd_sc_hd__nor2_1 U16022 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n13449), .Y(n12991) );
  sky130_fd_sc_hd__nand2_1 U16023 ( .A(n11209), .B(n12991), .Y(n13326) );
  sky130_fd_sc_hd__nor2_1 U16024 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .B(n14094), .Y(n15093) );
  sky130_fd_sc_hd__nand2_1 U16025 ( .A(n15093), .B(n15017), .Y(n13171) );
  sky130_fd_sc_hd__nor2_1 U16026 ( .A(n13449), .B(n13171), .Y(n13434) );
  sky130_fd_sc_hd__nand2_1 U16027 ( .A(n13326), .B(n13492), .Y(n11211) );
  sky130_fd_sc_hd__nor3_1 U16028 ( .A(n11232), .B(n13107), .C(n11211), .Y(
        n13415) );
  sky130_fd_sc_hd__nor2_1 U16029 ( .A(j202_soc_core_bootrom_00_address_w[7]), 
        .B(n15017), .Y(n14456) );
  sky130_fd_sc_hd__nand2_1 U16030 ( .A(n14456), .B(n14983), .Y(n14113) );
  sky130_fd_sc_hd__nor2_1 U16031 ( .A(n15149), .B(n14113), .Y(n13123) );
  sky130_fd_sc_hd__nand2_1 U16032 ( .A(n13123), .B(n13014), .Y(n13472) );
  sky130_fd_sc_hd__nor2_1 U16033 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(j202_soc_core_bootrom_00_address_w[3]), .Y(n13483) );
  sky130_fd_sc_hd__a31oi_1 U16034 ( .A1(n11210), .A2(n13415), .A3(n13472), 
        .B1(n17730), .Y(n11223) );
  sky130_fd_sc_hd__nand2_1 U16035 ( .A(n13014), .B(
        j202_soc_core_bootrom_00_address_w[4]), .Y(n14099) );
  sky130_fd_sc_hd__nor2_1 U16036 ( .A(n15017), .B(n14099), .Y(n17533) );
  sky130_fd_sc_hd__nand2_1 U16037 ( .A(n17533), .B(n14096), .Y(n13212) );
  sky130_fd_sc_hd__nor2_1 U16038 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .B(n13212), .Y(n11280) );
  sky130_fd_sc_hd__nor2_1 U16039 ( .A(n11280), .B(n13332), .Y(n11218) );
  sky130_fd_sc_hd__nand2_1 U16040 ( .A(n14111), .B(n11211), .Y(n13417) );
  sky130_fd_sc_hd__nand2_1 U16041 ( .A(n14098), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n12994) );
  sky130_fd_sc_hd__nand2_1 U16042 ( .A(n14613), .B(n15017), .Y(n13448) );
  sky130_fd_sc_hd__nor2_1 U16043 ( .A(n12994), .B(n13448), .Y(n13416) );
  sky130_fd_sc_hd__nand2_1 U16044 ( .A(n13589), .B(n14094), .Y(n13172) );
  sky130_fd_sc_hd__nor2_1 U16045 ( .A(n13416), .B(n13485), .Y(n11266) );
  sky130_fd_sc_hd__nor2_1 U16046 ( .A(j202_soc_core_bootrom_00_address_w[7]), 
        .B(j202_soc_core_bootrom_00_address_w[10]), .Y(n14236) );
  sky130_fd_sc_hd__nand2_1 U16047 ( .A(n17533), .B(n14236), .Y(n14777) );
  sky130_fd_sc_hd__nor2_1 U16048 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .B(n14777), .Y(n13452) );
  sky130_fd_sc_hd__nor2_1 U16049 ( .A(n14619), .B(n14120), .Y(n13440) );
  sky130_fd_sc_hd__or4_1 U16050 ( .A(n13308), .B(n13411), .C(n13452), .D(
        n13463), .X(n11212) );
  sky130_fd_sc_hd__nor2b_1 U16051 ( .B_N(n13417), .A(n11212), .Y(n13301) );
  sky130_fd_sc_hd__nor2_1 U16052 ( .A(n14094), .B(n14777), .Y(n11264) );
  sky130_fd_sc_hd__nand2_1 U16053 ( .A(n14352), .B(n15017), .Y(n11340) );
  sky130_fd_sc_hd__nor2_1 U16054 ( .A(n11340), .B(n12994), .Y(n13136) );
  sky130_fd_sc_hd__nor2_1 U16055 ( .A(n11264), .B(n13136), .Y(n13488) );
  sky130_fd_sc_hd__nand2_1 U16056 ( .A(n13334), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n13493) );
  sky130_fd_sc_hd__nand2_1 U16057 ( .A(n14613), .B(
        j202_soc_core_bootrom_00_address_w[11]), .Y(n11362) );
  sky130_fd_sc_hd__nor2_1 U16058 ( .A(n11362), .B(n11213), .Y(n13431) );
  sky130_fd_sc_hd__nand2_1 U16059 ( .A(n18250), .B(
        j202_soc_core_bootrom_00_address_w[7]), .Y(n13109) );
  sky130_fd_sc_hd__nand2_1 U16060 ( .A(n14236), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n13006) );
  sky130_fd_sc_hd__nand2_1 U16061 ( .A(n13374), .B(n13413), .Y(n13454) );
  sky130_fd_sc_hd__nand2_1 U16062 ( .A(n13109), .B(n13454), .Y(n13420) );
  sky130_fd_sc_hd__nor4b_1 U16063 ( .D_N(n13488), .A(n13435), .B(n13431), .C(
        n13420), .Y(n11214) );
  sky130_fd_sc_hd__nor2_1 U16064 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(n14100), .Y(n13489) );
  sky130_fd_sc_hd__a31oi_1 U16065 ( .A1(n11218), .A2(n13301), .A3(n11214), 
        .B1(n17468), .Y(n11222) );
  sky130_fd_sc_hd__nor2_1 U16066 ( .A(n11363), .B(n12994), .Y(n13333) );
  sky130_fd_sc_hd__nor2_1 U16067 ( .A(n11227), .B(n13333), .Y(n11217) );
  sky130_fd_sc_hd__nand2_1 U16068 ( .A(j202_soc_core_bootrom_00_address_w[3]), 
        .B(j202_soc_core_bootrom_00_address_w[6]), .Y(n13464) );
  sky130_fd_sc_hd__nand2_1 U16069 ( .A(n14236), .B(n13014), .Y(n11215) );
  sky130_fd_sc_hd__nor2_1 U16070 ( .A(n11215), .B(n11356), .Y(n13328) );
  sky130_fd_sc_hd__nor2_1 U16071 ( .A(n14631), .B(n18125), .Y(n13167) );
  sky130_fd_sc_hd__nor2_1 U16072 ( .A(n13328), .B(n13167), .Y(n13110) );
  sky130_fd_sc_hd__nand2_1 U16074 ( .A(n13454), .B(n13472), .Y(n13372) );
  sky130_fd_sc_hd__nor3b_1 U16075 ( .C_N(n13110), .A(n13421), .B(n13372), .Y(
        n11216) );
  sky130_fd_sc_hd__nor2_1 U16076 ( .A(j202_soc_core_bootrom_00_address_w[3]), 
        .B(n14998), .Y(n13121) );
  sky130_fd_sc_hd__o22ai_1 U16077 ( .A1(n11217), .A2(n13464), .B1(n11216), 
        .B2(n13500), .Y(n13303) );
  sky130_fd_sc_hd__nand2b_1 U16078 ( .A_N(n13171), .B(n13056), .Y(n13166) );
  sky130_fd_sc_hd__nand2_1 U16079 ( .A(n13166), .B(n13109), .Y(n13468) );
  sky130_fd_sc_hd__nand2_1 U16080 ( .A(n14348), .B(
        j202_soc_core_bootrom_00_address_w[11]), .Y(n11347) );
  sky130_fd_sc_hd__nand2_1 U16081 ( .A(n13412), .B(n13413), .Y(n13486) );
  sky130_fd_sc_hd__nand2_1 U16082 ( .A(n13434), .B(n13014), .Y(n13307) );
  sky130_fd_sc_hd__nand3_1 U16083 ( .A(n11218), .B(n13486), .C(n13307), .Y(
        n11219) );
  sky130_fd_sc_hd__a32oi_1 U16085 ( .A1(n13494), .A2(n11220), .A3(n11276), 
        .B1(n13464), .B2(n11220), .Y(n11221) );
  sky130_fd_sc_hd__nor4_1 U16086 ( .A(n11223), .B(n11222), .C(n13303), .D(
        n11221), .Y(n11332) );
  sky130_fd_sc_hd__nand2_1 U16087 ( .A(n13595), .B(
        j202_soc_core_bootrom_00_address_w[5]), .Y(n13365) );
  sky130_fd_sc_hd__nand2_1 U16088 ( .A(n11224), .B(n13365), .Y(n11230) );
  sky130_fd_sc_hd__nor2_1 U16089 ( .A(n11232), .B(n11280), .Y(n13502) );
  sky130_fd_sc_hd__nor2_1 U16090 ( .A(n13167), .B(n11258), .Y(n13424) );
  sky130_fd_sc_hd__nand2_1 U16091 ( .A(n13424), .B(n13454), .Y(n13120) );
  sky130_fd_sc_hd__nor2_1 U16092 ( .A(n11230), .B(n13120), .Y(n11228) );
  sky130_fd_sc_hd__nor2_1 U16093 ( .A(n11362), .B(n13006), .Y(n13299) );
  sky130_fd_sc_hd__nor2_1 U16094 ( .A(n13328), .B(n13299), .Y(n13460) );
  sky130_fd_sc_hd__nand2_1 U16095 ( .A(n15017), .B(n13014), .Y(n16741) );
  sky130_fd_sc_hd__nand3_1 U16096 ( .A(n11225), .B(n14098), .C(n14613), .Y(
        n13165) );
  sky130_fd_sc_hd__nor4_1 U16097 ( .A(n18250), .B(n13435), .C(n13433), .D(
        n13452), .Y(n11226) );
  sky130_fd_sc_hd__a31oi_1 U16098 ( .A1(n11228), .A2(n13460), .A3(n11226), 
        .B1(n13500), .Y(n13323) );
  sky130_fd_sc_hd__nor2_1 U16099 ( .A(n11347), .B(n14604), .Y(n13439) );
  sky130_fd_sc_hd__nor4_1 U16100 ( .A(n13416), .B(n13136), .C(n13439), .D(
        n13463), .Y(n13133) );
  sky130_fd_sc_hd__nor2_1 U16101 ( .A(n11227), .B(n13299), .Y(n11278) );
  sky130_fd_sc_hd__nand2_1 U16102 ( .A(n11278), .B(n13124), .Y(n11281) );
  sky130_fd_sc_hd__nor2_1 U16103 ( .A(n11264), .B(n11281), .Y(n13175) );
  sky130_fd_sc_hd__and3_1 U16104 ( .A(n11228), .B(n13133), .C(n13175), .X(
        n11229) );
  sky130_fd_sc_hd__a31oi_1 U16105 ( .A1(n11229), .A2(n13492), .A3(n13109), 
        .B1(n13464), .Y(n11238) );
  sky130_fd_sc_hd__nor2_1 U16106 ( .A(n13332), .B(n11230), .Y(n13418) );
  sky130_fd_sc_hd__nor2_1 U16107 ( .A(n11264), .B(n11280), .Y(n11257) );
  sky130_fd_sc_hd__nand2_1 U16108 ( .A(n13170), .B(n13166), .Y(n11261) );
  sky130_fd_sc_hd__nor2_1 U16109 ( .A(n13299), .B(n13439), .Y(n13129) );
  sky130_fd_sc_hd__nand3b_1 U16110 ( .A_N(n11261), .B(n13129), .C(n11234), .Y(
        n13317) );
  sky130_fd_sc_hd__nor2_1 U16111 ( .A(n13440), .B(n13317), .Y(n11231) );
  sky130_fd_sc_hd__a31oi_1 U16112 ( .A1(n13418), .A2(n11257), .A3(n11231), 
        .B1(n17730), .Y(n11237) );
  sky130_fd_sc_hd__nand2b_1 U16113 ( .A_N(n11232), .B(n11257), .Y(n13469) );
  sky130_fd_sc_hd__nor2_1 U16114 ( .A(n13300), .B(n13469), .Y(n13441) );
  sky130_fd_sc_hd__nand2_1 U16115 ( .A(n13441), .B(n13307), .Y(n13316) );
  sky130_fd_sc_hd__nor2_1 U16116 ( .A(n11340), .B(n11233), .Y(n11265) );
  sky130_fd_sc_hd__nor2_1 U16117 ( .A(n13433), .B(n11265), .Y(n13474) );
  sky130_fd_sc_hd__nand3b_1 U16118 ( .A_N(n13452), .B(n13474), .C(n11234), .Y(
        n11262) );
  sky130_fd_sc_hd__nor4_1 U16119 ( .A(n13114), .B(n13299), .C(n13316), .D(
        n11262), .Y(n11235) );
  sky130_fd_sc_hd__a21oi_1 U16120 ( .A1(n11235), .A2(n13109), .B1(n17468), .Y(
        n11236) );
  sky130_fd_sc_hd__nor4_1 U16121 ( .A(n13323), .B(n11238), .C(n11237), .D(
        n11236), .Y(n11240) );
  sky130_fd_sc_hd__nand2_1 U16122 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .B(j202_soc_core_bootrom_00_address_w[9]), .Y(n11239) );
  sky130_fd_sc_hd__nand2b_1 U16123 ( .A_N(n11240), .B(n18610), .Y(n11331) );
  sky130_fd_sc_hd__nand2_1 U16124 ( .A(n11242), .B(n11241), .Y(n18306) );
  sky130_fd_sc_hd__nand2_1 U16125 ( .A(n11428), .B(n18288), .Y(n11243) );
  sky130_fd_sc_hd__nor2_1 U16126 ( .A(n11243), .B(n18306), .Y(n11245) );
  sky130_fd_sc_hd__nand2_1 U16127 ( .A(n11245), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[3]), .Y(n17717) );
  sky130_fd_sc_hd__a22oi_1 U16128 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[21]), .B1(n18379), .B2(
        j202_soc_core_uart_div1[5]), .Y(n11275) );
  sky130_fd_sc_hd__nand2_1 U16129 ( .A(n18277), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[1]), .Y(n11246) );
  sky130_fd_sc_hd__nand2_1 U16130 ( .A(n11245), .B(n18283), .Y(n11410) );
  sky130_fd_sc_hd__a22oi_1 U16131 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[85]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[53]), .Y(n11274) );
  sky130_fd_sc_hd__nor2_1 U16132 ( .A(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[0]), .B(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[1]), .Y(n21227) );
  sky130_fd_sc_hd__nand3_1 U16133 ( .A(n21228), .B(n21227), .C(n11247), .Y(
        n15063) );
  sky130_fd_sc_hd__nor2_1 U16134 ( .A(j202_soc_core_aquc_ADR__2_), .B(n15063), 
        .Y(n17716) );
  sky130_fd_sc_hd__mux2i_1 U16135 ( .A0(j202_soc_core_aquc_ADR__3_), .A1(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[3]), .S(n15063), 
        .Y(n19742) );
  sky130_fd_sc_hd__nor2_1 U16136 ( .A(j202_soc_core_aquc_ADR__1_), .B(
        j202_soc_core_aquc_ADR__0_), .Y(n11249) );
  sky130_fd_sc_hd__nor3_1 U16137 ( .A(j202_soc_core_aquc_ADR__5_), .B(
        j202_soc_core_aquc_ADR__7_), .C(j202_soc_core_aquc_ADR__6_), .Y(n11248) );
  sky130_fd_sc_hd__nand2_1 U16138 ( .A(n11249), .B(n11248), .Y(n11253) );
  sky130_fd_sc_hd__nor2_1 U16139 ( .A(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[1]), .B(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[0]), .Y(n11251) );
  sky130_fd_sc_hd__nor3_1 U16140 ( .A(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[7]), .B(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[6]), .C(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[5]), .Y(n11250) );
  sky130_fd_sc_hd__a21oi_1 U16141 ( .A1(n11251), .A2(n11250), .B1(n25245), .Y(
        n11252) );
  sky130_fd_sc_hd__a21oi_1 U16142 ( .A1(n11253), .A2(n25245), .B1(n11252), .Y(
        n17709) );
  sky130_fd_sc_hd__nand2_1 U16143 ( .A(n15063), .B(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[4]), .Y(n11254) );
  sky130_fd_sc_hd__o21a_1 U16144 ( .A1(n11255), .A2(n15063), .B1(n11254), .X(
        n17710) );
  sky130_fd_sc_hd__nand2_1 U16145 ( .A(n17709), .B(n17710), .Y(n15065) );
  sky130_fd_sc_hd__nand2_1 U16146 ( .A(n19742), .B(n11256), .Y(n20496) );
  sky130_fd_sc_hd__nand2_1 U16147 ( .A(n17716), .B(n20430), .Y(n18282) );
  sky130_fd_sc_hd__nor2b_1 U16148 ( .B_N(n13109), .A(n13485), .Y(n13168) );
  sky130_fd_sc_hd__nand3_1 U16149 ( .A(n11257), .B(n13129), .C(n13168), .Y(
        n13313) );
  sky130_fd_sc_hd__nor3_1 U16150 ( .A(n13328), .B(n13300), .C(n11258), .Y(
        n13436) );
  sky130_fd_sc_hd__nor2_1 U16151 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n13465), .Y(n13422) );
  sky130_fd_sc_hd__a31oi_1 U16152 ( .A1(n13436), .A2(n13380), .A3(n11259), 
        .B1(n13464), .Y(n11260) );
  sky130_fd_sc_hd__a221oi_1 U16153 ( .A1(n11261), .A2(n13483), .B1(n13313), 
        .B2(n13483), .C1(n11260), .Y(n11271) );
  sky130_fd_sc_hd__o31ai_1 U16154 ( .A1(n13434), .A2(n13372), .A3(n11262), 
        .B1(n13121), .Y(n11270) );
  sky130_fd_sc_hd__nand2_1 U16155 ( .A(n13487), .B(n11263), .Y(n13458) );
  sky130_fd_sc_hd__nand2_1 U16156 ( .A(n13312), .B(n13112), .Y(n13381) );
  sky130_fd_sc_hd__nand2b_1 U16157 ( .A_N(n13381), .B(n13456), .Y(n13127) );
  sky130_fd_sc_hd__nor2_1 U16158 ( .A(n13299), .B(n13127), .Y(n13336) );
  sky130_fd_sc_hd__nand4_1 U16159 ( .A(n11266), .B(n13336), .C(n13326), .D(
        n13454), .Y(n11267) );
  sky130_fd_sc_hd__o21ai_1 U16160 ( .A1(n13458), .A2(n11267), .B1(n13489), .Y(
        n11269) );
  sky130_fd_sc_hd__nand2_1 U16161 ( .A(n13231), .B(
        j202_soc_core_bootrom_00_address_w[9]), .Y(n11268) );
  sky130_fd_sc_hd__a31oi_1 U16162 ( .A1(n11271), .A2(n11270), .A3(n11269), 
        .B1(n18552), .Y(n11272) );
  sky130_fd_sc_hd__a21oi_1 U16163 ( .A1(j202_soc_core_bldc_core_00_pwm_duty[9]), .A2(n18629), .B1(n11272), .Y(n11273) );
  sky130_fd_sc_hd__nand3_1 U16164 ( .A(n11275), .B(n11274), .C(n11273), .Y(
        n11329) );
  sky130_fd_sc_hd__nor3_1 U16165 ( .A(n13014), .B(n15149), .C(n14120), .Y(
        n13325) );
  sky130_fd_sc_hd__nor2_1 U16166 ( .A(n13325), .B(n13314), .Y(n13106) );
  sky130_fd_sc_hd__a211oi_1 U16167 ( .A1(n13056), .A2(n13412), .B1(n13114), 
        .C1(n13434), .Y(n13366) );
  sky130_fd_sc_hd__nand3_1 U16168 ( .A(n13480), .B(n13486), .C(n11276), .Y(
        n13457) );
  sky130_fd_sc_hd__a31oi_1 U16169 ( .A1(n13106), .A2(n13366), .A3(n11277), 
        .B1(n17468), .Y(n11286) );
  sky130_fd_sc_hd__a21oi_1 U16170 ( .A1(n13412), .A2(n13413), .B1(n13469), .Y(
        n13125) );
  sky130_fd_sc_hd__nor3_1 U16171 ( .A(n13411), .B(n13422), .C(n13314), .Y(
        n13331) );
  sky130_fd_sc_hd__nand2_1 U16172 ( .A(n13125), .B(n13331), .Y(n13173) );
  sky130_fd_sc_hd__a21oi_1 U16173 ( .A1(n13374), .A2(n13056), .B1(n13173), .Y(
        n13481) );
  sky130_fd_sc_hd__nand2_1 U16174 ( .A(n14399), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n13373) );
  sky130_fd_sc_hd__a21oi_1 U16175 ( .A1(n11356), .A2(n13171), .B1(n13373), .Y(
        n13367) );
  sky130_fd_sc_hd__nor3_1 U16176 ( .A(n13123), .B(n13367), .C(n13126), .Y(
        n11279) );
  sky130_fd_sc_hd__a21oi_1 U16177 ( .A1(n13481), .A2(n11279), .B1(n17730), .Y(
        n11285) );
  sky130_fd_sc_hd__nor3_1 U16179 ( .A(n11280), .B(n13136), .C(n13135), .Y(
        n11283) );
  sky130_fd_sc_hd__nand2_1 U16180 ( .A(n13326), .B(n13365), .Y(n13315) );
  sky130_fd_sc_hd__nor3_1 U16183 ( .A(n11286), .B(n11285), .C(n11284), .Y(
        n11327) );
  sky130_fd_sc_hd__nor2_1 U16184 ( .A(j202_soc_core_memory0_ram_dout0_sel[14]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[13]), .Y(n11302) );
  sky130_fd_sc_hd__nand2_1 U16185 ( .A(n11302), .B(n11289), .Y(n11295) );
  sky130_fd_sc_hd__nor2_1 U16186 ( .A(j202_soc_core_memory0_ram_dout0_sel[11]), 
        .B(n11295), .Y(n11299) );
  sky130_fd_sc_hd__nand2_1 U16187 ( .A(n11299), .B(n11290), .Y(n11297) );
  sky130_fd_sc_hd__nand2_1 U16188 ( .A(n11298), .B(n11291), .Y(n11292) );
  sky130_fd_sc_hd__nor2_1 U16189 ( .A(j202_soc_core_memory0_ram_dout0_sel[7]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[6]), .Y(n11315) );
  sky130_fd_sc_hd__nand2_1 U16190 ( .A(n11315), .B(n11293), .Y(n11316) );
  sky130_fd_sc_hd__nor2_1 U16191 ( .A(j202_soc_core_memory0_ram_dout0_sel[4]), 
        .B(n11316), .Y(n11313) );
  sky130_fd_sc_hd__nor2_1 U16192 ( .A(j202_soc_core_memory0_ram_dout0_sel[2]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[3]), .Y(n11294) );
  sky130_fd_sc_hd__nand3_1 U16193 ( .A(n11313), .B(
        j202_soc_core_memory0_ram_dout0_sel[1]), .C(n11294), .Y(n11389) );
  sky130_fd_sc_hd__nor2_1 U16194 ( .A(n18736), .B(n11389), .Y(n18739) );
  sky130_fd_sc_hd__a22oi_1 U16195 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[277]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[53]), .Y(n11324) );
  sky130_fd_sc_hd__nor2_1 U16196 ( .A(n11296), .B(n11295), .Y(n18743) );
  sky130_fd_sc_hd__nor2_1 U16197 ( .A(n11298), .B(n11297), .Y(n18741) );
  sky130_fd_sc_hd__a22o_1 U16198 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[309]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[341]), .X(n11300) );
  sky130_fd_sc_hd__a21oi_1 U16199 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[373]), .B1(n11300), .Y(n11323) );
  sky130_fd_sc_hd__nor2_1 U16200 ( .A(j202_soc_core_memory0_ram_dout0_sel[7]), 
        .B(n11301), .Y(n18360) );
  sky130_fd_sc_hd__nand2_1 U16201 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[245]), .Y(n11307) );
  sky130_fd_sc_hd__a21oi_1 U16202 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[469]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n11306) );
  sky130_fd_sc_hd__nand2_1 U16203 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[405]), .Y(n11305) );
  sky130_fd_sc_hd__nor2_1 U16204 ( .A(j202_soc_core_memory0_ram_dout0_sel[14]), 
        .B(n11303), .Y(n18746) );
  sky130_fd_sc_hd__nand2_1 U16205 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[437]), .Y(n11304) );
  sky130_fd_sc_hd__nand4_1 U16206 ( .A(n11307), .B(n11306), .C(n11305), .D(
        n11304), .Y(n11308) );
  sky130_fd_sc_hd__a21oi_1 U16207 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[213]), .B1(n11308), .Y(n11322) );
  sky130_fd_sc_hd__clkinv_1 U16208 ( .A(n11313), .Y(n11310) );
  sky130_fd_sc_hd__nor2_1 U16209 ( .A(n11312), .B(n11310), .Y(n18733) );
  sky130_fd_sc_hd__nand2_1 U16210 ( .A(n11309), .B(
        j202_soc_core_memory0_ram_dout0_sel[0]), .Y(n11311) );
  sky130_fd_sc_hd__nor4_1 U16211 ( .A(j202_soc_core_memory0_ram_dout0_sel[3]), 
        .B(j202_soc_core_memory0_ram_dout0_sel[1]), .C(n11311), .D(n11310), 
        .Y(n18367) );
  sky130_fd_sc_hd__clkbuf_1 U16212 ( .A(n18367), .X(n18731) );
  sky130_fd_sc_hd__and3_1 U16213 ( .A(n11313), .B(
        j202_soc_core_memory0_ram_dout0_sel[2]), .C(n11312), .X(n18730) );
  sky130_fd_sc_hd__a22o_1 U16214 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[21]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[85]), .X(n11314) );
  sky130_fd_sc_hd__a21oi_1 U16215 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[117]), .B1(n11314), .Y(n11319) );
  sky130_fd_sc_hd__nor2_1 U16216 ( .A(n11317), .B(n11316), .Y(n18734) );
  sky130_fd_sc_hd__a22oi_1 U16217 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[181]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[149]), .Y(n11318) );
  sky130_fd_sc_hd__nand2_1 U16218 ( .A(n11319), .B(n11318), .Y(n11320) );
  sky130_fd_sc_hd__nand2_1 U16219 ( .A(n11320), .B(n17639), .Y(n11321) );
  sky130_fd_sc_hd__nand4_1 U16220 ( .A(n11324), .B(n11323), .C(n11322), .D(
        n11321), .Y(n11325) );
  sky130_fd_sc_hd__o211ai_1 U16221 ( .A1(j202_soc_core_memory0_ram_dout0[501]), 
        .A2(n18758), .B1(n14906), .C1(n11325), .Y(n11326) );
  sky130_fd_sc_hd__o21ai_1 U16222 ( .A1(n18722), .A2(n11327), .B1(n11326), .Y(
        n11328) );
  sky130_fd_sc_hd__nor2_1 U16223 ( .A(n11329), .B(n11328), .Y(n11330) );
  sky130_fd_sc_hd__o211a_2 U16224 ( .A1(n18720), .A2(n11332), .B1(n11331), 
        .C1(n11330), .X(n22526) );
  sky130_fd_sc_hd__or3_1 U16225 ( .A(j202_soc_core_j22_cpu_id_op2_v_), .B(
        j202_soc_core_j22_cpu_id_opn_v_), .C(n22807), .X(n11333) );
  sky130_fd_sc_hd__nand2b_1 U16226 ( .A_N(n22526), .B(n19089), .Y(n11423) );
  sky130_fd_sc_hd__nand2_1 U16227 ( .A(j202_soc_core_bootrom_00_address_w[7]), 
        .B(j202_soc_core_bootrom_00_address_w[6]), .Y(n18792) );
  sky130_fd_sc_hd__nand2_1 U16228 ( .A(n18250), .B(n14100), .Y(n16925) );
  sky130_fd_sc_hd__nor2_1 U16229 ( .A(j202_soc_core_bootrom_00_address_w[3]), 
        .B(n14983), .Y(n14980) );
  sky130_fd_sc_hd__nor2_1 U16230 ( .A(n11339), .B(n13171), .Y(n11383) );
  sky130_fd_sc_hd__nand2_1 U16231 ( .A(n11383), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n18675) );
  sky130_fd_sc_hd__nor2_1 U16232 ( .A(n18770), .B(n15153), .Y(n18266) );
  sky130_fd_sc_hd__nand2_1 U16233 ( .A(n14352), .B(n14983), .Y(n11338) );
  sky130_fd_sc_hd__nand2_1 U16234 ( .A(j202_soc_core_bootrom_00_address_w[11]), 
        .B(j202_soc_core_bootrom_00_address_w[3]), .Y(n11336) );
  sky130_fd_sc_hd__nand2_1 U16235 ( .A(n14095), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n18296) );
  sky130_fd_sc_hd__nor2b_1 U16236 ( .B_N(n11334), .A(n18296), .Y(n16968) );
  sky130_fd_sc_hd__nand2_1 U16237 ( .A(n14100), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n11335) );
  sky130_fd_sc_hd__nand2_1 U16238 ( .A(n14613), .B(
        j202_soc_core_bootrom_00_address_w[10]), .Y(n11354) );
  sky130_fd_sc_hd__nand2b_1 U16239 ( .A_N(n11354), .B(n15017), .Y(n16985) );
  sky130_fd_sc_hd__nor2_1 U16240 ( .A(n11335), .B(n16985), .Y(n18710) );
  sky130_fd_sc_hd__nor2_1 U16241 ( .A(n16968), .B(n18710), .Y(n18264) );
  sky130_fd_sc_hd__nor2_1 U16242 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n11336), .Y(n11348) );
  sky130_fd_sc_hd__nor2_1 U16243 ( .A(n11338), .B(n11337), .Y(n18557) );
  sky130_fd_sc_hd__nor2_1 U16244 ( .A(n14100), .B(n16741), .Y(n11346) );
  sky130_fd_sc_hd__nand2_1 U16245 ( .A(n14352), .B(
        j202_soc_core_bootrom_00_address_w[10]), .Y(n18295) );
  sky130_fd_sc_hd__nor2b_1 U16246 ( .B_N(n11346), .A(n18295), .Y(n18585) );
  sky130_fd_sc_hd__nor2_1 U16247 ( .A(n18557), .B(n18585), .Y(n16929) );
  sky130_fd_sc_hd__nand2_1 U16248 ( .A(n14983), .B(
        j202_soc_core_bootrom_00_address_w[3]), .Y(n14108) );
  sky130_fd_sc_hd__nor3_1 U16249 ( .A(n14094), .B(n15017), .C(n14108), .Y(
        n18534) );
  sky130_fd_sc_hd__nand2_1 U16250 ( .A(n14472), .B(n18534), .Y(n18555) );
  sky130_fd_sc_hd__nor2_1 U16251 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n16985), .Y(n18543) );
  sky130_fd_sc_hd__nand2_1 U16252 ( .A(n15093), .B(
        j202_soc_core_bootrom_00_address_w[10]), .Y(n15090) );
  sky130_fd_sc_hd__nand2_1 U16253 ( .A(n15017), .B(
        j202_soc_core_bootrom_00_address_w[3]), .Y(n14989) );
  sky130_fd_sc_hd__nand2_1 U16254 ( .A(n14473), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n11355) );
  sky130_fd_sc_hd__nor2_1 U16255 ( .A(n15090), .B(n11355), .Y(n15121) );
  sky130_fd_sc_hd__nand2_1 U16256 ( .A(n14983), .B(n14100), .Y(n14978) );
  sky130_fd_sc_hd__nand2b_1 U16257 ( .A_N(n11356), .B(n14982), .Y(n16975) );
  sky130_fd_sc_hd__nor2_1 U16258 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n16975), .Y(n18673) );
  sky130_fd_sc_hd__nand2_1 U16259 ( .A(n14348), .B(
        j202_soc_core_bootrom_00_address_w[10]), .Y(n11342) );
  sky130_fd_sc_hd__nand2b_1 U16260 ( .A_N(n11342), .B(n11346), .Y(n18588) );
  sky130_fd_sc_hd__nor2_1 U16261 ( .A(n11340), .B(n11339), .Y(n15186) );
  sky130_fd_sc_hd__nand2_1 U16262 ( .A(n15186), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n16990) );
  sky130_fd_sc_hd__nor2_1 U16263 ( .A(n11354), .B(n11355), .Y(n15194) );
  sky130_fd_sc_hd__nor2_1 U16264 ( .A(n18645), .B(n15194), .Y(n18556) );
  sky130_fd_sc_hd__nand3_1 U16265 ( .A(n18713), .B(n18588), .C(n18556), .Y(
        n16926) );
  sky130_fd_sc_hd__nor4b_1 U16266 ( .D_N(n18555), .A(n18543), .B(n15121), .C(
        n16926), .Y(n11341) );
  sky130_fd_sc_hd__nand4_1 U16267 ( .A(n18266), .B(n18264), .C(n16929), .D(
        n11341), .Y(n11345) );
  sky130_fd_sc_hd__nor2_1 U16268 ( .A(n11342), .B(n11355), .Y(n18584) );
  sky130_fd_sc_hd__nand2_1 U16269 ( .A(n16974), .B(n18569), .Y(n18775) );
  sky130_fd_sc_hd__nor4_1 U16270 ( .A(n18645), .B(n18710), .C(n18775), .D(
        n16908), .Y(n11343) );
  sky130_fd_sc_hd__nor2_1 U16271 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(n14999), .Y(n18513) );
  sky130_fd_sc_hd__nand2_1 U16272 ( .A(n18543), .B(n14100), .Y(n18554) );
  sky130_fd_sc_hd__nor2_1 U16273 ( .A(n14978), .B(n17442), .Y(n17604) );
  sky130_fd_sc_hd__nand2_1 U16274 ( .A(n17604), .B(
        j202_soc_core_bootrom_00_address_w[5]), .Y(n18593) );
  sky130_fd_sc_hd__nand2_1 U16275 ( .A(n15186), .B(n13014), .Y(n15122) );
  sky130_fd_sc_hd__nand2_1 U16276 ( .A(n18593), .B(n15122), .Y(n15181) );
  sky130_fd_sc_hd__o21ai_1 U16278 ( .A1(n11343), .A2(n18783), .B1(n16918), .Y(
        n11344) );
  sky130_fd_sc_hd__a21oi_1 U16279 ( .A1(n18651), .A2(n11345), .B1(n11344), .Y(
        n11352) );
  sky130_fd_sc_hd__nor2_1 U16280 ( .A(j202_soc_core_bootrom_00_address_w[11]), 
        .B(n14099), .Y(n17777) );
  sky130_fd_sc_hd__nand2_1 U16281 ( .A(n17777), .B(n14980), .Y(n17799) );
  sky130_fd_sc_hd__nor2_1 U16282 ( .A(n18248), .B(n18645), .Y(n18292) );
  sky130_fd_sc_hd__nor2b_1 U16283 ( .B_N(n11346), .A(n15090), .Y(n18674) );
  sky130_fd_sc_hd__nand2_1 U16284 ( .A(n17533), .B(n14986), .Y(n17768) );
  sky130_fd_sc_hd__nor2_1 U16285 ( .A(n14094), .B(n17768), .Y(n18703) );
  sky130_fd_sc_hd__nand3_1 U16286 ( .A(n18292), .B(n18559), .C(n18558), .Y(
        n17000) );
  sky130_fd_sc_hd__nor2_1 U16287 ( .A(n14978), .B(n11347), .Y(n18704) );
  sky130_fd_sc_hd__nand2_1 U16288 ( .A(n18704), .B(n13014), .Y(n16916) );
  sky130_fd_sc_hd__nand2_1 U16289 ( .A(n11348), .B(n14348), .Y(n15140) );
  sky130_fd_sc_hd__nor2_1 U16290 ( .A(j202_soc_core_bootrom_00_address_w[10]), 
        .B(n15140), .Y(n18253) );
  sky130_fd_sc_hd__nand2_1 U16291 ( .A(n16916), .B(n18291), .Y(n18777) );
  sky130_fd_sc_hd__nor3_1 U16292 ( .A(n18673), .B(n18777), .C(n16908), .Y(
        n18663) );
  sky130_fd_sc_hd__nor2_1 U16293 ( .A(j202_soc_core_bootrom_00_address_w[7]), 
        .B(n14998), .Y(n18664) );
  sky130_fd_sc_hd__o21ai_1 U16294 ( .A1(n17000), .A2(n11349), .B1(n18664), .Y(
        n11351) );
  sky130_fd_sc_hd__nand2_1 U16295 ( .A(n18250), .B(
        j202_soc_core_bootrom_00_address_w[3]), .Y(n18289) );
  sky130_fd_sc_hd__nand4_1 U16296 ( .A(n18559), .B(n18558), .C(n18662), .D(
        n18289), .Y(n18525) );
  sky130_fd_sc_hd__nand2_1 U16297 ( .A(n18289), .B(n15122), .Y(n11357) );
  sky130_fd_sc_hd__nand2b_1 U16298 ( .A_N(n17604), .B(n18595), .Y(n15197) );
  sky130_fd_sc_hd__nor2_1 U16299 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(j202_soc_core_bootrom_00_address_w[7]), .Y(n18655) );
  sky130_fd_sc_hd__a31oi_1 U16301 ( .A1(n11352), .A2(n11351), .A3(n11350), 
        .B1(n18720), .Y(n11409) );
  sky130_fd_sc_hd__nand2_1 U16302 ( .A(n14472), .B(n14983), .Y(n13200) );
  sky130_fd_sc_hd__nand2b_1 U16303 ( .A_N(n13200), .B(n14095), .Y(n18519) );
  sky130_fd_sc_hd__nor2_1 U16304 ( .A(n14631), .B(n18519), .Y(n15182) );
  sky130_fd_sc_hd__nand2_1 U16305 ( .A(n16925), .B(n18592), .Y(n15096) );
  sky130_fd_sc_hd__nor3_1 U16306 ( .A(n18703), .B(n18766), .C(n15096), .Y(
        n11353) );
  sky130_fd_sc_hd__nor2_1 U16308 ( .A(n18295), .B(n11355), .Y(n18524) );
  sky130_fd_sc_hd__nand2_1 U16309 ( .A(n15189), .B(n18681), .Y(n18568) );
  sky130_fd_sc_hd__nor3_1 U16310 ( .A(j202_soc_core_bootrom_00_address_w[10]), 
        .B(n13014), .C(n11356), .Y(n18256) );
  sky130_fd_sc_hd__nand2_1 U16311 ( .A(n18256), .B(n14100), .Y(n18661) );
  sky130_fd_sc_hd__nand2_1 U16312 ( .A(n18704), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n16901) );
  sky130_fd_sc_hd__nand2_1 U16313 ( .A(n18661), .B(n16901), .Y(n15118) );
  sky130_fd_sc_hd__nor2_1 U16314 ( .A(n18253), .B(n15153), .Y(n16890) );
  sky130_fd_sc_hd__nand2_1 U16315 ( .A(n18533), .B(n16890), .Y(n18273) );
  sky130_fd_sc_hd__nor4_1 U16316 ( .A(n18527), .B(n18312), .C(n18568), .D(
        n18273), .Y(n11359) );
  sky130_fd_sc_hd__nand2_1 U16317 ( .A(n18593), .B(n18569), .Y(n16905) );
  sky130_fd_sc_hd__nor2_1 U16318 ( .A(n14978), .B(n11362), .Y(n16898) );
  sky130_fd_sc_hd__nand2_1 U16319 ( .A(n16898), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n18514) );
  sky130_fd_sc_hd__nand2_1 U16320 ( .A(n18543), .B(
        j202_soc_core_bootrom_00_address_w[3]), .Y(n16977) );
  sky130_fd_sc_hd__nand2_1 U16321 ( .A(n18514), .B(n16977), .Y(n18641) );
  sky130_fd_sc_hd__nor3_1 U16322 ( .A(n18641), .B(n16968), .C(n18644), .Y(
        n11381) );
  sky130_fd_sc_hd__nor3_1 U16323 ( .A(n11357), .B(n16905), .C(n11373), .Y(
        n11358) );
  sky130_fd_sc_hd__o22ai_1 U16324 ( .A1(n11359), .A2(n18792), .B1(n11358), 
        .B2(n18771), .Y(n11360) );
  sky130_fd_sc_hd__a21oi_1 U16325 ( .A1(n18513), .A2(n11361), .B1(n11360), .Y(
        n11366) );
  sky130_fd_sc_hd__nand2_1 U16326 ( .A(n16898), .B(n13014), .Y(n18680) );
  sky130_fd_sc_hd__nand2_1 U16327 ( .A(n18680), .B(n15122), .Y(n16986) );
  sky130_fd_sc_hd__nor2_1 U16328 ( .A(n14108), .B(n11362), .Y(n18638) );
  sky130_fd_sc_hd__nor2_1 U16329 ( .A(n15194), .B(n18638), .Y(n16907) );
  sky130_fd_sc_hd__nand2b_1 U16330 ( .A_N(n11363), .B(n14980), .Y(n15087) );
  sky130_fd_sc_hd__nor2_1 U16331 ( .A(n13014), .B(n15087), .Y(n18512) );
  sky130_fd_sc_hd__nand4_1 U16332 ( .A(n16907), .B(n18514), .C(n18291), .D(
        n18521), .Y(n11364) );
  sky130_fd_sc_hd__o21ai_1 U16333 ( .A1(n16986), .A2(n11364), .B1(n18655), .Y(
        n11365) );
  sky130_fd_sc_hd__a21oi_1 U16334 ( .A1(n11366), .A2(n11365), .B1(n18552), .Y(
        n11408) );
  sky130_fd_sc_hd__nor3_1 U16335 ( .A(n18704), .B(n18674), .C(n18253), .Y(
        n18252) );
  sky130_fd_sc_hd__nand2_1 U16336 ( .A(n15189), .B(n18593), .Y(n18540) );
  sky130_fd_sc_hd__nand2_1 U16337 ( .A(n16974), .B(n15122), .Y(n11367) );
  sky130_fd_sc_hd__nor2_1 U16338 ( .A(n11383), .B(n15194), .Y(n18314) );
  sky130_fd_sc_hd__nor2_1 U16339 ( .A(j202_soc_core_bootrom_00_address_w[10]), 
        .B(n14111), .Y(n13195) );
  sky130_fd_sc_hd__nand2_1 U16340 ( .A(n13195), .B(n14095), .Y(n14991) );
  sky130_fd_sc_hd__nor2_1 U16341 ( .A(n14094), .B(n14991), .Y(n16996) );
  sky130_fd_sc_hd__nand2_1 U16342 ( .A(n18314), .B(n18642), .Y(n16906) );
  sky130_fd_sc_hd__nor3_1 U16343 ( .A(n18540), .B(n11367), .C(n16906), .Y(
        n11368) );
  sky130_fd_sc_hd__nand4_1 U16344 ( .A(n18252), .B(n11368), .C(n18290), .D(
        n15199), .Y(n11371) );
  sky130_fd_sc_hd__nor3_1 U16345 ( .A(n18704), .B(n18703), .C(n16908), .Y(
        n16933) );
  sky130_fd_sc_hd__nor2_1 U16346 ( .A(n18674), .B(n15194), .Y(n18574) );
  sky130_fd_sc_hd__and3_1 U16347 ( .A(n18521), .B(n18660), .C(n18574), .X(
        n15204) );
  sky130_fd_sc_hd__nand2_1 U16348 ( .A(n18289), .B(n18592), .Y(n16976) );
  sky130_fd_sc_hd__nand2_1 U16349 ( .A(n18593), .B(n18555), .Y(n18263) );
  sky130_fd_sc_hd__nand2_1 U16350 ( .A(n16974), .B(n18661), .Y(n15085) );
  sky130_fd_sc_hd__nor2_1 U16351 ( .A(n18253), .B(n18643), .Y(n15151) );
  sky130_fd_sc_hd__nor4_1 U16352 ( .A(n16976), .B(n18263), .C(n15085), .D(
        n18255), .Y(n11369) );
  sky130_fd_sc_hd__a31oi_1 U16353 ( .A1(n16933), .A2(n15204), .A3(n11369), 
        .B1(n18792), .Y(n11370) );
  sky130_fd_sc_hd__a21oi_1 U16354 ( .A1(n18513), .A2(n11371), .B1(n11370), .Y(
        n11378) );
  sky130_fd_sc_hd__nor2_1 U16355 ( .A(n16996), .B(n18674), .Y(n18683) );
  sky130_fd_sc_hd__nand3_1 U16356 ( .A(n18558), .B(n18588), .C(n15151), .Y(
        n11375) );
  sky130_fd_sc_hd__nand4_1 U16357 ( .A(n18683), .B(n15191), .C(n16916), .D(
        n18555), .Y(n11372) );
  sky130_fd_sc_hd__o21ai_1 U16358 ( .A1(n11373), .A2(n11372), .B1(n18655), .Y(
        n11377) );
  sky130_fd_sc_hd__nand2_1 U16359 ( .A(n18554), .B(n18592), .Y(n18769) );
  sky130_fd_sc_hd__nor2_1 U16360 ( .A(n18687), .B(n18770), .Y(n11374) );
  sky130_fd_sc_hd__nand2_1 U16361 ( .A(n16974), .B(n18521), .Y(n15117) );
  sky130_fd_sc_hd__nor2_1 U16362 ( .A(n18568), .B(n15117), .Y(n16919) );
  sky130_fd_sc_hd__nand4_1 U16363 ( .A(n11374), .B(n16919), .C(n18555), .D(
        n16975), .Y(n18254) );
  sky130_fd_sc_hd__o31ai_1 U16364 ( .A1(n11375), .A2(n18769), .A3(n18254), 
        .B1(n18664), .Y(n11376) );
  sky130_fd_sc_hd__a31oi_1 U16365 ( .A1(n11378), .A2(n11377), .A3(n11376), 
        .B1(n18666), .Y(n11407) );
  sky130_fd_sc_hd__nor2_1 U16366 ( .A(n14983), .B(n15140), .Y(n16983) );
  sky130_fd_sc_hd__a21oi_1 U16367 ( .A1(n13374), .A2(n14980), .B1(n16983), .Y(
        n18594) );
  sky130_fd_sc_hd__nand2_1 U16368 ( .A(n18521), .B(n18660), .Y(n11379) );
  sky130_fd_sc_hd__nor4_1 U16369 ( .A(n16898), .B(n18263), .C(n16908), .D(
        n11379), .Y(n11380) );
  sky130_fd_sc_hd__a21oi_1 U16370 ( .A1(n18594), .A2(n11380), .B1(n18779), .Y(
        n11388) );
  sky130_fd_sc_hd__nand2_1 U16371 ( .A(n18698), .B(n18660), .Y(n18597) );
  sky130_fd_sc_hd__nor2_1 U16372 ( .A(n18673), .B(n18597), .Y(n15152) );
  sky130_fd_sc_hd__a31oi_1 U16373 ( .A1(n11381), .A2(n15152), .A3(n18593), 
        .B1(n18771), .Y(n11387) );
  sky130_fd_sc_hd__nand2_1 U16374 ( .A(n16916), .B(n18588), .Y(n11382) );
  sky130_fd_sc_hd__nor4_1 U16375 ( .A(n16898), .B(n18674), .C(n16976), .D(
        n11382), .Y(n11385) );
  sky130_fd_sc_hd__nor2_1 U16376 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .B(n17799), .Y(n18702) );
  sky130_fd_sc_hd__nand2_1 U16377 ( .A(n11383), .B(n13014), .Y(n18522) );
  sky130_fd_sc_hd__nor2_1 U16378 ( .A(n16968), .B(n16987), .Y(n18267) );
  sky130_fd_sc_hd__nand3_1 U16379 ( .A(n18267), .B(n16916), .C(n18588), .Y(
        n18294) );
  sky130_fd_sc_hd__nor4_1 U16380 ( .A(n18687), .B(n18674), .C(n18702), .D(
        n18294), .Y(n11384) );
  sky130_fd_sc_hd__o22ai_1 U16381 ( .A1(n11385), .A2(n18792), .B1(n11384), 
        .B2(n18783), .Y(n11386) );
  sky130_fd_sc_hd__nor3_1 U16382 ( .A(n11388), .B(n11387), .C(n11386), .Y(
        n11405) );
  sky130_fd_sc_hd__a22oi_1 U16383 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[229]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[197]), .Y(n11393) );
  sky130_fd_sc_hd__a22oi_1 U16384 ( .A1(n18734), .A2(
        j202_soc_core_memory0_ram_dout0[133]), .B1(n18733), .B2(
        j202_soc_core_memory0_ram_dout0[101]), .Y(n11392) );
  sky130_fd_sc_hd__a22oi_1 U16385 ( .A1(n18361), .A2(
        j202_soc_core_memory0_ram_dout0[37]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[69]), .Y(n11391) );
  sky130_fd_sc_hd__nand2_1 U16386 ( .A(n18735), .B(
        j202_soc_core_memory0_ram_dout0[165]), .Y(n11390) );
  sky130_fd_sc_hd__nand4_1 U16387 ( .A(n11393), .B(n11392), .C(n11391), .D(
        n11390), .Y(n11394) );
  sky130_fd_sc_hd__a21oi_1 U16388 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[5]), .B1(n11394), .Y(n11402) );
  sky130_fd_sc_hd__a22oi_1 U16389 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[293]), .B1(n18062), .B2(
        j202_soc_core_memory0_ram_dout0[261]), .Y(n11401) );
  sky130_fd_sc_hd__nand2_1 U16390 ( .A(n18743), .B(
        j202_soc_core_memory0_ram_dout0[357]), .Y(n11398) );
  sky130_fd_sc_hd__a21oi_1 U16391 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[453]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n11397) );
  sky130_fd_sc_hd__nand2_1 U16392 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[389]), .Y(n11396) );
  sky130_fd_sc_hd__nand2_1 U16393 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[421]), .Y(n11395) );
  sky130_fd_sc_hd__nand4_1 U16394 ( .A(n11398), .B(n11397), .C(n11396), .D(
        n11395), .Y(n11399) );
  sky130_fd_sc_hd__a21oi_1 U16395 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[325]), .B1(n11399), .Y(n11400) );
  sky130_fd_sc_hd__o211ai_1 U16396 ( .A1(n18736), .A2(n11402), .B1(n11401), 
        .C1(n11400), .Y(n11403) );
  sky130_fd_sc_hd__o21ai_1 U16397 ( .A1(j202_soc_core_memory0_ram_dout0[485]), 
        .A2(n18758), .B1(n11403), .Y(n11404) );
  sky130_fd_sc_hd__o22ai_1 U16398 ( .A1(n11405), .A2(n18722), .B1(n18761), 
        .B2(n11404), .Y(n11406) );
  sky130_fd_sc_hd__nor4_1 U16399 ( .A(n11409), .B(n11408), .C(n11407), .D(
        n11406), .Y(n11418) );
  sky130_fd_sc_hd__nand3_1 U16400 ( .A(n11430), .B(n18277), .C(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[0]), .Y(n18276) );
  sky130_fd_sc_hd__nor2_1 U16401 ( .A(n11410), .B(n18276), .Y(n18724) );
  sky130_fd_sc_hd__nor2_1 U16402 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[0]), 
        .B(n25203), .Y(n18242) );
  sky130_fd_sc_hd__nor2_1 U16403 ( .A(n25206), .B(n25203), .Y(n18243) );
  sky130_fd_sc_hd__a22oi_1 U16404 ( .A1(n18242), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[13]), .B1(n18243), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[5]), .Y(n11412) );
  sky130_fd_sc_hd__nand2_1 U16405 ( .A(n25203), .B(
        j202_soc_core_uart_TOP_rx_fifo_rp[0]), .Y(n25202) );
  sky130_fd_sc_hd__nor2_1 U16406 ( .A(j202_soc_core_uart_TOP_rx_fifo_rp[0]), 
        .B(j202_soc_core_uart_TOP_rx_fifo_rp[1]), .Y(n18241) );
  sky130_fd_sc_hd__a22oi_1 U16407 ( .A1(n18244), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[21]), .B1(n18241), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[29]), .Y(n11411) );
  sky130_fd_sc_hd__a21oi_1 U16408 ( .A1(n11412), .A2(n11411), .B1(n18245), .Y(
        n11413) );
  sky130_fd_sc_hd__a21oi_1 U16409 ( .A1(n18724), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[101]), .B1(n11413), .Y(
        n11416) );
  sky130_fd_sc_hd__a22oi_1 U16410 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[5]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[37]), .Y(n11415) );
  sky130_fd_sc_hd__a22oi_1 U16411 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[69]), .B1(n18629), .B2(
        j202_soc_core_bldc_core_00_pwm_period[5]), .Y(n11414) );
  sky130_fd_sc_hd__and3_1 U16412 ( .A(n11416), .B(n11415), .C(n11414), .X(
        n11417) );
  sky130_fd_sc_hd__nand2_1 U16413 ( .A(n11418), .B(n11417), .Y(n25255) );
  sky130_fd_sc_hd__nor2_1 U16414 ( .A(j202_soc_core_j22_cpu_id_op2_v_), .B(
        n22807), .Y(n11420) );
  sky130_fd_sc_hd__nand2_1 U16415 ( .A(n25255), .B(n19087), .Y(n11422) );
  sky130_fd_sc_hd__nor2b_1 U16416 ( .B_N(j202_soc_core_j22_cpu_id_opn_v_), .A(
        j202_soc_core_j22_cpu_id_op2_v_), .Y(n19088) );
  sky130_fd_sc_hd__a22oi_1 U16417 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__5_), .B1(n19088), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__5_), .Y(n11421) );
  sky130_fd_sc_hd__nand3_1 U16418 ( .A(n11423), .B(n11422), .C(n11421), .Y(
        n25382) );
  sky130_fd_sc_hd__clkinv_1 U16419 ( .A(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[1]), .Y(n20429) );
  sky130_fd_sc_hd__clkinv_1 U16420 ( .A(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[2]), .Y(n11425) );
  sky130_fd_sc_hd__o22ai_1 U16421 ( .A1(n20429), .A2(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[1]), .B1(n11425), 
        .B2(j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[2]), .Y(n11424) );
  sky130_fd_sc_hd__a221oi_1 U16422 ( .A1(n20429), .A2(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[1]), .B1(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[2]), .B2(n11425), 
        .C1(n11424), .Y(n11426) );
  sky130_fd_sc_hd__nand3_1 U16423 ( .A(n11426), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[0]), .C(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[0]), .Y(n25243) );
  sky130_fd_sc_hd__nor3b_1 U16424 ( .C_N(n11426), .A(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_1[0]), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[0]), .Y(n11427) );
  sky130_fd_sc_hd__o21ai_1 U16425 ( .A1(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[1]), .A2(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[2]), .B1(n11427), 
        .Y(n25241) );
  sky130_fd_sc_hd__nand2_1 U16426 ( .A(n25243), .B(n25241), .Y(n25406) );
  sky130_fd_sc_hd__nor2_1 U16427 ( .A(j202_soc_core_qspi_wb_ack), .B(n20103), 
        .Y(n23289) );
  sky130_fd_sc_hd__nor2_1 U16429 ( .A(j202_soc_core_ahb2apb_02_state[0]), .B(
        j202_soc_core_ahb2apb_02_state[1]), .Y(n21219) );
  sky130_fd_sc_hd__nand2_1 U16430 ( .A(n21219), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[2]), .Y(n11429) );
  sky130_fd_sc_hd__nand4_1 U16431 ( .A(n11429), .B(n18283), .C(n18288), .D(
        n11428), .Y(n11435) );
  sky130_fd_sc_hd__nand2_1 U16432 ( .A(n22767), .B(n22764), .Y(n22763) );
  sky130_fd_sc_hd__nand2_1 U16433 ( .A(n22763), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[0]), .Y(n11431) );
  sky130_fd_sc_hd__nand2_1 U16434 ( .A(n11431), .B(n11430), .Y(n11433) );
  sky130_fd_sc_hd__nor2_1 U16435 ( .A(j202_soc_core_ahb2apb_01_state[0]), .B(
        j202_soc_core_ahb2apb_01_state[1]), .Y(n21225) );
  sky130_fd_sc_hd__nand2_1 U16436 ( .A(n21225), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[1]), .Y(n11432) );
  sky130_fd_sc_hd__a21oi_1 U16437 ( .A1(n11433), .A2(n11432), .B1(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[2]), .Y(n11434) );
  sky130_fd_sc_hd__o22a_1 U16438 ( .A1(n10536), .A2(n18288), .B1(n11435), .B2(
        n11434), .X(n11437) );
  sky130_fd_sc_hd__nand2_1 U16439 ( .A(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[6]), .B(j202_soc_core_bootrom_00_sel_w), .Y(n11436) );
  sky130_fd_sc_hd__nand2_1 U16440 ( .A(n22715), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n12904) );
  sky130_fd_sc_hd__nand2_1 U16441 ( .A(n11438), .B(n22790), .Y(n12903) );
  sky130_fd_sc_hd__nor2_1 U16442 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[3]), 
        .B(n16652), .Y(n13093) );
  sky130_fd_sc_hd__nand2_1 U16443 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n22589) );
  sky130_fd_sc_hd__and3_1 U16444 ( .A(n12903), .B(n11439), .C(n22589), .X(
        n12113) );
  sky130_fd_sc_hd__nor2_1 U16445 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[2]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[4]), .Y(n22706) );
  sky130_fd_sc_hd__nand2_1 U16446 ( .A(n22706), .B(n16664), .Y(n22694) );
  sky130_fd_sc_hd__nand2_1 U16447 ( .A(n22706), .B(n22715), .Y(n11440) );
  sky130_fd_sc_hd__o21a_1 U16448 ( .A1(j202_soc_core_j22_cpu_exuop_EXU_[0]), 
        .A2(n22694), .B1(n11440), .X(n12112) );
  sky130_fd_sc_hd__nand2_1 U16449 ( .A(n22697), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[1]), .Y(n20836) );
  sky130_fd_sc_hd__nor2_1 U16450 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .B(n22790), .Y(n11441) );
  sky130_fd_sc_hd__nand3_1 U16451 ( .A(n16663), .B(n11441), .C(n22670), .Y(
        n12114) );
  sky130_fd_sc_hd__nand3_1 U16452 ( .A(n12113), .B(n12112), .C(n12114), .Y(
        n11511) );
  sky130_fd_sc_hd__nand3_1 U16453 ( .A(n16652), .B(n22790), .C(
        j202_soc_core_j22_cpu_exuop_EXU_[1]), .Y(n22691) );
  sky130_fd_sc_hd__nand2_1 U16454 ( .A(n22691), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[3]), .Y(n11442) );
  sky130_fd_sc_hd__o21ai_1 U16455 ( .A1(n22715), .A2(n22697), .B1(n11442), .Y(
        n11444) );
  sky130_fd_sc_hd__nor2_1 U16456 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .B(n22697), .Y(n22428) );
  sky130_fd_sc_hd__nand2_1 U16457 ( .A(n22428), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[0]), .Y(n11443) );
  sky130_fd_sc_hd__nand2_1 U16458 ( .A(n11443), .B(n22670), .Y(n12120) );
  sky130_fd_sc_hd__nor2_1 U16459 ( .A(n11444), .B(n12120), .Y(n11568) );
  sky130_fd_sc_hd__nor2_1 U16460 ( .A(j202_soc_core_j22_cpu_regop_Ra__1_), .B(
        n12971), .Y(n12920) );
  sky130_fd_sc_hd__nor2_1 U16461 ( .A(j202_soc_core_j22_cpu_regop_Rn__0_), .B(
        n11446), .Y(n11460) );
  sky130_fd_sc_hd__nor2_1 U16462 ( .A(j202_soc_core_j22_cpu_regop_Rn__3_), .B(
        n11447), .Y(n11474) );
  sky130_fd_sc_hd__nand2_1 U16463 ( .A(n11460), .B(n11474), .Y(n20297) );
  sky130_fd_sc_hd__nand2_1 U16464 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[214]), .Y(n11453) );
  sky130_fd_sc_hd__nor2_1 U16465 ( .A(j202_soc_core_j22_cpu_regop_Rn__2_), .B(
        j202_soc_core_j22_cpu_regop_Rn__3_), .Y(n11467) );
  sky130_fd_sc_hd__nand2_1 U16466 ( .A(n11461), .B(n11467), .Y(n20291) );
  sky130_fd_sc_hd__nand2_1 U16467 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[54]), .Y(n11452) );
  sky130_fd_sc_hd__nand2_1 U16468 ( .A(n11473), .B(n11467), .Y(n20294) );
  sky130_fd_sc_hd__nand2_1 U16469 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[118]), .Y(n11451) );
  sky130_fd_sc_hd__nor2_1 U16470 ( .A(j202_soc_core_j22_cpu_regop_Rn__2_), .B(
        n11449), .Y(n11462) );
  sky130_fd_sc_hd__nand2_1 U16471 ( .A(n11462), .B(n11473), .Y(n20280) );
  sky130_fd_sc_hd__nand2_1 U16472 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[374]), .Y(n11450) );
  sky130_fd_sc_hd__nand4_1 U16473 ( .A(n11453), .B(n11452), .C(n11451), .D(
        n11450), .Y(n11459) );
  sky130_fd_sc_hd__nand2_1 U16474 ( .A(n11460), .B(n11467), .Y(n20272) );
  sky130_fd_sc_hd__nand2_1 U16475 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[86]), .Y(n11457) );
  sky130_fd_sc_hd__nand2_1 U16476 ( .A(n11474), .B(n11461), .Y(n20302) );
  sky130_fd_sc_hd__nand2_1 U16477 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[182]), .Y(n11456) );
  sky130_fd_sc_hd__nor2_1 U16478 ( .A(j202_soc_core_j22_cpu_regop_Rn__1_), .B(
        j202_soc_core_j22_cpu_regop_Rn__0_), .Y(n11475) );
  sky130_fd_sc_hd__nand2_1 U16479 ( .A(n11474), .B(n11475), .Y(n20266) );
  sky130_fd_sc_hd__nand2_1 U16480 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[150]), .Y(n11455) );
  sky130_fd_sc_hd__nand2_1 U16481 ( .A(n11460), .B(n11476), .Y(n20289) );
  sky130_fd_sc_hd__nand2_1 U16482 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[470]), .Y(n11454) );
  sky130_fd_sc_hd__nand4_1 U16483 ( .A(n11457), .B(n11456), .C(n11455), .D(
        n11454), .Y(n11458) );
  sky130_fd_sc_hd__nor2_1 U16484 ( .A(n11459), .B(n11458), .Y(n11486) );
  sky130_fd_sc_hd__nand2_1 U16485 ( .A(n11462), .B(n11461), .Y(n20283) );
  sky130_fd_sc_hd__nand2_1 U16486 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[310]), .Y(n11466) );
  sky130_fd_sc_hd__nand2_1 U16487 ( .A(n11460), .B(n11462), .Y(n20305) );
  sky130_fd_sc_hd__nand2_1 U16488 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[342]), .Y(n11465) );
  sky130_fd_sc_hd__nand2_1 U16489 ( .A(n11461), .B(n11476), .Y(n20286) );
  sky130_fd_sc_hd__nand2_1 U16490 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[438]), .Y(n11464) );
  sky130_fd_sc_hd__nand2_1 U16491 ( .A(n11462), .B(n11475), .Y(n20258) );
  sky130_fd_sc_hd__nand2_1 U16492 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[278]), .Y(n11463) );
  sky130_fd_sc_hd__and4_1 U16493 ( .A(n11466), .B(n11465), .C(n11464), .D(
        n11463), .X(n11485) );
  sky130_fd_sc_hd__nand2_1 U16494 ( .A(n11475), .B(n11467), .Y(n20249) );
  sky130_fd_sc_hd__nand2_1 U16495 ( .A(n20249), .B(n12042), .Y(n11468) );
  sky130_fd_sc_hd__nor2_1 U16496 ( .A(n11469), .B(n13919), .Y(n11483) );
  sky130_fd_sc_hd__nand2_1 U16497 ( .A(n12042), .B(n21399), .Y(n11471) );
  sky130_fd_sc_hd__nand2_1 U16498 ( .A(n11471), .B(n12971), .Y(n12539) );
  sky130_fd_sc_hd__nor2_1 U16499 ( .A(n11472), .B(n12539), .Y(n13920) );
  sky130_fd_sc_hd__a21oi_1 U16500 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[22]), .B1(n13920), .Y(n11481) );
  sky130_fd_sc_hd__nand2_1 U16501 ( .A(n11476), .B(n11473), .Y(n20241) );
  sky130_fd_sc_hd__nand2_1 U16502 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[502]), .Y(n11480) );
  sky130_fd_sc_hd__nand2_1 U16503 ( .A(n11474), .B(n11473), .Y(n20299) );
  sky130_fd_sc_hd__nand2_1 U16504 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[246]), .Y(n11479) );
  sky130_fd_sc_hd__nand2_1 U16505 ( .A(n11476), .B(n11475), .Y(n20261) );
  sky130_fd_sc_hd__nand2_1 U16506 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[406]), .Y(n11478) );
  sky130_fd_sc_hd__nand4_1 U16507 ( .A(n11481), .B(n11480), .C(n11479), .D(
        n11478), .Y(n11482) );
  sky130_fd_sc_hd__nor2_1 U16508 ( .A(n11483), .B(n11482), .Y(n11484) );
  sky130_fd_sc_hd__nand3_1 U16509 ( .A(n11486), .B(n11485), .C(n11484), .Y(
        n21867) );
  sky130_fd_sc_hd__nand2_1 U16510 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[245]), .Y(n11490) );
  sky130_fd_sc_hd__nand2_1 U16511 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[53]), .Y(n11489) );
  sky130_fd_sc_hd__nand2_1 U16512 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[117]), .Y(n11488) );
  sky130_fd_sc_hd__nand2_1 U16513 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[501]), .Y(n11487) );
  sky130_fd_sc_hd__nand4_1 U16514 ( .A(n11490), .B(n11489), .C(n11488), .D(
        n11487), .Y(n11496) );
  sky130_fd_sc_hd__nand2_1 U16515 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[437]), .Y(n11494) );
  sky130_fd_sc_hd__nand2_1 U16516 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[341]), .Y(n11493) );
  sky130_fd_sc_hd__nand2_1 U16517 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[469]), .Y(n11492) );
  sky130_fd_sc_hd__nand2_1 U16518 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[277]), .Y(n11491) );
  sky130_fd_sc_hd__nand4_1 U16519 ( .A(n11494), .B(n11493), .C(n11492), .D(
        n11491), .Y(n11495) );
  sky130_fd_sc_hd__nor2_1 U16520 ( .A(n11496), .B(n11495), .Y(n11510) );
  sky130_fd_sc_hd__nor2_1 U16521 ( .A(n11497), .B(n13919), .Y(n11503) );
  sky130_fd_sc_hd__a21oi_1 U16522 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[21]), .B1(n13920), .Y(n11501) );
  sky130_fd_sc_hd__nand2_1 U16523 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[181]), .Y(n11500) );
  sky130_fd_sc_hd__nand2_1 U16524 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[149]), .Y(n11499) );
  sky130_fd_sc_hd__nand2_1 U16525 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[309]), .Y(n11498) );
  sky130_fd_sc_hd__nand4_1 U16526 ( .A(n11501), .B(n11500), .C(n11499), .D(
        n11498), .Y(n11502) );
  sky130_fd_sc_hd__nor2_1 U16527 ( .A(n11503), .B(n11502), .Y(n11509) );
  sky130_fd_sc_hd__nand2_1 U16528 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[213]), .Y(n11507) );
  sky130_fd_sc_hd__nand2_1 U16529 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[373]), .Y(n11506) );
  sky130_fd_sc_hd__nand2_1 U16530 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[405]), .Y(n11505) );
  sky130_fd_sc_hd__nand2_1 U16531 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[85]), .Y(n11504) );
  sky130_fd_sc_hd__and4_1 U16532 ( .A(n11507), .B(n11506), .C(n11505), .D(
        n11504), .X(n11508) );
  sky130_fd_sc_hd__nand3_1 U16533 ( .A(n11510), .B(n11509), .C(n11508), .Y(
        n22578) );
  sky130_fd_sc_hd__nand2_1 U16534 ( .A(n16652), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[3]), .Y(n14042) );
  sky130_fd_sc_hd__o22ai_1 U16535 ( .A1(n20677), .A2(n22567), .B1(n22600), 
        .B2(n14042), .Y(n12788) );
  sky130_fd_sc_hd__xor2_1 U16536 ( .A(j202_soc_core_j22_cpu_rfuo_sr__q_), .B(
        j202_soc_core_j22_cpu_rfuo_sr__m_), .X(n11566) );
  sky130_fd_sc_hd__nand2_1 U16537 ( .A(n11566), .B(n13681), .Y(n12111) );
  sky130_fd_sc_hd__nand2_1 U16538 ( .A(n11529), .B(
        j202_soc_core_j22_cpu_regop_Rm__0_), .Y(n11514) );
  sky130_fd_sc_hd__nor2_1 U16539 ( .A(j202_soc_core_j22_cpu_regop_Rm__3_), .B(
        n11520), .Y(n11535) );
  sky130_fd_sc_hd__nand2_1 U16541 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[182]), .Y(n11518) );
  sky130_fd_sc_hd__nand2_1 U16542 ( .A(j202_soc_core_j22_cpu_regop_Rm__0_), 
        .B(j202_soc_core_j22_cpu_regop_Rm__1_), .Y(n11513) );
  sky130_fd_sc_hd__nand2_1 U16543 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[246]), .Y(n11517) );
  sky130_fd_sc_hd__nand2_1 U16544 ( .A(j202_soc_core_j22_cpu_regop_Rm__2_), 
        .B(j202_soc_core_j22_cpu_regop_Rm__3_), .Y(n11522) );
  sky130_fd_sc_hd__nor2_1 U16545 ( .A(n11513), .B(n11522), .Y(n20238) );
  sky130_fd_sc_hd__nand2_1 U16546 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[502]), .Y(n11516) );
  sky130_fd_sc_hd__nand2_1 U16548 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[438]), .Y(n11515) );
  sky130_fd_sc_hd__nand4_1 U16549 ( .A(n11518), .B(n11517), .C(n11516), .D(
        n11515), .Y(n11528) );
  sky130_fd_sc_hd__nor2_1 U16550 ( .A(j202_soc_core_j22_cpu_regop_Rm__1_), .B(
        j202_soc_core_j22_cpu_regop_Rm__0_), .Y(n11541) );
  sky130_fd_sc_hd__nand2_1 U16551 ( .A(n11519), .B(n11541), .Y(n20260) );
  sky130_fd_sc_hd__nand2_1 U16552 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[406]), .Y(n11526) );
  sky130_fd_sc_hd__nor2_1 U16553 ( .A(j202_soc_core_j22_cpu_regop_Rm__3_), .B(
        j202_soc_core_j22_cpu_regop_Rm__2_), .Y(n11536) );
  sky130_fd_sc_hd__nand2_1 U16554 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[22]), .Y(n11525) );
  sky130_fd_sc_hd__nand2_1 U16555 ( .A(n11529), .B(n11538), .Y(n11521) );
  sky130_fd_sc_hd__nand2_1 U16556 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[54]), .Y(n11524) );
  sky130_fd_sc_hd__nand2_1 U16557 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[470]), .Y(n11523) );
  sky130_fd_sc_hd__nand4_1 U16558 ( .A(n11526), .B(n11525), .C(n11524), .D(
        n11523), .Y(n11527) );
  sky130_fd_sc_hd__nor2_1 U16559 ( .A(n11528), .B(n11527), .Y(n11550) );
  sky130_fd_sc_hd__nand2_1 U16560 ( .A(n11529), .B(
        j202_soc_core_j22_cpu_regop_Rm__3_), .Y(n11530) );
  sky130_fd_sc_hd__a22oi_1 U16562 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[310]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[214]), .Y(n11549) );
  sky130_fd_sc_hd__nand2_1 U16563 ( .A(j202_soc_core_j22_cpu_regop_Rm__1_), 
        .B(j202_soc_core_j22_cpu_regop_Rm__3_), .Y(n11532) );
  sky130_fd_sc_hd__nor2_1 U16565 ( .A(j202_soc_core_j22_cpu_regop_Rm__2_), .B(
        n11538), .Y(n11542) );
  sky130_fd_sc_hd__a22oi_1 U16566 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[374]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[342]), .Y(n11548) );
  sky130_fd_sc_hd__nand2_1 U16567 ( .A(n11535), .B(n11541), .Y(n20265) );
  sky130_fd_sc_hd__nand2_1 U16568 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[150]), .Y(n11546) );
  sky130_fd_sc_hd__nand2_1 U16569 ( .A(n11537), .B(n11536), .Y(n20270) );
  sky130_fd_sc_hd__nand2_1 U16570 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[86]), .Y(n11545) );
  sky130_fd_sc_hd__nand2_1 U16571 ( .A(n11538), .B(
        j202_soc_core_j22_cpu_regop_Rm__1_), .Y(n11540) );
  sky130_fd_sc_hd__nand2_1 U16572 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[118]), .Y(n11544) );
  sky130_fd_sc_hd__nand2_1 U16573 ( .A(n11542), .B(n11541), .Y(n20257) );
  sky130_fd_sc_hd__nand2_1 U16574 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[278]), .Y(n11543) );
  sky130_fd_sc_hd__and4_1 U16575 ( .A(n11546), .B(n11545), .C(n11544), .D(
        n11543), .X(n11547) );
  sky130_fd_sc_hd__nand4_1 U16576 ( .A(n11550), .B(n11549), .C(n11548), .D(
        n11547), .Y(n19544) );
  sky130_fd_sc_hd__nand2_1 U16577 ( .A(n19544), .B(n14086), .Y(n11565) );
  sky130_fd_sc_hd__nand2_1 U16578 ( .A(j202_soc_core_j22_cpu_regop_Rb__0_), 
        .B(j202_soc_core_j22_cpu_regop_Rb__1_), .Y(n11555) );
  sky130_fd_sc_hd__nor2_1 U16579 ( .A(j202_soc_core_j22_cpu_regop_other__0_), 
        .B(n12941), .Y(n12940) );
  sky130_fd_sc_hd__nand2_1 U16580 ( .A(n12940), .B(
        j202_soc_core_j22_cpu_regop_other__2_), .Y(n15213) );
  sky130_fd_sc_hd__nor2_1 U16581 ( .A(n11555), .B(n15213), .Y(n14069) );
  sky130_fd_sc_hd__nand2_1 U16582 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[22]), .Y(n11554) );
  sky130_fd_sc_hd__nand2_1 U16583 ( .A(j202_soc_core_j22_cpu_regop_other__2_), 
        .B(j202_soc_core_j22_cpu_regop_other__0_), .Y(n12019) );
  sky130_fd_sc_hd__nor2_1 U16584 ( .A(n12941), .B(n12019), .Y(n15219) );
  sky130_fd_sc_hd__nand2_1 U16585 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[22]), .Y(n11553) );
  sky130_fd_sc_hd__nor2_1 U16586 ( .A(j202_soc_core_j22_cpu_regop_Rb__0_), .B(
        n14086), .Y(n11551) );
  sky130_fd_sc_hd__nand2_1 U16587 ( .A(n11551), .B(
        j202_soc_core_j22_cpu_regop_imm__12_), .Y(n14022) );
  sky130_fd_sc_hd__nor2_1 U16588 ( .A(j202_soc_core_j22_cpu_regop_other__1_), 
        .B(j202_soc_core_j22_cpu_regop_other__0_), .Y(n15215) );
  sky130_fd_sc_hd__nand2_1 U16589 ( .A(n15215), .B(
        j202_soc_core_j22_cpu_regop_other__2_), .Y(n15221) );
  sky130_fd_sc_hd__nor2_1 U16590 ( .A(n11555), .B(n15221), .Y(n14072) );
  sky130_fd_sc_hd__nand2_1 U16591 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[502]), .Y(n11552) );
  sky130_fd_sc_hd__and4_1 U16592 ( .A(n11554), .B(n11553), .C(n14022), .D(
        n11552), .X(n11564) );
  sky130_fd_sc_hd__nor2_1 U16593 ( .A(j202_soc_core_j22_cpu_regop_other__2_), 
        .B(n11555), .Y(n11558) );
  sky130_fd_sc_hd__nand2_1 U16594 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[22]), .Y(n11562) );
  sky130_fd_sc_hd__nor2_1 U16595 ( .A(j202_soc_core_j22_cpu_regop_other__1_), 
        .B(n11556), .Y(n15212) );
  sky130_fd_sc_hd__nand2_1 U16596 ( .A(n14025), .B(
        j202_soc_core_j22_cpu_pc[22]), .Y(n11561) );
  sky130_fd_sc_hd__nand2_1 U16597 ( .A(j202_soc_core_j22_cpu_regop_other__0_), 
        .B(j202_soc_core_j22_cpu_regop_other__1_), .Y(n12916) );
  sky130_fd_sc_hd__nand2_1 U16598 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[22]), .Y(n11560) );
  sky130_fd_sc_hd__nand2_1 U16599 ( .A(n11558), .B(n15215), .Y(n14077) );
  sky130_fd_sc_hd__nand2_1 U16600 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[22]), .Y(n11559) );
  sky130_fd_sc_hd__and4_1 U16601 ( .A(n11562), .B(n11561), .C(n11560), .D(
        n11559), .X(n11563) );
  sky130_fd_sc_hd__nand3_1 U16602 ( .A(n11565), .B(n11564), .C(n11563), .Y(
        n23316) );
  sky130_fd_sc_hd__nand2_1 U16603 ( .A(n11567), .B(n13681), .Y(n12116) );
  sky130_fd_sc_hd__nand2_1 U16604 ( .A(n11568), .B(n12116), .Y(n14087) );
  sky130_fd_sc_hd__nand2_1 U16605 ( .A(n21878), .B(n14087), .Y(n11569) );
  sky130_fd_sc_hd__o21ai_1 U16606 ( .A1(n14089), .A2(n21878), .B1(n11569), .Y(
        n12789) );
  sky130_fd_sc_hd__nor2_1 U16607 ( .A(n12788), .B(n12789), .Y(n13293) );
  sky130_fd_sc_hd__nand2_1 U16608 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[243]), .Y(n11573) );
  sky130_fd_sc_hd__nand2_1 U16609 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[371]), .Y(n11572) );
  sky130_fd_sc_hd__nand2_1 U16610 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[115]), .Y(n11571) );
  sky130_fd_sc_hd__nand2_1 U16611 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[499]), .Y(n11570) );
  sky130_fd_sc_hd__nand4_1 U16612 ( .A(n11573), .B(n11572), .C(n11571), .D(
        n11570), .Y(n11579) );
  sky130_fd_sc_hd__nand2_1 U16613 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[147]), .Y(n11577) );
  sky130_fd_sc_hd__nand2_1 U16614 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[339]), .Y(n11576) );
  sky130_fd_sc_hd__nand2_1 U16615 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[467]), .Y(n11575) );
  sky130_fd_sc_hd__nand2_1 U16616 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[435]), .Y(n11574) );
  sky130_fd_sc_hd__nand4_1 U16617 ( .A(n11577), .B(n11576), .C(n11575), .D(
        n11574), .Y(n11578) );
  sky130_fd_sc_hd__nor2_1 U16618 ( .A(n11579), .B(n11578), .Y(n11593) );
  sky130_fd_sc_hd__nor2_1 U16619 ( .A(n11580), .B(n13919), .Y(n11586) );
  sky130_fd_sc_hd__a21oi_1 U16620 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[19]), .B1(n13920), .Y(n11584) );
  sky130_fd_sc_hd__nand2_1 U16621 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[179]), .Y(n11583) );
  sky130_fd_sc_hd__nand2_1 U16622 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[83]), .Y(n11582) );
  sky130_fd_sc_hd__nand2_1 U16623 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[51]), .Y(n11581) );
  sky130_fd_sc_hd__nand4_1 U16624 ( .A(n11584), .B(n11583), .C(n11582), .D(
        n11581), .Y(n11585) );
  sky130_fd_sc_hd__nor2_1 U16625 ( .A(n11586), .B(n11585), .Y(n11592) );
  sky130_fd_sc_hd__nand2_1 U16626 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[211]), .Y(n11590) );
  sky130_fd_sc_hd__nand2_1 U16627 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[307]), .Y(n11589) );
  sky130_fd_sc_hd__nand2_1 U16628 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[403]), .Y(n11588) );
  sky130_fd_sc_hd__nand2_1 U16629 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[275]), .Y(n11587) );
  sky130_fd_sc_hd__and4_1 U16630 ( .A(n11590), .B(n11589), .C(n11588), .D(
        n11587), .X(n11591) );
  sky130_fd_sc_hd__nand3_1 U16631 ( .A(n11593), .B(n11592), .C(n11591), .Y(
        n21963) );
  sky130_fd_sc_hd__nand2_1 U16632 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[148]), .Y(n11597) );
  sky130_fd_sc_hd__nand2_1 U16633 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[308]), .Y(n11596) );
  sky130_fd_sc_hd__nand2_1 U16634 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[276]), .Y(n11595) );
  sky130_fd_sc_hd__nand2_1 U16635 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[468]), .Y(n11594) );
  sky130_fd_sc_hd__nand4_1 U16636 ( .A(n11597), .B(n11596), .C(n11595), .D(
        n11594), .Y(n11603) );
  sky130_fd_sc_hd__nand2_1 U16637 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[244]), .Y(n11601) );
  sky130_fd_sc_hd__nand2_1 U16638 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[340]), .Y(n11600) );
  sky130_fd_sc_hd__nand2_1 U16639 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[52]), .Y(n11599) );
  sky130_fd_sc_hd__nand2_1 U16640 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[84]), .Y(n11598) );
  sky130_fd_sc_hd__nand4_1 U16641 ( .A(n11601), .B(n11600), .C(n11599), .D(
        n11598), .Y(n11602) );
  sky130_fd_sc_hd__nor2_1 U16642 ( .A(n11603), .B(n11602), .Y(n11617) );
  sky130_fd_sc_hd__nand2_1 U16643 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[212]), .Y(n11607) );
  sky130_fd_sc_hd__nand2_1 U16644 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[180]), .Y(n11606) );
  sky130_fd_sc_hd__nand2_1 U16645 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[404]), .Y(n11605) );
  sky130_fd_sc_hd__nand2_1 U16646 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[116]), .Y(n11604) );
  sky130_fd_sc_hd__and4_1 U16647 ( .A(n11607), .B(n11606), .C(n11605), .D(
        n11604), .X(n11616) );
  sky130_fd_sc_hd__nor2_1 U16648 ( .A(n11608), .B(n13919), .Y(n11614) );
  sky130_fd_sc_hd__a21oi_1 U16649 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[20]), .B1(n13920), .Y(n11612) );
  sky130_fd_sc_hd__nand2_1 U16650 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[372]), .Y(n11611) );
  sky130_fd_sc_hd__nand2_1 U16651 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[500]), .Y(n11610) );
  sky130_fd_sc_hd__nand2_1 U16652 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[436]), .Y(n11609) );
  sky130_fd_sc_hd__nand4_1 U16653 ( .A(n11612), .B(n11611), .C(n11610), .D(
        n11609), .Y(n11613) );
  sky130_fd_sc_hd__nor2_1 U16654 ( .A(n11614), .B(n11613), .Y(n11615) );
  sky130_fd_sc_hd__nand3_1 U16655 ( .A(n11617), .B(n11616), .C(n11615), .Y(
        n22577) );
  sky130_fd_sc_hd__o22ai_1 U16656 ( .A1(n14042), .A2(n22643), .B1(n22641), 
        .B2(n20677), .Y(n12754) );
  sky130_fd_sc_hd__nand2_1 U16657 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[180]), .Y(n11621) );
  sky130_fd_sc_hd__nand2_1 U16658 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[244]), .Y(n11620) );
  sky130_fd_sc_hd__nand2_1 U16659 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[500]), .Y(n11619) );
  sky130_fd_sc_hd__nand2_1 U16660 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[436]), .Y(n11618) );
  sky130_fd_sc_hd__nand4_1 U16661 ( .A(n11621), .B(n11620), .C(n11619), .D(
        n11618), .Y(n11627) );
  sky130_fd_sc_hd__nand2_1 U16662 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[404]), .Y(n11625) );
  sky130_fd_sc_hd__nand2_1 U16663 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[20]), .Y(n11624) );
  sky130_fd_sc_hd__nand2_1 U16664 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[52]), .Y(n11623) );
  sky130_fd_sc_hd__nand2_1 U16665 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[468]), .Y(n11622) );
  sky130_fd_sc_hd__nand4_1 U16666 ( .A(n11625), .B(n11624), .C(n11623), .D(
        n11622), .Y(n11626) );
  sky130_fd_sc_hd__nor2_1 U16667 ( .A(n11627), .B(n11626), .Y(n11635) );
  sky130_fd_sc_hd__a22oi_1 U16668 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[308]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[212]), .Y(n11634) );
  sky130_fd_sc_hd__a22oi_1 U16669 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[372]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[340]), .Y(n11633) );
  sky130_fd_sc_hd__nand2_1 U16670 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[148]), .Y(n11631) );
  sky130_fd_sc_hd__nand2_1 U16671 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[84]), .Y(n11630) );
  sky130_fd_sc_hd__nand2_1 U16672 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[116]), .Y(n11629) );
  sky130_fd_sc_hd__nand2_1 U16673 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[276]), .Y(n11628) );
  sky130_fd_sc_hd__and4_1 U16674 ( .A(n11631), .B(n11630), .C(n11629), .D(
        n11628), .X(n11632) );
  sky130_fd_sc_hd__nand4_1 U16675 ( .A(n11635), .B(n11634), .C(n11633), .D(
        n11632), .Y(n19417) );
  sky130_fd_sc_hd__nand2_1 U16676 ( .A(n19417), .B(n14086), .Y(n11645) );
  sky130_fd_sc_hd__nand2_1 U16677 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[20]), .Y(n11638) );
  sky130_fd_sc_hd__nand2_1 U16678 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[20]), .Y(n11637) );
  sky130_fd_sc_hd__nand2_1 U16679 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[500]), .Y(n11636) );
  sky130_fd_sc_hd__and4_1 U16680 ( .A(n11638), .B(n11637), .C(n14022), .D(
        n11636), .X(n11644) );
  sky130_fd_sc_hd__nand2_1 U16681 ( .A(n14025), .B(
        j202_soc_core_j22_cpu_pc[20]), .Y(n11642) );
  sky130_fd_sc_hd__nand2_1 U16682 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[20]), .Y(n11641) );
  sky130_fd_sc_hd__nand2_1 U16683 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[20]), .Y(n11640) );
  sky130_fd_sc_hd__nand2_1 U16684 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[20]), .Y(n11639) );
  sky130_fd_sc_hd__and4_1 U16685 ( .A(n11642), .B(n11641), .C(n11640), .D(
        n11639), .X(n11643) );
  sky130_fd_sc_hd__nand3_1 U16686 ( .A(n11645), .B(n11644), .C(n11643), .Y(
        n23310) );
  sky130_fd_sc_hd__nand2_1 U16687 ( .A(n22640), .B(n14087), .Y(n11646) );
  sky130_fd_sc_hd__nor2_1 U16689 ( .A(n12754), .B(n12755), .Y(n13403) );
  sky130_fd_sc_hd__nand2_1 U16690 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[338]), .Y(n11650) );
  sky130_fd_sc_hd__nand2_1 U16691 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[242]), .Y(n11649) );
  sky130_fd_sc_hd__nand2_1 U16692 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[498]), .Y(n11648) );
  sky130_fd_sc_hd__nand2_1 U16693 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[82]), .Y(n11647) );
  sky130_fd_sc_hd__nand4_1 U16694 ( .A(n11650), .B(n11649), .C(n11648), .D(
        n11647), .Y(n11656) );
  sky130_fd_sc_hd__nand2_1 U16695 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[210]), .Y(n11654) );
  sky130_fd_sc_hd__nand2_1 U16696 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[178]), .Y(n11653) );
  sky130_fd_sc_hd__nand2_1 U16697 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[146]), .Y(n11652) );
  sky130_fd_sc_hd__nand2_1 U16698 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[274]), .Y(n11651) );
  sky130_fd_sc_hd__nand4_1 U16699 ( .A(n11654), .B(n11653), .C(n11652), .D(
        n11651), .Y(n11655) );
  sky130_fd_sc_hd__nor2_1 U16700 ( .A(n11656), .B(n11655), .Y(n11670) );
  sky130_fd_sc_hd__nand2_1 U16701 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[306]), .Y(n11660) );
  sky130_fd_sc_hd__nand2_1 U16702 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[434]), .Y(n11659) );
  sky130_fd_sc_hd__nand2_1 U16703 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[114]), .Y(n11658) );
  sky130_fd_sc_hd__nand2_1 U16704 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[466]), .Y(n11657) );
  sky130_fd_sc_hd__and4_1 U16705 ( .A(n11660), .B(n11659), .C(n11658), .D(
        n11657), .X(n11669) );
  sky130_fd_sc_hd__nor2_1 U16706 ( .A(n11661), .B(n13919), .Y(n11667) );
  sky130_fd_sc_hd__a21oi_1 U16707 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[18]), .B1(n13920), .Y(n11665) );
  sky130_fd_sc_hd__nand2_1 U16708 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[370]), .Y(n11664) );
  sky130_fd_sc_hd__nand2_1 U16709 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[50]), .Y(n11663) );
  sky130_fd_sc_hd__nand2_1 U16710 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[402]), .Y(n11662) );
  sky130_fd_sc_hd__nand4_1 U16711 ( .A(n11665), .B(n11664), .C(n11663), .D(
        n11662), .Y(n11666) );
  sky130_fd_sc_hd__nor2_1 U16712 ( .A(n11667), .B(n11666), .Y(n11668) );
  sky130_fd_sc_hd__nand3_1 U16713 ( .A(n11670), .B(n11669), .C(n11668), .Y(
        n21775) );
  sky130_fd_sc_hd__nand2_1 U16714 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[177]), .Y(n11674) );
  sky130_fd_sc_hd__nand2_1 U16715 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[433]), .Y(n11673) );
  sky130_fd_sc_hd__nand2_1 U16716 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[497]), .Y(n11672) );
  sky130_fd_sc_hd__nand2_1 U16717 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[273]), .Y(n11671) );
  sky130_fd_sc_hd__nand4_1 U16718 ( .A(n11674), .B(n11673), .C(n11672), .D(
        n11671), .Y(n11680) );
  sky130_fd_sc_hd__nand2_1 U16719 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[337]), .Y(n11678) );
  sky130_fd_sc_hd__nand2_1 U16720 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[209]), .Y(n11677) );
  sky130_fd_sc_hd__nand2_1 U16721 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[369]), .Y(n11676) );
  sky130_fd_sc_hd__nand2_1 U16722 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[401]), .Y(n11675) );
  sky130_fd_sc_hd__nand4_1 U16723 ( .A(n11678), .B(n11677), .C(n11676), .D(
        n11675), .Y(n11679) );
  sky130_fd_sc_hd__nor2_1 U16724 ( .A(n11680), .B(n11679), .Y(n11694) );
  sky130_fd_sc_hd__nand2_1 U16725 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[305]), .Y(n11684) );
  sky130_fd_sc_hd__nand2_1 U16726 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[145]), .Y(n11683) );
  sky130_fd_sc_hd__nand2_1 U16727 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[113]), .Y(n11682) );
  sky130_fd_sc_hd__nand2_1 U16728 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[465]), .Y(n11681) );
  sky130_fd_sc_hd__and4_1 U16729 ( .A(n11684), .B(n11683), .C(n11682), .D(
        n11681), .X(n11693) );
  sky130_fd_sc_hd__nor2_1 U16730 ( .A(n11685), .B(n13919), .Y(n11691) );
  sky130_fd_sc_hd__a21oi_1 U16731 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[17]), .B1(n13920), .Y(n11689) );
  sky130_fd_sc_hd__nand2_1 U16732 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[49]), .Y(n11688) );
  sky130_fd_sc_hd__nand2_1 U16733 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[241]), .Y(n11687) );
  sky130_fd_sc_hd__nand2_1 U16734 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[81]), .Y(n11686) );
  sky130_fd_sc_hd__nand4_1 U16735 ( .A(n11689), .B(n11688), .C(n11687), .D(
        n11686), .Y(n11690) );
  sky130_fd_sc_hd__nor2_1 U16736 ( .A(n11691), .B(n11690), .Y(n11692) );
  sky130_fd_sc_hd__nand3_1 U16737 ( .A(n11694), .B(n11693), .C(n11692), .Y(
        n21683) );
  sky130_fd_sc_hd__o22ai_1 U16738 ( .A1(n20677), .A2(n22566), .B1(n22565), 
        .B2(n14042), .Y(n12720) );
  sky130_fd_sc_hd__nand2_1 U16739 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[178]), .Y(n11698) );
  sky130_fd_sc_hd__nand2_1 U16740 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[242]), .Y(n11697) );
  sky130_fd_sc_hd__nand2_1 U16741 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[498]), .Y(n11696) );
  sky130_fd_sc_hd__nand2_1 U16742 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[434]), .Y(n11695) );
  sky130_fd_sc_hd__nand4_1 U16743 ( .A(n11698), .B(n11697), .C(n11696), .D(
        n11695), .Y(n11704) );
  sky130_fd_sc_hd__nand2_1 U16744 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[402]), .Y(n11702) );
  sky130_fd_sc_hd__nand2_1 U16745 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[18]), .Y(n11701) );
  sky130_fd_sc_hd__nand2_1 U16746 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[50]), .Y(n11700) );
  sky130_fd_sc_hd__nand2_1 U16747 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[466]), .Y(n11699) );
  sky130_fd_sc_hd__nand4_1 U16748 ( .A(n11702), .B(n11701), .C(n11700), .D(
        n11699), .Y(n11703) );
  sky130_fd_sc_hd__nor2_1 U16749 ( .A(n11704), .B(n11703), .Y(n11712) );
  sky130_fd_sc_hd__a22oi_1 U16750 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[306]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[210]), .Y(n11711) );
  sky130_fd_sc_hd__a22oi_1 U16751 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[370]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[338]), .Y(n11710) );
  sky130_fd_sc_hd__nand2_1 U16752 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[146]), .Y(n11708) );
  sky130_fd_sc_hd__nand2_1 U16753 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[82]), .Y(n11707) );
  sky130_fd_sc_hd__nand2_1 U16754 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[114]), .Y(n11706) );
  sky130_fd_sc_hd__nand2_1 U16755 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[274]), .Y(n11705) );
  sky130_fd_sc_hd__and4_1 U16756 ( .A(n11708), .B(n11707), .C(n11706), .D(
        n11705), .X(n11709) );
  sky130_fd_sc_hd__nand4_1 U16757 ( .A(n11712), .B(n11711), .C(n11710), .D(
        n11709), .Y(n19460) );
  sky130_fd_sc_hd__nand2_1 U16758 ( .A(n19460), .B(n14086), .Y(n11722) );
  sky130_fd_sc_hd__nand2_1 U16759 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[18]), .Y(n11715) );
  sky130_fd_sc_hd__nand2_1 U16760 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[18]), .Y(n11714) );
  sky130_fd_sc_hd__nand2_1 U16761 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[498]), .Y(n11713) );
  sky130_fd_sc_hd__and4_1 U16762 ( .A(n11715), .B(n11714), .C(n14022), .D(
        n11713), .X(n11721) );
  sky130_fd_sc_hd__nand2_1 U16763 ( .A(n14025), .B(
        j202_soc_core_j22_cpu_pc[18]), .Y(n11719) );
  sky130_fd_sc_hd__nand2_1 U16764 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[18]), .Y(n11718) );
  sky130_fd_sc_hd__nand2_1 U16765 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[18]), .Y(n11717) );
  sky130_fd_sc_hd__nand2_1 U16766 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[18]), .Y(n11716) );
  sky130_fd_sc_hd__and4_1 U16767 ( .A(n11719), .B(n11718), .C(n11717), .D(
        n11716), .X(n11720) );
  sky130_fd_sc_hd__nand3_1 U16768 ( .A(n11722), .B(n11721), .C(n11720), .Y(
        n23304) );
  sky130_fd_sc_hd__nand2_1 U16769 ( .A(n21787), .B(n14087), .Y(n11723) );
  sky130_fd_sc_hd__nor2_1 U16771 ( .A(n12720), .B(n12721), .Y(n13541) );
  sky130_fd_sc_hd__nand2_1 U16772 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[240]), .Y(n11727) );
  sky130_fd_sc_hd__nand2_1 U16773 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[48]), .Y(n11726) );
  sky130_fd_sc_hd__nand2_1 U16774 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[112]), .Y(n11725) );
  sky130_fd_sc_hd__nand2_1 U16775 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[496]), .Y(n11724) );
  sky130_fd_sc_hd__nand4_1 U16776 ( .A(n11727), .B(n11726), .C(n11725), .D(
        n11724), .Y(n11733) );
  sky130_fd_sc_hd__nand2_1 U16777 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[144]), .Y(n11731) );
  sky130_fd_sc_hd__nand2_1 U16778 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[336]), .Y(n11730) );
  sky130_fd_sc_hd__nand2_1 U16779 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[272]), .Y(n11729) );
  sky130_fd_sc_hd__nand2_1 U16780 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[432]), .Y(n11728) );
  sky130_fd_sc_hd__nand4_1 U16781 ( .A(n11731), .B(n11730), .C(n11729), .D(
        n11728), .Y(n11732) );
  sky130_fd_sc_hd__nor2_1 U16782 ( .A(n11733), .B(n11732), .Y(n11747) );
  sky130_fd_sc_hd__nor2_1 U16783 ( .A(n11734), .B(n13919), .Y(n11740) );
  sky130_fd_sc_hd__a21oi_1 U16784 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[16]), .B1(n13920), .Y(n11738) );
  sky130_fd_sc_hd__nand2_1 U16785 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[176]), .Y(n11737) );
  sky130_fd_sc_hd__nand2_1 U16786 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[400]), .Y(n11736) );
  sky130_fd_sc_hd__nand2_1 U16787 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[80]), .Y(n11735) );
  sky130_fd_sc_hd__nand4_1 U16788 ( .A(n11738), .B(n11737), .C(n11736), .D(
        n11735), .Y(n11739) );
  sky130_fd_sc_hd__nor2_1 U16789 ( .A(n11740), .B(n11739), .Y(n11746) );
  sky130_fd_sc_hd__nand2_1 U16790 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[208]), .Y(n11744) );
  sky130_fd_sc_hd__nand2_1 U16791 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[304]), .Y(n11743) );
  sky130_fd_sc_hd__nand2_1 U16792 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[368]), .Y(n11742) );
  sky130_fd_sc_hd__nand2_1 U16793 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[464]), .Y(n11741) );
  sky130_fd_sc_hd__and4_1 U16794 ( .A(n11744), .B(n11743), .C(n11742), .D(
        n11741), .X(n11745) );
  sky130_fd_sc_hd__nand3_1 U16795 ( .A(n11747), .B(n11746), .C(n11745), .Y(
        n22133) );
  sky130_fd_sc_hd__nand2_1 U16796 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[239]), .Y(n11751) );
  sky130_fd_sc_hd__nand2_1 U16797 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[47]), .Y(n11750) );
  sky130_fd_sc_hd__nand2_1 U16798 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[111]), .Y(n11749) );
  sky130_fd_sc_hd__nand2_1 U16799 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[495]), .Y(n11748) );
  sky130_fd_sc_hd__nand4_1 U16800 ( .A(n11751), .B(n11750), .C(n11749), .D(
        n11748), .Y(n11757) );
  sky130_fd_sc_hd__nand2_1 U16801 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[207]), .Y(n11755) );
  sky130_fd_sc_hd__nand2_1 U16802 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[303]), .Y(n11754) );
  sky130_fd_sc_hd__nand2_1 U16803 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[431]), .Y(n11753) );
  sky130_fd_sc_hd__nand2_1 U16804 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[463]), .Y(n11752) );
  sky130_fd_sc_hd__nand4_1 U16805 ( .A(n11755), .B(n11754), .C(n11753), .D(
        n11752), .Y(n11756) );
  sky130_fd_sc_hd__nor2_1 U16806 ( .A(n11757), .B(n11756), .Y(n11770) );
  sky130_fd_sc_hd__nor2_1 U16807 ( .A(n12676), .B(n13919), .Y(n11763) );
  sky130_fd_sc_hd__a21oi_1 U16808 ( .A1(j202_soc_core_j22_cpu_rf_tmp[15]), 
        .A2(n11184), .B1(n13920), .Y(n11761) );
  sky130_fd_sc_hd__nand2_1 U16809 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[79]), .Y(n11760) );
  sky130_fd_sc_hd__nand2_1 U16810 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[367]), .Y(n11759) );
  sky130_fd_sc_hd__nand2_1 U16811 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[399]), .Y(n11758) );
  sky130_fd_sc_hd__nand4_1 U16812 ( .A(n11761), .B(n11760), .C(n11759), .D(
        n11758), .Y(n11762) );
  sky130_fd_sc_hd__nor2_1 U16813 ( .A(n11763), .B(n11762), .Y(n11769) );
  sky130_fd_sc_hd__nand2_1 U16814 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[175]), .Y(n11767) );
  sky130_fd_sc_hd__nand2_1 U16815 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[335]), .Y(n11766) );
  sky130_fd_sc_hd__nand2_1 U16816 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[143]), .Y(n11765) );
  sky130_fd_sc_hd__nand2_1 U16817 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[271]), .Y(n11764) );
  sky130_fd_sc_hd__and4_1 U16818 ( .A(n11767), .B(n11766), .C(n11765), .D(
        n11764), .X(n11768) );
  sky130_fd_sc_hd__nand3_1 U16819 ( .A(n11770), .B(n11769), .C(n11768), .Y(
        n22136) );
  sky130_fd_sc_hd__o22ai_1 U16820 ( .A1(n20677), .A2(n22563), .B1(n22556), 
        .B2(n14042), .Y(n12686) );
  sky130_fd_sc_hd__nand2_1 U16821 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[176]), .Y(n11774) );
  sky130_fd_sc_hd__nand2_1 U16822 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[240]), .Y(n11773) );
  sky130_fd_sc_hd__nand2_1 U16823 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[496]), .Y(n11772) );
  sky130_fd_sc_hd__nand2_1 U16824 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[432]), .Y(n11771) );
  sky130_fd_sc_hd__nand4_1 U16825 ( .A(n11774), .B(n11773), .C(n11772), .D(
        n11771), .Y(n11780) );
  sky130_fd_sc_hd__nand2_1 U16826 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[400]), .Y(n11778) );
  sky130_fd_sc_hd__nand2_1 U16827 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[16]), .Y(n11777) );
  sky130_fd_sc_hd__nand2_1 U16828 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[48]), .Y(n11776) );
  sky130_fd_sc_hd__nand2_1 U16829 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[464]), .Y(n11775) );
  sky130_fd_sc_hd__nand4_1 U16830 ( .A(n11778), .B(n11777), .C(n11776), .D(
        n11775), .Y(n11779) );
  sky130_fd_sc_hd__nor2_1 U16831 ( .A(n11780), .B(n11779), .Y(n11788) );
  sky130_fd_sc_hd__a22oi_1 U16832 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[304]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[208]), .Y(n11787) );
  sky130_fd_sc_hd__a22oi_1 U16833 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[368]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[336]), .Y(n11786) );
  sky130_fd_sc_hd__nand2_1 U16834 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[144]), .Y(n11784) );
  sky130_fd_sc_hd__nand2_1 U16835 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[80]), .Y(n11783) );
  sky130_fd_sc_hd__nand2_1 U16836 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[112]), .Y(n11782) );
  sky130_fd_sc_hd__nand2_1 U16837 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[272]), .Y(n11781) );
  sky130_fd_sc_hd__and4_1 U16838 ( .A(n11784), .B(n11783), .C(n11782), .D(
        n11781), .X(n11785) );
  sky130_fd_sc_hd__nand4_1 U16839 ( .A(n11788), .B(n11787), .C(n11786), .D(
        n11785), .Y(n19684) );
  sky130_fd_sc_hd__nand2_1 U16840 ( .A(n19684), .B(n14086), .Y(n11798) );
  sky130_fd_sc_hd__nand2_1 U16841 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[16]), .Y(n11791) );
  sky130_fd_sc_hd__nand2_1 U16842 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[16]), .Y(n11790) );
  sky130_fd_sc_hd__nand2_1 U16843 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[496]), .Y(n11789) );
  sky130_fd_sc_hd__and4_1 U16844 ( .A(n11791), .B(n11790), .C(n14022), .D(
        n11789), .X(n11797) );
  sky130_fd_sc_hd__nand2_1 U16845 ( .A(n14025), .B(
        j202_soc_core_j22_cpu_pc[16]), .Y(n11795) );
  sky130_fd_sc_hd__nand2_1 U16846 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[16]), .Y(n11794) );
  sky130_fd_sc_hd__nand2_1 U16847 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[16]), .Y(n11793) );
  sky130_fd_sc_hd__nand2_1 U16848 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[16]), .Y(n11792) );
  sky130_fd_sc_hd__and4_1 U16849 ( .A(n11795), .B(n11794), .C(n11793), .D(
        n11792), .X(n11796) );
  sky130_fd_sc_hd__nand3_1 U16850 ( .A(n11798), .B(n11797), .C(n11796), .Y(
        n23298) );
  sky130_fd_sc_hd__nand2_1 U16851 ( .A(n22375), .B(n14087), .Y(n11799) );
  sky130_fd_sc_hd__o21ai_1 U16852 ( .A1(n14089), .A2(n22375), .B1(n11799), .Y(
        n12687) );
  sky130_fd_sc_hd__nor2_1 U16853 ( .A(n12686), .B(n12687), .Y(n18481) );
  sky130_fd_sc_hd__nand2_1 U16854 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[430]), .Y(n11803) );
  sky130_fd_sc_hd__nand2_1 U16855 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[462]), .Y(n11802) );
  sky130_fd_sc_hd__nand2_1 U16856 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[110]), .Y(n11801) );
  sky130_fd_sc_hd__nand2_1 U16857 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[46]), .Y(n11800) );
  sky130_fd_sc_hd__nand4_1 U16858 ( .A(n11803), .B(n11802), .C(n11801), .D(
        n11800), .Y(n11809) );
  sky130_fd_sc_hd__nand2_1 U16859 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[174]), .Y(n11807) );
  sky130_fd_sc_hd__nand2_1 U16860 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[302]), .Y(n11806) );
  sky130_fd_sc_hd__nand2_1 U16861 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[238]), .Y(n11805) );
  sky130_fd_sc_hd__nand2_1 U16862 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[142]), .Y(n11804) );
  sky130_fd_sc_hd__nand4_1 U16863 ( .A(n11807), .B(n11806), .C(n11805), .D(
        n11804), .Y(n11808) );
  sky130_fd_sc_hd__nor2_1 U16864 ( .A(n11809), .B(n11808), .Y(n11823) );
  sky130_fd_sc_hd__nand2_1 U16865 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[206]), .Y(n11813) );
  sky130_fd_sc_hd__nand2_1 U16866 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[78]), .Y(n11812) );
  sky130_fd_sc_hd__nand2_1 U16867 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[494]), .Y(n11811) );
  sky130_fd_sc_hd__nand2_1 U16868 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[270]), .Y(n11810) );
  sky130_fd_sc_hd__and4_1 U16869 ( .A(n11813), .B(n11812), .C(n11811), .D(
        n11810), .X(n11822) );
  sky130_fd_sc_hd__nand2_1 U16870 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[366]), .Y(n11818) );
  sky130_fd_sc_hd__nand2_1 U16871 ( .A(n11184), .B(
        j202_soc_core_j22_cpu_rf_tmp[14]), .Y(n11816) );
  sky130_fd_sc_hd__nand2_1 U16872 ( .A(n11814), .B(
        j202_soc_core_j22_cpu_rf_gpr[14]), .Y(n11815) );
  sky130_fd_sc_hd__nand4_1 U16873 ( .A(n11818), .B(n11817), .C(n11816), .D(
        n11815), .Y(n11820) );
  sky130_fd_sc_hd__a22o_1 U16874 ( .A1(n13913), .A2(
        j202_soc_core_j22_cpu_rf_gpr[398]), .B1(n13902), .B2(
        j202_soc_core_j22_cpu_rf_gpr[334]), .X(n11819) );
  sky130_fd_sc_hd__nor2_1 U16875 ( .A(n11820), .B(n11819), .Y(n11821) );
  sky130_fd_sc_hd__nand3_1 U16876 ( .A(n11823), .B(n11822), .C(n11821), .Y(
        n21152) );
  sky130_fd_sc_hd__nand2_1 U16877 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[365]), .Y(n11827) );
  sky130_fd_sc_hd__nand2_1 U16878 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[173]), .Y(n11826) );
  sky130_fd_sc_hd__nand2_1 U16879 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[269]), .Y(n11825) );
  sky130_fd_sc_hd__nand2_1 U16880 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[461]), .Y(n11824) );
  sky130_fd_sc_hd__nand4_1 U16881 ( .A(n11827), .B(n11826), .C(n11825), .D(
        n11824), .Y(n11833) );
  sky130_fd_sc_hd__nand2_1 U16882 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[333]), .Y(n11831) );
  sky130_fd_sc_hd__nand2_1 U16883 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[205]), .Y(n11830) );
  sky130_fd_sc_hd__nand2_1 U16884 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[45]), .Y(n11829) );
  sky130_fd_sc_hd__nand2_1 U16885 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[77]), .Y(n11828) );
  sky130_fd_sc_hd__nand4_1 U16886 ( .A(n11831), .B(n11830), .C(n11829), .D(
        n11828), .Y(n11832) );
  sky130_fd_sc_hd__nor2_1 U16887 ( .A(n11833), .B(n11832), .Y(n11846) );
  sky130_fd_sc_hd__nand2_1 U16888 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[301]), .Y(n11837) );
  sky130_fd_sc_hd__nand2_1 U16889 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[429]), .Y(n11836) );
  sky130_fd_sc_hd__nand2_1 U16890 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[109]), .Y(n11835) );
  sky130_fd_sc_hd__nand2_1 U16891 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[141]), .Y(n11834) );
  sky130_fd_sc_hd__and4_1 U16892 ( .A(n11837), .B(n11836), .C(n11835), .D(
        n11834), .X(n11845) );
  sky130_fd_sc_hd__nor2_1 U16893 ( .A(n12642), .B(n13919), .Y(n11843) );
  sky130_fd_sc_hd__a21oi_1 U16894 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[13]), .B1(n13920), .Y(n11841) );
  sky130_fd_sc_hd__nand2_1 U16895 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[493]), .Y(n11840) );
  sky130_fd_sc_hd__nand2_1 U16896 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[237]), .Y(n11839) );
  sky130_fd_sc_hd__nand2_1 U16897 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[397]), .Y(n11838) );
  sky130_fd_sc_hd__nand4_1 U16898 ( .A(n11841), .B(n11840), .C(n11839), .D(
        n11838), .Y(n11842) );
  sky130_fd_sc_hd__nor2_1 U16899 ( .A(n11843), .B(n11842), .Y(n11844) );
  sky130_fd_sc_hd__nand3_1 U16900 ( .A(n11846), .B(n11845), .C(n11844), .Y(
        n20648) );
  sky130_fd_sc_hd__o22ai_1 U16901 ( .A1(n20677), .A2(n22562), .B1(n22561), 
        .B2(n14042), .Y(n12652) );
  sky130_fd_sc_hd__nand2_1 U16902 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[174]), .Y(n11850) );
  sky130_fd_sc_hd__nand2_1 U16903 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[238]), .Y(n11849) );
  sky130_fd_sc_hd__nand2_1 U16904 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[494]), .Y(n11848) );
  sky130_fd_sc_hd__nand2_1 U16905 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[430]), .Y(n11847) );
  sky130_fd_sc_hd__nand4_1 U16906 ( .A(n11850), .B(n11849), .C(n11848), .D(
        n11847), .Y(n11856) );
  sky130_fd_sc_hd__nand2_1 U16907 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[398]), .Y(n11854) );
  sky130_fd_sc_hd__nand2_1 U16908 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[14]), .Y(n11853) );
  sky130_fd_sc_hd__nand2_1 U16909 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[46]), .Y(n11852) );
  sky130_fd_sc_hd__nand2_1 U16910 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[462]), .Y(n11851) );
  sky130_fd_sc_hd__nand4_1 U16911 ( .A(n11854), .B(n11853), .C(n11852), .D(
        n11851), .Y(n11855) );
  sky130_fd_sc_hd__nor2_1 U16912 ( .A(n11856), .B(n11855), .Y(n11864) );
  sky130_fd_sc_hd__a22oi_1 U16913 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[302]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[206]), .Y(n11863) );
  sky130_fd_sc_hd__a22oi_1 U16914 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[366]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[334]), .Y(n11862) );
  sky130_fd_sc_hd__nand2_1 U16915 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[142]), .Y(n11860) );
  sky130_fd_sc_hd__nand2_1 U16916 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[78]), .Y(n11859) );
  sky130_fd_sc_hd__nand2_1 U16917 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[110]), .Y(n11858) );
  sky130_fd_sc_hd__nand2_1 U16918 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[270]), .Y(n11857) );
  sky130_fd_sc_hd__and4_1 U16919 ( .A(n11860), .B(n11859), .C(n11858), .D(
        n11857), .X(n11861) );
  sky130_fd_sc_hd__nand4_1 U16920 ( .A(n11864), .B(n11863), .C(n11862), .D(
        n11861), .Y(n18962) );
  sky130_fd_sc_hd__nand2_1 U16921 ( .A(n18962), .B(n14086), .Y(n11874) );
  sky130_fd_sc_hd__nand2_1 U16922 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[14]), .Y(n11867) );
  sky130_fd_sc_hd__nand2_1 U16923 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[14]), .Y(n11866) );
  sky130_fd_sc_hd__nand2_1 U16924 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[494]), .Y(n11865) );
  sky130_fd_sc_hd__and4_1 U16925 ( .A(n11867), .B(n11866), .C(n14022), .D(
        n11865), .X(n11873) );
  sky130_fd_sc_hd__nand2_1 U16926 ( .A(n14025), .B(
        j202_soc_core_j22_cpu_pc[14]), .Y(n11871) );
  sky130_fd_sc_hd__nand2_1 U16927 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[14]), .Y(n11870) );
  sky130_fd_sc_hd__nand2_1 U16928 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[14]), .Y(n11869) );
  sky130_fd_sc_hd__nand2_1 U16929 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[14]), .Y(n11868) );
  sky130_fd_sc_hd__and4_1 U16930 ( .A(n11871), .B(n11870), .C(n11869), .D(
        n11868), .X(n11872) );
  sky130_fd_sc_hd__nand3_1 U16931 ( .A(n11874), .B(n11873), .C(n11872), .Y(
        n22156) );
  sky130_fd_sc_hd__nand2_1 U16932 ( .A(n21862), .B(n14087), .Y(n11875) );
  sky130_fd_sc_hd__nor2_1 U16934 ( .A(n12652), .B(n12653), .Y(n18805) );
  sky130_fd_sc_hd__nand2_1 U16935 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[427]), .Y(n11879) );
  sky130_fd_sc_hd__nand2_1 U16936 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[267]), .Y(n11878) );
  sky130_fd_sc_hd__nand2_1 U16937 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[395]), .Y(n11877) );
  sky130_fd_sc_hd__nand2_1 U16938 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[491]), .Y(n11876) );
  sky130_fd_sc_hd__nand4_1 U16939 ( .A(n11879), .B(n11878), .C(n11877), .D(
        n11876), .Y(n11885) );
  sky130_fd_sc_hd__nand2_1 U16940 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[203]), .Y(n11883) );
  sky130_fd_sc_hd__nand2_1 U16941 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[171]), .Y(n11882) );
  sky130_fd_sc_hd__nand2_1 U16942 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[139]), .Y(n11881) );
  sky130_fd_sc_hd__nand2_1 U16943 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[43]), .Y(n11880) );
  sky130_fd_sc_hd__nand4_1 U16944 ( .A(n11883), .B(n11882), .C(n11881), .D(
        n11880), .Y(n11884) );
  sky130_fd_sc_hd__nor2_1 U16945 ( .A(n11885), .B(n11884), .Y(n11899) );
  sky130_fd_sc_hd__nand2_1 U16946 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[299]), .Y(n11889) );
  sky130_fd_sc_hd__nand2_1 U16947 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[331]), .Y(n11888) );
  sky130_fd_sc_hd__nand2_1 U16948 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[107]), .Y(n11887) );
  sky130_fd_sc_hd__nand2_1 U16949 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[459]), .Y(n11886) );
  sky130_fd_sc_hd__and4_1 U16950 ( .A(n11889), .B(n11888), .C(n11887), .D(
        n11886), .X(n11898) );
  sky130_fd_sc_hd__nor2_1 U16951 ( .A(n12406), .B(n13919), .Y(n11896) );
  sky130_fd_sc_hd__nand2_1 U16952 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[363]), .Y(n11894) );
  sky130_fd_sc_hd__nand2_1 U16953 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[235]), .Y(n11893) );
  sky130_fd_sc_hd__nand2_1 U16954 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[75]), .Y(n11891) );
  sky130_fd_sc_hd__nand4_1 U16955 ( .A(n11894), .B(n11893), .C(n11892), .D(
        n11891), .Y(n11895) );
  sky130_fd_sc_hd__nor2_1 U16956 ( .A(n11896), .B(n11895), .Y(n11897) );
  sky130_fd_sc_hd__nand3_1 U16957 ( .A(n11899), .B(n11898), .C(n11897), .Y(
        n20689) );
  sky130_fd_sc_hd__nand2_1 U16958 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[364]), .Y(n11903) );
  sky130_fd_sc_hd__nand2_1 U16959 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[76]), .Y(n11902) );
  sky130_fd_sc_hd__nand2_1 U16960 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[108]), .Y(n11901) );
  sky130_fd_sc_hd__nand2_1 U16961 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[396]), .Y(n11900) );
  sky130_fd_sc_hd__nand4_1 U16962 ( .A(n11903), .B(n11902), .C(n11901), .D(
        n11900), .Y(n11909) );
  sky130_fd_sc_hd__nand2_1 U16963 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[332]), .Y(n11907) );
  sky130_fd_sc_hd__nand2_1 U16964 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[268]), .Y(n11906) );
  sky130_fd_sc_hd__nand2_1 U16965 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[492]), .Y(n11905) );
  sky130_fd_sc_hd__nand2_1 U16966 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[140]), .Y(n11904) );
  sky130_fd_sc_hd__nand4_1 U16967 ( .A(n11907), .B(n11906), .C(n11905), .D(
        n11904), .Y(n11908) );
  sky130_fd_sc_hd__nor2_1 U16968 ( .A(n11909), .B(n11908), .Y(n11922) );
  sky130_fd_sc_hd__nor2_1 U16969 ( .A(n11944), .B(n13919), .Y(n11915) );
  sky130_fd_sc_hd__a21oi_1 U16970 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[12]), .B1(n13920), .Y(n11913) );
  sky130_fd_sc_hd__nand2_1 U16971 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[204]), .Y(n11912) );
  sky130_fd_sc_hd__nand2_1 U16972 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[44]), .Y(n11911) );
  sky130_fd_sc_hd__nand2_1 U16973 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[236]), .Y(n11910) );
  sky130_fd_sc_hd__nand4_1 U16974 ( .A(n11913), .B(n11912), .C(n11911), .D(
        n11910), .Y(n11914) );
  sky130_fd_sc_hd__nor2_1 U16975 ( .A(n11915), .B(n11914), .Y(n11921) );
  sky130_fd_sc_hd__nand2_1 U16976 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[172]), .Y(n11919) );
  sky130_fd_sc_hd__nand2_1 U16977 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[300]), .Y(n11918) );
  sky130_fd_sc_hd__nand2_1 U16978 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[428]), .Y(n11917) );
  sky130_fd_sc_hd__nand2_1 U16979 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[460]), .Y(n11916) );
  sky130_fd_sc_hd__and4_1 U16980 ( .A(n11919), .B(n11918), .C(n11917), .D(
        n11916), .X(n11920) );
  sky130_fd_sc_hd__nand3_1 U16981 ( .A(n11922), .B(n11921), .C(n11920), .Y(
        n20720) );
  sky130_fd_sc_hd__o22ai_1 U16982 ( .A1(n14042), .A2(n22564), .B1(n22560), 
        .B2(n20677), .Y(n12619) );
  sky130_fd_sc_hd__nand2_1 U16983 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[172]), .Y(n11926) );
  sky130_fd_sc_hd__nand2_1 U16984 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[236]), .Y(n11925) );
  sky130_fd_sc_hd__nand2_1 U16985 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[492]), .Y(n11924) );
  sky130_fd_sc_hd__nand2_1 U16986 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[428]), .Y(n11923) );
  sky130_fd_sc_hd__nand4_1 U16987 ( .A(n11926), .B(n11925), .C(n11924), .D(
        n11923), .Y(n11932) );
  sky130_fd_sc_hd__nand2_1 U16988 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[396]), .Y(n11930) );
  sky130_fd_sc_hd__nand2_1 U16989 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[12]), .Y(n11929) );
  sky130_fd_sc_hd__nand2_1 U16990 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[44]), .Y(n11928) );
  sky130_fd_sc_hd__nand2_1 U16991 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[460]), .Y(n11927) );
  sky130_fd_sc_hd__nand4_1 U16992 ( .A(n11930), .B(n11929), .C(n11928), .D(
        n11927), .Y(n11931) );
  sky130_fd_sc_hd__nor2_1 U16993 ( .A(n11932), .B(n11931), .Y(n11943) );
  sky130_fd_sc_hd__nand2_1 U16994 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[332]), .Y(n11936) );
  sky130_fd_sc_hd__nand2_1 U16995 ( .A(n11191), .B(
        j202_soc_core_j22_cpu_rf_gpr[204]), .Y(n11935) );
  sky130_fd_sc_hd__nand2_1 U16996 ( .A(n20285), .B(
        j202_soc_core_j22_cpu_rf_gpr[300]), .Y(n11934) );
  sky130_fd_sc_hd__nand2_1 U16997 ( .A(n20282), .B(
        j202_soc_core_j22_cpu_rf_gpr[364]), .Y(n11933) );
  sky130_fd_sc_hd__and4_1 U16998 ( .A(n11936), .B(n11935), .C(n11934), .D(
        n11933), .X(n11942) );
  sky130_fd_sc_hd__nand2_1 U16999 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[140]), .Y(n11940) );
  sky130_fd_sc_hd__nand2_1 U17000 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[76]), .Y(n11939) );
  sky130_fd_sc_hd__nand2_1 U17001 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[108]), .Y(n11938) );
  sky130_fd_sc_hd__nand2_1 U17002 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[268]), .Y(n11937) );
  sky130_fd_sc_hd__and4_1 U17003 ( .A(n11940), .B(n11939), .C(n11938), .D(
        n11937), .X(n11941) );
  sky130_fd_sc_hd__nand3_1 U17004 ( .A(n11943), .B(n11942), .C(n11941), .Y(
        n17051) );
  sky130_fd_sc_hd__a21oi_1 U17005 ( .A1(n14069), .A2(
        j202_soc_core_j22_cpu_rf_vbr[12]), .B1(n14068), .Y(n11948) );
  sky130_fd_sc_hd__a2bb2oi_1 U17006 ( .B1(j202_soc_core_j22_cpu_rf_gpr[492]), 
        .B2(n14072), .A1_N(n14071), .A2_N(n17057), .Y(n11947) );
  sky130_fd_sc_hd__o22a_1 U17007 ( .A1(n11944), .A2(n14075), .B1(n17053), .B2(
        n14073), .X(n11946) );
  sky130_fd_sc_hd__o22a_1 U17008 ( .A1(n17052), .A2(n14079), .B1(n17056), .B2(
        n14077), .X(n11945) );
  sky130_fd_sc_hd__nand4_1 U17009 ( .A(n11948), .B(n11947), .C(n11946), .D(
        n11945), .Y(n11949) );
  sky130_fd_sc_hd__nand2_1 U17010 ( .A(n22064), .B(n14087), .Y(n11950) );
  sky130_fd_sc_hd__nor2_1 U17012 ( .A(n12619), .B(n12620), .Y(n18817) );
  sky130_fd_sc_hd__nor2_1 U17013 ( .A(n12022), .B(n13919), .Y(n11957) );
  sky130_fd_sc_hd__nand2_1 U17014 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[225]), .Y(n11955) );
  sky130_fd_sc_hd__nand2_1 U17015 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[481]), .Y(n11954) );
  sky130_fd_sc_hd__a2bb2oi_1 U17016 ( .B1(j202_soc_core_j22_cpu_rf_tmp[1]), 
        .B2(n11184), .A1_N(n12539), .A2_N(n11951), .Y(n11953) );
  sky130_fd_sc_hd__nand2_1 U17017 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[385]), .Y(n11952) );
  sky130_fd_sc_hd__nand4_1 U17018 ( .A(n11955), .B(n11954), .C(n11953), .D(
        n11952), .Y(n11956) );
  sky130_fd_sc_hd__nor2_1 U17019 ( .A(n11957), .B(n11956), .Y(n11972) );
  sky130_fd_sc_hd__nand2_1 U17020 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[193]), .Y(n11961) );
  sky130_fd_sc_hd__nand2_1 U17021 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[161]), .Y(n11960) );
  sky130_fd_sc_hd__nand2_1 U17022 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[129]), .Y(n11959) );
  sky130_fd_sc_hd__nand2_1 U17023 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[321]), .Y(n11958) );
  sky130_fd_sc_hd__nand2_1 U17024 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[33]), .Y(n11965) );
  sky130_fd_sc_hd__nand2_1 U17025 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[353]), .Y(n11964) );
  sky130_fd_sc_hd__nand2_1 U17026 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[97]), .Y(n11963) );
  sky130_fd_sc_hd__nand2_1 U17027 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[65]), .Y(n11962) );
  sky130_fd_sc_hd__and4_1 U17028 ( .A(n11965), .B(n11964), .C(n11963), .D(
        n11962), .X(n11971) );
  sky130_fd_sc_hd__nand2_1 U17029 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[417]), .Y(n11969) );
  sky130_fd_sc_hd__nand2_1 U17030 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[289]), .Y(n11968) );
  sky130_fd_sc_hd__nand2_1 U17031 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[449]), .Y(n11967) );
  sky130_fd_sc_hd__nand2_1 U17032 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[257]), .Y(n11966) );
  sky130_fd_sc_hd__and4_1 U17033 ( .A(n11969), .B(n11968), .C(n11967), .D(
        n11966), .X(n11970) );
  sky130_fd_sc_hd__nand4_1 U17034 ( .A(n11972), .B(n11197), .C(n11971), .D(
        n11970), .Y(n22141) );
  sky130_fd_sc_hd__nand2_1 U17035 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[192]), .Y(n11976) );
  sky130_fd_sc_hd__nand2_1 U17036 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[64]), .Y(n11975) );
  sky130_fd_sc_hd__nand2_1 U17037 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[480]), .Y(n11974) );
  sky130_fd_sc_hd__nand2_1 U17038 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[128]), .Y(n11973) );
  sky130_fd_sc_hd__nand4_1 U17039 ( .A(n11976), .B(n11975), .C(n11974), .D(
        n11973), .Y(n11982) );
  sky130_fd_sc_hd__nand2_1 U17040 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[160]), .Y(n11980) );
  sky130_fd_sc_hd__nand2_1 U17041 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[416]), .Y(n11979) );
  sky130_fd_sc_hd__nand2_1 U17042 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[384]), .Y(n11978) );
  sky130_fd_sc_hd__nand2_1 U17043 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[256]), .Y(n11977) );
  sky130_fd_sc_hd__nand4_1 U17044 ( .A(n11980), .B(n11979), .C(n11978), .D(
        n11977), .Y(n11981) );
  sky130_fd_sc_hd__nor2_1 U17045 ( .A(n11982), .B(n11981), .Y(n11996) );
  sky130_fd_sc_hd__nand2_1 U17046 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[288]), .Y(n11986) );
  sky130_fd_sc_hd__nand2_1 U17047 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[320]), .Y(n11985) );
  sky130_fd_sc_hd__nand2_1 U17048 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[96]), .Y(n11984) );
  sky130_fd_sc_hd__nand2_1 U17049 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[448]), .Y(n11983) );
  sky130_fd_sc_hd__and4_1 U17050 ( .A(n11986), .B(n11985), .C(n11984), .D(
        n11983), .X(n11995) );
  sky130_fd_sc_hd__nor2_1 U17051 ( .A(n19278), .B(n13919), .Y(n11993) );
  sky130_fd_sc_hd__nand2_1 U17052 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[32]), .Y(n11991) );
  sky130_fd_sc_hd__nand2_1 U17053 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[224]), .Y(n11990) );
  sky130_fd_sc_hd__a2bb2oi_1 U17054 ( .B1(j202_soc_core_j22_cpu_rf_tmp[0]), 
        .B2(n11184), .A1_N(n12539), .A2_N(n11987), .Y(n11989) );
  sky130_fd_sc_hd__nand2_1 U17055 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[352]), .Y(n11988) );
  sky130_fd_sc_hd__nand4_1 U17056 ( .A(n11991), .B(n11990), .C(n11989), .D(
        n11988), .Y(n11992) );
  sky130_fd_sc_hd__nor2_1 U17057 ( .A(n11993), .B(n11992), .Y(n11994) );
  sky130_fd_sc_hd__nand3_1 U17058 ( .A(n11996), .B(n11995), .C(n11994), .Y(
        n22584) );
  sky130_fd_sc_hd__o22ai_1 U17059 ( .A1(n20677), .A2(n20805), .B1(n22146), 
        .B2(n14042), .Y(n12125) );
  sky130_fd_sc_hd__nand2_1 U17060 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[161]), .Y(n12000) );
  sky130_fd_sc_hd__nand2_1 U17061 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[225]), .Y(n11999) );
  sky130_fd_sc_hd__nand2_1 U17062 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[481]), .Y(n11998) );
  sky130_fd_sc_hd__nand2_1 U17063 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[417]), .Y(n11997) );
  sky130_fd_sc_hd__nand4_1 U17064 ( .A(n12000), .B(n11999), .C(n11998), .D(
        n11997), .Y(n12006) );
  sky130_fd_sc_hd__nand2_1 U17065 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[385]), .Y(n12004) );
  sky130_fd_sc_hd__nand2_1 U17066 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[1]), .Y(n12003) );
  sky130_fd_sc_hd__nand2_1 U17067 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[33]), .Y(n12002) );
  sky130_fd_sc_hd__nand2_1 U17068 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[449]), .Y(n12001) );
  sky130_fd_sc_hd__nand4_1 U17069 ( .A(n12004), .B(n12003), .C(n12002), .D(
        n12001), .Y(n12005) );
  sky130_fd_sc_hd__nor2_1 U17070 ( .A(n12006), .B(n12005), .Y(n12014) );
  sky130_fd_sc_hd__a22oi_1 U17071 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[289]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[193]), .Y(n12013) );
  sky130_fd_sc_hd__a22oi_1 U17072 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[353]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[321]), .Y(n12012) );
  sky130_fd_sc_hd__nand2_1 U17073 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[129]), .Y(n12010) );
  sky130_fd_sc_hd__nand2_1 U17074 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[65]), .Y(n12009) );
  sky130_fd_sc_hd__nand2_1 U17075 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[97]), .Y(n12008) );
  sky130_fd_sc_hd__nand2_1 U17076 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[257]), .Y(n12007) );
  sky130_fd_sc_hd__and4_1 U17077 ( .A(n12010), .B(n12009), .C(n12008), .D(
        n12007), .X(n12011) );
  sky130_fd_sc_hd__nand4_1 U17078 ( .A(n12014), .B(n12013), .C(n12012), .D(
        n12011), .Y(n19849) );
  sky130_fd_sc_hd__nand2_1 U17079 ( .A(n19849), .B(n14086), .Y(n12027) );
  sky130_fd_sc_hd__nand2_1 U17080 ( .A(n14025), .B(j202_soc_core_j22_cpu_pc[1]), .Y(n12018) );
  sky130_fd_sc_hd__nand2_1 U17081 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[1]), .Y(n12017) );
  sky130_fd_sc_hd__nand2_1 U17082 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[481]), .Y(n12016) );
  sky130_fd_sc_hd__nand2_1 U17083 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[1]), .Y(n12015) );
  sky130_fd_sc_hd__and4_1 U17084 ( .A(n12018), .B(n12017), .C(n12016), .D(
        n12015), .X(n12026) );
  sky130_fd_sc_hd__nand3_1 U17085 ( .A(n12020), .B(n12942), .C(n12941), .Y(
        n12943) );
  sky130_fd_sc_hd__a2bb2oi_1 U17086 ( .B1(n11551), .B2(
        j202_soc_core_j22_cpu_regop_imm__1_), .A1_N(n21653), .A2_N(n12943), 
        .Y(n12021) );
  sky130_fd_sc_hd__o22ai_1 U17088 ( .A1(n12022), .A2(n14075), .B1(n14079), 
        .B2(n19837), .Y(n12023) );
  sky130_fd_sc_hd__nor2_1 U17089 ( .A(n12024), .B(n12023), .Y(n12025) );
  sky130_fd_sc_hd__nand2_1 U17090 ( .A(n22754), .B(n14087), .Y(n12028) );
  sky130_fd_sc_hd__o21ai_1 U17091 ( .A1(n14089), .A2(n22754), .B1(n12028), .Y(
        n12126) );
  sky130_fd_sc_hd__nor2_1 U17092 ( .A(n12125), .B(n12126), .Y(n17824) );
  sky130_fd_sc_hd__nand2_1 U17093 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[290]), .Y(n12032) );
  sky130_fd_sc_hd__nand2_1 U17094 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[34]), .Y(n12031) );
  sky130_fd_sc_hd__nand2_1 U17095 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[98]), .Y(n12030) );
  sky130_fd_sc_hd__nand2_1 U17096 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[66]), .Y(n12029) );
  sky130_fd_sc_hd__nand4_1 U17097 ( .A(n12032), .B(n12031), .C(n12030), .D(
        n12029), .Y(n12038) );
  sky130_fd_sc_hd__nand2_1 U17098 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[418]), .Y(n12036) );
  sky130_fd_sc_hd__nand2_1 U17099 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[162]), .Y(n12035) );
  sky130_fd_sc_hd__nand2_1 U17100 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[450]), .Y(n12034) );
  sky130_fd_sc_hd__nand2_1 U17101 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[226]), .Y(n12033) );
  sky130_fd_sc_hd__nand4_1 U17102 ( .A(n12036), .B(n12035), .C(n12034), .D(
        n12033), .Y(n12037) );
  sky130_fd_sc_hd__nor2_1 U17103 ( .A(n12038), .B(n12037), .Y(n12054) );
  sky130_fd_sc_hd__nand2_1 U17104 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[194]), .Y(n12040) );
  sky130_fd_sc_hd__nand2_1 U17105 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[258]), .Y(n12039) );
  sky130_fd_sc_hd__o211a_2 U17106 ( .A1(n12041), .A2(n13919), .B1(n12040), 
        .C1(n12039), .X(n12053) );
  sky130_fd_sc_hd__nand3_1 U17107 ( .A(n12042), .B(n12971), .C(
        j202_soc_core_intr_req_), .Y(n12280) );
  sky130_fd_sc_hd__a21oi_1 U17108 ( .A1(n12426), .A2(
        j202_soc_core_intr_vec__0_), .B1(j202_soc_core_j22_cpu_regop_imm__2_), 
        .Y(n12045) );
  sky130_fd_sc_hd__nand2_1 U17109 ( .A(n11184), .B(
        j202_soc_core_j22_cpu_rf_tmp[2]), .Y(n12044) );
  sky130_fd_sc_hd__nand2_1 U17110 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[322]), .Y(n12043) );
  sky130_fd_sc_hd__o211ai_1 U17111 ( .A1(n12045), .A2(n12539), .B1(n12044), 
        .C1(n12043), .Y(n12051) );
  sky130_fd_sc_hd__nand2_1 U17112 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[354]), .Y(n12049) );
  sky130_fd_sc_hd__nand2_1 U17113 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[130]), .Y(n12048) );
  sky130_fd_sc_hd__nand2_1 U17114 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[386]), .Y(n12047) );
  sky130_fd_sc_hd__nand2_1 U17115 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[482]), .Y(n12046) );
  sky130_fd_sc_hd__nand4_1 U17116 ( .A(n12049), .B(n12048), .C(n12047), .D(
        n12046), .Y(n12050) );
  sky130_fd_sc_hd__nor2_1 U17117 ( .A(n12051), .B(n12050), .Y(n12052) );
  sky130_fd_sc_hd__nand3_1 U17118 ( .A(n12054), .B(n12053), .C(n12052), .Y(
        n21019) );
  sky130_fd_sc_hd__o22ai_1 U17119 ( .A1(n14042), .A2(n20805), .B1(n22487), 
        .B2(n20677), .Y(n12127) );
  sky130_fd_sc_hd__nand2_1 U17120 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[162]), .Y(n12058) );
  sky130_fd_sc_hd__nand2_1 U17121 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[226]), .Y(n12057) );
  sky130_fd_sc_hd__nand2_1 U17122 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[482]), .Y(n12056) );
  sky130_fd_sc_hd__nand2_1 U17123 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[418]), .Y(n12055) );
  sky130_fd_sc_hd__nand4_1 U17124 ( .A(n12058), .B(n12057), .C(n12056), .D(
        n12055), .Y(n12064) );
  sky130_fd_sc_hd__nand2_1 U17125 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[386]), .Y(n12062) );
  sky130_fd_sc_hd__nand2_1 U17126 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[2]), .Y(n12061) );
  sky130_fd_sc_hd__nand2_1 U17127 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[34]), .Y(n12060) );
  sky130_fd_sc_hd__nand2_1 U17128 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[450]), .Y(n12059) );
  sky130_fd_sc_hd__nand4_1 U17129 ( .A(n12062), .B(n12061), .C(n12060), .D(
        n12059), .Y(n12063) );
  sky130_fd_sc_hd__nor2_1 U17130 ( .A(n12064), .B(n12063), .Y(n12072) );
  sky130_fd_sc_hd__a22oi_1 U17131 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[290]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[194]), .Y(n12071) );
  sky130_fd_sc_hd__a22oi_1 U17132 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[354]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[322]), .Y(n12070) );
  sky130_fd_sc_hd__nand2_1 U17133 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[130]), .Y(n12068) );
  sky130_fd_sc_hd__nand2_1 U17134 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[66]), .Y(n12067) );
  sky130_fd_sc_hd__nand2_1 U17135 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[98]), .Y(n12066) );
  sky130_fd_sc_hd__nand2_1 U17136 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[258]), .Y(n12065) );
  sky130_fd_sc_hd__and4_1 U17137 ( .A(n12068), .B(n12067), .C(n12066), .D(
        n12065), .X(n12069) );
  sky130_fd_sc_hd__nand4_1 U17138 ( .A(n12072), .B(n12071), .C(n12070), .D(
        n12069), .Y(n16821) );
  sky130_fd_sc_hd__nand2_1 U17139 ( .A(n16821), .B(n14086), .Y(n12083) );
  sky130_fd_sc_hd__nand2_1 U17140 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[2]), .Y(n12076) );
  sky130_fd_sc_hd__nand2_1 U17141 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[2]), .Y(n12075) );
  sky130_fd_sc_hd__nand2_1 U17142 ( .A(n11551), .B(
        j202_soc_core_j22_cpu_regop_imm__2_), .Y(n12074) );
  sky130_fd_sc_hd__nand2_1 U17143 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[482]), .Y(n12073) );
  sky130_fd_sc_hd__and4_1 U17144 ( .A(n12076), .B(n12075), .C(n12074), .D(
        n12073), .X(n12082) );
  sky130_fd_sc_hd__nand2_1 U17145 ( .A(n14025), .B(j202_soc_core_j22_cpu_pc[2]), .Y(n12080) );
  sky130_fd_sc_hd__nand2_1 U17146 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[2]), .Y(n12079) );
  sky130_fd_sc_hd__nand2_1 U17147 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[2]), .Y(n12078) );
  sky130_fd_sc_hd__nand2_1 U17148 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[2]), .Y(n12077) );
  sky130_fd_sc_hd__and4_1 U17149 ( .A(n12080), .B(n12079), .C(n12078), .D(
        n12077), .X(n12081) );
  sky130_fd_sc_hd__nand3_1 U17150 ( .A(n12083), .B(n12082), .C(n12081), .Y(
        n22181) );
  sky130_fd_sc_hd__nand2_1 U17151 ( .A(n22264), .B(n14087), .Y(n12084) );
  sky130_fd_sc_hd__o21ai_1 U17152 ( .A1(n14089), .A2(n22264), .B1(n12084), .Y(
        n12128) );
  sky130_fd_sc_hd__nor2_1 U17153 ( .A(n17824), .B(n15073), .Y(n12130) );
  sky130_fd_sc_hd__nand2_1 U17154 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[160]), .Y(n12088) );
  sky130_fd_sc_hd__nand2_1 U17155 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[224]), .Y(n12087) );
  sky130_fd_sc_hd__nand2_1 U17156 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[480]), .Y(n12086) );
  sky130_fd_sc_hd__nand2_1 U17157 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[416]), .Y(n12085) );
  sky130_fd_sc_hd__nand4_1 U17158 ( .A(n12088), .B(n12087), .C(n12086), .D(
        n12085), .Y(n12094) );
  sky130_fd_sc_hd__nand2_1 U17159 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[384]), .Y(n12092) );
  sky130_fd_sc_hd__nand2_1 U17160 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[0]), .Y(n12091) );
  sky130_fd_sc_hd__nand2_1 U17161 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[32]), .Y(n12090) );
  sky130_fd_sc_hd__nand2_1 U17162 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[448]), .Y(n12089) );
  sky130_fd_sc_hd__nand4_1 U17163 ( .A(n12092), .B(n12091), .C(n12090), .D(
        n12089), .Y(n12093) );
  sky130_fd_sc_hd__nor2_1 U17164 ( .A(n12094), .B(n12093), .Y(n12102) );
  sky130_fd_sc_hd__a22oi_1 U17165 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[288]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[192]), .Y(n12101) );
  sky130_fd_sc_hd__a22oi_1 U17166 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[352]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[320]), .Y(n12100) );
  sky130_fd_sc_hd__nand2_1 U17167 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[128]), .Y(n12098) );
  sky130_fd_sc_hd__nand2_1 U17168 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[64]), .Y(n12097) );
  sky130_fd_sc_hd__nand2_1 U17169 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[96]), .Y(n12096) );
  sky130_fd_sc_hd__nand2_1 U17170 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[256]), .Y(n12095) );
  sky130_fd_sc_hd__and4_1 U17171 ( .A(n12098), .B(n12097), .C(n12096), .D(
        n12095), .X(n12099) );
  sky130_fd_sc_hd__nand4_1 U17172 ( .A(n12102), .B(n12101), .C(n12100), .D(
        n12099), .Y(n19272) );
  sky130_fd_sc_hd__nand2_1 U17173 ( .A(n19272), .B(n14086), .Y(n12110) );
  sky130_fd_sc_hd__o22ai_1 U17174 ( .A1(n19277), .A2(n14071), .B1(n14073), 
        .B2(n21630), .Y(n12104) );
  sky130_fd_sc_hd__a22o_1 U17175 ( .A1(n14072), .A2(
        j202_soc_core_j22_cpu_rf_gpr[480]), .B1(n14069), .B2(
        j202_soc_core_j22_cpu_rf_vbr[0]), .X(n12103) );
  sky130_fd_sc_hd__nor2_1 U17176 ( .A(n12104), .B(n12103), .Y(n12109) );
  sky130_fd_sc_hd__a2bb2oi_1 U17177 ( .B1(n11551), .B2(
        j202_soc_core_j22_cpu_regop_imm__0_), .A1_N(n11202), .A2_N(n12943), 
        .Y(n12105) );
  sky130_fd_sc_hd__o22ai_1 U17179 ( .A1(n19278), .A2(n14075), .B1(n14079), 
        .B2(n19273), .Y(n12106) );
  sky130_fd_sc_hd__nor2_1 U17180 ( .A(n12107), .B(n12106), .Y(n12108) );
  sky130_fd_sc_hd__a21oi_1 U17181 ( .A1(n12112), .A2(n12111), .B1(n21627), .Y(
        n12115) );
  sky130_fd_sc_hd__o21ai_1 U17182 ( .A1(n12114), .A2(n22754), .B1(n12113), .Y(
        n12118) );
  sky130_fd_sc_hd__a211o_1 U17183 ( .A1(n21627), .A2(n14087), .B1(n12115), 
        .C1(n12118), .X(n19247) );
  sky130_fd_sc_hd__o22ai_1 U17184 ( .A1(n11202), .A2(n14042), .B1(n20677), 
        .B2(n22146), .Y(n12122) );
  sky130_fd_sc_hd__nand2_1 U17185 ( .A(n22715), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[0]), .Y(n22695) );
  sky130_fd_sc_hd__nand2_1 U17186 ( .A(n22510), .B(
        j202_soc_core_j22_cpu_rfuo_sr__t_), .Y(n12905) );
  sky130_fd_sc_hd__o211ai_1 U17187 ( .A1(j202_soc_core_j22_cpu_exuop_EXU_[1]), 
        .A2(n16664), .B1(n12905), .C1(n12117), .Y(n12119) );
  sky130_fd_sc_hd__or4_1 U17188 ( .A(n12121), .B(n12120), .C(n12119), .D(
        n12118), .X(n12123) );
  sky130_fd_sc_hd__nor2_1 U17189 ( .A(n12122), .B(n12123), .Y(n19243) );
  sky130_fd_sc_hd__nand2_1 U17190 ( .A(n12123), .B(n12122), .Y(n19244) );
  sky130_fd_sc_hd__nand2_1 U17192 ( .A(n12126), .B(n12125), .Y(n17825) );
  sky130_fd_sc_hd__nand2_1 U17193 ( .A(n12128), .B(n12127), .Y(n15074) );
  sky130_fd_sc_hd__o21ai_1 U17194 ( .A1(n17825), .A2(n15073), .B1(n15074), .Y(
        n12129) );
  sky130_fd_sc_hd__a21oi_1 U17195 ( .A1(n12130), .A2(n15076), .B1(n12129), .Y(
        n17122) );
  sky130_fd_sc_hd__nand2_1 U17196 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[198]), .Y(n12134) );
  sky130_fd_sc_hd__nand2_1 U17197 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[70]), .Y(n12133) );
  sky130_fd_sc_hd__nand2_1 U17198 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[390]), .Y(n12132) );
  sky130_fd_sc_hd__nand2_1 U17199 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[134]), .Y(n12131) );
  sky130_fd_sc_hd__nand4_1 U17200 ( .A(n12134), .B(n12133), .C(n12132), .D(
        n12131), .Y(n12140) );
  sky130_fd_sc_hd__nand2_1 U17201 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[166]), .Y(n12138) );
  sky130_fd_sc_hd__nand2_1 U17202 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[294]), .Y(n12137) );
  sky130_fd_sc_hd__nand2_1 U17203 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[422]), .Y(n12136) );
  sky130_fd_sc_hd__nand2_1 U17204 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[454]), .Y(n12135) );
  sky130_fd_sc_hd__nand4_1 U17205 ( .A(n12138), .B(n12137), .C(n12136), .D(
        n12135), .Y(n12139) );
  sky130_fd_sc_hd__nor2_1 U17206 ( .A(n12140), .B(n12139), .Y(n12155) );
  sky130_fd_sc_hd__nand2_1 U17207 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[262]), .Y(n12142) );
  sky130_fd_sc_hd__nand2_1 U17208 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[326]), .Y(n12141) );
  sky130_fd_sc_hd__o211a_2 U17209 ( .A1(n12204), .A2(n13919), .B1(n12142), 
        .C1(n12141), .X(n12154) );
  sky130_fd_sc_hd__o22ai_1 U17210 ( .A1(n12280), .A2(n22900), .B1(n12143), 
        .B2(n12539), .Y(n12144) );
  sky130_fd_sc_hd__a21oi_1 U17211 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[6]), .B1(n12144), .Y(n12146) );
  sky130_fd_sc_hd__nand2_1 U17212 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[102]), .Y(n12145) );
  sky130_fd_sc_hd__nand2_1 U17213 ( .A(n12146), .B(n12145), .Y(n12152) );
  sky130_fd_sc_hd__nand2_1 U17214 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[38]), .Y(n12150) );
  sky130_fd_sc_hd__nand2_1 U17215 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[230]), .Y(n12149) );
  sky130_fd_sc_hd__nand2_1 U17216 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[486]), .Y(n12148) );
  sky130_fd_sc_hd__nand2_1 U17217 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[358]), .Y(n12147) );
  sky130_fd_sc_hd__nand4_1 U17218 ( .A(n12150), .B(n12149), .C(n12148), .D(
        n12147), .Y(n12151) );
  sky130_fd_sc_hd__nor2_1 U17219 ( .A(n12152), .B(n12151), .Y(n12153) );
  sky130_fd_sc_hd__nand3_1 U17220 ( .A(n12155), .B(n12154), .C(n12153), .Y(
        n20530) );
  sky130_fd_sc_hd__nand2_1 U17221 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[293]), .Y(n12159) );
  sky130_fd_sc_hd__nand2_1 U17222 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[229]), .Y(n12158) );
  sky130_fd_sc_hd__nand2_1 U17223 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[389]), .Y(n12157) );
  sky130_fd_sc_hd__nand2_1 U17224 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[261]), .Y(n12156) );
  sky130_fd_sc_hd__nand4_1 U17225 ( .A(n12159), .B(n12158), .C(n12157), .D(
        n12156), .Y(n12165) );
  sky130_fd_sc_hd__nand2_1 U17226 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[165]), .Y(n12163) );
  sky130_fd_sc_hd__nand2_1 U17227 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[197]), .Y(n12162) );
  sky130_fd_sc_hd__nand2_1 U17228 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[69]), .Y(n12161) );
  sky130_fd_sc_hd__nand2_1 U17229 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[453]), .Y(n12160) );
  sky130_fd_sc_hd__nand4_1 U17230 ( .A(n12163), .B(n12162), .C(n12161), .D(
        n12160), .Y(n12164) );
  sky130_fd_sc_hd__nor2_1 U17231 ( .A(n12165), .B(n12164), .Y(n12180) );
  sky130_fd_sc_hd__nand2_1 U17232 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[421]), .Y(n12167) );
  sky130_fd_sc_hd__nand2_1 U17233 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[325]), .Y(n12166) );
  sky130_fd_sc_hd__o211a_2 U17234 ( .A1(n12259), .A2(n13919), .B1(n12167), 
        .C1(n12166), .X(n12179) );
  sky130_fd_sc_hd__o22ai_1 U17235 ( .A1(n12280), .A2(n22905), .B1(n12168), 
        .B2(n12539), .Y(n12169) );
  sky130_fd_sc_hd__a21oi_1 U17236 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[5]), .B1(n12169), .Y(n12171) );
  sky130_fd_sc_hd__nand2_1 U17237 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[101]), .Y(n12170) );
  sky130_fd_sc_hd__nand2_1 U17238 ( .A(n12171), .B(n12170), .Y(n12177) );
  sky130_fd_sc_hd__nand2_1 U17239 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[37]), .Y(n12175) );
  sky130_fd_sc_hd__nand2_1 U17240 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[357]), .Y(n12174) );
  sky130_fd_sc_hd__nand2_1 U17241 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[485]), .Y(n12173) );
  sky130_fd_sc_hd__nand2_1 U17242 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[133]), .Y(n12172) );
  sky130_fd_sc_hd__nand4_1 U17243 ( .A(n12175), .B(n12174), .C(n12173), .D(
        n12172), .Y(n12176) );
  sky130_fd_sc_hd__nor2_1 U17244 ( .A(n12177), .B(n12176), .Y(n12178) );
  sky130_fd_sc_hd__nand3_1 U17245 ( .A(n12180), .B(n12179), .C(n12178), .Y(
        n19173) );
  sky130_fd_sc_hd__o22ai_1 U17246 ( .A1(n20677), .A2(n22612), .B1(n22580), 
        .B2(n14042), .Y(n12356) );
  sky130_fd_sc_hd__nand2_1 U17247 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[166]), .Y(n12184) );
  sky130_fd_sc_hd__nand2_1 U17248 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[230]), .Y(n12183) );
  sky130_fd_sc_hd__nand2_1 U17249 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[486]), .Y(n12182) );
  sky130_fd_sc_hd__nand2_1 U17250 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[422]), .Y(n12181) );
  sky130_fd_sc_hd__nand4_1 U17251 ( .A(n12184), .B(n12183), .C(n12182), .D(
        n12181), .Y(n12190) );
  sky130_fd_sc_hd__nand2_1 U17252 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[390]), .Y(n12188) );
  sky130_fd_sc_hd__nand2_1 U17253 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[6]), .Y(n12187) );
  sky130_fd_sc_hd__nand2_1 U17254 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[38]), .Y(n12186) );
  sky130_fd_sc_hd__nand2_1 U17255 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[454]), .Y(n12185) );
  sky130_fd_sc_hd__nand4_1 U17256 ( .A(n12188), .B(n12187), .C(n12186), .D(
        n12185), .Y(n12189) );
  sky130_fd_sc_hd__nor2_1 U17257 ( .A(n12190), .B(n12189), .Y(n12198) );
  sky130_fd_sc_hd__a22oi_1 U17258 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[294]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[198]), .Y(n12197) );
  sky130_fd_sc_hd__a22oi_1 U17259 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[358]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[326]), .Y(n12196) );
  sky130_fd_sc_hd__nand2_1 U17260 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[134]), .Y(n12194) );
  sky130_fd_sc_hd__nand2_1 U17261 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[70]), .Y(n12193) );
  sky130_fd_sc_hd__nand2_1 U17262 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[102]), .Y(n12192) );
  sky130_fd_sc_hd__nand2_1 U17263 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[262]), .Y(n12191) );
  sky130_fd_sc_hd__and4_1 U17264 ( .A(n12194), .B(n12193), .C(n12192), .D(
        n12191), .X(n12195) );
  sky130_fd_sc_hd__nand4_1 U17265 ( .A(n12198), .B(n12197), .C(n12196), .D(
        n12195), .Y(n19063) );
  sky130_fd_sc_hd__nand2_1 U17266 ( .A(n19063), .B(n14086), .Y(n12209) );
  sky130_fd_sc_hd__nand2_1 U17267 ( .A(n14025), .B(j202_soc_core_j22_cpu_pc[6]), .Y(n12202) );
  sky130_fd_sc_hd__nand2_1 U17268 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[6]), .Y(n12201) );
  sky130_fd_sc_hd__nand2_1 U17269 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[486]), .Y(n12200) );
  sky130_fd_sc_hd__nand2_1 U17270 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[6]), .Y(n12199) );
  sky130_fd_sc_hd__and4_1 U17271 ( .A(n12202), .B(n12201), .C(n12200), .D(
        n12199), .X(n12208) );
  sky130_fd_sc_hd__a2bb2oi_1 U17272 ( .B1(n11551), .B2(
        j202_soc_core_j22_cpu_regop_imm__6_), .A1_N(n19052), .A2_N(n12943), 
        .Y(n12203) );
  sky130_fd_sc_hd__o22ai_1 U17274 ( .A1(n12204), .A2(n14075), .B1(n14079), 
        .B2(n19051), .Y(n12205) );
  sky130_fd_sc_hd__nor2_1 U17275 ( .A(n12206), .B(n12205), .Y(n12207) );
  sky130_fd_sc_hd__nand3_1 U17276 ( .A(n12209), .B(n12208), .C(n12207), .Y(
        n22708) );
  sky130_fd_sc_hd__nand2_1 U17277 ( .A(n22611), .B(n14087), .Y(n12210) );
  sky130_fd_sc_hd__o21ai_1 U17278 ( .A1(n14089), .A2(n22611), .B1(n12210), .Y(
        n12357) );
  sky130_fd_sc_hd__nor2_1 U17279 ( .A(n12356), .B(n12357), .Y(n19040) );
  sky130_fd_sc_hd__nand2_1 U17280 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[196]), .Y(n12214) );
  sky130_fd_sc_hd__nand2_1 U17281 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[68]), .Y(n12213) );
  sky130_fd_sc_hd__nand2_1 U17282 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[388]), .Y(n12212) );
  sky130_fd_sc_hd__nand2_1 U17283 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[132]), .Y(n12211) );
  sky130_fd_sc_hd__nand4_1 U17284 ( .A(n12214), .B(n12213), .C(n12212), .D(
        n12211), .Y(n12220) );
  sky130_fd_sc_hd__nand2_1 U17285 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[164]), .Y(n12218) );
  sky130_fd_sc_hd__nand2_1 U17286 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[292]), .Y(n12217) );
  sky130_fd_sc_hd__nand2_1 U17287 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[420]), .Y(n12216) );
  sky130_fd_sc_hd__nand2_1 U17288 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[452]), .Y(n12215) );
  sky130_fd_sc_hd__nand4_1 U17289 ( .A(n12218), .B(n12217), .C(n12216), .D(
        n12215), .Y(n12219) );
  sky130_fd_sc_hd__nor2_1 U17290 ( .A(n12220), .B(n12219), .Y(n12235) );
  sky130_fd_sc_hd__nand2_1 U17291 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[260]), .Y(n12222) );
  sky130_fd_sc_hd__nand2_1 U17292 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[324]), .Y(n12221) );
  sky130_fd_sc_hd__o211a_2 U17293 ( .A1(n12343), .A2(n13919), .B1(n12222), 
        .C1(n12221), .X(n12234) );
  sky130_fd_sc_hd__o22ai_1 U17294 ( .A1(n12280), .A2(n22903), .B1(n12223), 
        .B2(n12539), .Y(n12224) );
  sky130_fd_sc_hd__a21oi_1 U17295 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[4]), .B1(n12224), .Y(n12226) );
  sky130_fd_sc_hd__nand2_1 U17296 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[100]), .Y(n12225) );
  sky130_fd_sc_hd__nand2_1 U17297 ( .A(n12226), .B(n12225), .Y(n12232) );
  sky130_fd_sc_hd__nand2_1 U17298 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[36]), .Y(n12230) );
  sky130_fd_sc_hd__nand2_1 U17299 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[228]), .Y(n12229) );
  sky130_fd_sc_hd__nand2_1 U17300 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[484]), .Y(n12228) );
  sky130_fd_sc_hd__nand2_1 U17301 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[356]), .Y(n12227) );
  sky130_fd_sc_hd__nand4_1 U17302 ( .A(n12230), .B(n12229), .C(n12228), .D(
        n12227), .Y(n12231) );
  sky130_fd_sc_hd__nor2_1 U17303 ( .A(n12232), .B(n12231), .Y(n12233) );
  sky130_fd_sc_hd__nand3_1 U17304 ( .A(n12235), .B(n12234), .C(n12233), .Y(
        n22483) );
  sky130_fd_sc_hd__o22ai_1 U17305 ( .A1(n20677), .A2(n22580), .B1(n22647), 
        .B2(n14042), .Y(n12354) );
  sky130_fd_sc_hd__nand2_1 U17306 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[165]), .Y(n12239) );
  sky130_fd_sc_hd__nand2_1 U17307 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[229]), .Y(n12238) );
  sky130_fd_sc_hd__nand2_1 U17308 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[485]), .Y(n12237) );
  sky130_fd_sc_hd__nand2_1 U17309 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[421]), .Y(n12236) );
  sky130_fd_sc_hd__nand4_1 U17310 ( .A(n12239), .B(n12238), .C(n12237), .D(
        n12236), .Y(n12245) );
  sky130_fd_sc_hd__nand2_1 U17311 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[389]), .Y(n12243) );
  sky130_fd_sc_hd__nand2_1 U17312 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[5]), .Y(n12242) );
  sky130_fd_sc_hd__nand2_1 U17313 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[37]), .Y(n12241) );
  sky130_fd_sc_hd__nand2_1 U17314 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[453]), .Y(n12240) );
  sky130_fd_sc_hd__nand4_1 U17315 ( .A(n12243), .B(n12242), .C(n12241), .D(
        n12240), .Y(n12244) );
  sky130_fd_sc_hd__nor2_1 U17316 ( .A(n12245), .B(n12244), .Y(n12253) );
  sky130_fd_sc_hd__a22oi_1 U17317 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[293]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[197]), .Y(n12252) );
  sky130_fd_sc_hd__a22oi_1 U17318 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[357]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[325]), .Y(n12251) );
  sky130_fd_sc_hd__nand2_1 U17319 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[133]), .Y(n12249) );
  sky130_fd_sc_hd__nand2_1 U17320 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[69]), .Y(n12248) );
  sky130_fd_sc_hd__nand2_1 U17321 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[101]), .Y(n12247) );
  sky130_fd_sc_hd__nand2_1 U17322 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[261]), .Y(n12246) );
  sky130_fd_sc_hd__and4_1 U17323 ( .A(n12249), .B(n12248), .C(n12247), .D(
        n12246), .X(n12250) );
  sky130_fd_sc_hd__nand4_1 U17324 ( .A(n12253), .B(n12252), .C(n12251), .D(
        n12250), .Y(n19191) );
  sky130_fd_sc_hd__nand2_1 U17325 ( .A(n19191), .B(n14086), .Y(n12264) );
  sky130_fd_sc_hd__nand2_1 U17326 ( .A(n14025), .B(j202_soc_core_j22_cpu_pc[5]), .Y(n12257) );
  sky130_fd_sc_hd__nand2_1 U17327 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[5]), .Y(n12256) );
  sky130_fd_sc_hd__nand2_1 U17328 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[485]), .Y(n12255) );
  sky130_fd_sc_hd__nand2_1 U17329 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[5]), .Y(n12254) );
  sky130_fd_sc_hd__and4_1 U17330 ( .A(n12257), .B(n12256), .C(n12255), .D(
        n12254), .X(n12263) );
  sky130_fd_sc_hd__a2bb2oi_1 U17331 ( .B1(n11551), .B2(
        j202_soc_core_j22_cpu_regop_imm__5_), .A1_N(n19180), .A2_N(n12943), 
        .Y(n12258) );
  sky130_fd_sc_hd__o22ai_1 U17333 ( .A1(n12259), .A2(n14075), .B1(n14079), 
        .B2(n19179), .Y(n12260) );
  sky130_fd_sc_hd__nor2_1 U17334 ( .A(n12261), .B(n12260), .Y(n12262) );
  sky130_fd_sc_hd__nand3_1 U17335 ( .A(n12264), .B(n12263), .C(n12262), .Y(
        n22176) );
  sky130_fd_sc_hd__nand2_1 U17336 ( .A(n22037), .B(n14087), .Y(n12265) );
  sky130_fd_sc_hd__nor2_1 U17338 ( .A(n12354), .B(n12355), .Y(n19072) );
  sky130_fd_sc_hd__nor2_1 U17339 ( .A(n19040), .B(n19072), .Y(n12359) );
  sky130_fd_sc_hd__nand2_1 U17340 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[163]), .Y(n12269) );
  sky130_fd_sc_hd__nand2_1 U17341 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[451]), .Y(n12268) );
  sky130_fd_sc_hd__nand2_1 U17342 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[99]), .Y(n12267) );
  sky130_fd_sc_hd__nand2_1 U17343 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[227]), .Y(n12266) );
  sky130_fd_sc_hd__nand4_1 U17344 ( .A(n12269), .B(n12268), .C(n12267), .D(
        n12266), .Y(n12275) );
  sky130_fd_sc_hd__nand2_1 U17345 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[195]), .Y(n12273) );
  sky130_fd_sc_hd__nand2_1 U17346 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[291]), .Y(n12272) );
  sky130_fd_sc_hd__nand2_1 U17347 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[355]), .Y(n12271) );
  sky130_fd_sc_hd__nand2_1 U17348 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[483]), .Y(n12270) );
  sky130_fd_sc_hd__nand4_1 U17349 ( .A(n12273), .B(n12272), .C(n12271), .D(
        n12270), .Y(n12274) );
  sky130_fd_sc_hd__nor2_1 U17350 ( .A(n12275), .B(n12274), .Y(n12292) );
  sky130_fd_sc_hd__nand2b_1 U17351 ( .A_N(n13919), .B(
        j202_soc_core_j22_cpu_rf_gpr[3]), .Y(n12278) );
  sky130_fd_sc_hd__nand2_1 U17352 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[387]), .Y(n12277) );
  sky130_fd_sc_hd__nand2_1 U17353 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[259]), .Y(n12276) );
  sky130_fd_sc_hd__and3_1 U17354 ( .A(n12278), .B(n12277), .C(n12276), .X(
        n12291) );
  sky130_fd_sc_hd__nand2_1 U17355 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[323]), .Y(n12283) );
  sky130_fd_sc_hd__o22ai_1 U17356 ( .A1(n12280), .A2(n22899), .B1(n12279), 
        .B2(n12539), .Y(n12281) );
  sky130_fd_sc_hd__a21oi_1 U17357 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[3]), .B1(n12281), .Y(n12282) );
  sky130_fd_sc_hd__nand2_1 U17358 ( .A(n12283), .B(n12282), .Y(n12289) );
  sky130_fd_sc_hd__nand2_1 U17359 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[35]), .Y(n12287) );
  sky130_fd_sc_hd__nand2_1 U17360 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[131]), .Y(n12286) );
  sky130_fd_sc_hd__nand2_1 U17361 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[67]), .Y(n12285) );
  sky130_fd_sc_hd__nand2_1 U17362 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[419]), .Y(n12284) );
  sky130_fd_sc_hd__nand4_1 U17363 ( .A(n12287), .B(n12286), .C(n12285), .D(
        n12284), .Y(n12288) );
  sky130_fd_sc_hd__nor2_1 U17364 ( .A(n12289), .B(n12288), .Y(n12290) );
  sky130_fd_sc_hd__nand3_1 U17365 ( .A(n12292), .B(n12291), .C(n12290), .Y(
        n22583) );
  sky130_fd_sc_hd__o22ai_1 U17366 ( .A1(n20677), .A2(n22488), .B1(n22487), 
        .B2(n14042), .Y(n12350) );
  sky130_fd_sc_hd__nand2_1 U17367 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[163]), .Y(n12296) );
  sky130_fd_sc_hd__nand2_1 U17368 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[227]), .Y(n12295) );
  sky130_fd_sc_hd__nand2_1 U17369 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[483]), .Y(n12294) );
  sky130_fd_sc_hd__nand2_1 U17370 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[419]), .Y(n12293) );
  sky130_fd_sc_hd__nand4_1 U17371 ( .A(n12296), .B(n12295), .C(n12294), .D(
        n12293), .Y(n12302) );
  sky130_fd_sc_hd__nand2_1 U17372 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[387]), .Y(n12300) );
  sky130_fd_sc_hd__nand2_1 U17373 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[3]), .Y(n12299) );
  sky130_fd_sc_hd__nand2_1 U17374 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[35]), .Y(n12298) );
  sky130_fd_sc_hd__nand2_1 U17375 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[451]), .Y(n12297) );
  sky130_fd_sc_hd__nand4_1 U17376 ( .A(n12300), .B(n12299), .C(n12298), .D(
        n12297), .Y(n12301) );
  sky130_fd_sc_hd__nor2_1 U17377 ( .A(n12302), .B(n12301), .Y(n12312) );
  sky130_fd_sc_hd__nand2_1 U17378 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[323]), .Y(n12306) );
  sky130_fd_sc_hd__nand2_1 U17379 ( .A(n11191), .B(
        j202_soc_core_j22_cpu_rf_gpr[195]), .Y(n12305) );
  sky130_fd_sc_hd__nand2_1 U17380 ( .A(n20285), .B(
        j202_soc_core_j22_cpu_rf_gpr[291]), .Y(n12304) );
  sky130_fd_sc_hd__nand2_1 U17381 ( .A(n20282), .B(
        j202_soc_core_j22_cpu_rf_gpr[355]), .Y(n12303) );
  sky130_fd_sc_hd__nand2_1 U17382 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[131]), .Y(n12310) );
  sky130_fd_sc_hd__nand2_1 U17383 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[67]), .Y(n12309) );
  sky130_fd_sc_hd__nand2_1 U17384 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[99]), .Y(n12308) );
  sky130_fd_sc_hd__nand2_1 U17385 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[259]), .Y(n12307) );
  sky130_fd_sc_hd__and4_1 U17386 ( .A(n12310), .B(n12309), .C(n12308), .D(
        n12307), .X(n12311) );
  sky130_fd_sc_hd__nand3_1 U17387 ( .A(n12312), .B(n11187), .C(n12311), .Y(
        n18912) );
  sky130_fd_sc_hd__a22oi_1 U17388 ( .A1(n11551), .A2(
        j202_soc_core_j22_cpu_regop_imm__3_), .B1(n14069), .B2(
        j202_soc_core_j22_cpu_rf_vbr[3]), .Y(n12317) );
  sky130_fd_sc_hd__a2bb2oi_1 U17389 ( .B1(j202_soc_core_j22_cpu_rf_gpr[483]), 
        .B2(n14072), .A1_N(n14071), .A2_N(n18917), .Y(n12316) );
  sky130_fd_sc_hd__o22a_1 U17390 ( .A1(n18914), .A2(n14079), .B1(n18918), .B2(
        n14073), .X(n12315) );
  sky130_fd_sc_hd__o22a_1 U17391 ( .A1(n12313), .A2(n14075), .B1(n18913), .B2(
        n14077), .X(n12314) );
  sky130_fd_sc_hd__nand4_1 U17392 ( .A(n12317), .B(n12316), .C(n12315), .D(
        n12314), .Y(n12318) );
  sky130_fd_sc_hd__nand2_1 U17393 ( .A(n22711), .B(n14087), .Y(n12319) );
  sky130_fd_sc_hd__o21ai_1 U17394 ( .A1(n14089), .A2(n22711), .B1(n12319), .Y(
        n12351) );
  sky130_fd_sc_hd__nor2_1 U17395 ( .A(n12350), .B(n12351), .Y(n17123) );
  sky130_fd_sc_hd__o22ai_1 U17396 ( .A1(n20677), .A2(n22647), .B1(n22488), 
        .B2(n14042), .Y(n12352) );
  sky130_fd_sc_hd__nand2_1 U17397 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[164]), .Y(n12323) );
  sky130_fd_sc_hd__nand2_1 U17398 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[228]), .Y(n12322) );
  sky130_fd_sc_hd__nand2_1 U17399 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[484]), .Y(n12321) );
  sky130_fd_sc_hd__nand2_1 U17400 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[420]), .Y(n12320) );
  sky130_fd_sc_hd__nand4_1 U17401 ( .A(n12323), .B(n12322), .C(n12321), .D(
        n12320), .Y(n12329) );
  sky130_fd_sc_hd__nand2_1 U17402 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[388]), .Y(n12327) );
  sky130_fd_sc_hd__nand2_1 U17403 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[4]), .Y(n12326) );
  sky130_fd_sc_hd__nand2_1 U17404 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[36]), .Y(n12325) );
  sky130_fd_sc_hd__nand2_1 U17405 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[452]), .Y(n12324) );
  sky130_fd_sc_hd__nand4_1 U17406 ( .A(n12327), .B(n12326), .C(n12325), .D(
        n12324), .Y(n12328) );
  sky130_fd_sc_hd__nor2_1 U17407 ( .A(n12329), .B(n12328), .Y(n12337) );
  sky130_fd_sc_hd__a22oi_1 U17408 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[292]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[196]), .Y(n12336) );
  sky130_fd_sc_hd__a22oi_1 U17409 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[356]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[324]), .Y(n12335) );
  sky130_fd_sc_hd__nand2_1 U17410 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[132]), .Y(n12333) );
  sky130_fd_sc_hd__nand2_1 U17411 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[68]), .Y(n12332) );
  sky130_fd_sc_hd__nand2_1 U17412 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[100]), .Y(n12331) );
  sky130_fd_sc_hd__nand2_1 U17413 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[260]), .Y(n12330) );
  sky130_fd_sc_hd__and4_1 U17414 ( .A(n12333), .B(n12332), .C(n12331), .D(
        n12330), .X(n12334) );
  sky130_fd_sc_hd__nand4_1 U17415 ( .A(n12337), .B(n12336), .C(n12335), .D(
        n12334), .Y(n17075) );
  sky130_fd_sc_hd__nand2_1 U17416 ( .A(n17075), .B(n14086), .Y(n12348) );
  sky130_fd_sc_hd__nand2_1 U17417 ( .A(n14025), .B(j202_soc_core_j22_cpu_pc[4]), .Y(n12341) );
  sky130_fd_sc_hd__nand2_1 U17418 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[4]), .Y(n12340) );
  sky130_fd_sc_hd__nand2_1 U17419 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[484]), .Y(n12339) );
  sky130_fd_sc_hd__nand2_1 U17420 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[4]), .Y(n12338) );
  sky130_fd_sc_hd__and4_1 U17421 ( .A(n12341), .B(n12340), .C(n12339), .D(
        n12338), .X(n12347) );
  sky130_fd_sc_hd__a2bb2oi_1 U17422 ( .B1(n11551), .B2(
        j202_soc_core_j22_cpu_regop_imm__4_), .A1_N(n17064), .A2_N(n12943), 
        .Y(n12342) );
  sky130_fd_sc_hd__o22ai_1 U17424 ( .A1(n12343), .A2(n14075), .B1(n14079), 
        .B2(n17063), .Y(n12344) );
  sky130_fd_sc_hd__nor2_1 U17425 ( .A(n12345), .B(n12344), .Y(n12346) );
  sky130_fd_sc_hd__nand3_1 U17426 ( .A(n12348), .B(n12347), .C(n12346), .Y(
        n22705) );
  sky130_fd_sc_hd__nand2_1 U17427 ( .A(n22646), .B(n14087), .Y(n12349) );
  sky130_fd_sc_hd__nor2_1 U17429 ( .A(n12352), .B(n12353), .Y(n17125) );
  sky130_fd_sc_hd__nor2_1 U17430 ( .A(n17123), .B(n17125), .Y(n19044) );
  sky130_fd_sc_hd__nand2_1 U17431 ( .A(n12359), .B(n19044), .Y(n12361) );
  sky130_fd_sc_hd__nand2_1 U17432 ( .A(n12351), .B(n12350), .Y(n17833) );
  sky130_fd_sc_hd__nand2_1 U17433 ( .A(n12353), .B(n12352), .Y(n17126) );
  sky130_fd_sc_hd__nand2_1 U17435 ( .A(n12355), .B(n12354), .Y(n19073) );
  sky130_fd_sc_hd__nand2_1 U17436 ( .A(n12357), .B(n12356), .Y(n19041) );
  sky130_fd_sc_hd__a21oi_1 U17438 ( .A1(n12359), .A2(n19043), .B1(n12358), .Y(
        n12360) );
  sky130_fd_sc_hd__o21ai_1 U17439 ( .A1(n17122), .A2(n12361), .B1(n12360), .Y(
        n16679) );
  sky130_fd_sc_hd__nor2_1 U17440 ( .A(n12570), .B(n13919), .Y(n12368) );
  sky130_fd_sc_hd__nand2_1 U17441 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[42]), .Y(n12366) );
  sky130_fd_sc_hd__nand2_1 U17442 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[74]), .Y(n12365) );
  sky130_fd_sc_hd__a2bb2oi_1 U17443 ( .B1(j202_soc_core_j22_cpu_rf_tmp[10]), 
        .B2(n11184), .A1_N(n12539), .A2_N(n12362), .Y(n12364) );
  sky130_fd_sc_hd__nand2_1 U17444 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[490]), .Y(n12363) );
  sky130_fd_sc_hd__nand4_1 U17445 ( .A(n12366), .B(n12365), .C(n12364), .D(
        n12363), .Y(n12367) );
  sky130_fd_sc_hd__nor2_1 U17446 ( .A(n12368), .B(n12367), .Y(n12384) );
  sky130_fd_sc_hd__nand2_1 U17447 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[362]), .Y(n12372) );
  sky130_fd_sc_hd__nand2_1 U17448 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[266]), .Y(n12371) );
  sky130_fd_sc_hd__nand2_1 U17449 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[138]), .Y(n12370) );
  sky130_fd_sc_hd__nand2_1 U17450 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[458]), .Y(n12369) );
  sky130_fd_sc_hd__and4_1 U17451 ( .A(n12372), .B(n12371), .C(n12370), .D(
        n12369), .X(n12383) );
  sky130_fd_sc_hd__nand2_1 U17452 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[202]), .Y(n12376) );
  sky130_fd_sc_hd__nand2_1 U17453 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[170]), .Y(n12375) );
  sky130_fd_sc_hd__nand2_1 U17454 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[106]), .Y(n12374) );
  sky130_fd_sc_hd__nand2_1 U17455 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[234]), .Y(n12373) );
  sky130_fd_sc_hd__and4_1 U17456 ( .A(n12376), .B(n12375), .C(n12374), .D(
        n12373), .X(n12382) );
  sky130_fd_sc_hd__nand2_1 U17457 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[330]), .Y(n12380) );
  sky130_fd_sc_hd__nand2_1 U17458 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[298]), .Y(n12379) );
  sky130_fd_sc_hd__nand2_1 U17459 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[394]), .Y(n12378) );
  sky130_fd_sc_hd__nand2_1 U17460 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[426]), .Y(n12377) );
  sky130_fd_sc_hd__and4_1 U17461 ( .A(n12380), .B(n12379), .C(n12378), .D(
        n12377), .X(n12381) );
  sky130_fd_sc_hd__nand4_1 U17462 ( .A(n12384), .B(n12383), .C(n12382), .D(
        n12381), .Y(n20935) );
  sky130_fd_sc_hd__o22ai_1 U17463 ( .A1(n20677), .A2(n22564), .B1(n22557), 
        .B2(n14042), .Y(n12615) );
  sky130_fd_sc_hd__nand2_1 U17464 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[171]), .Y(n12388) );
  sky130_fd_sc_hd__nand2_1 U17465 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[235]), .Y(n12387) );
  sky130_fd_sc_hd__nand2_1 U17466 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[491]), .Y(n12386) );
  sky130_fd_sc_hd__nand2_1 U17467 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[427]), .Y(n12385) );
  sky130_fd_sc_hd__nand4_1 U17468 ( .A(n12388), .B(n12387), .C(n12386), .D(
        n12385), .Y(n12394) );
  sky130_fd_sc_hd__nand2_1 U17469 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[395]), .Y(n12392) );
  sky130_fd_sc_hd__nand2_1 U17470 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[11]), .Y(n12391) );
  sky130_fd_sc_hd__nand2_1 U17471 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[43]), .Y(n12390) );
  sky130_fd_sc_hd__nand2_1 U17472 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[459]), .Y(n12389) );
  sky130_fd_sc_hd__nand4_1 U17473 ( .A(n12392), .B(n12391), .C(n12390), .D(
        n12389), .Y(n12393) );
  sky130_fd_sc_hd__nor2_1 U17474 ( .A(n12394), .B(n12393), .Y(n12405) );
  sky130_fd_sc_hd__nand2_1 U17475 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[331]), .Y(n12398) );
  sky130_fd_sc_hd__nand2_1 U17476 ( .A(n11191), .B(
        j202_soc_core_j22_cpu_rf_gpr[203]), .Y(n12397) );
  sky130_fd_sc_hd__nand2_1 U17477 ( .A(n20285), .B(
        j202_soc_core_j22_cpu_rf_gpr[299]), .Y(n12396) );
  sky130_fd_sc_hd__nand2_1 U17478 ( .A(n20282), .B(
        j202_soc_core_j22_cpu_rf_gpr[363]), .Y(n12395) );
  sky130_fd_sc_hd__and4_1 U17479 ( .A(n12398), .B(n12397), .C(n12396), .D(
        n12395), .X(n12404) );
  sky130_fd_sc_hd__nand2_1 U17480 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[139]), .Y(n12402) );
  sky130_fd_sc_hd__nand2_1 U17481 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[75]), .Y(n12401) );
  sky130_fd_sc_hd__nand2_1 U17482 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[107]), .Y(n12400) );
  sky130_fd_sc_hd__nand2_1 U17483 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[267]), .Y(n12399) );
  sky130_fd_sc_hd__and4_1 U17484 ( .A(n12402), .B(n12401), .C(n12400), .D(
        n12399), .X(n12403) );
  sky130_fd_sc_hd__nand3_1 U17485 ( .A(n12405), .B(n12404), .C(n12403), .Y(
        n18925) );
  sky130_fd_sc_hd__a22oi_1 U17486 ( .A1(n11551), .A2(
        j202_soc_core_j22_cpu_regop_imm__11_), .B1(n14069), .B2(
        j202_soc_core_j22_cpu_rf_vbr[11]), .Y(n12410) );
  sky130_fd_sc_hd__a2bb2oi_1 U17487 ( .B1(j202_soc_core_j22_cpu_rf_gpr[491]), 
        .B2(n14072), .A1_N(n14071), .A2_N(n18931), .Y(n12409) );
  sky130_fd_sc_hd__o22a_1 U17488 ( .A1(n12406), .A2(n14075), .B1(n18927), .B2(
        n14073), .X(n12408) );
  sky130_fd_sc_hd__o22a_1 U17489 ( .A1(n18926), .A2(n14079), .B1(n18930), .B2(
        n14077), .X(n12407) );
  sky130_fd_sc_hd__nand4_1 U17490 ( .A(n12410), .B(n12409), .C(n12408), .D(
        n12407), .Y(n12411) );
  sky130_fd_sc_hd__a21oi_1 U17491 ( .A1(n18925), .A2(n14086), .B1(n12411), .Y(
        n22351) );
  sky130_fd_sc_hd__nand2_1 U17492 ( .A(n22351), .B(n14087), .Y(n12412) );
  sky130_fd_sc_hd__nor2_1 U17494 ( .A(n12615), .B(n12616), .Y(n18837) );
  sky130_fd_sc_hd__nand2_1 U17495 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[264]), .Y(n12416) );
  sky130_fd_sc_hd__nand2_1 U17496 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[232]), .Y(n12415) );
  sky130_fd_sc_hd__nand2_1 U17497 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[392]), .Y(n12414) );
  sky130_fd_sc_hd__nand2_1 U17498 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[456]), .Y(n12413) );
  sky130_fd_sc_hd__nand4_1 U17499 ( .A(n12416), .B(n12415), .C(n12414), .D(
        n12413), .Y(n12422) );
  sky130_fd_sc_hd__nand2_1 U17500 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[296]), .Y(n12420) );
  sky130_fd_sc_hd__nand2_1 U17501 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[40]), .Y(n12419) );
  sky130_fd_sc_hd__nand2_1 U17502 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[488]), .Y(n12418) );
  sky130_fd_sc_hd__nand2_1 U17503 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[136]), .Y(n12417) );
  sky130_fd_sc_hd__nand4_1 U17504 ( .A(n12420), .B(n12419), .C(n12418), .D(
        n12417), .Y(n12421) );
  sky130_fd_sc_hd__nor2_1 U17505 ( .A(n12422), .B(n12421), .Y(n12439) );
  sky130_fd_sc_hd__nand2_1 U17506 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[168]), .Y(n12424) );
  sky130_fd_sc_hd__nand2_1 U17507 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[328]), .Y(n12423) );
  sky130_fd_sc_hd__o211a_2 U17508 ( .A1(n12487), .A2(n13919), .B1(n12424), 
        .C1(n12423), .X(n12438) );
  sky130_fd_sc_hd__nand2_1 U17509 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[104]), .Y(n12430) );
  sky130_fd_sc_hd__nand2_1 U17510 ( .A(n11184), .B(
        j202_soc_core_j22_cpu_rf_tmp[8]), .Y(n12429) );
  sky130_fd_sc_hd__nand2_1 U17511 ( .A(n12425), .B(
        j202_soc_core_j22_cpu_regop_imm__8_), .Y(n12428) );
  sky130_fd_sc_hd__nand2_1 U17512 ( .A(n12426), .B(j202_soc_core_intr_vec__6_), 
        .Y(n12427) );
  sky130_fd_sc_hd__nand4_1 U17513 ( .A(n12430), .B(n12429), .C(n12428), .D(
        n12427), .Y(n12436) );
  sky130_fd_sc_hd__nand2_1 U17514 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[360]), .Y(n12434) );
  sky130_fd_sc_hd__nand2_1 U17515 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[200]), .Y(n12433) );
  sky130_fd_sc_hd__nand2_1 U17516 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[72]), .Y(n12432) );
  sky130_fd_sc_hd__nand2_1 U17517 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[424]), .Y(n12431) );
  sky130_fd_sc_hd__nand4_1 U17518 ( .A(n12434), .B(n12433), .C(n12432), .D(
        n12431), .Y(n12435) );
  sky130_fd_sc_hd__nor2_1 U17519 ( .A(n12436), .B(n12435), .Y(n12437) );
  sky130_fd_sc_hd__nand3_1 U17520 ( .A(n12439), .B(n12438), .C(n12437), .Y(
        n20721) );
  sky130_fd_sc_hd__nand2_1 U17521 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[199]), .Y(n12443) );
  sky130_fd_sc_hd__nand2_1 U17522 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[71]), .Y(n12442) );
  sky130_fd_sc_hd__nand2_1 U17523 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[487]), .Y(n12441) );
  sky130_fd_sc_hd__nand2_1 U17524 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[135]), .Y(n12440) );
  sky130_fd_sc_hd__nand4_1 U17525 ( .A(n12443), .B(n12442), .C(n12441), .D(
        n12440), .Y(n12449) );
  sky130_fd_sc_hd__nand2_1 U17526 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[167]), .Y(n12447) );
  sky130_fd_sc_hd__nand2_1 U17527 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[423]), .Y(n12446) );
  sky130_fd_sc_hd__nand2_1 U17528 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[391]), .Y(n12445) );
  sky130_fd_sc_hd__nand2_1 U17529 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[263]), .Y(n12444) );
  sky130_fd_sc_hd__nand4_1 U17530 ( .A(n12447), .B(n12446), .C(n12445), .D(
        n12444), .Y(n12448) );
  sky130_fd_sc_hd__nor2_1 U17531 ( .A(n12449), .B(n12448), .Y(n12463) );
  sky130_fd_sc_hd__nand2_1 U17532 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[295]), .Y(n12453) );
  sky130_fd_sc_hd__nand2_1 U17533 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[327]), .Y(n12452) );
  sky130_fd_sc_hd__nand2_1 U17534 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[103]), .Y(n12451) );
  sky130_fd_sc_hd__nand2_1 U17535 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[455]), .Y(n12450) );
  sky130_fd_sc_hd__and4_1 U17536 ( .A(n12453), .B(n12452), .C(n12451), .D(
        n12450), .X(n12462) );
  sky130_fd_sc_hd__nor2_1 U17537 ( .A(n12517), .B(n13919), .Y(n12460) );
  sky130_fd_sc_hd__nand2_1 U17538 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[39]), .Y(n12458) );
  sky130_fd_sc_hd__nand2_1 U17539 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[231]), .Y(n12457) );
  sky130_fd_sc_hd__a2bb2oi_1 U17540 ( .B1(j202_soc_core_j22_cpu_rf_tmp[7]), 
        .B2(n11184), .A1_N(n12539), .A2_N(n12454), .Y(n12456) );
  sky130_fd_sc_hd__nand2_1 U17541 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[359]), .Y(n12455) );
  sky130_fd_sc_hd__nand4_1 U17542 ( .A(n12458), .B(n12457), .C(n12456), .D(
        n12455), .Y(n12459) );
  sky130_fd_sc_hd__nor2_1 U17543 ( .A(n12460), .B(n12459), .Y(n12461) );
  sky130_fd_sc_hd__nand3_1 U17544 ( .A(n12463), .B(n12462), .C(n12461), .Y(
        n22496) );
  sky130_fd_sc_hd__o22ai_1 U17545 ( .A1(n20677), .A2(n22558), .B1(n22645), 
        .B2(n14042), .Y(n12607) );
  sky130_fd_sc_hd__nand2_1 U17546 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[168]), .Y(n12467) );
  sky130_fd_sc_hd__nand2_1 U17547 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[232]), .Y(n12466) );
  sky130_fd_sc_hd__nand2_1 U17548 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[488]), .Y(n12465) );
  sky130_fd_sc_hd__nand2_1 U17549 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[424]), .Y(n12464) );
  sky130_fd_sc_hd__nand4_1 U17550 ( .A(n12467), .B(n12466), .C(n12465), .D(
        n12464), .Y(n12473) );
  sky130_fd_sc_hd__nand2_1 U17551 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[392]), .Y(n12471) );
  sky130_fd_sc_hd__nand2_1 U17552 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[8]), .Y(n12470) );
  sky130_fd_sc_hd__nand2_1 U17553 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[40]), .Y(n12469) );
  sky130_fd_sc_hd__nand2_1 U17554 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[456]), .Y(n12468) );
  sky130_fd_sc_hd__nand4_1 U17555 ( .A(n12471), .B(n12470), .C(n12469), .D(
        n12468), .Y(n12472) );
  sky130_fd_sc_hd__nor2_1 U17556 ( .A(n12473), .B(n12472), .Y(n12481) );
  sky130_fd_sc_hd__a22oi_1 U17557 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[296]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[200]), .Y(n12480) );
  sky130_fd_sc_hd__a22oi_1 U17558 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[360]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[328]), .Y(n12479) );
  sky130_fd_sc_hd__nand2_1 U17559 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[136]), .Y(n12477) );
  sky130_fd_sc_hd__nand2_1 U17560 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[72]), .Y(n12476) );
  sky130_fd_sc_hd__nand2_1 U17561 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[104]), .Y(n12475) );
  sky130_fd_sc_hd__nand2_1 U17562 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[264]), .Y(n12474) );
  sky130_fd_sc_hd__and4_1 U17563 ( .A(n12477), .B(n12476), .C(n12475), .D(
        n12474), .X(n12478) );
  sky130_fd_sc_hd__nand4_1 U17564 ( .A(n12481), .B(n12480), .C(n12479), .D(
        n12478), .Y(n19212) );
  sky130_fd_sc_hd__nand2_1 U17565 ( .A(n19212), .B(n14086), .Y(n12492) );
  sky130_fd_sc_hd__nand2_1 U17566 ( .A(n14025), .B(j202_soc_core_j22_cpu_pc[8]), .Y(n12485) );
  sky130_fd_sc_hd__nand2_1 U17567 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[8]), .Y(n12484) );
  sky130_fd_sc_hd__nand2_1 U17568 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[488]), .Y(n12483) );
  sky130_fd_sc_hd__nand2_1 U17569 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[8]), .Y(n12482) );
  sky130_fd_sc_hd__and4_1 U17570 ( .A(n12485), .B(n12484), .C(n12483), .D(
        n12482), .X(n12491) );
  sky130_fd_sc_hd__a2bb2oi_1 U17571 ( .B1(n11551), .B2(
        j202_soc_core_j22_cpu_regop_imm__8_), .A1_N(n19201), .A2_N(n12943), 
        .Y(n12486) );
  sky130_fd_sc_hd__o22ai_1 U17573 ( .A1(n12487), .A2(n14075), .B1(n14079), 
        .B2(n19200), .Y(n12488) );
  sky130_fd_sc_hd__nor2_1 U17574 ( .A(n12489), .B(n12488), .Y(n12490) );
  sky130_fd_sc_hd__nand3_1 U17575 ( .A(n12492), .B(n12491), .C(n12490), .Y(
        n22171) );
  sky130_fd_sc_hd__nand2_1 U17576 ( .A(n21929), .B(n14087), .Y(n12493) );
  sky130_fd_sc_hd__nor2_1 U17578 ( .A(n12607), .B(n12608), .Y(n19721) );
  sky130_fd_sc_hd__o22ai_1 U17579 ( .A1(n20677), .A2(n22645), .B1(n22612), 
        .B2(n14042), .Y(n12605) );
  sky130_fd_sc_hd__nand2_1 U17580 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[167]), .Y(n12497) );
  sky130_fd_sc_hd__nand2_1 U17581 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[231]), .Y(n12496) );
  sky130_fd_sc_hd__nand2_1 U17582 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[487]), .Y(n12495) );
  sky130_fd_sc_hd__nand2_1 U17583 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[423]), .Y(n12494) );
  sky130_fd_sc_hd__nand4_1 U17584 ( .A(n12497), .B(n12496), .C(n12495), .D(
        n12494), .Y(n12503) );
  sky130_fd_sc_hd__nand2_1 U17585 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[391]), .Y(n12501) );
  sky130_fd_sc_hd__nand2_1 U17586 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[7]), .Y(n12500) );
  sky130_fd_sc_hd__nand2_1 U17587 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[39]), .Y(n12499) );
  sky130_fd_sc_hd__nand2_1 U17588 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[455]), .Y(n12498) );
  sky130_fd_sc_hd__nand4_1 U17589 ( .A(n12501), .B(n12500), .C(n12499), .D(
        n12498), .Y(n12502) );
  sky130_fd_sc_hd__nor2_1 U17590 ( .A(n12503), .B(n12502), .Y(n12511) );
  sky130_fd_sc_hd__a22oi_1 U17591 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[295]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[199]), .Y(n12510) );
  sky130_fd_sc_hd__a22oi_1 U17592 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[359]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[327]), .Y(n12509) );
  sky130_fd_sc_hd__nand2_1 U17593 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[135]), .Y(n12507) );
  sky130_fd_sc_hd__nand2_1 U17594 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[71]), .Y(n12506) );
  sky130_fd_sc_hd__nand2_1 U17595 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[103]), .Y(n12505) );
  sky130_fd_sc_hd__nand2_1 U17596 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[263]), .Y(n12504) );
  sky130_fd_sc_hd__and4_1 U17597 ( .A(n12507), .B(n12506), .C(n12505), .D(
        n12504), .X(n12508) );
  sky130_fd_sc_hd__nand4_1 U17598 ( .A(n12511), .B(n12510), .C(n12509), .D(
        n12508), .Y(n16703) );
  sky130_fd_sc_hd__nand2_1 U17599 ( .A(n16703), .B(n14086), .Y(n12522) );
  sky130_fd_sc_hd__nand2_1 U17600 ( .A(n14025), .B(j202_soc_core_j22_cpu_pc[7]), .Y(n12515) );
  sky130_fd_sc_hd__nand2_1 U17601 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[7]), .Y(n12514) );
  sky130_fd_sc_hd__nand2_1 U17602 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[487]), .Y(n12513) );
  sky130_fd_sc_hd__nand2_1 U17603 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[7]), .Y(n12512) );
  sky130_fd_sc_hd__and4_1 U17604 ( .A(n12515), .B(n12514), .C(n12513), .D(
        n12512), .X(n12521) );
  sky130_fd_sc_hd__a2bb2oi_1 U17605 ( .B1(n11551), .B2(
        j202_soc_core_j22_cpu_regop_imm__7_), .A1_N(n16692), .A2_N(n12943), 
        .Y(n12516) );
  sky130_fd_sc_hd__o22ai_1 U17607 ( .A1(n12517), .A2(n14075), .B1(n14079), 
        .B2(n16691), .Y(n12518) );
  sky130_fd_sc_hd__nor2_1 U17608 ( .A(n12519), .B(n12518), .Y(n12520) );
  sky130_fd_sc_hd__nand3_1 U17609 ( .A(n12522), .B(n12521), .C(n12520), .Y(
        n22704) );
  sky130_fd_sc_hd__nand2_1 U17610 ( .A(n22644), .B(n14087), .Y(n12523) );
  sky130_fd_sc_hd__nor2_1 U17612 ( .A(n12605), .B(n12606), .Y(n19726) );
  sky130_fd_sc_hd__nor2_1 U17613 ( .A(n19721), .B(n19726), .Y(n18940) );
  sky130_fd_sc_hd__nand2_1 U17614 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[233]), .Y(n12527) );
  sky130_fd_sc_hd__nand2_1 U17615 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[361]), .Y(n12526) );
  sky130_fd_sc_hd__nand2_1 U17616 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[105]), .Y(n12525) );
  sky130_fd_sc_hd__nand2_1 U17617 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[137]), .Y(n12524) );
  sky130_fd_sc_hd__nand4_1 U17618 ( .A(n12527), .B(n12526), .C(n12525), .D(
        n12524), .Y(n12533) );
  sky130_fd_sc_hd__nand2_1 U17619 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[73]), .Y(n12531) );
  sky130_fd_sc_hd__nand2_1 U17620 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[297]), .Y(n12530) );
  sky130_fd_sc_hd__nand2_1 U17621 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[425]), .Y(n12529) );
  sky130_fd_sc_hd__nand2_1 U17622 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[265]), .Y(n12528) );
  sky130_fd_sc_hd__nand4_1 U17623 ( .A(n12531), .B(n12530), .C(n12529), .D(
        n12528), .Y(n12532) );
  sky130_fd_sc_hd__nor2_1 U17624 ( .A(n12533), .B(n12532), .Y(n12548) );
  sky130_fd_sc_hd__nand2_1 U17625 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[169]), .Y(n12537) );
  sky130_fd_sc_hd__nand2_1 U17626 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[329]), .Y(n12536) );
  sky130_fd_sc_hd__nand2_1 U17627 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[393]), .Y(n12535) );
  sky130_fd_sc_hd__nand2_1 U17628 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[457]), .Y(n12534) );
  sky130_fd_sc_hd__and4_1 U17629 ( .A(n12537), .B(n12536), .C(n12535), .D(
        n12534), .X(n12547) );
  sky130_fd_sc_hd__nor2_1 U17630 ( .A(n19984), .B(n13919), .Y(n12545) );
  sky130_fd_sc_hd__nand2_1 U17631 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[201]), .Y(n12543) );
  sky130_fd_sc_hd__nand2_1 U17632 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[41]), .Y(n12542) );
  sky130_fd_sc_hd__nand2_1 U17634 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[489]), .Y(n12540) );
  sky130_fd_sc_hd__nand4_1 U17635 ( .A(n12543), .B(n12542), .C(n12541), .D(
        n12540), .Y(n12544) );
  sky130_fd_sc_hd__nor2_1 U17636 ( .A(n12545), .B(n12544), .Y(n12546) );
  sky130_fd_sc_hd__nand3_1 U17637 ( .A(n12548), .B(n12547), .C(n12546), .Y(
        n20699) );
  sky130_fd_sc_hd__o22ai_1 U17638 ( .A1(n20677), .A2(n22557), .B1(n22559), 
        .B2(n14042), .Y(n12611) );
  sky130_fd_sc_hd__nand2_1 U17639 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[170]), .Y(n12552) );
  sky130_fd_sc_hd__nand2_1 U17640 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[234]), .Y(n12551) );
  sky130_fd_sc_hd__nand2_1 U17641 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[490]), .Y(n12550) );
  sky130_fd_sc_hd__nand2_1 U17642 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[426]), .Y(n12549) );
  sky130_fd_sc_hd__nand4_1 U17643 ( .A(n12552), .B(n12551), .C(n12550), .D(
        n12549), .Y(n12558) );
  sky130_fd_sc_hd__nand2_1 U17644 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[394]), .Y(n12556) );
  sky130_fd_sc_hd__nand2_1 U17645 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[10]), .Y(n12555) );
  sky130_fd_sc_hd__nand2_1 U17646 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[42]), .Y(n12554) );
  sky130_fd_sc_hd__nand2_1 U17647 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[458]), .Y(n12553) );
  sky130_fd_sc_hd__nand4_1 U17648 ( .A(n12556), .B(n12555), .C(n12554), .D(
        n12553), .Y(n12557) );
  sky130_fd_sc_hd__nor2_1 U17649 ( .A(n12558), .B(n12557), .Y(n12569) );
  sky130_fd_sc_hd__nand2_1 U17650 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[330]), .Y(n12562) );
  sky130_fd_sc_hd__nand2_1 U17651 ( .A(n11191), .B(
        j202_soc_core_j22_cpu_rf_gpr[202]), .Y(n12561) );
  sky130_fd_sc_hd__nand2_1 U17652 ( .A(n20285), .B(
        j202_soc_core_j22_cpu_rf_gpr[298]), .Y(n12560) );
  sky130_fd_sc_hd__nand2_1 U17653 ( .A(n20282), .B(
        j202_soc_core_j22_cpu_rf_gpr[362]), .Y(n12559) );
  sky130_fd_sc_hd__and4_1 U17654 ( .A(n12562), .B(n12561), .C(n12560), .D(
        n12559), .X(n12568) );
  sky130_fd_sc_hd__nand2_1 U17655 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[138]), .Y(n12566) );
  sky130_fd_sc_hd__nand2_1 U17656 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[74]), .Y(n12565) );
  sky130_fd_sc_hd__nand2_1 U17657 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[106]), .Y(n12564) );
  sky130_fd_sc_hd__nand2_1 U17658 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[266]), .Y(n12563) );
  sky130_fd_sc_hd__and4_1 U17659 ( .A(n12566), .B(n12565), .C(n12564), .D(
        n12563), .X(n12567) );
  sky130_fd_sc_hd__nand3_1 U17660 ( .A(n12569), .B(n12568), .C(n12567), .Y(
        n16875) );
  sky130_fd_sc_hd__a22oi_1 U17661 ( .A1(n11551), .A2(
        j202_soc_core_j22_cpu_regop_imm__10_), .B1(n14069), .B2(
        j202_soc_core_j22_cpu_rf_vbr[10]), .Y(n12574) );
  sky130_fd_sc_hd__a2bb2oi_1 U17662 ( .B1(j202_soc_core_j22_cpu_rf_gpr[490]), 
        .B2(n14072), .A1_N(n14071), .A2_N(n16881), .Y(n12573) );
  sky130_fd_sc_hd__o22a_1 U17663 ( .A1(n12570), .A2(n14075), .B1(n16877), .B2(
        n14073), .X(n12572) );
  sky130_fd_sc_hd__o22a_1 U17664 ( .A1(n16876), .A2(n14079), .B1(n16880), .B2(
        n14077), .X(n12571) );
  sky130_fd_sc_hd__nand4_1 U17665 ( .A(n12574), .B(n12573), .C(n12572), .D(
        n12571), .Y(n12575) );
  sky130_fd_sc_hd__a21oi_1 U17666 ( .A1(n16875), .A2(n14086), .B1(n12575), .Y(
        n21807) );
  sky130_fd_sc_hd__nand2_1 U17667 ( .A(n21807), .B(n14087), .Y(n12576) );
  sky130_fd_sc_hd__nor2_1 U17669 ( .A(n12611), .B(n12612), .Y(n19511) );
  sky130_fd_sc_hd__o22ai_1 U17670 ( .A1(n20677), .A2(n22559), .B1(n22558), 
        .B2(n14042), .Y(n12609) );
  sky130_fd_sc_hd__nand2_1 U17671 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[169]), .Y(n12580) );
  sky130_fd_sc_hd__nand2_1 U17672 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[233]), .Y(n12579) );
  sky130_fd_sc_hd__nand2_1 U17673 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[489]), .Y(n12578) );
  sky130_fd_sc_hd__nand2_1 U17674 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[425]), .Y(n12577) );
  sky130_fd_sc_hd__nand4_1 U17675 ( .A(n12580), .B(n12579), .C(n12578), .D(
        n12577), .Y(n12586) );
  sky130_fd_sc_hd__nand2_1 U17676 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[393]), .Y(n12584) );
  sky130_fd_sc_hd__nand2_1 U17677 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[9]), .Y(n12583) );
  sky130_fd_sc_hd__nand2_1 U17678 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[41]), .Y(n12582) );
  sky130_fd_sc_hd__nand2_1 U17679 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[457]), .Y(n12581) );
  sky130_fd_sc_hd__nand4_1 U17680 ( .A(n12584), .B(n12583), .C(n12582), .D(
        n12581), .Y(n12585) );
  sky130_fd_sc_hd__nor2_1 U17681 ( .A(n12586), .B(n12585), .Y(n12597) );
  sky130_fd_sc_hd__nand2_1 U17682 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[329]), .Y(n12590) );
  sky130_fd_sc_hd__nand2_1 U17683 ( .A(n11191), .B(
        j202_soc_core_j22_cpu_rf_gpr[201]), .Y(n12589) );
  sky130_fd_sc_hd__nand2_1 U17684 ( .A(n20285), .B(
        j202_soc_core_j22_cpu_rf_gpr[297]), .Y(n12588) );
  sky130_fd_sc_hd__nand2_1 U17685 ( .A(n20282), .B(
        j202_soc_core_j22_cpu_rf_gpr[361]), .Y(n12587) );
  sky130_fd_sc_hd__and4_1 U17686 ( .A(n12590), .B(n12589), .C(n12588), .D(
        n12587), .X(n12596) );
  sky130_fd_sc_hd__nand2_1 U17687 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[137]), .Y(n12594) );
  sky130_fd_sc_hd__nand2_1 U17688 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[73]), .Y(n12593) );
  sky130_fd_sc_hd__nand2_1 U17689 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[105]), .Y(n12592) );
  sky130_fd_sc_hd__nand2_1 U17690 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[265]), .Y(n12591) );
  sky130_fd_sc_hd__and4_1 U17691 ( .A(n12594), .B(n12593), .C(n12592), .D(
        n12591), .X(n12595) );
  sky130_fd_sc_hd__nand3_1 U17692 ( .A(n12597), .B(n12596), .C(n12595), .Y(
        n19970) );
  sky130_fd_sc_hd__a22oi_1 U17693 ( .A1(n14072), .A2(
        j202_soc_core_j22_cpu_rf_gpr[489]), .B1(n14069), .B2(
        j202_soc_core_j22_cpu_rf_vbr[9]), .Y(n12602) );
  sky130_fd_sc_hd__o2bb2ai_1 U17694 ( .B1(n19974), .B2(n12943), .A1_N(n11551), 
        .A2_N(j202_soc_core_j22_cpu_regop_imm__9_), .Y(n12598) );
  sky130_fd_sc_hd__a21oi_1 U17695 ( .A1(n14028), .A2(
        j202_soc_core_j22_cpu_rf_gbr[9]), .B1(n12598), .Y(n12601) );
  sky130_fd_sc_hd__o22a_1 U17696 ( .A1(n19978), .A2(n14073), .B1(n14071), .B2(
        n19982), .X(n12600) );
  sky130_fd_sc_hd__o22a_1 U17697 ( .A1(n19984), .A2(n14075), .B1(n19972), .B2(
        n14079), .X(n12599) );
  sky130_fd_sc_hd__nand4_1 U17698 ( .A(n12602), .B(n12601), .C(n12600), .D(
        n12599), .Y(n12603) );
  sky130_fd_sc_hd__a21oi_1 U17699 ( .A1(n19970), .A2(n14086), .B1(n12603), .Y(
        n22314) );
  sky130_fd_sc_hd__nand2_1 U17700 ( .A(n22314), .B(n14087), .Y(n12604) );
  sky130_fd_sc_hd__o21ai_1 U17701 ( .A1(n14089), .A2(n22314), .B1(n12604), .Y(
        n12610) );
  sky130_fd_sc_hd__nor2_1 U17702 ( .A(n12609), .B(n12610), .Y(n18939) );
  sky130_fd_sc_hd__nor2_1 U17703 ( .A(n19511), .B(n18939), .Y(n12614) );
  sky130_fd_sc_hd__nand2_1 U17704 ( .A(n18940), .B(n12614), .Y(n18841) );
  sky130_fd_sc_hd__nor2_1 U17705 ( .A(n18837), .B(n18841), .Y(n12618) );
  sky130_fd_sc_hd__nand2_1 U17706 ( .A(n12606), .B(n12605), .Y(n19724) );
  sky130_fd_sc_hd__nand2_1 U17707 ( .A(n12608), .B(n12607), .Y(n19722) );
  sky130_fd_sc_hd__nand2_1 U17709 ( .A(n12610), .B(n12609), .Y(n19507) );
  sky130_fd_sc_hd__nand2_1 U17710 ( .A(n12612), .B(n12611), .Y(n19512) );
  sky130_fd_sc_hd__a21oi_1 U17712 ( .A1(n12614), .A2(n18941), .B1(n12613), .Y(
        n18840) );
  sky130_fd_sc_hd__nand2_1 U17713 ( .A(n12616), .B(n12615), .Y(n18838) );
  sky130_fd_sc_hd__a21oi_1 U17715 ( .A1(n16679), .A2(n12618), .B1(n12617), .Y(
        n18821) );
  sky130_fd_sc_hd__nand2_1 U17716 ( .A(n12620), .B(n12619), .Y(n18818) );
  sky130_fd_sc_hd__o21ai_1 U17717 ( .A1(n18817), .A2(n18821), .B1(n18818), .Y(
        n18829) );
  sky130_fd_sc_hd__o22ai_1 U17718 ( .A1(n14042), .A2(n22560), .B1(n22561), 
        .B2(n20677), .Y(n12649) );
  sky130_fd_sc_hd__nand2_1 U17719 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[173]), .Y(n12624) );
  sky130_fd_sc_hd__nand2_1 U17720 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[237]), .Y(n12623) );
  sky130_fd_sc_hd__nand2_1 U17721 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[493]), .Y(n12622) );
  sky130_fd_sc_hd__nand2_1 U17722 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[429]), .Y(n12621) );
  sky130_fd_sc_hd__nand4_1 U17723 ( .A(n12624), .B(n12623), .C(n12622), .D(
        n12621), .Y(n12630) );
  sky130_fd_sc_hd__nand2_1 U17724 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[397]), .Y(n12628) );
  sky130_fd_sc_hd__nand2_1 U17725 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[13]), .Y(n12627) );
  sky130_fd_sc_hd__nand2_1 U17726 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[45]), .Y(n12626) );
  sky130_fd_sc_hd__nand2_1 U17727 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[461]), .Y(n12625) );
  sky130_fd_sc_hd__nand4_1 U17728 ( .A(n12628), .B(n12627), .C(n12626), .D(
        n12625), .Y(n12629) );
  sky130_fd_sc_hd__nor2_1 U17729 ( .A(n12630), .B(n12629), .Y(n12641) );
  sky130_fd_sc_hd__nand2_1 U17730 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[333]), .Y(n12634) );
  sky130_fd_sc_hd__nand2_1 U17731 ( .A(n11191), .B(
        j202_soc_core_j22_cpu_rf_gpr[205]), .Y(n12633) );
  sky130_fd_sc_hd__nand2_1 U17732 ( .A(n20285), .B(
        j202_soc_core_j22_cpu_rf_gpr[301]), .Y(n12632) );
  sky130_fd_sc_hd__nand2_1 U17733 ( .A(n20282), .B(
        j202_soc_core_j22_cpu_rf_gpr[365]), .Y(n12631) );
  sky130_fd_sc_hd__and4_1 U17734 ( .A(n12634), .B(n12633), .C(n12632), .D(
        n12631), .X(n12640) );
  sky130_fd_sc_hd__nand2_1 U17735 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[141]), .Y(n12638) );
  sky130_fd_sc_hd__nand2_1 U17736 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[77]), .Y(n12637) );
  sky130_fd_sc_hd__nand2_1 U17737 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[109]), .Y(n12636) );
  sky130_fd_sc_hd__nand2_1 U17738 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[269]), .Y(n12635) );
  sky130_fd_sc_hd__and4_1 U17739 ( .A(n12638), .B(n12637), .C(n12636), .D(
        n12635), .X(n12639) );
  sky130_fd_sc_hd__nand3_1 U17740 ( .A(n12641), .B(n12640), .C(n12639), .Y(
        n19115) );
  sky130_fd_sc_hd__a21oi_1 U17741 ( .A1(n14069), .A2(
        j202_soc_core_j22_cpu_rf_vbr[13]), .B1(n14068), .Y(n12646) );
  sky130_fd_sc_hd__a2bb2oi_1 U17742 ( .B1(j202_soc_core_j22_cpu_rf_gpr[493]), 
        .B2(n14072), .A1_N(n14071), .A2_N(n19120), .Y(n12645) );
  sky130_fd_sc_hd__o22a_1 U17743 ( .A1(n19117), .A2(n14079), .B1(n19121), .B2(
        n14073), .X(n12644) );
  sky130_fd_sc_hd__o22a_1 U17744 ( .A1(n12642), .A2(n14075), .B1(n19116), .B2(
        n14077), .X(n12643) );
  sky130_fd_sc_hd__nand4_1 U17745 ( .A(n12646), .B(n12645), .C(n12644), .D(
        n12643), .Y(n12647) );
  sky130_fd_sc_hd__nand2_1 U17746 ( .A(n22300), .B(n14087), .Y(n12648) );
  sky130_fd_sc_hd__o21ai_1 U17747 ( .A1(n14089), .A2(n22300), .B1(n12648), .Y(
        n12650) );
  sky130_fd_sc_hd__nand2_1 U17748 ( .A(n12650), .B(n12649), .Y(n18828) );
  sky130_fd_sc_hd__nand2_1 U17749 ( .A(n12653), .B(n12652), .Y(n18806) );
  sky130_fd_sc_hd__o21ai_1 U17750 ( .A1(n18805), .A2(n18809), .B1(n18806), .Y(
        n19654) );
  sky130_fd_sc_hd__o22ai_1 U17751 ( .A1(n20677), .A2(n22556), .B1(n22562), 
        .B2(n14042), .Y(n12683) );
  sky130_fd_sc_hd__nand2_1 U17752 ( .A(n11191), .B(
        j202_soc_core_j22_cpu_rf_gpr[207]), .Y(n12657) );
  sky130_fd_sc_hd__nand2_1 U17753 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[335]), .Y(n12656) );
  sky130_fd_sc_hd__nand2_1 U17754 ( .A(n20285), .B(
        j202_soc_core_j22_cpu_rf_gpr[303]), .Y(n12655) );
  sky130_fd_sc_hd__nand2_1 U17755 ( .A(n20282), .B(
        j202_soc_core_j22_cpu_rf_gpr[367]), .Y(n12654) );
  sky130_fd_sc_hd__nand4_1 U17756 ( .A(n12657), .B(n12656), .C(n12655), .D(
        n12654), .Y(n12663) );
  sky130_fd_sc_hd__nand2_1 U17757 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[143]), .Y(n12661) );
  sky130_fd_sc_hd__nand2_1 U17758 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[79]), .Y(n12660) );
  sky130_fd_sc_hd__nand2_1 U17759 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[111]), .Y(n12659) );
  sky130_fd_sc_hd__nand2_1 U17760 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[271]), .Y(n12658) );
  sky130_fd_sc_hd__nand4_1 U17761 ( .A(n12661), .B(n12660), .C(n12659), .D(
        n12658), .Y(n12662) );
  sky130_fd_sc_hd__nor2_1 U17762 ( .A(n12663), .B(n12662), .Y(n12671) );
  sky130_fd_sc_hd__a22oi_1 U17763 ( .A1(n20301), .A2(
        j202_soc_core_j22_cpu_rf_gpr[239]), .B1(n20304), .B2(
        j202_soc_core_j22_cpu_rf_gpr[175]), .Y(n12670) );
  sky130_fd_sc_hd__a22oi_1 U17764 ( .A1(n20238), .A2(
        j202_soc_core_j22_cpu_rf_gpr[495]), .B1(n20288), .B2(
        j202_soc_core_j22_cpu_rf_gpr[431]), .Y(n12669) );
  sky130_fd_sc_hd__nand2_1 U17765 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[399]), .Y(n12667) );
  sky130_fd_sc_hd__nand2_1 U17766 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[15]), .Y(n12666) );
  sky130_fd_sc_hd__nand2_1 U17767 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[47]), .Y(n12665) );
  sky130_fd_sc_hd__nand2_1 U17768 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[463]), .Y(n12664) );
  sky130_fd_sc_hd__and4_1 U17769 ( .A(n12667), .B(n12666), .C(n12665), .D(
        n12664), .X(n12668) );
  sky130_fd_sc_hd__nand4_1 U17770 ( .A(n12671), .B(n12670), .C(n12669), .D(
        n12668), .Y(n15228) );
  sky130_fd_sc_hd__nand2_1 U17771 ( .A(n15228), .B(n14086), .Y(n12681) );
  sky130_fd_sc_hd__nand2_1 U17772 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[15]), .Y(n12674) );
  sky130_fd_sc_hd__nand2_1 U17773 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[15]), .Y(n12673) );
  sky130_fd_sc_hd__nand2_1 U17774 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[495]), .Y(n12672) );
  sky130_fd_sc_hd__and4_1 U17775 ( .A(n12674), .B(n12673), .C(n14022), .D(
        n12672), .X(n12680) );
  sky130_fd_sc_hd__o22ai_1 U17776 ( .A1(n12676), .A2(n14075), .B1(n14073), 
        .B2(n12675), .Y(n12678) );
  sky130_fd_sc_hd__o22ai_1 U17777 ( .A1(n15218), .A2(n14079), .B1(n14077), 
        .B2(n15217), .Y(n12677) );
  sky130_fd_sc_hd__nor2_1 U17778 ( .A(n12678), .B(n12677), .Y(n12679) );
  sky130_fd_sc_hd__nand3_1 U17779 ( .A(n12681), .B(n12680), .C(n12679), .Y(
        n22154) );
  sky130_fd_sc_hd__nand2_1 U17780 ( .A(n22275), .B(n14087), .Y(n12682) );
  sky130_fd_sc_hd__o21ai_1 U17781 ( .A1(n14089), .A2(n22275), .B1(n12682), .Y(
        n12684) );
  sky130_fd_sc_hd__nand2_1 U17782 ( .A(n12684), .B(n12683), .Y(n19653) );
  sky130_fd_sc_hd__a21oi_1 U17783 ( .A1(n19654), .A2(n11186), .B1(n12685), .Y(
        n18485) );
  sky130_fd_sc_hd__nand2_1 U17784 ( .A(n12687), .B(n12686), .Y(n18482) );
  sky130_fd_sc_hd__o22ai_1 U17786 ( .A1(n14042), .A2(n22563), .B1(n22565), 
        .B2(n20677), .Y(n12717) );
  sky130_fd_sc_hd__nand2_1 U17787 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[177]), .Y(n12691) );
  sky130_fd_sc_hd__nand2_1 U17788 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[241]), .Y(n12690) );
  sky130_fd_sc_hd__nand2_1 U17789 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[497]), .Y(n12689) );
  sky130_fd_sc_hd__nand2_1 U17790 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[433]), .Y(n12688) );
  sky130_fd_sc_hd__nand4_1 U17791 ( .A(n12691), .B(n12690), .C(n12689), .D(
        n12688), .Y(n12697) );
  sky130_fd_sc_hd__nand2_1 U17792 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[401]), .Y(n12695) );
  sky130_fd_sc_hd__nand2_1 U17793 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[17]), .Y(n12694) );
  sky130_fd_sc_hd__nand2_1 U17794 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[49]), .Y(n12693) );
  sky130_fd_sc_hd__nand2_1 U17795 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[465]), .Y(n12692) );
  sky130_fd_sc_hd__nand4_1 U17796 ( .A(n12695), .B(n12694), .C(n12693), .D(
        n12692), .Y(n12696) );
  sky130_fd_sc_hd__nor2_1 U17797 ( .A(n12697), .B(n12696), .Y(n12705) );
  sky130_fd_sc_hd__a22oi_1 U17798 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[305]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[209]), .Y(n12704) );
  sky130_fd_sc_hd__a22oi_1 U17799 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[369]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[337]), .Y(n12703) );
  sky130_fd_sc_hd__nand2_1 U17800 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[145]), .Y(n12701) );
  sky130_fd_sc_hd__nand2_1 U17801 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[81]), .Y(n12700) );
  sky130_fd_sc_hd__nand2_1 U17802 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[113]), .Y(n12699) );
  sky130_fd_sc_hd__nand2_1 U17803 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[273]), .Y(n12698) );
  sky130_fd_sc_hd__and4_1 U17804 ( .A(n12701), .B(n12700), .C(n12699), .D(
        n12698), .X(n12702) );
  sky130_fd_sc_hd__nand4_1 U17805 ( .A(n12705), .B(n12704), .C(n12703), .D(
        n12702), .Y(n19915) );
  sky130_fd_sc_hd__nand2_1 U17806 ( .A(n19915), .B(n14086), .Y(n12715) );
  sky130_fd_sc_hd__nand2_1 U17807 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[17]), .Y(n12708) );
  sky130_fd_sc_hd__nand2_1 U17808 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[17]), .Y(n12707) );
  sky130_fd_sc_hd__nand2_1 U17809 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[497]), .Y(n12706) );
  sky130_fd_sc_hd__and4_1 U17810 ( .A(n12708), .B(n12707), .C(n14022), .D(
        n12706), .X(n12714) );
  sky130_fd_sc_hd__nand2_1 U17811 ( .A(n14025), .B(
        j202_soc_core_j22_cpu_pc[17]), .Y(n12712) );
  sky130_fd_sc_hd__nand2_1 U17812 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[17]), .Y(n12711) );
  sky130_fd_sc_hd__nand2_1 U17813 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[17]), .Y(n12710) );
  sky130_fd_sc_hd__nand2_1 U17814 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[17]), .Y(n12709) );
  sky130_fd_sc_hd__and4_1 U17815 ( .A(n12712), .B(n12711), .C(n12710), .D(
        n12709), .X(n12713) );
  sky130_fd_sc_hd__nand3_1 U17816 ( .A(n12715), .B(n12714), .C(n12713), .Y(
        n23301) );
  sky130_fd_sc_hd__nand2_1 U17817 ( .A(n22116), .B(n14087), .Y(n12716) );
  sky130_fd_sc_hd__o21ai_1 U17818 ( .A1(n14089), .A2(n22116), .B1(n12716), .Y(
        n12718) );
  sky130_fd_sc_hd__nand2_1 U17819 ( .A(n12718), .B(n12717), .Y(n18493) );
  sky130_fd_sc_hd__nand2_1 U17820 ( .A(n12721), .B(n12720), .Y(n13542) );
  sky130_fd_sc_hd__o22ai_1 U17822 ( .A1(n20677), .A2(n22643), .B1(n22566), 
        .B2(n14042), .Y(n12751) );
  sky130_fd_sc_hd__nand2_1 U17823 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[179]), .Y(n12725) );
  sky130_fd_sc_hd__nand2_1 U17824 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[243]), .Y(n12724) );
  sky130_fd_sc_hd__nand2_1 U17825 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[499]), .Y(n12723) );
  sky130_fd_sc_hd__nand2_1 U17826 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[435]), .Y(n12722) );
  sky130_fd_sc_hd__nand4_1 U17827 ( .A(n12725), .B(n12724), .C(n12723), .D(
        n12722), .Y(n12731) );
  sky130_fd_sc_hd__nand2_1 U17828 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[403]), .Y(n12729) );
  sky130_fd_sc_hd__nand2_1 U17829 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[19]), .Y(n12728) );
  sky130_fd_sc_hd__nand2_1 U17830 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[51]), .Y(n12727) );
  sky130_fd_sc_hd__nand2_1 U17831 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[467]), .Y(n12726) );
  sky130_fd_sc_hd__nand4_1 U17832 ( .A(n12729), .B(n12728), .C(n12727), .D(
        n12726), .Y(n12730) );
  sky130_fd_sc_hd__nor2_1 U17833 ( .A(n12731), .B(n12730), .Y(n12739) );
  sky130_fd_sc_hd__a22oi_1 U17834 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[307]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[211]), .Y(n12738) );
  sky130_fd_sc_hd__a22oi_1 U17835 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[371]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[339]), .Y(n12737) );
  sky130_fd_sc_hd__nand2_1 U17836 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[147]), .Y(n12735) );
  sky130_fd_sc_hd__nand2_1 U17837 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[83]), .Y(n12734) );
  sky130_fd_sc_hd__nand2_1 U17838 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[115]), .Y(n12733) );
  sky130_fd_sc_hd__nand2_1 U17839 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[275]), .Y(n12732) );
  sky130_fd_sc_hd__and4_1 U17840 ( .A(n12735), .B(n12734), .C(n12733), .D(
        n12732), .X(n12736) );
  sky130_fd_sc_hd__nand4_1 U17841 ( .A(n12739), .B(n12738), .C(n12737), .D(
        n12736), .Y(n20054) );
  sky130_fd_sc_hd__nand2_1 U17842 ( .A(n20054), .B(n14086), .Y(n12749) );
  sky130_fd_sc_hd__nand2_1 U17843 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[19]), .Y(n12742) );
  sky130_fd_sc_hd__nand2_1 U17844 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[19]), .Y(n12741) );
  sky130_fd_sc_hd__nand2_1 U17845 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[499]), .Y(n12740) );
  sky130_fd_sc_hd__and4_1 U17846 ( .A(n12742), .B(n12741), .C(n14022), .D(
        n12740), .X(n12748) );
  sky130_fd_sc_hd__nand2_1 U17847 ( .A(n14025), .B(
        j202_soc_core_j22_cpu_pc[19]), .Y(n12746) );
  sky130_fd_sc_hd__nand2_1 U17848 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[19]), .Y(n12745) );
  sky130_fd_sc_hd__nand2_1 U17849 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[19]), .Y(n12744) );
  sky130_fd_sc_hd__nand2_1 U17850 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[19]), .Y(n12743) );
  sky130_fd_sc_hd__and4_1 U17851 ( .A(n12746), .B(n12745), .C(n12744), .D(
        n12743), .X(n12747) );
  sky130_fd_sc_hd__nand3_1 U17852 ( .A(n12749), .B(n12748), .C(n12747), .Y(
        n23307) );
  sky130_fd_sc_hd__nand2_1 U17853 ( .A(n22642), .B(n14087), .Y(n12750) );
  sky130_fd_sc_hd__o21ai_1 U17854 ( .A1(n14089), .A2(n22642), .B1(n12750), .Y(
        n12752) );
  sky130_fd_sc_hd__nand2_1 U17855 ( .A(n12752), .B(n12751), .Y(n13188) );
  sky130_fd_sc_hd__a21oi_1 U17856 ( .A1(n13189), .A2(n11192), .B1(n12753), .Y(
        n13407) );
  sky130_fd_sc_hd__nand2_1 U17857 ( .A(n12755), .B(n12754), .Y(n13404) );
  sky130_fd_sc_hd__o21ai_1 U17858 ( .A1(n13403), .A2(n13407), .B1(n13404), .Y(
        n13396) );
  sky130_fd_sc_hd__o22ai_1 U17859 ( .A1(n20677), .A2(n22600), .B1(n22641), 
        .B2(n14042), .Y(n12785) );
  sky130_fd_sc_hd__nand2_1 U17860 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[181]), .Y(n12759) );
  sky130_fd_sc_hd__nand2_1 U17861 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[245]), .Y(n12758) );
  sky130_fd_sc_hd__nand2_1 U17862 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[501]), .Y(n12757) );
  sky130_fd_sc_hd__nand2_1 U17863 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[437]), .Y(n12756) );
  sky130_fd_sc_hd__nand4_1 U17864 ( .A(n12759), .B(n12758), .C(n12757), .D(
        n12756), .Y(n12765) );
  sky130_fd_sc_hd__nand2_1 U17865 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[405]), .Y(n12763) );
  sky130_fd_sc_hd__nand2_1 U17866 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[21]), .Y(n12762) );
  sky130_fd_sc_hd__nand2_1 U17867 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[53]), .Y(n12761) );
  sky130_fd_sc_hd__nand2_1 U17868 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[469]), .Y(n12760) );
  sky130_fd_sc_hd__nand4_1 U17869 ( .A(n12763), .B(n12762), .C(n12761), .D(
        n12760), .Y(n12764) );
  sky130_fd_sc_hd__nor2_1 U17870 ( .A(n12765), .B(n12764), .Y(n12773) );
  sky130_fd_sc_hd__a22oi_1 U17871 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[309]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[213]), .Y(n12772) );
  sky130_fd_sc_hd__a22oi_1 U17872 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[373]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[341]), .Y(n12771) );
  sky130_fd_sc_hd__nand2_1 U17873 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[149]), .Y(n12769) );
  sky130_fd_sc_hd__nand2_1 U17874 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[85]), .Y(n12768) );
  sky130_fd_sc_hd__nand2_1 U17875 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[117]), .Y(n12767) );
  sky130_fd_sc_hd__nand2_1 U17876 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[277]), .Y(n12766) );
  sky130_fd_sc_hd__and4_1 U17877 ( .A(n12769), .B(n12768), .C(n12767), .D(
        n12766), .X(n12770) );
  sky130_fd_sc_hd__nand4_1 U17878 ( .A(n12773), .B(n12772), .C(n12771), .D(
        n12770), .Y(n19408) );
  sky130_fd_sc_hd__nand2_1 U17879 ( .A(n19408), .B(n14086), .Y(n12783) );
  sky130_fd_sc_hd__nand2_1 U17880 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[21]), .Y(n12776) );
  sky130_fd_sc_hd__nand2_1 U17881 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[21]), .Y(n12775) );
  sky130_fd_sc_hd__nand2_1 U17882 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[501]), .Y(n12774) );
  sky130_fd_sc_hd__and4_1 U17883 ( .A(n12776), .B(n12775), .C(n14022), .D(
        n12774), .X(n12782) );
  sky130_fd_sc_hd__nand2_1 U17884 ( .A(n14025), .B(
        j202_soc_core_j22_cpu_pc[21]), .Y(n12780) );
  sky130_fd_sc_hd__nand2_1 U17885 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[21]), .Y(n12779) );
  sky130_fd_sc_hd__nand2_1 U17886 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[21]), .Y(n12778) );
  sky130_fd_sc_hd__nand2_1 U17887 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[21]), .Y(n12777) );
  sky130_fd_sc_hd__and4_1 U17888 ( .A(n12780), .B(n12779), .C(n12778), .D(
        n12777), .X(n12781) );
  sky130_fd_sc_hd__nand3_1 U17889 ( .A(n12783), .B(n12782), .C(n12781), .Y(
        n23313) );
  sky130_fd_sc_hd__nand2_1 U17890 ( .A(n22599), .B(n14087), .Y(n12784) );
  sky130_fd_sc_hd__nand2_1 U17892 ( .A(n12786), .B(n12785), .Y(n13395) );
  sky130_fd_sc_hd__a21oi_1 U17893 ( .A1(n13396), .A2(n11188), .B1(n12787), .Y(
        n13297) );
  sky130_fd_sc_hd__nand2_1 U17894 ( .A(n12789), .B(n12788), .Y(n13294) );
  sky130_fd_sc_hd__o21ai_1 U17895 ( .A1(n13293), .A2(n13297), .B1(n13294), .Y(
        n13103) );
  sky130_fd_sc_hd__nand2_1 U17896 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[183]), .Y(n12793) );
  sky130_fd_sc_hd__nand2_1 U17897 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[439]), .Y(n12792) );
  sky130_fd_sc_hd__nand2_1 U17898 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[407]), .Y(n12791) );
  sky130_fd_sc_hd__nand2_1 U17899 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[503]), .Y(n12790) );
  sky130_fd_sc_hd__nand4_1 U17900 ( .A(n12793), .B(n12792), .C(n12791), .D(
        n12790), .Y(n12799) );
  sky130_fd_sc_hd__nand2_1 U17901 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[343]), .Y(n12797) );
  sky130_fd_sc_hd__nand2_1 U17902 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[215]), .Y(n12796) );
  sky130_fd_sc_hd__nand2_1 U17903 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[375]), .Y(n12795) );
  sky130_fd_sc_hd__nand2_1 U17904 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[151]), .Y(n12794) );
  sky130_fd_sc_hd__nand4_1 U17905 ( .A(n12797), .B(n12796), .C(n12795), .D(
        n12794), .Y(n12798) );
  sky130_fd_sc_hd__nor2_1 U17906 ( .A(n12799), .B(n12798), .Y(n12813) );
  sky130_fd_sc_hd__nor2_1 U17907 ( .A(n12800), .B(n13919), .Y(n12806) );
  sky130_fd_sc_hd__a21oi_1 U17908 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[23]), .B1(n13920), .Y(n12804) );
  sky130_fd_sc_hd__nand2_1 U17909 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[55]), .Y(n12803) );
  sky130_fd_sc_hd__nand2_1 U17910 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[247]), .Y(n12802) );
  sky130_fd_sc_hd__nand2_1 U17911 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[87]), .Y(n12801) );
  sky130_fd_sc_hd__nand4_1 U17912 ( .A(n12804), .B(n12803), .C(n12802), .D(
        n12801), .Y(n12805) );
  sky130_fd_sc_hd__nor2_1 U17913 ( .A(n12806), .B(n12805), .Y(n12812) );
  sky130_fd_sc_hd__nand2_1 U17914 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[311]), .Y(n12810) );
  sky130_fd_sc_hd__nand2_1 U17915 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[279]), .Y(n12809) );
  sky130_fd_sc_hd__nand2_1 U17916 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[119]), .Y(n12808) );
  sky130_fd_sc_hd__nand2_1 U17917 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[471]), .Y(n12807) );
  sky130_fd_sc_hd__and4_1 U17918 ( .A(n12810), .B(n12809), .C(n12808), .D(
        n12807), .X(n12811) );
  sky130_fd_sc_hd__nand3_1 U17919 ( .A(n12813), .B(n12812), .C(n12811), .Y(
        n21828) );
  sky130_fd_sc_hd__o22ai_1 U17920 ( .A1(n20677), .A2(n22614), .B1(n22567), 
        .B2(n14042), .Y(n12843) );
  sky130_fd_sc_hd__nand2_1 U17921 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[183]), .Y(n12817) );
  sky130_fd_sc_hd__nand2_1 U17922 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[247]), .Y(n12816) );
  sky130_fd_sc_hd__nand2_1 U17923 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[503]), .Y(n12815) );
  sky130_fd_sc_hd__nand2_1 U17924 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[439]), .Y(n12814) );
  sky130_fd_sc_hd__nand4_1 U17925 ( .A(n12817), .B(n12816), .C(n12815), .D(
        n12814), .Y(n12823) );
  sky130_fd_sc_hd__nand2_1 U17926 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[407]), .Y(n12821) );
  sky130_fd_sc_hd__nand2_1 U17927 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[23]), .Y(n12820) );
  sky130_fd_sc_hd__nand2_1 U17928 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[55]), .Y(n12819) );
  sky130_fd_sc_hd__nand2_1 U17929 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[471]), .Y(n12818) );
  sky130_fd_sc_hd__nand4_1 U17930 ( .A(n12821), .B(n12820), .C(n12819), .D(
        n12818), .Y(n12822) );
  sky130_fd_sc_hd__nor2_1 U17931 ( .A(n12823), .B(n12822), .Y(n12831) );
  sky130_fd_sc_hd__a22oi_1 U17932 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[311]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[215]), .Y(n12830) );
  sky130_fd_sc_hd__a22oi_1 U17933 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[375]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[343]), .Y(n12829) );
  sky130_fd_sc_hd__nand2_1 U17934 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[151]), .Y(n12827) );
  sky130_fd_sc_hd__nand2_1 U17935 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[87]), .Y(n12826) );
  sky130_fd_sc_hd__nand2_1 U17936 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[119]), .Y(n12825) );
  sky130_fd_sc_hd__nand2_1 U17937 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[279]), .Y(n12824) );
  sky130_fd_sc_hd__and4_1 U17938 ( .A(n12827), .B(n12826), .C(n12825), .D(
        n12824), .X(n12828) );
  sky130_fd_sc_hd__nand4_1 U17939 ( .A(n12831), .B(n12830), .C(n12829), .D(
        n12828), .Y(n19386) );
  sky130_fd_sc_hd__nand2_1 U17940 ( .A(n19386), .B(n14086), .Y(n12841) );
  sky130_fd_sc_hd__nand2_1 U17941 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[23]), .Y(n12834) );
  sky130_fd_sc_hd__nand2_1 U17942 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[23]), .Y(n12833) );
  sky130_fd_sc_hd__nand2_1 U17943 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[503]), .Y(n12832) );
  sky130_fd_sc_hd__and4_1 U17944 ( .A(n12834), .B(n12833), .C(n14022), .D(
        n12832), .X(n12840) );
  sky130_fd_sc_hd__nand2_1 U17945 ( .A(n14025), .B(
        j202_soc_core_j22_cpu_pc[23]), .Y(n12838) );
  sky130_fd_sc_hd__nand2_1 U17946 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[23]), .Y(n12837) );
  sky130_fd_sc_hd__nand2_1 U17947 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[23]), .Y(n12836) );
  sky130_fd_sc_hd__nand2_1 U17948 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[23]), .Y(n12835) );
  sky130_fd_sc_hd__and4_1 U17949 ( .A(n12838), .B(n12837), .C(n12836), .D(
        n12835), .X(n12839) );
  sky130_fd_sc_hd__nand3_1 U17950 ( .A(n12841), .B(n12840), .C(n12839), .Y(
        n23319) );
  sky130_fd_sc_hd__nand2_1 U17951 ( .A(n22613), .B(n14087), .Y(n12842) );
  sky130_fd_sc_hd__o21ai_1 U17952 ( .A1(n14089), .A2(n22613), .B1(n12842), .Y(
        n12844) );
  sky130_fd_sc_hd__nand2_1 U17953 ( .A(n12844), .B(n12843), .Y(n13102) );
  sky130_fd_sc_hd__a21oi_1 U17954 ( .A1(n13103), .A2(n11190), .B1(n12845), .Y(
        n13966) );
  sky130_fd_sc_hd__nand2_1 U17955 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[184]), .Y(n12849) );
  sky130_fd_sc_hd__nand2_1 U17956 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[248]), .Y(n12848) );
  sky130_fd_sc_hd__nand2_1 U17957 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[120]), .Y(n12847) );
  sky130_fd_sc_hd__nand2_1 U17958 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[408]), .Y(n12846) );
  sky130_fd_sc_hd__nand4_1 U17959 ( .A(n12849), .B(n12848), .C(n12847), .D(
        n12846), .Y(n12855) );
  sky130_fd_sc_hd__nand2_1 U17960 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[216]), .Y(n12853) );
  sky130_fd_sc_hd__nand2_1 U17961 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[344]), .Y(n12852) );
  sky130_fd_sc_hd__nand2_1 U17962 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[376]), .Y(n12851) );
  sky130_fd_sc_hd__nand2_1 U17963 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[152]), .Y(n12850) );
  sky130_fd_sc_hd__nand4_1 U17964 ( .A(n12853), .B(n12852), .C(n12851), .D(
        n12850), .Y(n12854) );
  sky130_fd_sc_hd__nor2_1 U17965 ( .A(n12855), .B(n12854), .Y(n12869) );
  sky130_fd_sc_hd__nor2_1 U17966 ( .A(n12856), .B(n13919), .Y(n12862) );
  sky130_fd_sc_hd__a21oi_1 U17967 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[24]), .B1(n13920), .Y(n12860) );
  sky130_fd_sc_hd__nand2_1 U17968 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[504]), .Y(n12859) );
  sky130_fd_sc_hd__nand2_1 U17969 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[56]), .Y(n12858) );
  sky130_fd_sc_hd__nand2_1 U17970 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[88]), .Y(n12857) );
  sky130_fd_sc_hd__nand4_1 U17971 ( .A(n12860), .B(n12859), .C(n12858), .D(
        n12857), .Y(n12861) );
  sky130_fd_sc_hd__nor2_1 U17972 ( .A(n12862), .B(n12861), .Y(n12868) );
  sky130_fd_sc_hd__nand2_1 U17973 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[312]), .Y(n12866) );
  sky130_fd_sc_hd__nand2_1 U17974 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[440]), .Y(n12865) );
  sky130_fd_sc_hd__nand2_1 U17975 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[280]), .Y(n12864) );
  sky130_fd_sc_hd__nand2_1 U17976 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[472]), .Y(n12863) );
  sky130_fd_sc_hd__and4_1 U17977 ( .A(n12866), .B(n12865), .C(n12864), .D(
        n12863), .X(n12867) );
  sky130_fd_sc_hd__nand3_1 U17978 ( .A(n12869), .B(n12868), .C(n12867), .Y(
        n21935) );
  sky130_fd_sc_hd__o22ai_1 U17979 ( .A1(n20677), .A2(n22568), .B1(n22614), 
        .B2(n14042), .Y(n12899) );
  sky130_fd_sc_hd__nand2_1 U17980 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[184]), .Y(n12873) );
  sky130_fd_sc_hd__nand2_1 U17981 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[248]), .Y(n12872) );
  sky130_fd_sc_hd__nand2_1 U17982 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[504]), .Y(n12871) );
  sky130_fd_sc_hd__nand2_1 U17983 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[440]), .Y(n12870) );
  sky130_fd_sc_hd__nand4_1 U17984 ( .A(n12873), .B(n12872), .C(n12871), .D(
        n12870), .Y(n12879) );
  sky130_fd_sc_hd__nand2_1 U17985 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[408]), .Y(n12877) );
  sky130_fd_sc_hd__nand2_1 U17986 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[24]), .Y(n12876) );
  sky130_fd_sc_hd__nand2_1 U17987 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[56]), .Y(n12875) );
  sky130_fd_sc_hd__nand2_1 U17988 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[472]), .Y(n12874) );
  sky130_fd_sc_hd__nand4_1 U17989 ( .A(n12877), .B(n12876), .C(n12875), .D(
        n12874), .Y(n12878) );
  sky130_fd_sc_hd__nor2_1 U17990 ( .A(n12879), .B(n12878), .Y(n12887) );
  sky130_fd_sc_hd__a22oi_1 U17991 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[312]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[216]), .Y(n12886) );
  sky130_fd_sc_hd__a22oi_1 U17992 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[376]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[344]), .Y(n12885) );
  sky130_fd_sc_hd__nand2_1 U17993 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[152]), .Y(n12883) );
  sky130_fd_sc_hd__nand2_1 U17994 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[88]), .Y(n12882) );
  sky130_fd_sc_hd__nand2_1 U17995 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[120]), .Y(n12881) );
  sky130_fd_sc_hd__nand2_1 U17996 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[280]), .Y(n12880) );
  sky130_fd_sc_hd__and4_1 U17997 ( .A(n12883), .B(n12882), .C(n12881), .D(
        n12880), .X(n12884) );
  sky130_fd_sc_hd__nand4_1 U17998 ( .A(n12887), .B(n12886), .C(n12885), .D(
        n12884), .Y(n19715) );
  sky130_fd_sc_hd__nand2_1 U17999 ( .A(n19715), .B(n14086), .Y(n12897) );
  sky130_fd_sc_hd__nand2_1 U18000 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[24]), .Y(n12890) );
  sky130_fd_sc_hd__nand2_1 U18001 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[24]), .Y(n12889) );
  sky130_fd_sc_hd__nand2_1 U18002 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[504]), .Y(n12888) );
  sky130_fd_sc_hd__and4_1 U18003 ( .A(n12890), .B(n12889), .C(n14022), .D(
        n12888), .X(n12896) );
  sky130_fd_sc_hd__nand2_1 U18004 ( .A(n14025), .B(
        j202_soc_core_j22_cpu_pc[24]), .Y(n12894) );
  sky130_fd_sc_hd__nand2_1 U18005 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[24]), .Y(n12893) );
  sky130_fd_sc_hd__nand2_1 U18006 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[24]), .Y(n12892) );
  sky130_fd_sc_hd__nand2_1 U18007 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[24]), .Y(n12891) );
  sky130_fd_sc_hd__and4_1 U18008 ( .A(n12894), .B(n12893), .C(n12892), .D(
        n12891), .X(n12895) );
  sky130_fd_sc_hd__nand3_1 U18009 ( .A(n12897), .B(n12896), .C(n12895), .Y(
        n23322) );
  sky130_fd_sc_hd__nand2_1 U18010 ( .A(n21840), .B(n14087), .Y(n12898) );
  sky130_fd_sc_hd__o21ai_1 U18011 ( .A1(n14089), .A2(n21840), .B1(n12898), .Y(
        n12900) );
  sky130_fd_sc_hd__nor2_1 U18012 ( .A(n12899), .B(n12900), .Y(n13967) );
  sky130_fd_sc_hd__nand2_1 U18013 ( .A(n12900), .B(n12899), .Y(n13965) );
  sky130_fd_sc_hd__nand2_1 U18014 ( .A(n12901), .B(n13965), .Y(n12902) );
  sky130_fd_sc_hd__xor2_1 U18015 ( .A(n13966), .B(n12902), .X(n21839) );
  sky130_fd_sc_hd__nor2_1 U18016 ( .A(n11202), .B(n12903), .Y(n12908) );
  sky130_fd_sc_hd__nand2_1 U18017 ( .A(n22687), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[4]), .Y(n22429) );
  sky130_fd_sc_hd__a21oi_1 U18018 ( .A1(n12904), .A2(n20836), .B1(n22429), .Y(
        n22791) );
  sky130_fd_sc_hd__nand2_1 U18019 ( .A(n12905), .B(n20836), .Y(n12906) );
  sky130_fd_sc_hd__nand2_1 U18020 ( .A(n22697), .B(
        j202_soc_core_j22_cpu_rfuo_sr__t_), .Y(n19253) );
  sky130_fd_sc_hd__nand2_1 U18021 ( .A(n12906), .B(n19253), .Y(n12907) );
  sky130_fd_sc_hd__nand2_1 U18022 ( .A(n22791), .B(n12907), .Y(n12986) );
  sky130_fd_sc_hd__nor2_1 U18023 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[2]), .B(
        j202_soc_core_j22_cpu_ma_M_MEM[3]), .Y(n12966) );
  sky130_fd_sc_hd__nand3_1 U18024 ( .A(n16643), .B(n12966), .C(n20352), .Y(
        n12909) );
  sky130_fd_sc_hd__nand2_1 U18025 ( .A(n21657), .B(
        j202_soc_core_j22_cpu_ifetchl), .Y(n20221) );
  sky130_fd_sc_hd__nand2_1 U18026 ( .A(n20506), .B(
        j202_soc_core_j22_cpu_regop_We__2_), .Y(n12910) );
  sky130_fd_sc_hd__nor2_1 U18027 ( .A(j202_soc_core_j22_cpu_regop_We__3_), .B(
        n12910), .Y(n20276) );
  sky130_fd_sc_hd__nand2_1 U18028 ( .A(n20276), .B(
        j202_soc_core_j22_cpu_regop_We__1_), .Y(n20239) );
  sky130_fd_sc_hd__nor2_1 U18029 ( .A(j202_soc_core_j22_cpu_memop_MEM__2_), 
        .B(j202_soc_core_j22_cpu_memop_MEM__1_), .Y(n13654) );
  sky130_fd_sc_hd__nand2_1 U18030 ( .A(n13654), .B(n23245), .Y(n14943) );
  sky130_fd_sc_hd__nand2b_1 U18031 ( .A_N(n14943), .B(
        j202_soc_core_j22_cpu_memop_MEM__0_), .Y(n22789) );
  sky130_fd_sc_hd__nand2_1 U18032 ( .A(n23245), .B(n23240), .Y(n21220) );
  sky130_fd_sc_hd__nand2_1 U18033 ( .A(n23243), .B(
        j202_soc_core_j22_cpu_memop_MEM__1_), .Y(n13652) );
  sky130_fd_sc_hd__o22a_1 U18034 ( .A1(n20479), .A2(n12910), .B1(n21220), .B2(
        n13652), .X(n12911) );
  sky130_fd_sc_hd__nand3_1 U18035 ( .A(n20239), .B(n22789), .C(n12911), .Y(
        n12912) );
  sky130_fd_sc_hd__nor2_1 U18036 ( .A(j202_soc_core_j22_cpu_opst[2]), .B(
        n22418), .Y(n21604) );
  sky130_fd_sc_hd__nand2_1 U18037 ( .A(n12912), .B(n21604), .Y(n12913) );
  sky130_fd_sc_hd__or3_1 U18038 ( .A(j202_soc_core_j22_cpu_opst[3]), .B(
        j202_soc_core_j22_cpu_opst[1]), .C(j202_soc_core_j22_cpu_opst[4]), .X(
        n21329) );
  sky130_fd_sc_hd__nor2_1 U18039 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__1_), 
        .B(j202_soc_core_j22_cpu_regop_M_Rn__0_), .Y(n20245) );
  sky130_fd_sc_hd__nor2_1 U18040 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__2_), 
        .B(j202_soc_core_j22_cpu_regop_M_Rn__3_), .Y(n20246) );
  sky130_fd_sc_hd__nand2_1 U18041 ( .A(n20245), .B(n20246), .Y(n12937) );
  sky130_fd_sc_hd__nand2_1 U18042 ( .A(n21657), .B(n12915), .Y(n12972) );
  sky130_fd_sc_hd__o21ai_1 U18043 ( .A1(j202_soc_core_j22_cpu_regop_other__2_), 
        .A2(n12916), .B1(j202_soc_core_j22_cpu_regop_Rs__0_), .Y(n12917) );
  sky130_fd_sc_hd__nand2_1 U18044 ( .A(n12917), .B(
        j202_soc_core_j22_cpu_regop_Rs__1_), .Y(n19983) );
  sky130_fd_sc_hd__nand2_1 U18045 ( .A(j202_soc_core_j22_cpu_regop_Ra__0_), 
        .B(j202_soc_core_j22_cpu_regop_Ra__1_), .Y(n12918) );
  sky130_fd_sc_hd__nand3_1 U18046 ( .A(n14075), .B(n19983), .C(n12918), .Y(
        n12919) );
  sky130_fd_sc_hd__o21ba_2 U18047 ( .A1(j202_soc_core_j22_cpu_regop_We__1_), 
        .A2(n12972), .B1_N(n12919), .X(n12976) );
  sky130_fd_sc_hd__a21oi_1 U18048 ( .A1(n21657), .A2(n20309), .B1(n12920), .Y(
        n12935) );
  sky130_fd_sc_hd__xnor2_1 U18049 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__1_), 
        .B(j202_soc_core_j22_cpu_regop_Rn__1_), .Y(n12924) );
  sky130_fd_sc_hd__xnor2_1 U18050 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__0_), 
        .B(j202_soc_core_j22_cpu_regop_Rn__0_), .Y(n12923) );
  sky130_fd_sc_hd__xnor2_1 U18051 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__2_), 
        .B(j202_soc_core_j22_cpu_regop_Rn__2_), .Y(n12922) );
  sky130_fd_sc_hd__xnor2_1 U18052 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__3_), 
        .B(j202_soc_core_j22_cpu_regop_Rn__3_), .Y(n12921) );
  sky130_fd_sc_hd__nand4_1 U18053 ( .A(n12924), .B(n12923), .C(n12922), .D(
        n12921), .Y(n12934) );
  sky130_fd_sc_hd__xnor2_1 U18054 ( .A(j202_soc_core_j22_cpu_regop_Rm__2_), 
        .B(j202_soc_core_j22_cpu_regop_M_Rn__2_), .Y(n12928) );
  sky130_fd_sc_hd__xnor2_1 U18055 ( .A(j202_soc_core_j22_cpu_regop_Rm__0_), 
        .B(j202_soc_core_j22_cpu_regop_M_Rn__0_), .Y(n12927) );
  sky130_fd_sc_hd__xnor2_1 U18056 ( .A(j202_soc_core_j22_cpu_regop_Rm__1_), 
        .B(j202_soc_core_j22_cpu_regop_M_Rn__1_), .Y(n12926) );
  sky130_fd_sc_hd__xnor2_1 U18057 ( .A(j202_soc_core_j22_cpu_regop_Rm__3_), 
        .B(j202_soc_core_j22_cpu_regop_M_Rn__3_), .Y(n12925) );
  sky130_fd_sc_hd__nand4_1 U18058 ( .A(n12928), .B(n12927), .C(n12926), .D(
        n12925), .Y(n12933) );
  sky130_fd_sc_hd__nand2_1 U18059 ( .A(n20506), .B(n20478), .Y(n12929) );
  sky130_fd_sc_hd__o22ai_1 U18060 ( .A1(j202_soc_core_j22_cpu_regop_Rs__1_), 
        .A2(n12931), .B1(j202_soc_core_j22_cpu_regop_Rb__1_), .B2(n12930), .Y(
        n12932) );
  sky130_fd_sc_hd__a21oi_1 U18061 ( .A1(n21657), .A2(n20256), .B1(n12932), .Y(
        n12970) );
  sky130_fd_sc_hd__o22a_1 U18062 ( .A1(n12935), .A2(n12934), .B1(n12933), .B2(
        n12970), .X(n12936) );
  sky130_fd_sc_hd__nor2_1 U18064 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__3_), 
        .B(j202_soc_core_j22_cpu_regop_M_Wm__0_), .Y(n23234) );
  sky130_fd_sc_hd__nand3_1 U18065 ( .A(n23234), .B(
        j202_soc_core_j22_cpu_regop_M_Wm__2_), .C(
        j202_soc_core_j22_cpu_regop_M_Wm__1_), .Y(n20234) );
  sky130_fd_sc_hd__nand2_1 U18066 ( .A(n12939), .B(n12938), .Y(n12982) );
  sky130_fd_sc_hd__nand2_1 U18067 ( .A(n20487), .B(
        j202_soc_core_j22_cpu_regop_M_Wm__0_), .Y(n20231) );
  sky130_fd_sc_hd__nand2_1 U18068 ( .A(j202_soc_core_j22_cpu_regop_Rs__1_), 
        .B(j202_soc_core_j22_cpu_regop_Rs__0_), .Y(n15214) );
  sky130_fd_sc_hd__nor2_1 U18069 ( .A(j202_soc_core_j22_cpu_regop_other__2_), 
        .B(n15214), .Y(n15216) );
  sky130_fd_sc_hd__nand2_1 U18070 ( .A(n15216), .B(n12940), .Y(n19971) );
  sky130_fd_sc_hd__nand2_1 U18071 ( .A(n14079), .B(n19971), .Y(n12945) );
  sky130_fd_sc_hd__nor2_1 U18072 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__2_), 
        .B(n20235), .Y(n20274) );
  sky130_fd_sc_hd__nand3_1 U18073 ( .A(n12942), .B(n15220), .C(n12941), .Y(
        n19973) );
  sky130_fd_sc_hd__nand2_1 U18074 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__2_), 
        .B(j202_soc_core_j22_cpu_regop_M_Wm__1_), .Y(n20482) );
  sky130_fd_sc_hd__a21oi_1 U18075 ( .A1(n12943), .A2(n19973), .B1(n20482), .Y(
        n12944) );
  sky130_fd_sc_hd__a21oi_1 U18076 ( .A1(n12945), .A2(n20274), .B1(n12944), .Y(
        n12962) );
  sky130_fd_sc_hd__nor4_1 U18077 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__3_), 
        .B(j202_soc_core_j22_cpu_regop_M_Wm__0_), .C(
        j202_soc_core_j22_cpu_regop_M_Wm__2_), .D(n20235), .Y(n20225) );
  sky130_fd_sc_hd__nand2b_1 U18078 ( .A_N(n14073), .B(n20225), .Y(n14939) );
  sky130_fd_sc_hd__nor2_1 U18079 ( .A(n12947), .B(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[4]), .Y(n12952) );
  sky130_fd_sc_hd__a21oi_1 U18080 ( .A1(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]), .A2(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[3]), .B1(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .Y(n12946) );
  sky130_fd_sc_hd__nor2b_1 U18081 ( .B_N(n12952), .A(n12946), .Y(n20098) );
  sky130_fd_sc_hd__nand3_1 U18082 ( .A(n15241), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .C(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .Y(n21664) );
  sky130_fd_sc_hd__nand3_1 U18083 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[4]), .B(n12947), .C(n22128), .Y(
        n20099) );
  sky130_fd_sc_hd__a21oi_1 U18084 ( .A1(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]), .A2(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .B1(n20099), .Y(n22147) );
  sky130_fd_sc_hd__nand3_1 U18085 ( .A(n12949), .B(n21664), .C(n12948), .Y(
        n21671) );
  sky130_fd_sc_hd__nand2_1 U18086 ( .A(j202_soc_core_j22_cpu_macop_MAC_[3]), 
        .B(j202_soc_core_j22_cpu_macop_MAC_[1]), .Y(n21654) );
  sky130_fd_sc_hd__nand2_1 U18087 ( .A(j202_soc_core_j22_cpu_macop_MAC_[0]), 
        .B(n21679), .Y(n21676) );
  sky130_fd_sc_hd__a21oi_1 U18088 ( .A1(j202_soc_core_j22_cpu_macop_MAC_[3]), 
        .A2(j202_soc_core_j22_cpu_macop_MAC_[0]), .B1(
        j202_soc_core_j22_cpu_macop_MAC_[1]), .Y(n21678) );
  sky130_fd_sc_hd__nand3_1 U18089 ( .A(n12950), .B(
        j202_soc_core_j22_cpu_macop_MAC_[2]), .C(n23247), .Y(n20085) );
  sky130_fd_sc_hd__nor2_1 U18090 ( .A(j202_soc_core_j22_cpu_macop_MAC_[2]), 
        .B(j202_soc_core_j22_cpu_macop_MAC_[3]), .Y(n21675) );
  sky130_fd_sc_hd__nand3_1 U18091 ( .A(n21675), .B(
        j202_soc_core_j22_cpu_macop_MAC_[4]), .C(n22923), .Y(n21650) );
  sky130_fd_sc_hd__nand2_1 U18093 ( .A(n21671), .B(n21656), .Y(n12954) );
  sky130_fd_sc_hd__nor2_1 U18094 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .B(n21659), .Y(n15234) );
  sky130_fd_sc_hd__nand2_1 U18095 ( .A(n15234), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .Y(n16594) );
  sky130_fd_sc_hd__nor2_1 U18096 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .B(j202_soc_core_j22_cpu_ml_X_macop_MAC_[0]), .Y(n15237) );
  sky130_fd_sc_hd__nand2_1 U18097 ( .A(n15241), .B(n15237), .Y(n21665) );
  sky130_fd_sc_hd__o21a_1 U18098 ( .A1(n16596), .A2(n16594), .B1(n21665), .X(
        n20089) );
  sky130_fd_sc_hd__nand2_1 U18099 ( .A(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .B(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[3]), .Y(n20097) );
  sky130_fd_sc_hd__nand2_1 U18100 ( .A(n12953), .B(n12952), .Y(n23347) );
  sky130_fd_sc_hd__nand3_1 U18101 ( .A(n12954), .B(n20089), .C(n23347), .Y(
        n12961) );
  sky130_fd_sc_hd__nand2_1 U18102 ( .A(n22923), .B(n22125), .Y(n12955) );
  sky130_fd_sc_hd__nor2_1 U18103 ( .A(n12955), .B(
        j202_soc_core_j22_cpu_macop_MAC_[4]), .Y(n12956) );
  sky130_fd_sc_hd__nand2_1 U18104 ( .A(n21675), .B(n12956), .Y(n12960) );
  sky130_fd_sc_hd__nand2_1 U18105 ( .A(n15232), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .Y(n21723) );
  sky130_fd_sc_hd__nand2_1 U18106 ( .A(n15232), .B(n15234), .Y(n15233) );
  sky130_fd_sc_hd__nand4_1 U18107 ( .A(n16594), .B(n21675), .C(
        j202_soc_core_j22_cpu_macop_MAC_[1]), .D(n23247), .Y(n12958) );
  sky130_fd_sc_hd__a21oi_1 U18108 ( .A1(n21723), .A2(n15233), .B1(n12958), .Y(
        n12959) );
  sky130_fd_sc_hd__a21oi_1 U18109 ( .A1(n12961), .A2(n12960), .B1(n12959), .Y(
        n21652) );
  sky130_fd_sc_hd__o211ai_1 U18110 ( .A1(n20231), .A2(n12962), .B1(n14939), 
        .C1(n21652), .Y(n12969) );
  sky130_fd_sc_hd__nor3_1 U18111 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[2]), 
        .B(n22695), .C(n22429), .Y(n12965) );
  sky130_fd_sc_hd__nand3_1 U18112 ( .A(n22670), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[0]), .C(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n12963) );
  sky130_fd_sc_hd__nor2_1 U18113 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[3]), 
        .B(n22670), .Y(n19254) );
  sky130_fd_sc_hd__nand2_1 U18114 ( .A(n19254), .B(n22428), .Y(n22688) );
  sky130_fd_sc_hd__o22ai_1 U18115 ( .A1(n12963), .A2(n14042), .B1(
        j202_soc_core_j22_cpu_exuop_EXU_[0]), .B2(n22688), .Y(n12964) );
  sky130_fd_sc_hd__nor2_1 U18116 ( .A(n12965), .B(n12964), .Y(n12968) );
  sky130_fd_sc_hd__nand2_1 U18117 ( .A(n22530), .B(n12966), .Y(n12967) );
  sky130_fd_sc_hd__nor2_1 U18118 ( .A(n12968), .B(n23235), .Y(n22801) );
  sky130_fd_sc_hd__nand2_1 U18119 ( .A(n12972), .B(n12971), .Y(n12974) );
  sky130_fd_sc_hd__a22oi_1 U18120 ( .A1(n12975), .A2(n20250), .B1(n12974), 
        .B2(n12973), .Y(n12977) );
  sky130_fd_sc_hd__nand2_1 U18121 ( .A(n12977), .B(n12976), .Y(n12979) );
  sky130_fd_sc_hd__nand2_1 U18122 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__2_), 
        .B(n23234), .Y(n12978) );
  sky130_fd_sc_hd__nor2_1 U18123 ( .A(j202_soc_core_j22_cpu_regop_M_Wm__1_), 
        .B(n12978), .Y(n20247) );
  sky130_fd_sc_hd__nand2_1 U18124 ( .A(n12979), .B(n20247), .Y(n12980) );
  sky130_fd_sc_hd__nand2b_1 U18125 ( .A_N(n14943), .B(n23240), .Y(n21213) );
  sky130_fd_sc_hd__nand2_1 U18126 ( .A(n23239), .B(n21213), .Y(n12985) );
  sky130_fd_sc_hd__nand2b_1 U18127 ( .A_N(n23235), .B(n21215), .Y(n12984) );
  sky130_fd_sc_hd__nand2_1 U18128 ( .A(n21839), .B(n19729), .Y(n13101) );
  sky130_fd_sc_hd__nor2_1 U18129 ( .A(n22790), .B(n12986), .Y(n21616) );
  sky130_fd_sc_hd__nand2b_1 U18130 ( .A_N(n13095), .B(n21616), .Y(n19734) );
  sky130_fd_sc_hd__nand2_1 U18131 ( .A(j202_soc_core_bootrom_00_address_w[10]), 
        .B(j202_soc_core_bootrom_00_address_w[3]), .Y(n17778) );
  sky130_fd_sc_hd__nor2_1 U18132 ( .A(n14999), .B(n17778), .Y(n14141) );
  sky130_fd_sc_hd__nand2_1 U18133 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .B(j202_soc_core_bootrom_00_address_w[6]), .Y(n14605) );
  sky130_fd_sc_hd__nand2_1 U18134 ( .A(n14141), .B(n12989), .Y(n14219) );
  sky130_fd_sc_hd__nor2_1 U18135 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n14219), .Y(n14624) );
  sky130_fd_sc_hd__nor2_1 U18136 ( .A(j202_soc_core_bootrom_00_address_w[7]), 
        .B(n17778), .Y(n14102) );
  sky130_fd_sc_hd__nor2_1 U18137 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(n13210), .Y(n14292) );
  sky130_fd_sc_hd__nand2_1 U18138 ( .A(n14292), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n13008) );
  sky130_fd_sc_hd__nor2_1 U18139 ( .A(n14575), .B(n13008), .Y(n14636) );
  sky130_fd_sc_hd__nand2_1 U18140 ( .A(n14292), .B(n13014), .Y(n13016) );
  sky130_fd_sc_hd__nand2_1 U18141 ( .A(n14235), .B(n14141), .Y(n14566) );
  sky130_fd_sc_hd__nand2_1 U18142 ( .A(n14980), .B(
        j202_soc_core_bootrom_00_address_w[7]), .Y(n14296) );
  sky130_fd_sc_hd__nand2_1 U18143 ( .A(n13031), .B(n14104), .Y(n14580) );
  sky130_fd_sc_hd__nand2_1 U18144 ( .A(n14566), .B(n14580), .Y(n13055) );
  sky130_fd_sc_hd__nor3_1 U18145 ( .A(n14624), .B(n14636), .C(n13055), .Y(
        n14218) );
  sky130_fd_sc_hd__nor2_1 U18146 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(j202_soc_core_bootrom_00_address_w[9]), .Y(n14313) );
  sky130_fd_sc_hd__nand2_1 U18147 ( .A(n14313), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n13015) );
  sky130_fd_sc_hd__nor2_1 U18148 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(j202_soc_core_bootrom_00_address_w[9]), .Y(n13025) );
  sky130_fd_sc_hd__nand2_1 U18149 ( .A(n13025), .B(n14998), .Y(n14310) );
  sky130_fd_sc_hd__o21a_1 U18151 ( .A1(n14296), .A2(n13015), .B1(n14186), .X(
        n14286) );
  sky130_fd_sc_hd__nand2_1 U18152 ( .A(n14399), .B(n14100), .Y(n14293) );
  sky130_fd_sc_hd__nor2_1 U18153 ( .A(n13014), .B(n14605), .Y(n13005) );
  sky130_fd_sc_hd__nand2_1 U18154 ( .A(n14571), .B(n13005), .Y(n14567) );
  sky130_fd_sc_hd__nor2_1 U18155 ( .A(n13014), .B(n14219), .Y(n14278) );
  sky130_fd_sc_hd__nor2_1 U18156 ( .A(n13016), .B(n14296), .Y(n14630) );
  sky130_fd_sc_hd__nor2_1 U18157 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .B(n14998), .Y(n14201) );
  sky130_fd_sc_hd__nor2_1 U18158 ( .A(n12987), .B(n14296), .Y(n14188) );
  sky130_fd_sc_hd__nand2_1 U18159 ( .A(n14188), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n14185) );
  sky130_fd_sc_hd__nand2_1 U18160 ( .A(n14201), .B(n13014), .Y(n14576) );
  sky130_fd_sc_hd__nand2_1 U18161 ( .A(n14571), .B(n13028), .Y(n14637) );
  sky130_fd_sc_hd__nand2_1 U18162 ( .A(n14185), .B(n14637), .Y(n14585) );
  sky130_fd_sc_hd__nor4_1 U18163 ( .A(n14579), .B(n14278), .C(n14630), .D(
        n14585), .Y(n12988) );
  sky130_fd_sc_hd__a31oi_1 U18164 ( .A1(n14218), .A2(n14286), .A3(n12988), 
        .B1(n14639), .Y(n13000) );
  sky130_fd_sc_hd__nor2_1 U18165 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n14605), .Y(n13018) );
  sky130_fd_sc_hd__nand2_1 U18166 ( .A(n13018), .B(n14571), .Y(n14625) );
  sky130_fd_sc_hd__nand2_1 U18167 ( .A(n13018), .B(n14102), .Y(n14287) );
  sky130_fd_sc_hd__nand2_1 U18168 ( .A(n14287), .B(n14186), .Y(n14577) );
  sky130_fd_sc_hd__nor4b_1 U18169 ( .D_N(n12988), .A(n14565), .B(n14277), .C(
        n14577), .Y(n12990) );
  sky130_fd_sc_hd__nand2_1 U18170 ( .A(n14104), .B(n12989), .Y(n14288) );
  sky130_fd_sc_hd__nand2_1 U18171 ( .A(n13027), .B(n14141), .Y(n13054) );
  sky130_fd_sc_hd__a31oi_1 U18172 ( .A1(n12990), .A2(n14288), .A3(n13054), 
        .B1(n14631), .Y(n12999) );
  sky130_fd_sc_hd__nand2_1 U18173 ( .A(n14549), .B(n14141), .Y(n13063) );
  sky130_fd_sc_hd__nor2_1 U18174 ( .A(n13015), .B(n14296), .Y(n12992) );
  sky130_fd_sc_hd__nand2_1 U18175 ( .A(n12991), .B(n14201), .Y(n14184) );
  sky130_fd_sc_hd__nand2_1 U18176 ( .A(n13031), .B(n14141), .Y(n14632) );
  sky130_fd_sc_hd__nand2_1 U18177 ( .A(n14201), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n13017) );
  sky130_fd_sc_hd__nor2_1 U18178 ( .A(n17778), .B(n13017), .Y(n14570) );
  sky130_fd_sc_hd__nand2_1 U18179 ( .A(n14570), .B(n14999), .Y(n14280) );
  sky130_fd_sc_hd__nand2_1 U18180 ( .A(n14571), .B(n13031), .Y(n14332) );
  sky130_fd_sc_hd__nand3_1 U18181 ( .A(n14632), .B(n14280), .C(n14332), .Y(
        n14618) );
  sky130_fd_sc_hd__nor4b_1 U18182 ( .D_N(n13063), .A(n12992), .B(n14283), .C(
        n14618), .Y(n12993) );
  sky130_fd_sc_hd__a21oi_1 U18183 ( .A1(n12993), .A2(n14625), .B1(n15149), .Y(
        n12998) );
  sky130_fd_sc_hd__a21oi_1 U18185 ( .A1(n14201), .A2(n14571), .B1(n13058), .Y(
        n12996) );
  sky130_fd_sc_hd__a31oi_1 U18186 ( .A1(n12996), .A2(n13063), .A3(n14632), 
        .B1(n14619), .Y(n12997) );
  sky130_fd_sc_hd__nor4_1 U18187 ( .A(n13000), .B(n12999), .C(n12998), .D(
        n12997), .Y(n13003) );
  sky130_fd_sc_hd__nor2_1 U18188 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n14288), .Y(n13066) );
  sky130_fd_sc_hd__nor2_1 U18189 ( .A(n13066), .B(n14579), .Y(n14621) );
  sky130_fd_sc_hd__nand2_1 U18190 ( .A(n13027), .B(n14571), .Y(n14279) );
  sky130_fd_sc_hd__nand2_1 U18191 ( .A(n13056), .B(n14313), .Y(n13001) );
  sky130_fd_sc_hd__nand2_1 U18192 ( .A(n13027), .B(n14102), .Y(n14627) );
  sky130_fd_sc_hd__nand2_1 U18193 ( .A(n14102), .B(n14292), .Y(n13065) );
  sky130_fd_sc_hd__nand2b_1 U18194 ( .A_N(n13065), .B(n13014), .Y(n14333) );
  sky130_fd_sc_hd__nand4_1 U18195 ( .A(n14583), .B(n13001), .C(n14627), .D(
        n14333), .Y(n14291) );
  sky130_fd_sc_hd__a21oi_1 U18196 ( .A1(j202_soc_core_bootrom_00_address_w[7]), 
        .A2(n14570), .B1(n14291), .Y(n14569) );
  sky130_fd_sc_hd__nand4b_1 U18197 ( .A_N(n14585), .B(n14621), .C(n14569), .D(
        n14287), .Y(n13002) );
  sky130_fd_sc_hd__nor2_1 U18198 ( .A(n13066), .B(n14300), .Y(n14574) );
  sky130_fd_sc_hd__nor2_1 U18199 ( .A(n14295), .B(n14575), .Y(n14284) );
  sky130_fd_sc_hd__a21oi_1 U18200 ( .A1(n14574), .A2(n14330), .B1(n14619), .Y(
        n14307) );
  sky130_fd_sc_hd__a21oi_1 U18201 ( .A1(n15093), .A2(n13002), .B1(n14307), .Y(
        n14190) );
  sky130_fd_sc_hd__nand2_1 U18202 ( .A(n13003), .B(n14190), .Y(n13004) );
  sky130_fd_sc_hd__nor2_1 U18203 ( .A(j202_soc_core_bootrom_00_address_w[11]), 
        .B(j202_soc_core_bootrom_00_address_w[8]), .Y(n14308) );
  sky130_fd_sc_hd__nand2_1 U18204 ( .A(n13004), .B(n14308), .Y(n13071) );
  sky130_fd_sc_hd__nor2_1 U18205 ( .A(j202_soc_core_bootrom_00_address_w[7]), 
        .B(n14978), .Y(n14723) );
  sky130_fd_sc_hd__nand2_1 U18206 ( .A(n14723), .B(n14201), .Y(n13013) );
  sky130_fd_sc_hd__nor2_1 U18207 ( .A(j202_soc_core_bootrom_00_address_w[2]), 
        .B(n13013), .Y(n13042) );
  sky130_fd_sc_hd__nor2_1 U18208 ( .A(j202_soc_core_bootrom_00_address_w[7]), 
        .B(n14108), .Y(n14314) );
  sky130_fd_sc_hd__nor2_1 U18209 ( .A(n14110), .B(n14310), .Y(n14607) );
  sky130_fd_sc_hd__nand2b_1 U18210 ( .A_N(n13016), .B(n14096), .Y(n14200) );
  sky130_fd_sc_hd__nor2_1 U18211 ( .A(j202_soc_core_bootrom_00_address_w[3]), 
        .B(n14200), .Y(n14211) );
  sky130_fd_sc_hd__nor2_1 U18212 ( .A(n14999), .B(n14978), .Y(n14404) );
  sky130_fd_sc_hd__nand2_1 U18213 ( .A(n14404), .B(n13018), .Y(n14342) );
  sky130_fd_sc_hd__nor2_1 U18214 ( .A(n14999), .B(n14108), .Y(n13032) );
  sky130_fd_sc_hd__nand2_1 U18215 ( .A(n13032), .B(n13005), .Y(n13033) );
  sky130_fd_sc_hd__nand2_1 U18216 ( .A(n14342), .B(n13033), .Y(n14230) );
  sky130_fd_sc_hd__nor2_1 U18217 ( .A(n14211), .B(n14230), .Y(n14552) );
  sky130_fd_sc_hd__nor2_1 U18218 ( .A(n14605), .B(n13006), .Y(n14196) );
  sky130_fd_sc_hd__nand2_1 U18219 ( .A(n14196), .B(
        j202_soc_core_bootrom_00_address_w[3]), .Y(n14344) );
  sky130_fd_sc_hd__nand2_1 U18220 ( .A(n14552), .B(n14344), .Y(n14600) );
  sky130_fd_sc_hd__nand2_1 U18221 ( .A(n13031), .B(n14236), .Y(n13041) );
  sky130_fd_sc_hd__nand2_1 U18222 ( .A(n13007), .B(n14100), .Y(n14591) );
  sky130_fd_sc_hd__nor4_1 U18224 ( .A(n13042), .B(n14607), .C(n14600), .D(
        n14343), .Y(n13011) );
  sky130_fd_sc_hd__nor2_1 U18225 ( .A(n14103), .B(n13008), .Y(n14232) );
  sky130_fd_sc_hd__nor2_1 U18226 ( .A(n13016), .B(n14309), .Y(n13009) );
  sky130_fd_sc_hd__nor2_1 U18227 ( .A(n14100), .B(n14200), .Y(n14553) );
  sky130_fd_sc_hd__nor2_1 U18228 ( .A(n13012), .B(n14309), .Y(n14537) );
  sky130_fd_sc_hd__nand3_1 U18229 ( .A(n14314), .B(
        j202_soc_core_bootrom_00_address_w[9]), .C(n13014), .Y(n14209) );
  sky130_fd_sc_hd__nand2_1 U18230 ( .A(n14572), .B(n14314), .Y(n14227) );
  sky130_fd_sc_hd__nand2_1 U18231 ( .A(n13032), .B(n13027), .Y(n13044) );
  sky130_fd_sc_hd__nand4b_1 U18232 ( .A_N(n14537), .B(n14209), .C(n14227), .D(
        n13044), .Y(n13034) );
  sky130_fd_sc_hd__nor4_1 U18233 ( .A(n14232), .B(n13009), .C(n14553), .D(
        n13034), .Y(n13010) );
  sky130_fd_sc_hd__a21oi_1 U18234 ( .A1(n13011), .A2(n13010), .B1(n14631), .Y(
        n13024) );
  sky130_fd_sc_hd__nor2_1 U18235 ( .A(n14161), .B(n13012), .Y(n14597) );
  sky130_fd_sc_hd__a21oi_1 U18236 ( .A1(n13032), .A2(n14572), .B1(n14537), .Y(
        n14546) );
  sky130_fd_sc_hd__nand2_1 U18237 ( .A(n14196), .B(n14100), .Y(n14550) );
  sky130_fd_sc_hd__nand3_1 U18238 ( .A(n14542), .B(n14546), .C(n14550), .Y(
        n14354) );
  sky130_fd_sc_hd__nor2_1 U18239 ( .A(n14597), .B(n14354), .Y(n14557) );
  sky130_fd_sc_hd__nand2_1 U18240 ( .A(n13027), .B(n14982), .Y(n14205) );
  sky130_fd_sc_hd__a21oi_1 U18241 ( .A1(n14557), .A2(n14205), .B1(n14619), .Y(
        n13023) );
  sky130_fd_sc_hd__nand2_1 U18242 ( .A(n14161), .B(n14309), .Y(n14548) );
  sky130_fd_sc_hd__nand2_1 U18243 ( .A(n13033), .B(n14592), .Y(n14543) );
  sky130_fd_sc_hd__a21oi_1 U18244 ( .A1(n13025), .A2(n14548), .B1(n14543), .Y(
        n13021) );
  sky130_fd_sc_hd__nor2_1 U18245 ( .A(n13014), .B(n13013), .Y(n14229) );
  sky130_fd_sc_hd__nor2_1 U18246 ( .A(n14110), .B(n13015), .Y(n13046) );
  sky130_fd_sc_hd__o21bai_1 U18247 ( .A1(n14604), .A2(n13016), .B1_N(n13046), 
        .Y(n14601) );
  sky130_fd_sc_hd__nor2b_1 U18248 ( .B_N(n14342), .A(n14601), .Y(n14603) );
  sky130_fd_sc_hd__nor2_1 U18249 ( .A(n14604), .B(n14310), .Y(n14207) );
  sky130_fd_sc_hd__nor2_1 U18250 ( .A(j202_soc_core_bootrom_00_address_w[7]), 
        .B(n14205), .Y(n14539) );
  sky130_fd_sc_hd__nor2_1 U18251 ( .A(n14207), .B(n14539), .Y(n14593) );
  sky130_fd_sc_hd__nand2_1 U18252 ( .A(n14603), .B(n14593), .Y(n14199) );
  sky130_fd_sc_hd__nor2_1 U18253 ( .A(n14103), .B(n14576), .Y(n14311) );
  sky130_fd_sc_hd__nand2_1 U18254 ( .A(n13032), .B(n13028), .Y(n14350) );
  sky130_fd_sc_hd__nor2_1 U18256 ( .A(n14311), .B(n14325), .Y(n14198) );
  sky130_fd_sc_hd__nand2_1 U18257 ( .A(n14314), .B(n13018), .Y(n14202) );
  sky130_fd_sc_hd__nor2b_1 U18258 ( .B_N(n14202), .A(n14232), .Y(n14351) );
  sky130_fd_sc_hd__nand2_1 U18259 ( .A(n13032), .B(n14549), .Y(n13040) );
  sky130_fd_sc_hd__nand4_1 U18260 ( .A(n14198), .B(n14351), .C(n13041), .D(
        n13040), .Y(n13019) );
  sky130_fd_sc_hd__nor4_1 U18261 ( .A(n14229), .B(n14554), .C(n14199), .D(
        n13019), .Y(n13020) );
  sky130_fd_sc_hd__o22ai_1 U18262 ( .A1(n13021), .A2(n15149), .B1(n13020), 
        .B2(n14639), .Y(n13022) );
  sky130_fd_sc_hd__nor3_1 U18263 ( .A(n13024), .B(n13023), .C(n13022), .Y(
        n13053) );
  sky130_fd_sc_hd__nand2_1 U18264 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .B(j202_soc_core_bootrom_00_address_w[11]), .Y(n14562) );
  sky130_fd_sc_hd__nand2_1 U18265 ( .A(n13231), .B(
        j202_soc_core_bootrom_00_address_w[11]), .Y(n14615) );
  sky130_fd_sc_hd__o21ai_1 U18266 ( .A1(n13025), .A2(n13027), .B1(n14404), .Y(
        n14555) );
  sky130_fd_sc_hd__nand2_1 U18268 ( .A(n14208), .B(n13044), .Y(n14544) );
  sky130_fd_sc_hd__nor2b_1 U18269 ( .B_N(n14555), .A(n14544), .Y(n14594) );
  sky130_fd_sc_hd__nand2_1 U18270 ( .A(n14572), .B(n13032), .Y(n13026) );
  sky130_fd_sc_hd__nand2_1 U18271 ( .A(n14314), .B(n14235), .Y(n14315) );
  sky130_fd_sc_hd__nand4b_1 U18272 ( .A_N(n14232), .B(n14594), .C(n13026), .D(
        n14315), .Y(n14322) );
  sky130_fd_sc_hd__nand2_1 U18274 ( .A(n14572), .B(n14404), .Y(n13029) );
  sky130_fd_sc_hd__nand3_1 U18275 ( .A(n13036), .B(n13029), .C(n13041), .Y(
        n13030) );
  sky130_fd_sc_hd__nor3_1 U18276 ( .A(n14211), .B(n14322), .C(n13030), .Y(
        n14228) );
  sky130_fd_sc_hd__nand2_1 U18277 ( .A(n13032), .B(n13031), .Y(n14349) );
  sky130_fd_sc_hd__a31oi_1 U18279 ( .A1(n14228), .A2(n14345), .A3(n14202), 
        .B1(n14639), .Y(n13051) );
  sky130_fd_sc_hd__nand2_1 U18280 ( .A(n14200), .B(n14344), .Y(n13039) );
  sky130_fd_sc_hd__nand2_1 U18281 ( .A(n14404), .B(n14549), .Y(n14540) );
  sky130_fd_sc_hd__nand2_1 U18282 ( .A(n14540), .B(n13033), .Y(n14206) );
  sky130_fd_sc_hd__nor2_1 U18283 ( .A(n14103), .B(n14295), .Y(n14598) );
  sky130_fd_sc_hd__nor2_1 U18284 ( .A(n14538), .B(n14598), .Y(n13035) );
  sky130_fd_sc_hd__nor2_1 U18285 ( .A(n14358), .B(n13034), .Y(n14319) );
  sky130_fd_sc_hd__nand3_1 U18286 ( .A(n13036), .B(n13035), .C(n14319), .Y(
        n14231) );
  sky130_fd_sc_hd__nor3_1 U18287 ( .A(n13039), .B(n14206), .C(n14231), .Y(
        n13038) );
  sky130_fd_sc_hd__a31oi_1 U18288 ( .A1(n13038), .A2(n14349), .A3(n13037), 
        .B1(n15149), .Y(n13050) );
  sky130_fd_sc_hd__nor2_1 U18289 ( .A(n14310), .B(n14575), .Y(n14602) );
  sky130_fd_sc_hd__nor3b_1 U18290 ( .C_N(n13044), .A(n14602), .B(n13039), .Y(
        n14317) );
  sky130_fd_sc_hd__nand2_1 U18291 ( .A(n14317), .B(n14540), .Y(n14234) );
  sky130_fd_sc_hd__nor4b_1 U18292 ( .D_N(n14227), .A(n14325), .B(n14199), .C(
        n14234), .Y(n13048) );
  sky130_fd_sc_hd__nand2_1 U18293 ( .A(n14205), .B(n13040), .Y(n14204) );
  sky130_fd_sc_hd__nor2_1 U18294 ( .A(n14100), .B(n13041), .Y(n14357) );
  sky130_fd_sc_hd__nand2_1 U18295 ( .A(n13043), .B(n14227), .Y(n14194) );
  sky130_fd_sc_hd__nand4_1 U18296 ( .A(n13044), .B(n14200), .C(n14202), .D(
        n14627), .Y(n13045) );
  sky130_fd_sc_hd__nor3_1 U18297 ( .A(n14357), .B(n14194), .C(n13045), .Y(
        n14596) );
  sky130_fd_sc_hd__nand2_1 U18298 ( .A(n14596), .B(n14279), .Y(n14326) );
  sky130_fd_sc_hd__nor4_1 U18299 ( .A(n13046), .B(n14204), .C(n14230), .D(
        n14326), .Y(n13047) );
  sky130_fd_sc_hd__o22ai_1 U18300 ( .A1(n13048), .A2(n14631), .B1(n13047), 
        .B2(n14619), .Y(n13049) );
  sky130_fd_sc_hd__nor3_1 U18301 ( .A(n13051), .B(n13050), .C(n13049), .Y(
        n13052) );
  sky130_fd_sc_hd__o22a_1 U18302 ( .A1(n13053), .A2(n14562), .B1(n14615), .B2(
        n13052), .X(n13070) );
  sky130_fd_sc_hd__nand2b_1 U18303 ( .A_N(n13055), .B(n13054), .Y(n13057) );
  sky130_fd_sc_hd__a21oi_1 U18304 ( .A1(n13056), .A2(n14292), .B1(n13057), .Y(
        n14331) );
  sky130_fd_sc_hd__nor2_1 U18305 ( .A(n14602), .B(n14278), .Y(n14337) );
  sky130_fd_sc_hd__a31oi_1 U18306 ( .A1(n14331), .A2(n14337), .A3(n14632), 
        .B1(n14639), .Y(n14638) );
  sky130_fd_sc_hd__nor3_1 U18307 ( .A(n14602), .B(n14284), .C(n13057), .Y(
        n14620) );
  sky130_fd_sc_hd__a31oi_1 U18308 ( .A1(n14620), .A2(n14219), .A3(n13063), 
        .B1(n14619), .Y(n13062) );
  sky130_fd_sc_hd__nand2_1 U18309 ( .A(n14571), .B(n14235), .Y(n14289) );
  sky130_fd_sc_hd__nor2_1 U18310 ( .A(n14310), .B(n14296), .Y(n13064) );
  sky130_fd_sc_hd__nor2_1 U18311 ( .A(n13064), .B(n13058), .Y(n13059) );
  sky130_fd_sc_hd__nand2_1 U18312 ( .A(n14289), .B(n13059), .Y(n14623) );
  sky130_fd_sc_hd__a31oi_1 U18313 ( .A1(n14102), .A2(n13210), .A3(n14576), 
        .B1(n14623), .Y(n13060) );
  sky130_fd_sc_hd__a21oi_1 U18314 ( .A1(n13060), .A2(n14566), .B1(n15149), .Y(
        n13061) );
  sky130_fd_sc_hd__nor3_1 U18315 ( .A(n14638), .B(n13062), .C(n13061), .Y(
        n14220) );
  sky130_fd_sc_hd__nand2_1 U18316 ( .A(n14287), .B(n13063), .Y(n14298) );
  sky130_fd_sc_hd__nor4_1 U18317 ( .A(n14188), .B(n14570), .C(n13064), .D(
        n14298), .Y(n14634) );
  sky130_fd_sc_hd__nand2_1 U18318 ( .A(n14634), .B(n14637), .Y(n14217) );
  sky130_fd_sc_hd__nand2b_1 U18319 ( .A_N(n14578), .B(n14566), .Y(n14282) );
  sky130_fd_sc_hd__o31ai_1 U18320 ( .A1(n13066), .A2(n14217), .A3(n14282), 
        .B1(n14348), .Y(n13067) );
  sky130_fd_sc_hd__nand2_1 U18321 ( .A(n14220), .B(n13067), .Y(n13068) );
  sky130_fd_sc_hd__nand2_1 U18322 ( .A(n15017), .B(
        j202_soc_core_bootrom_00_address_w[8]), .Y(n14339) );
  sky130_fd_sc_hd__nand2_1 U18323 ( .A(n13068), .B(n14645), .Y(n13069) );
  sky130_fd_sc_hd__nand3_1 U18324 ( .A(n13071), .B(n13070), .C(n13069), .Y(
        n13072) );
  sky130_fd_sc_hd__nand2_1 U18325 ( .A(n13072), .B(n14668), .Y(n13091) );
  sky130_fd_sc_hd__nand2_1 U18326 ( .A(n18379), .B(j202_soc_core_uart_div0[0]), 
        .Y(n13076) );
  sky130_fd_sc_hd__nand2_1 U18327 ( .A(n18727), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[88]), .Y(n13075) );
  sky130_fd_sc_hd__nand2_1 U18328 ( .A(n18725), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[24]), .Y(n13074) );
  sky130_fd_sc_hd__nand2_1 U18329 ( .A(n18726), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[56]), .Y(n13073) );
  sky130_fd_sc_hd__and4_1 U18330 ( .A(n13076), .B(n13075), .C(n13074), .D(
        n13073), .X(n13090) );
  sky130_fd_sc_hd__a22oi_1 U18331 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[184]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[152]), .Y(n13080) );
  sky130_fd_sc_hd__a22oi_1 U18332 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[248]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[216]), .Y(n13079) );
  sky130_fd_sc_hd__a22o_1 U18333 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[24]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[88]), .X(n13077) );
  sky130_fd_sc_hd__a21oi_1 U18334 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[120]), .B1(n13077), .Y(n13078) );
  sky130_fd_sc_hd__a31oi_1 U18335 ( .A1(n13080), .A2(n13079), .A3(n13078), 
        .B1(n18736), .Y(n13085) );
  sky130_fd_sc_hd__a22oi_1 U18336 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[472]), .B1(n18745), .B2(
        j202_soc_core_memory0_ram_dout0[408]), .Y(n13083) );
  sky130_fd_sc_hd__a21oi_1 U18337 ( .A1(n18746), .A2(
        j202_soc_core_memory0_ram_dout0[440]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n13082) );
  sky130_fd_sc_hd__a22oi_1 U18338 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[344]), .B1(n18743), .B2(
        j202_soc_core_memory0_ram_dout0[376]), .Y(n13081) );
  sky130_fd_sc_hd__nand3_1 U18339 ( .A(n13083), .B(n13082), .C(n13081), .Y(
        n13084) );
  sky130_fd_sc_hd__a211oi_1 U18340 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[312]), .B1(n13085), .C1(n13084), .Y(
        n13087) );
  sky130_fd_sc_hd__a22oi_1 U18341 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[280]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[56]), .Y(n13086) );
  sky130_fd_sc_hd__nand2_1 U18342 ( .A(n13087), .B(n13086), .Y(n13088) );
  sky130_fd_sc_hd__o211ai_1 U18343 ( .A1(j202_soc_core_memory0_ram_dout0[504]), 
        .A2(n18758), .B1(n14906), .C1(n13088), .Y(n13089) );
  sky130_fd_sc_hd__nand3_1 U18344 ( .A(n13091), .B(n13090), .C(n13089), .Y(
        n22524) );
  sky130_fd_sc_hd__nand2_1 U18345 ( .A(n22524), .B(n19737), .Y(n13098) );
  sky130_fd_sc_hd__nand3_1 U18346 ( .A(n19078), .B(
        j202_soc_core_j22_cpu_memop_Ma__0_), .C(n13092), .Y(n19731) );
  sky130_fd_sc_hd__nand2_1 U18347 ( .A(n13093), .B(n22790), .Y(n20835) );
  sky130_fd_sc_hd__nor2_1 U18348 ( .A(n20835), .B(n13094), .Y(n21621) );
  sky130_fd_sc_hd__nand3_1 U18350 ( .A(n19078), .B(
        j202_soc_core_j22_cpu_memop_Ma__1_), .C(n13096), .Y(n18948) );
  sky130_fd_sc_hd__a22oi_1 U18351 ( .A1(n19657), .A2(n21935), .B1(n19736), 
        .B2(n23322), .Y(n13097) );
  sky130_fd_sc_hd__nand2_1 U18352 ( .A(n13098), .B(n13097), .Y(n13099) );
  sky130_fd_sc_hd__a21oi_1 U18353 ( .A1(n21842), .A2(n19661), .B1(n13099), .Y(
        n13100) );
  sky130_fd_sc_hd__nand2_1 U18354 ( .A(n13101), .B(n13100), .Y(n25257) );
  sky130_fd_sc_hd__nand2_1 U18355 ( .A(n11190), .B(n13102), .Y(n13104) );
  sky130_fd_sc_hd__xnor2_1 U18356 ( .A(n13104), .B(n13103), .Y(n21823) );
  sky130_fd_sc_hd__nand2_1 U18357 ( .A(n21823), .B(n19729), .Y(n13187) );
  sky130_fd_sc_hd__ha_1 U18358 ( .A(j202_soc_core_j22_cpu_pc[23]), .B(n13105), 
        .COUT(n14175), .SUM(n21825) );
  sky130_fd_sc_hd__a31oi_1 U18359 ( .A1(n13415), .A2(n13106), .A3(n13112), 
        .B1(n17730), .Y(n13305) );
  sky130_fd_sc_hd__nor3_1 U18360 ( .A(n13333), .B(n13463), .C(n13107), .Y(
        n13410) );
  sky130_fd_sc_hd__nand2_1 U18361 ( .A(n13413), .B(n14724), .Y(n17988) );
  sky130_fd_sc_hd__nor2_1 U18362 ( .A(n14680), .B(n13332), .Y(n13108) );
  sky130_fd_sc_hd__o22ai_1 U18363 ( .A1(n13410), .A2(n13464), .B1(n13108), 
        .B2(n17730), .Y(n13118) );
  sky130_fd_sc_hd__nand2_1 U18364 ( .A(n13110), .B(n13109), .Y(n13364) );
  sky130_fd_sc_hd__nor4_1 U18365 ( .A(n13411), .B(n13314), .C(n13421), .D(
        n13364), .Y(n13116) );
  sky130_fd_sc_hd__nand4_1 U18366 ( .A(n13301), .B(n13124), .C(n13112), .D(
        n13111), .Y(n13113) );
  sky130_fd_sc_hd__nor3_1 U18367 ( .A(n13114), .B(n13299), .C(n13113), .Y(
        n13115) );
  sky130_fd_sc_hd__o22ai_1 U18368 ( .A1(n13116), .A2(n13500), .B1(n13115), 
        .B2(n17468), .Y(n13117) );
  sky130_fd_sc_hd__nor3_1 U18369 ( .A(n13305), .B(n13118), .C(n13117), .Y(
        n13119) );
  sky130_fd_sc_hd__nand2b_1 U18370 ( .A_N(n13119), .B(n17609), .Y(n13182) );
  sky130_fd_sc_hd__nor2_1 U18371 ( .A(j202_soc_core_bootrom_00_address_w[11]), 
        .B(n14111), .Y(n17469) );
  sky130_fd_sc_hd__nand2_1 U18372 ( .A(n17469), .B(n14098), .Y(n14155) );
  sky130_fd_sc_hd__or4_1 U18373 ( .A(n13433), .B(n13485), .C(n14683), .D(
        n13120), .X(n13122) );
  sky130_fd_sc_hd__nand3_1 U18375 ( .A(n13125), .B(n13380), .C(n13124), .Y(
        n13371) );
  sky130_fd_sc_hd__nor3_1 U18376 ( .A(n13372), .B(n13127), .C(n13126), .Y(
        n13128) );
  sky130_fd_sc_hd__o22ai_1 U18377 ( .A1(n13129), .A2(n17730), .B1(n13128), 
        .B2(n17468), .Y(n13130) );
  sky130_fd_sc_hd__a21oi_1 U18378 ( .A1(n13496), .A2(n13371), .B1(n13130), .Y(
        n13131) );
  sky130_fd_sc_hd__nand2_1 U18379 ( .A(n13132), .B(n13131), .Y(n13164) );
  sky130_fd_sc_hd__a31oi_1 U18380 ( .A1(n13133), .A2(n13134), .A3(n13166), 
        .B1(n17730), .Y(n13141) );
  sky130_fd_sc_hd__a31oi_1 U18381 ( .A1(n13492), .A2(n13134), .A3(n13165), 
        .B1(n13500), .Y(n13140) );
  sky130_fd_sc_hd__nor3_1 U18382 ( .A(n13333), .B(n13452), .C(n13135), .Y(
        n13138) );
  sky130_fd_sc_hd__nand2_1 U18383 ( .A(n13480), .B(n13311), .Y(n13370) );
  sky130_fd_sc_hd__nand2_1 U18384 ( .A(n13380), .B(n13329), .Y(n13309) );
  sky130_fd_sc_hd__nor3_1 U18385 ( .A(n13434), .B(n13370), .C(n13309), .Y(
        n13137) );
  sky130_fd_sc_hd__o22ai_1 U18386 ( .A1(n13138), .A2(n17468), .B1(n13137), 
        .B2(n13464), .Y(n13139) );
  sky130_fd_sc_hd__nor3_1 U18387 ( .A(n13141), .B(n13140), .C(n13139), .Y(
        n13162) );
  sky130_fd_sc_hd__a22oi_1 U18388 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[247]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[215]), .Y(n13145) );
  sky130_fd_sc_hd__a22oi_1 U18389 ( .A1(n18734), .A2(
        j202_soc_core_memory0_ram_dout0[151]), .B1(n18733), .B2(
        j202_soc_core_memory0_ram_dout0[119]), .Y(n13144) );
  sky130_fd_sc_hd__a22oi_1 U18390 ( .A1(n18361), .A2(
        j202_soc_core_memory0_ram_dout0[55]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[87]), .Y(n13143) );
  sky130_fd_sc_hd__nand2_1 U18391 ( .A(n18735), .B(
        j202_soc_core_memory0_ram_dout0[183]), .Y(n13142) );
  sky130_fd_sc_hd__nand4_1 U18392 ( .A(n13145), .B(n13144), .C(n13143), .D(
        n13142), .Y(n13146) );
  sky130_fd_sc_hd__a21oi_1 U18393 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[23]), .B1(n13146), .Y(n13147) );
  sky130_fd_sc_hd__nand2b_1 U18394 ( .A_N(n13147), .B(n17639), .Y(n13155) );
  sky130_fd_sc_hd__a22oi_1 U18395 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[311]), .B1(n18062), .B2(
        j202_soc_core_memory0_ram_dout0[279]), .Y(n13154) );
  sky130_fd_sc_hd__nand2_1 U18396 ( .A(n18743), .B(
        j202_soc_core_memory0_ram_dout0[375]), .Y(n13151) );
  sky130_fd_sc_hd__a21oi_1 U18397 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[471]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n13150) );
  sky130_fd_sc_hd__nand2_1 U18398 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[407]), .Y(n13149) );
  sky130_fd_sc_hd__nand2_1 U18399 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[439]), .Y(n13148) );
  sky130_fd_sc_hd__nand4_1 U18400 ( .A(n13151), .B(n13150), .C(n13149), .D(
        n13148), .Y(n13152) );
  sky130_fd_sc_hd__a21oi_1 U18401 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[343]), .B1(n13152), .Y(n13153) );
  sky130_fd_sc_hd__nand3_1 U18402 ( .A(n13155), .B(n13154), .C(n13153), .Y(
        n13156) );
  sky130_fd_sc_hd__o211ai_1 U18403 ( .A1(j202_soc_core_memory0_ram_dout0[503]), 
        .A2(n18758), .B1(n14906), .C1(n13156), .Y(n13160) );
  sky130_fd_sc_hd__a22oi_1 U18404 ( .A1(n18726), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[55]), .B1(n18379), .B2(
        j202_soc_core_uart_div1[7]), .Y(n13159) );
  sky130_fd_sc_hd__a22oi_1 U18405 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[23]), .B1(n18727), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[87]), .Y(n13158) );
  sky130_fd_sc_hd__nand2_1 U18406 ( .A(n18629), .B(
        j202_soc_core_bldc_core_00_pwm_duty[11]), .Y(n13157) );
  sky130_fd_sc_hd__nand4_1 U18407 ( .A(n13160), .B(n13159), .C(n13158), .D(
        n13157), .Y(n13161) );
  sky130_fd_sc_hd__o21bai_1 U18408 ( .A1(n13162), .A2(n18666), .B1_N(n13161), 
        .Y(n13163) );
  sky130_fd_sc_hd__a21oi_1 U18409 ( .A1(n13164), .A2(n18798), .B1(n13163), .Y(
        n13181) );
  sky130_fd_sc_hd__nand2_1 U18410 ( .A(n13166), .B(n13165), .Y(n13324) );
  sky130_fd_sc_hd__nor2_1 U18411 ( .A(n13325), .B(n13167), .Y(n13461) );
  sky130_fd_sc_hd__nand4_1 U18412 ( .A(n13366), .B(n13369), .C(n13168), .D(
        n13461), .Y(n13178) );
  sky130_fd_sc_hd__a21oi_1 U18413 ( .A1(n13169), .A2(n13329), .B1(n13464), .Y(
        n13177) );
  sky130_fd_sc_hd__nand2_1 U18415 ( .A(n13365), .B(n13172), .Y(n13432) );
  sky130_fd_sc_hd__nor3_1 U18416 ( .A(n13378), .B(n13432), .C(n13173), .Y(
        n13174) );
  sky130_fd_sc_hd__o22ai_1 U18417 ( .A1(n13175), .A2(n13500), .B1(n13174), 
        .B2(n17730), .Y(n13176) );
  sky130_fd_sc_hd__a211oi_1 U18418 ( .A1(n13489), .A2(n13178), .B1(n13177), 
        .C1(n13176), .Y(n13179) );
  sky130_fd_sc_hd__nand2b_1 U18419 ( .A_N(n13179), .B(n18605), .Y(n13180) );
  sky130_fd_sc_hd__nand2_1 U18420 ( .A(n22531), .B(n19737), .Y(n13184) );
  sky130_fd_sc_hd__a22oi_1 U18421 ( .A1(n19657), .A2(n21828), .B1(n19736), 
        .B2(n23319), .Y(n13183) );
  sky130_fd_sc_hd__nand2_1 U18422 ( .A(n13184), .B(n13183), .Y(n13185) );
  sky130_fd_sc_hd__a21oi_1 U18423 ( .A1(n21825), .A2(n19661), .B1(n13185), .Y(
        n13186) );
  sky130_fd_sc_hd__nand2_1 U18424 ( .A(n13187), .B(n13186), .Y(n25280) );
  sky130_fd_sc_hd__nand2_1 U18425 ( .A(n11192), .B(n13188), .Y(n13190) );
  sky130_fd_sc_hd__xnor2_1 U18426 ( .A(n13190), .B(n13189), .Y(n21756) );
  sky130_fd_sc_hd__nand2_1 U18427 ( .A(n21756), .B(n19729), .Y(n13292) );
  sky130_fd_sc_hd__ha_1 U18428 ( .A(j202_soc_core_j22_cpu_pc[19]), .B(n13191), 
        .COUT(n13408), .SUM(n21758) );
  sky130_fd_sc_hd__nor2_1 U18429 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .B(n14100), .Y(n18161) );
  sky130_fd_sc_hd__nand2_1 U18430 ( .A(n14456), .B(n13210), .Y(n13596) );
  sky130_fd_sc_hd__nor2_1 U18431 ( .A(n13213), .B(n13596), .Y(n18045) );
  sky130_fd_sc_hd__nand2_1 U18432 ( .A(n15017), .B(
        j202_soc_core_bootrom_00_address_w[9]), .Y(n13246) );
  sky130_fd_sc_hd__nor2_1 U18433 ( .A(n13449), .B(n13246), .Y(n13194) );
  sky130_fd_sc_hd__nand2_1 U18434 ( .A(n13194), .B(n14472), .Y(n18007) );
  sky130_fd_sc_hd__nor2_1 U18435 ( .A(n18045), .B(n18041), .Y(n18144) );
  sky130_fd_sc_hd__nand2_1 U18436 ( .A(n13192), .B(
        j202_soc_core_bootrom_00_address_w[10]), .Y(n13222) );
  sky130_fd_sc_hd__nor2_1 U18437 ( .A(n13246), .B(n13222), .Y(n18006) );
  sky130_fd_sc_hd__nand2_1 U18438 ( .A(n18006), .B(
        j202_soc_core_bootrom_00_address_w[7]), .Y(n13234) );
  sky130_fd_sc_hd__nor2_1 U18439 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .B(n14777), .Y(n13608) );
  sky130_fd_sc_hd__nand2_1 U18440 ( .A(n13234), .B(n18086), .Y(n18024) );
  sky130_fd_sc_hd__nand2_1 U18441 ( .A(n13193), .B(n14399), .Y(n13197) );
  sky130_fd_sc_hd__nor2_1 U18442 ( .A(n14101), .B(n13197), .Y(n18031) );
  sky130_fd_sc_hd__nand2_1 U18443 ( .A(n13194), .B(n13198), .Y(n13223) );
  sky130_fd_sc_hd__or3_1 U18444 ( .A(n18024), .B(n18031), .C(n17991), .X(
        n18098) );
  sky130_fd_sc_hd__nor2_1 U18445 ( .A(n18114), .B(n18098), .Y(n17983) );
  sky130_fd_sc_hd__nand2_1 U18446 ( .A(n13195), .B(n13199), .Y(n13581) );
  sky130_fd_sc_hd__nand2_1 U18447 ( .A(n13196), .B(n13210), .Y(n13236) );
  sky130_fd_sc_hd__nand2_1 U18448 ( .A(n15016), .B(n13255), .Y(n13240) );
  sky130_fd_sc_hd__nor2_1 U18449 ( .A(n13553), .B(n18044), .Y(n18154) );
  sky130_fd_sc_hd__nand2b_1 U18450 ( .A_N(n18125), .B(n13210), .Y(n13235) );
  sky130_fd_sc_hd__nor2_1 U18451 ( .A(n13222), .B(n13596), .Y(n18132) );
  sky130_fd_sc_hd__nor2_1 U18452 ( .A(n18101), .B(n18132), .Y(n13610) );
  sky130_fd_sc_hd__nand2_1 U18453 ( .A(n15016), .B(
        j202_soc_core_bootrom_00_address_w[10]), .Y(n14988) );
  sky130_fd_sc_hd__nor2_1 U18454 ( .A(n13246), .B(n14988), .Y(n17990) );
  sky130_fd_sc_hd__nand2_1 U18455 ( .A(n17990), .B(
        j202_soc_core_bootrom_00_address_w[7]), .Y(n18180) );
  sky130_fd_sc_hd__nor2_1 U18456 ( .A(n15016), .B(n13236), .Y(n18124) );
  sky130_fd_sc_hd__nor2_1 U18457 ( .A(n17975), .B(n18124), .Y(n17971) );
  sky130_fd_sc_hd__nor2b_1 U18458 ( .B_N(n18180), .A(n18039), .Y(n18174) );
  sky130_fd_sc_hd__nand4_1 U18459 ( .A(n17983), .B(n18154), .C(n13610), .D(
        n18174), .Y(n13207) );
  sky130_fd_sc_hd__nor2_1 U18460 ( .A(n14111), .B(n13197), .Y(n17963) );
  sky130_fd_sc_hd__nor2_1 U18461 ( .A(n17975), .B(n17963), .Y(n18136) );
  sky130_fd_sc_hd__nand2_1 U18462 ( .A(n17990), .B(n14999), .Y(n13237) );
  sky130_fd_sc_hd__nor2_1 U18463 ( .A(n18043), .B(n18034), .Y(n18029) );
  sky130_fd_sc_hd__nand3_1 U18464 ( .A(n13210), .B(n15017), .C(
        j202_soc_core_bootrom_00_address_w[7]), .Y(n13221) );
  sky130_fd_sc_hd__nor2_1 U18465 ( .A(n14988), .B(n13221), .Y(n17968) );
  sky130_fd_sc_hd__nand2_1 U18466 ( .A(n14472), .B(n13255), .Y(n18134) );
  sky130_fd_sc_hd__nor2_1 U18467 ( .A(n17968), .B(n13208), .Y(n13549) );
  sky130_fd_sc_hd__nand2_1 U18468 ( .A(n15016), .B(n14983), .Y(n13201) );
  sky130_fd_sc_hd__nand3_1 U18469 ( .A(n13210), .B(
        j202_soc_core_bootrom_00_address_w[7]), .C(
        j202_soc_core_bootrom_00_address_w[11]), .Y(n13214) );
  sky130_fd_sc_hd__nor2_1 U18470 ( .A(n13201), .B(n13214), .Y(n18092) );
  sky130_fd_sc_hd__nor2_1 U18471 ( .A(n18045), .B(n18092), .Y(n18181) );
  sky130_fd_sc_hd__nand2_1 U18472 ( .A(n13549), .B(n18181), .Y(n18099) );
  sky130_fd_sc_hd__nor2_1 U18473 ( .A(n13218), .B(n18099), .Y(n17959) );
  sky130_fd_sc_hd__nor2_1 U18474 ( .A(n13210), .B(n13212), .Y(n17984) );
  sky130_fd_sc_hd__nor2_1 U18475 ( .A(j202_soc_core_bootrom_00_address_w[11]), 
        .B(n14101), .Y(n14977) );
  sky130_fd_sc_hd__nand3_1 U18476 ( .A(n14977), .B(
        j202_soc_core_bootrom_00_address_w[10]), .C(n13210), .Y(n13583) );
  sky130_fd_sc_hd__nor2_1 U18477 ( .A(n14999), .B(n13583), .Y(n13567) );
  sky130_fd_sc_hd__nand2_1 U18478 ( .A(n13241), .B(n18180), .Y(n17962) );
  sky130_fd_sc_hd__nor2_1 U18479 ( .A(n17984), .B(n17962), .Y(n13216) );
  sky130_fd_sc_hd__nand2_1 U18480 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .B(j202_soc_core_bootrom_00_address_w[3]), .Y(n18147) );
  sky130_fd_sc_hd__a21oi_1 U18481 ( .A1(n17959), .A2(n13216), .B1(n18147), .Y(
        n13206) );
  sky130_fd_sc_hd__nor2_1 U18482 ( .A(n14099), .B(n13236), .Y(n13215) );
  sky130_fd_sc_hd__nand2_1 U18483 ( .A(n18154), .B(n18102), .Y(n18012) );
  sky130_fd_sc_hd__nand2_1 U18484 ( .A(n13198), .B(
        j202_soc_core_bootrom_00_address_w[10]), .Y(n13245) );
  sky130_fd_sc_hd__nor2b_1 U18485 ( .B_N(n13199), .A(n13200), .Y(n18100) );
  sky130_fd_sc_hd__nand2_1 U18486 ( .A(n13253), .B(n18133), .Y(n18117) );
  sky130_fd_sc_hd__nor2_1 U18487 ( .A(n17991), .B(n18117), .Y(n18170) );
  sky130_fd_sc_hd__nor4_1 U18489 ( .A(n17975), .B(n18101), .C(n18012), .D(
        n18017), .Y(n13204) );
  sky130_fd_sc_hd__nor2_1 U18490 ( .A(j202_soc_core_bootrom_00_address_w[3]), 
        .B(j202_soc_core_bootrom_00_address_w[5]), .Y(n18189) );
  sky130_fd_sc_hd__nor3_1 U18491 ( .A(n17991), .B(n18045), .C(n13215), .Y(
        n13566) );
  sky130_fd_sc_hd__nand2b_1 U18492 ( .A_N(n13201), .B(n13199), .Y(n18173) );
  sky130_fd_sc_hd__nor3_1 U18493 ( .A(n13608), .B(n18040), .C(n13567), .Y(
        n18135) );
  sky130_fd_sc_hd__nor2_1 U18494 ( .A(n13200), .B(n13596), .Y(n18091) );
  sky130_fd_sc_hd__nor2_1 U18495 ( .A(n13210), .B(n18125), .Y(n13256) );
  sky130_fd_sc_hd__nor2_1 U18496 ( .A(n13201), .B(n13596), .Y(n17960) );
  sky130_fd_sc_hd__nor2_1 U18497 ( .A(n13256), .B(n17960), .Y(n17972) );
  sky130_fd_sc_hd__nand2_1 U18498 ( .A(n18081), .B(n17972), .Y(n13584) );
  sky130_fd_sc_hd__nand2_1 U18499 ( .A(n14983), .B(
        j202_soc_core_bootrom_00_address_w[9]), .Y(n13202) );
  sky130_fd_sc_hd__nor2_1 U18500 ( .A(n13202), .B(n15009), .Y(n18010) );
  sky130_fd_sc_hd__nand2_1 U18501 ( .A(n18010), .B(
        j202_soc_core_bootrom_00_address_w[7]), .Y(n18168) );
  sky130_fd_sc_hd__nand2_1 U18502 ( .A(n13224), .B(n18168), .Y(n13601) );
  sky130_fd_sc_hd__nor4b_1 U18503 ( .D_N(n13566), .A(n13220), .B(n13584), .C(
        n13601), .Y(n13203) );
  sky130_fd_sc_hd__nor2_1 U18504 ( .A(j202_soc_core_bootrom_00_address_w[3]), 
        .B(n14094), .Y(n18155) );
  sky130_fd_sc_hd__o22ai_1 U18505 ( .A1(n13204), .A2(n18047), .B1(n13203), 
        .B2(n18172), .Y(n13205) );
  sky130_fd_sc_hd__a211oi_1 U18506 ( .A1(n18161), .A2(n13207), .B1(n13206), 
        .C1(n13205), .Y(n13233) );
  sky130_fd_sc_hd__nand2_1 U18507 ( .A(n13231), .B(n14998), .Y(n18139) );
  sky130_fd_sc_hd__nor2_1 U18508 ( .A(n13553), .B(n13208), .Y(n17981) );
  sky130_fd_sc_hd__nand2_1 U18509 ( .A(n18006), .B(n14999), .Y(n13257) );
  sky130_fd_sc_hd__nand2_1 U18510 ( .A(n13223), .B(n13257), .Y(n17996) );
  sky130_fd_sc_hd__nor2_1 U18511 ( .A(n18101), .B(n17996), .Y(n18182) );
  sky130_fd_sc_hd__nand2_1 U18512 ( .A(n18182), .B(n13234), .Y(n17956) );
  sky130_fd_sc_hd__nor4_1 U18513 ( .A(n18044), .B(n18092), .C(n13554), .D(
        n17956), .Y(n13209) );
  sky130_fd_sc_hd__a31oi_1 U18514 ( .A1(n17981), .A2(n13209), .A3(n13237), 
        .B1(n18183), .Y(n13230) );
  sky130_fd_sc_hd__nor2_1 U18515 ( .A(n13210), .B(n14777), .Y(n13568) );
  sky130_fd_sc_hd__nor2_1 U18516 ( .A(n13568), .B(n13256), .Y(n13600) );
  sky130_fd_sc_hd__nor2_1 U18517 ( .A(n17984), .B(n18100), .Y(n13605) );
  sky130_fd_sc_hd__nand2_1 U18518 ( .A(n13605), .B(n13257), .Y(n13557) );
  sky130_fd_sc_hd__nand2_1 U18519 ( .A(n13234), .B(n13587), .Y(n13569) );
  sky130_fd_sc_hd__nor4_1 U18520 ( .A(n17975), .B(n17990), .C(n13557), .D(
        n13569), .Y(n13211) );
  sky130_fd_sc_hd__a31oi_1 U18521 ( .A1(n13549), .A2(n13600), .A3(n13211), 
        .B1(n18172), .Y(n13229) );
  sky130_fd_sc_hd__nand2_1 U18522 ( .A(n13235), .B(n13240), .Y(n13219) );
  sky130_fd_sc_hd__nor2_1 U18523 ( .A(n14111), .B(n13236), .Y(n13586) );
  sky130_fd_sc_hd__nand2_1 U18524 ( .A(n17958), .B(n13253), .Y(n13611) );
  sky130_fd_sc_hd__nor2_1 U18525 ( .A(j202_soc_core_bootrom_00_address_w[9]), 
        .B(n13212), .Y(n17997) );
  sky130_fd_sc_hd__nand2_1 U18526 ( .A(n18118), .B(n18032), .Y(n18112) );
  sky130_fd_sc_hd__nor2_1 U18527 ( .A(n13221), .B(n13245), .Y(n18005) );
  sky130_fd_sc_hd__nor2_1 U18528 ( .A(n17960), .B(n18005), .Y(n18104) );
  sky130_fd_sc_hd__nor2_1 U18529 ( .A(n18040), .B(n13215), .Y(n18093) );
  sky130_fd_sc_hd__nand4_1 U18530 ( .A(n18143), .B(n18104), .C(n13216), .D(
        n18093), .Y(n13217) );
  sky130_fd_sc_hd__nor4_1 U18531 ( .A(n13219), .B(n13218), .C(n13611), .D(
        n13217), .Y(n13227) );
  sky130_fd_sc_hd__nor2_1 U18532 ( .A(n13553), .B(n13220), .Y(n18145) );
  sky130_fd_sc_hd__nor2_1 U18533 ( .A(n13222), .B(n13221), .Y(n13607) );
  sky130_fd_sc_hd__nor2_1 U18534 ( .A(n17968), .B(n18005), .Y(n18037) );
  sky130_fd_sc_hd__nor2_1 U18535 ( .A(n13607), .B(n13247), .Y(n13239) );
  sky130_fd_sc_hd__nand3_1 U18536 ( .A(n18145), .B(n13239), .C(n13223), .Y(
        n18131) );
  sky130_fd_sc_hd__nor2_1 U18537 ( .A(n17984), .B(n18026), .Y(n13571) );
  sky130_fd_sc_hd__nand2_1 U18538 ( .A(n13571), .B(n13224), .Y(n17957) );
  sky130_fd_sc_hd__nor2_1 U18539 ( .A(n13568), .B(n18041), .Y(n18185) );
  sky130_fd_sc_hd__nand2_1 U18540 ( .A(n18185), .B(n18134), .Y(n17989) );
  sky130_fd_sc_hd__nand2_1 U18541 ( .A(n18032), .B(n18180), .Y(n13225) );
  sky130_fd_sc_hd__nor4_1 U18542 ( .A(n18131), .B(n17957), .C(n17989), .D(
        n13225), .Y(n13226) );
  sky130_fd_sc_hd__o22ai_1 U18543 ( .A1(n13227), .A2(n18147), .B1(n13226), 
        .B2(n18047), .Y(n13228) );
  sky130_fd_sc_hd__nor3_1 U18544 ( .A(n13230), .B(n13229), .C(n13228), .Y(
        n13232) );
  sky130_fd_sc_hd__nand2_1 U18545 ( .A(n13231), .B(
        j202_soc_core_bootrom_00_address_w[6]), .Y(n18164) );
  sky130_fd_sc_hd__o22ai_1 U18546 ( .A1(n13233), .A2(n18139), .B1(n13232), 
        .B2(n18164), .Y(n13267) );
  sky130_fd_sc_hd__nor2_1 U18548 ( .A(n17969), .B(n18113), .Y(n17961) );
  sky130_fd_sc_hd__nand2_1 U18549 ( .A(n13257), .B(n18102), .Y(n13578) );
  sky130_fd_sc_hd__nor2_1 U18550 ( .A(n17960), .B(n13578), .Y(n17993) );
  sky130_fd_sc_hd__nand2_1 U18551 ( .A(n17993), .B(n13237), .Y(n18009) );
  sky130_fd_sc_hd__nor3_1 U18552 ( .A(n18031), .B(n18026), .C(n18009), .Y(
        n13238) );
  sky130_fd_sc_hd__a31oi_1 U18553 ( .A1(n13239), .A2(n17961), .A3(n13238), 
        .B1(n18047), .Y(n13252) );
  sky130_fd_sc_hd__nor2_1 U18554 ( .A(n13568), .B(n17990), .Y(n18095) );
  sky130_fd_sc_hd__nand2_1 U18555 ( .A(n13240), .B(n18102), .Y(n13243) );
  sky130_fd_sc_hd__nand2b_1 U18556 ( .A_N(n13243), .B(n18136), .Y(n17995) );
  sky130_fd_sc_hd__nor2b_1 U18557 ( .B_N(n18095), .A(n17995), .Y(n18169) );
  sky130_fd_sc_hd__nand3_1 U18558 ( .A(n13241), .B(n18032), .C(n18180), .Y(
        n13254) );
  sky130_fd_sc_hd__a31oi_1 U18559 ( .A1(n18169), .A2(n18003), .A3(n13242), 
        .B1(n18147), .Y(n13251) );
  sky130_fd_sc_hd__nand2_1 U18560 ( .A(n18143), .B(n13555), .Y(n13550) );
  sky130_fd_sc_hd__nor4_1 U18561 ( .A(n13585), .B(n13243), .C(n18130), .D(
        n13550), .Y(n13244) );
  sky130_fd_sc_hd__a31oi_1 U18562 ( .A1(n18037), .A2(n13244), .A3(n18086), 
        .B1(n18183), .Y(n13250) );
  sky130_fd_sc_hd__nor2_1 U18563 ( .A(n13246), .B(n13245), .Y(n18004) );
  sky130_fd_sc_hd__nor2_1 U18564 ( .A(n13608), .B(n18034), .Y(n18121) );
  sky130_fd_sc_hd__nand2_1 U18565 ( .A(n18115), .B(n18121), .Y(n18030) );
  sky130_fd_sc_hd__nor4_1 U18566 ( .A(n13568), .B(n18004), .C(n13247), .D(
        n18030), .Y(n13248) );
  sky130_fd_sc_hd__nand2_1 U18567 ( .A(n18124), .B(n14099), .Y(n18158) );
  sky130_fd_sc_hd__a21oi_1 U18568 ( .A1(n13248), .A2(n18158), .B1(n18172), .Y(
        n13249) );
  sky130_fd_sc_hd__nor4_1 U18569 ( .A(n13252), .B(n13251), .C(n13250), .D(
        n13249), .Y(n13265) );
  sky130_fd_sc_hd__nand2_1 U18570 ( .A(n14998), .B(
        j202_soc_core_bootrom_00_address_w[8]), .Y(n18107) );
  sky130_fd_sc_hd__nor2_1 U18571 ( .A(n18044), .B(n18010), .Y(n17992) );
  sky130_fd_sc_hd__nand4_1 U18572 ( .A(n17992), .B(n18104), .C(n18158), .D(
        n18007), .Y(n13263) );
  sky130_fd_sc_hd__nand2_1 U18573 ( .A(n18179), .B(n13253), .Y(n13602) );
  sky130_fd_sc_hd__nor2_1 U18574 ( .A(n18039), .B(n13602), .Y(n18033) );
  sky130_fd_sc_hd__nor3_1 U18575 ( .A(n18034), .B(n18123), .C(n18112), .Y(
        n13564) );
  sky130_fd_sc_hd__a31oi_1 U18576 ( .A1(n18033), .A2(n17992), .A3(n13564), 
        .B1(n18147), .Y(n13262) );
  sky130_fd_sc_hd__nor2_1 U18577 ( .A(n17997), .B(n17963), .Y(n17982) );
  sky130_fd_sc_hd__nand3_1 U18578 ( .A(n17982), .B(n13253), .C(n18081), .Y(
        n18084) );
  sky130_fd_sc_hd__nor4_1 U18579 ( .A(n13568), .B(n13553), .C(n13254), .D(
        n18084), .Y(n13260) );
  sky130_fd_sc_hd__nor2_1 U18580 ( .A(n13256), .B(n13255), .Y(n17985) );
  sky130_fd_sc_hd__nand2_1 U18581 ( .A(n14977), .B(n14098), .Y(n17970) );
  sky130_fd_sc_hd__nand4_1 U18582 ( .A(n17985), .B(n17970), .C(n13555), .D(
        n13257), .Y(n13258) );
  sky130_fd_sc_hd__a211oi_1 U18585 ( .A1(n18155), .A2(n13263), .B1(n13262), 
        .C1(n13261), .Y(n13264) );
  sky130_fd_sc_hd__nand2_1 U18586 ( .A(j202_soc_core_bootrom_00_address_w[8]), 
        .B(j202_soc_core_bootrom_00_address_w[6]), .Y(n18190) );
  sky130_fd_sc_hd__o22ai_1 U18587 ( .A1(n13265), .A2(n18107), .B1(n13264), 
        .B2(n18190), .Y(n13266) );
  sky130_fd_sc_hd__nor2_1 U18588 ( .A(n13267), .B(n13266), .Y(n13288) );
  sky130_fd_sc_hd__a22oi_1 U18589 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[275]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[51]), .Y(n13281) );
  sky130_fd_sc_hd__a22o_1 U18590 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[307]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[339]), .X(n13268) );
  sky130_fd_sc_hd__a21oi_1 U18591 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[371]), .B1(n13268), .Y(n13280) );
  sky130_fd_sc_hd__nand2_1 U18592 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[243]), .Y(n13272) );
  sky130_fd_sc_hd__a21oi_1 U18593 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[467]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n13271) );
  sky130_fd_sc_hd__nand2_1 U18594 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[403]), .Y(n13270) );
  sky130_fd_sc_hd__nand2_1 U18595 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[435]), .Y(n13269) );
  sky130_fd_sc_hd__nand4_1 U18596 ( .A(n13272), .B(n13271), .C(n13270), .D(
        n13269), .Y(n13273) );
  sky130_fd_sc_hd__a21oi_1 U18597 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[211]), .B1(n13273), .Y(n13279) );
  sky130_fd_sc_hd__a22o_1 U18598 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[19]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[83]), .X(n13274) );
  sky130_fd_sc_hd__a21oi_1 U18599 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[115]), .B1(n13274), .Y(n13276) );
  sky130_fd_sc_hd__a22oi_1 U18600 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[179]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[147]), .Y(n13275) );
  sky130_fd_sc_hd__nand2_1 U18601 ( .A(n13276), .B(n13275), .Y(n13277) );
  sky130_fd_sc_hd__nand2_1 U18602 ( .A(n13277), .B(n17639), .Y(n13278) );
  sky130_fd_sc_hd__nand4_1 U18603 ( .A(n13281), .B(n13280), .C(n13279), .D(
        n13278), .Y(n13282) );
  sky130_fd_sc_hd__o211ai_1 U18604 ( .A1(j202_soc_core_memory0_ram_dout0[499]), 
        .A2(n18758), .B1(n14906), .C1(n13282), .Y(n13286) );
  sky130_fd_sc_hd__a22oi_1 U18605 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[83]), .B1(n18379), .B2(
        j202_soc_core_uart_div1[3]), .Y(n13285) );
  sky130_fd_sc_hd__a22oi_1 U18606 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[19]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[51]), .Y(n13284) );
  sky130_fd_sc_hd__nand2_1 U18607 ( .A(n18629), .B(
        j202_soc_core_bldc_core_00_pwm_duty[7]), .Y(n13283) );
  sky130_fd_sc_hd__nand4_1 U18608 ( .A(n13286), .B(n13285), .C(n13284), .D(
        n13283), .Y(n13287) );
  sky130_fd_sc_hd__o21ba_2 U18609 ( .A1(n18212), .A2(n13288), .B1_N(n13287), 
        .X(n20778) );
  sky130_fd_sc_hd__a22oi_1 U18610 ( .A1(n19657), .A2(n21963), .B1(n19736), 
        .B2(n23307), .Y(n13289) );
  sky130_fd_sc_hd__a21oi_1 U18612 ( .A1(n21758), .A2(n19661), .B1(n13290), .Y(
        n13291) );
  sky130_fd_sc_hd__nand2_1 U18613 ( .A(n13292), .B(n13291), .Y(n25252) );
  sky130_fd_sc_hd__nand2_1 U18614 ( .A(n13295), .B(n13294), .Y(n13296) );
  sky130_fd_sc_hd__xor2_1 U18615 ( .A(n13297), .B(n13296), .X(n21877) );
  sky130_fd_sc_hd__nand2_1 U18616 ( .A(n21877), .B(n19729), .Y(n13394) );
  sky130_fd_sc_hd__ha_1 U18617 ( .A(j202_soc_core_j22_cpu_pc[22]), .B(n13298), 
        .COUT(n13105), .SUM(n21880) );
  sky130_fd_sc_hd__nand2b_1 U18618 ( .A_N(n13299), .B(n13329), .Y(n13462) );
  sky130_fd_sc_hd__nor2_1 U18619 ( .A(n13300), .B(n13462), .Y(n13302) );
  sky130_fd_sc_hd__a21oi_1 U18620 ( .A1(n13302), .A2(n13301), .B1(n17468), .Y(
        n13304) );
  sky130_fd_sc_hd__nor3_1 U18621 ( .A(n13305), .B(n13304), .C(n13303), .Y(
        n13306) );
  sky130_fd_sc_hd__nand2b_1 U18622 ( .A_N(n13306), .B(n17609), .Y(n13389) );
  sky130_fd_sc_hd__nor2_1 U18623 ( .A(n13452), .B(n13453), .Y(n13310) );
  sky130_fd_sc_hd__nor2_1 U18624 ( .A(n13309), .B(n13308), .Y(n13495) );
  sky130_fd_sc_hd__a31oi_1 U18625 ( .A1(n13310), .A2(n13441), .A3(n13495), 
        .B1(n17468), .Y(n13322) );
  sky130_fd_sc_hd__a21oi_1 U18626 ( .A1(n13488), .A2(n13311), .B1(n13500), .Y(
        n13321) );
  sky130_fd_sc_hd__nand2_1 U18627 ( .A(n13312), .B(n13492), .Y(n13430) );
  sky130_fd_sc_hd__nor3_1 U18628 ( .A(n13314), .B(n13430), .C(n13313), .Y(
        n13319) );
  sky130_fd_sc_hd__nor4_1 U18629 ( .A(n13463), .B(n13317), .C(n13316), .D(
        n13315), .Y(n13318) );
  sky130_fd_sc_hd__o22ai_1 U18630 ( .A1(n13319), .A2(n13464), .B1(n13318), 
        .B2(n17730), .Y(n13320) );
  sky130_fd_sc_hd__nor4_1 U18631 ( .A(n13323), .B(n13322), .C(n13321), .D(
        n13320), .Y(n13363) );
  sky130_fd_sc_hd__nor3_1 U18632 ( .A(n13325), .B(n13435), .C(n13324), .Y(
        n13327) );
  sky130_fd_sc_hd__a31oi_1 U18633 ( .A1(n13327), .A2(n17988), .A3(n13326), 
        .B1(n17730), .Y(n13340) );
  sky130_fd_sc_hd__nor3_1 U18634 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .B(j202_soc_core_bootrom_00_address_w[2]), .C(n14120), .Y(n13450) );
  sky130_fd_sc_hd__nor2_1 U18635 ( .A(n13328), .B(n13450), .Y(n13379) );
  sky130_fd_sc_hd__a31oi_1 U18636 ( .A1(n13379), .A2(n13480), .A3(n13329), 
        .B1(n13464), .Y(n13339) );
  sky130_fd_sc_hd__nor2_1 U18637 ( .A(n13330), .B(n14683), .Y(n13482) );
  sky130_fd_sc_hd__a31oi_1 U18638 ( .A1(n13331), .A2(n13369), .A3(n13482), 
        .B1(n13500), .Y(n13338) );
  sky130_fd_sc_hd__nor4_1 U18639 ( .A(n13334), .B(n13333), .C(n13433), .D(
        n13332), .Y(n13335) );
  sky130_fd_sc_hd__a21oi_1 U18640 ( .A1(n13336), .A2(n13335), .B1(n17468), .Y(
        n13337) );
  sky130_fd_sc_hd__nor4_1 U18641 ( .A(n13340), .B(n13339), .C(n13338), .D(
        n13337), .Y(n13361) );
  sky130_fd_sc_hd__a22oi_1 U18642 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[22]), .B1(n18379), .B2(
        j202_soc_core_uart_div1[6]), .Y(n13342) );
  sky130_fd_sc_hd__a22oi_1 U18643 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[86]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[54]), .Y(n13341) );
  sky130_fd_sc_hd__nand2_1 U18644 ( .A(n13342), .B(n13341), .Y(n13343) );
  sky130_fd_sc_hd__a21oi_1 U18645 ( .A1(n18629), .A2(
        j202_soc_core_bldc_core_00_pwm_duty[10]), .B1(n13343), .Y(n13360) );
  sky130_fd_sc_hd__a22oi_1 U18646 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[246]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[214]), .Y(n13347) );
  sky130_fd_sc_hd__a22oi_1 U18647 ( .A1(n18734), .A2(
        j202_soc_core_memory0_ram_dout0[150]), .B1(n18733), .B2(
        j202_soc_core_memory0_ram_dout0[118]), .Y(n13346) );
  sky130_fd_sc_hd__a22oi_1 U18648 ( .A1(n18361), .A2(
        j202_soc_core_memory0_ram_dout0[54]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[86]), .Y(n13345) );
  sky130_fd_sc_hd__nand2_1 U18649 ( .A(n18735), .B(
        j202_soc_core_memory0_ram_dout0[182]), .Y(n13344) );
  sky130_fd_sc_hd__nand4_1 U18650 ( .A(n13347), .B(n13346), .C(n13345), .D(
        n13344), .Y(n13348) );
  sky130_fd_sc_hd__a21oi_1 U18651 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[22]), .B1(n13348), .Y(n13349) );
  sky130_fd_sc_hd__nand2b_1 U18652 ( .A_N(n13349), .B(n17639), .Y(n13357) );
  sky130_fd_sc_hd__a22oi_1 U18653 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[310]), .B1(n18062), .B2(
        j202_soc_core_memory0_ram_dout0[278]), .Y(n13356) );
  sky130_fd_sc_hd__nand2_1 U18654 ( .A(n18743), .B(
        j202_soc_core_memory0_ram_dout0[374]), .Y(n13353) );
  sky130_fd_sc_hd__a21oi_1 U18655 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[470]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n13352) );
  sky130_fd_sc_hd__nand2_1 U18656 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[406]), .Y(n13351) );
  sky130_fd_sc_hd__nand2_1 U18657 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[438]), .Y(n13350) );
  sky130_fd_sc_hd__nand4_1 U18658 ( .A(n13353), .B(n13352), .C(n13351), .D(
        n13350), .Y(n13354) );
  sky130_fd_sc_hd__a21oi_1 U18659 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[342]), .B1(n13354), .Y(n13355) );
  sky130_fd_sc_hd__nand3_1 U18660 ( .A(n13357), .B(n13356), .C(n13355), .Y(
        n13358) );
  sky130_fd_sc_hd__o211ai_1 U18661 ( .A1(j202_soc_core_memory0_ram_dout0[502]), 
        .A2(n18758), .B1(n14906), .C1(n13358), .Y(n13359) );
  sky130_fd_sc_hd__o211a_2 U18662 ( .A1(n18552), .A2(n13361), .B1(n13360), 
        .C1(n13359), .X(n13362) );
  sky130_fd_sc_hd__o21a_1 U18663 ( .A1(n18666), .A2(n13363), .B1(n13362), .X(
        n13388) );
  sky130_fd_sc_hd__nor2_1 U18664 ( .A(n13411), .B(n13364), .Y(n13467) );
  sky130_fd_sc_hd__nand2_1 U18665 ( .A(n13366), .B(n13365), .Y(n13490) );
  sky130_fd_sc_hd__nor3_1 U18666 ( .A(n13416), .B(n13490), .C(n13367), .Y(
        n13368) );
  sky130_fd_sc_hd__a31oi_1 U18667 ( .A1(n13369), .A2(n13467), .A3(n13368), 
        .B1(n17468), .Y(n13385) );
  sky130_fd_sc_hd__nor4_1 U18668 ( .A(n13372), .B(n13371), .C(n13462), .D(
        n13370), .Y(n13377) );
  sky130_fd_sc_hd__nand2_1 U18669 ( .A(n13375), .B(n13374), .Y(n13376) );
  sky130_fd_sc_hd__a31oi_1 U18670 ( .A1(n13377), .A2(n13487), .A3(n13376), 
        .B1(n17730), .Y(n13384) );
  sky130_fd_sc_hd__nor3b_1 U18671 ( .C_N(n13379), .A(n13411), .B(n13378), .Y(
        n13501) );
  sky130_fd_sc_hd__nor2_1 U18672 ( .A(n16741), .B(n18295), .Y(n18268) );
  sky130_fd_sc_hd__nand2_1 U18673 ( .A(n13380), .B(n13493), .Y(n13470) );
  sky130_fd_sc_hd__nor4_1 U18674 ( .A(n18268), .B(n13421), .C(n13470), .D(
        n13381), .Y(n13382) );
  sky130_fd_sc_hd__o22ai_1 U18675 ( .A1(n13501), .A2(n13500), .B1(n13382), 
        .B2(n13464), .Y(n13383) );
  sky130_fd_sc_hd__nor3_1 U18676 ( .A(n13385), .B(n13384), .C(n13383), .Y(
        n13386) );
  sky130_fd_sc_hd__nand2b_1 U18677 ( .A_N(n13386), .B(n18605), .Y(n13387) );
  sky130_fd_sc_hd__nand3_1 U18678 ( .A(n13389), .B(n13388), .C(n13387), .Y(
        n21135) );
  sky130_fd_sc_hd__nand2_1 U18679 ( .A(n21135), .B(n19737), .Y(n13391) );
  sky130_fd_sc_hd__a22oi_1 U18680 ( .A1(n19657), .A2(n21867), .B1(n19736), 
        .B2(n23316), .Y(n13390) );
  sky130_fd_sc_hd__nand2_1 U18681 ( .A(n13391), .B(n13390), .Y(n13392) );
  sky130_fd_sc_hd__a21oi_1 U18682 ( .A1(n21880), .A2(n19661), .B1(n13392), .Y(
        n13393) );
  sky130_fd_sc_hd__nand2_1 U18683 ( .A(n13394), .B(n13393), .Y(n25277) );
  sky130_fd_sc_hd__nand2_1 U18684 ( .A(n11188), .B(n13395), .Y(n13397) );
  sky130_fd_sc_hd__xnor2_1 U18685 ( .A(n13397), .B(n13396), .Y(n21974) );
  sky130_fd_sc_hd__nand2_1 U18686 ( .A(n21974), .B(n19729), .Y(n13402) );
  sky130_fd_sc_hd__ha_1 U18687 ( .A(j202_soc_core_j22_cpu_pc[21]), .B(n13398), 
        .COUT(n13298), .SUM(n21976) );
  sky130_fd_sc_hd__a22oi_1 U18688 ( .A1(n19657), .A2(n22578), .B1(n19736), 
        .B2(n23313), .Y(n13399) );
  sky130_fd_sc_hd__a21oi_1 U18690 ( .A1(n21976), .A2(n19661), .B1(n13400), .Y(
        n13401) );
  sky130_fd_sc_hd__nand2_1 U18691 ( .A(n13402), .B(n13401), .Y(n25281) );
  sky130_fd_sc_hd__nand2_1 U18692 ( .A(n13405), .B(n13404), .Y(n13406) );
  sky130_fd_sc_hd__xor2_1 U18693 ( .A(n13407), .B(n13406), .X(n22020) );
  sky130_fd_sc_hd__nand2_1 U18694 ( .A(n22020), .B(n19729), .Y(n13536) );
  sky130_fd_sc_hd__ha_1 U18695 ( .A(j202_soc_core_j22_cpu_pc[20]), .B(n13408), 
        .COUT(n13398), .SUM(n22022) );
  sky130_fd_sc_hd__nor4_1 U18696 ( .A(n13422), .B(n13439), .C(n13432), .D(
        n13458), .Y(n13409) );
  sky130_fd_sc_hd__a21oi_1 U18697 ( .A1(n13410), .A2(n13409), .B1(n13464), .Y(
        n13428) );
  sky130_fd_sc_hd__a21oi_1 U18698 ( .A1(n13413), .A2(n13412), .B1(n13411), .Y(
        n13414) );
  sky130_fd_sc_hd__a31oi_1 U18699 ( .A1(n13461), .A2(n13415), .A3(n13414), 
        .B1(n17730), .Y(n13427) );
  sky130_fd_sc_hd__nor2_1 U18700 ( .A(n13416), .B(n13439), .Y(n13419) );
  sky130_fd_sc_hd__a31oi_1 U18701 ( .A1(n13419), .A2(n13418), .A3(n13417), 
        .B1(n17468), .Y(n13426) );
  sky130_fd_sc_hd__nor4_1 U18702 ( .A(n14680), .B(n13422), .C(n13421), .D(
        n13420), .Y(n13423) );
  sky130_fd_sc_hd__a21oi_1 U18703 ( .A1(n13424), .A2(n13423), .B1(n13500), .Y(
        n13425) );
  sky130_fd_sc_hd__nor4_1 U18704 ( .A(n13428), .B(n13427), .C(n13426), .D(
        n13425), .Y(n13429) );
  sky130_fd_sc_hd__nand2b_1 U18705 ( .A_N(n13429), .B(n17609), .Y(n13531) );
  sky130_fd_sc_hd__nor4_1 U18706 ( .A(n13589), .B(n13431), .C(n13462), .D(
        n13430), .Y(n13471) );
  sky130_fd_sc_hd__a31oi_1 U18707 ( .A1(n13471), .A2(n14777), .A3(n13480), 
        .B1(n13464), .Y(n13446) );
  sky130_fd_sc_hd__nor3_1 U18708 ( .A(n13435), .B(n13434), .C(n13433), .Y(
        n13437) );
  sky130_fd_sc_hd__a31oi_1 U18709 ( .A1(n13438), .A2(n13437), .A3(n13436), 
        .B1(n13500), .Y(n13445) );
  sky130_fd_sc_hd__nor4b_1 U18710 ( .D_N(n13441), .A(n13551), .B(n13440), .C(
        n13439), .Y(n13443) );
  sky130_fd_sc_hd__nor3_1 U18711 ( .A(n13452), .B(n13453), .C(n13450), .Y(
        n13442) );
  sky130_fd_sc_hd__o22ai_1 U18712 ( .A1(n13443), .A2(n17730), .B1(n13442), 
        .B2(n17468), .Y(n13444) );
  sky130_fd_sc_hd__nor3_1 U18713 ( .A(n13446), .B(n13445), .C(n13444), .Y(
        n13447) );
  sky130_fd_sc_hd__nand2b_1 U18714 ( .A_N(n13447), .B(n18610), .Y(n13530) );
  sky130_fd_sc_hd__nor2_1 U18715 ( .A(n13449), .B(n13448), .Y(n13451) );
  sky130_fd_sc_hd__nor4_1 U18716 ( .A(n13453), .B(n13452), .C(n13451), .D(
        n13450), .Y(n13455) );
  sky130_fd_sc_hd__a31oi_1 U18717 ( .A1(n13456), .A2(n13455), .A3(n13454), 
        .B1(n13500), .Y(n13478) );
  sky130_fd_sc_hd__nor2_1 U18718 ( .A(n13458), .B(n13457), .Y(n13459) );
  sky130_fd_sc_hd__a31oi_1 U18719 ( .A1(n13461), .A2(n13460), .A3(n13459), 
        .B1(n17730), .Y(n13477) );
  sky130_fd_sc_hd__nor2_1 U18720 ( .A(n13463), .B(n13462), .Y(n13466) );
  sky130_fd_sc_hd__a31oi_1 U18721 ( .A1(n13467), .A2(n13466), .A3(n13465), 
        .B1(n13464), .Y(n13476) );
  sky130_fd_sc_hd__nor4b_1 U18722 ( .D_N(n13471), .A(n13470), .B(n13469), .C(
        n13468), .Y(n13473) );
  sky130_fd_sc_hd__a31oi_1 U18723 ( .A1(n13474), .A2(n13473), .A3(n13472), 
        .B1(n17468), .Y(n13475) );
  sky130_fd_sc_hd__nor4_1 U18724 ( .A(n13478), .B(n13477), .C(n13476), .D(
        n13475), .Y(n13479) );
  sky130_fd_sc_hd__nand2b_1 U18725 ( .A_N(n13479), .B(n18798), .Y(n13529) );
  sky130_fd_sc_hd__nand4_1 U18726 ( .A(n13482), .B(n13481), .C(n13480), .D(
        n13493), .Y(n13484) );
  sky130_fd_sc_hd__nand2_1 U18728 ( .A(n14098), .B(n15017), .Y(n14097) );
  sky130_fd_sc_hd__nor2_1 U18729 ( .A(n14099), .B(n14097), .Y(n14447) );
  sky130_fd_sc_hd__nand4_1 U18730 ( .A(n13488), .B(n13487), .C(n13486), .D(
        n14828), .Y(n13491) );
  sky130_fd_sc_hd__nand4_1 U18732 ( .A(n13495), .B(n13494), .C(n13493), .D(
        n13492), .Y(n13497) );
  sky130_fd_sc_hd__nand2_1 U18733 ( .A(n13497), .B(n13496), .Y(n13498) );
  sky130_fd_sc_hd__nand2_1 U18734 ( .A(n13499), .B(n13498), .Y(n13504) );
  sky130_fd_sc_hd__a31oi_1 U18735 ( .A1(n13502), .A2(n13501), .A3(n14828), 
        .B1(n13500), .Y(n13503) );
  sky130_fd_sc_hd__nor2_1 U18736 ( .A(n13504), .B(n13503), .Y(n13505) );
  sky130_fd_sc_hd__nand2_1 U18737 ( .A(n13506), .B(n13505), .Y(n13527) );
  sky130_fd_sc_hd__a22oi_1 U18738 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[276]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[52]), .Y(n13520) );
  sky130_fd_sc_hd__a22o_1 U18739 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[308]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[340]), .X(n13507) );
  sky130_fd_sc_hd__a21oi_1 U18740 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[372]), .B1(n13507), .Y(n13519) );
  sky130_fd_sc_hd__nand2_1 U18741 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[244]), .Y(n13511) );
  sky130_fd_sc_hd__a21oi_1 U18742 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[468]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n13510) );
  sky130_fd_sc_hd__nand2_1 U18743 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[404]), .Y(n13509) );
  sky130_fd_sc_hd__nand2_1 U18744 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[436]), .Y(n13508) );
  sky130_fd_sc_hd__nand4_1 U18745 ( .A(n13511), .B(n13510), .C(n13509), .D(
        n13508), .Y(n13512) );
  sky130_fd_sc_hd__a21oi_1 U18746 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[212]), .B1(n13512), .Y(n13518) );
  sky130_fd_sc_hd__a22o_1 U18747 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[20]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[84]), .X(n13513) );
  sky130_fd_sc_hd__a21oi_1 U18748 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[116]), .B1(n13513), .Y(n13515) );
  sky130_fd_sc_hd__a22oi_1 U18749 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[180]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[148]), .Y(n13514) );
  sky130_fd_sc_hd__nand2_1 U18750 ( .A(n13515), .B(n13514), .Y(n13516) );
  sky130_fd_sc_hd__nand2_1 U18751 ( .A(n13516), .B(n17639), .Y(n13517) );
  sky130_fd_sc_hd__nand4_1 U18752 ( .A(n13520), .B(n13519), .C(n13518), .D(
        n13517), .Y(n13521) );
  sky130_fd_sc_hd__o211ai_1 U18753 ( .A1(j202_soc_core_memory0_ram_dout0[500]), 
        .A2(n18758), .B1(n14906), .C1(n13521), .Y(n13525) );
  sky130_fd_sc_hd__a22oi_1 U18754 ( .A1(n18726), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[52]), .B1(n18379), .B2(
        j202_soc_core_uart_div1[4]), .Y(n13524) );
  sky130_fd_sc_hd__a22oi_1 U18755 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[20]), .B1(n18727), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[84]), .Y(n13523) );
  sky130_fd_sc_hd__nand2_1 U18756 ( .A(n18629), .B(
        j202_soc_core_bldc_core_00_pwm_duty[8]), .Y(n13522) );
  sky130_fd_sc_hd__nand4_1 U18757 ( .A(n13525), .B(n13524), .C(n13523), .D(
        n13522), .Y(n13526) );
  sky130_fd_sc_hd__a21oi_1 U18758 ( .A1(n13527), .A2(n18605), .B1(n13526), .Y(
        n13528) );
  sky130_fd_sc_hd__nand4_1 U18759 ( .A(n13531), .B(n13530), .C(n13529), .D(
        n13528), .Y(n22540) );
  sky130_fd_sc_hd__nand2_1 U18760 ( .A(n22540), .B(n19737), .Y(n13533) );
  sky130_fd_sc_hd__a22oi_1 U18761 ( .A1(n19657), .A2(n22577), .B1(n19736), 
        .B2(n23310), .Y(n13532) );
  sky130_fd_sc_hd__nand2_1 U18762 ( .A(n13533), .B(n13532), .Y(n13534) );
  sky130_fd_sc_hd__a21oi_1 U18763 ( .A1(n22022), .A2(n19661), .B1(n13534), .Y(
        n13535) );
  sky130_fd_sc_hd__nand2_1 U18764 ( .A(n13536), .B(n13535), .Y(n25250) );
  sky130_fd_sc_hd__nor2_1 U18765 ( .A(n13538), .B(j202_soc_core_j22_cpu_istall), .Y(n20220) );
  sky130_fd_sc_hd__nand2_1 U18767 ( .A(n23239), .B(
        j202_soc_core_j22_cpu_pc_hold), .Y(n22800) );
  sky130_fd_sc_hd__nor3_1 U18768 ( .A(j202_soc_core_j22_cpu_opst[4]), .B(
        n20773), .C(n22417), .Y(n20348) );
  sky130_fd_sc_hd__nor2_1 U18769 ( .A(j202_soc_core_j22_cpu_opst[2]), .B(
        j202_soc_core_j22_cpu_opst[0]), .Y(n21328) );
  sky130_fd_sc_hd__nand3_1 U18770 ( .A(n20773), .B(
        j202_soc_core_j22_cpu_opst[4]), .C(n21328), .Y(n22804) );
  sky130_fd_sc_hd__nand2b_1 U18771 ( .A_N(n24878), .B(n22804), .Y(n22788) );
  sky130_fd_sc_hd__nor2b_1 U18772 ( .B_N(n22788), .A(n21441), .Y(n24897) );
  sky130_fd_sc_hd__nor2_1 U18773 ( .A(n20348), .B(n24897), .Y(n21338) );
  sky130_fd_sc_hd__nor2_1 U18774 ( .A(j202_soc_core_j22_cpu_opst[4]), .B(
        n21441), .Y(n20774) );
  sky130_fd_sc_hd__nand3_1 U18775 ( .A(j202_soc_core_j22_cpu_opst[3]), .B(
        n21604), .C(n20774), .Y(n21408) );
  sky130_fd_sc_hd__nand4b_1 U18776 ( .A_N(n22800), .B(n21338), .C(n21408), .D(
        n22789), .Y(n13539) );
  sky130_fd_sc_hd__nand2_1 U18777 ( .A(n13540), .B(n13539), .Y(n25299) );
  sky130_fd_sc_hd__nand2_1 U18778 ( .A(j202_soc_core_ahbcs_6__HREADY_), .B(
        n25734), .Y(n23250) );
  sky130_fd_sc_hd__nand2_1 U18779 ( .A(n13543), .B(n13542), .Y(n13544) );
  sky130_fd_sc_hd__xor2_1 U18780 ( .A(n13545), .B(n13544), .X(n21786) );
  sky130_fd_sc_hd__nand2_1 U18781 ( .A(n21786), .B(n19729), .Y(n13650) );
  sky130_fd_sc_hd__ha_1 U18782 ( .A(j202_soc_core_j22_cpu_pc[18]), .B(n13546), 
        .COUT(n13191), .SUM(n21789) );
  sky130_fd_sc_hd__nor2b_1 U18783 ( .B_N(n17970), .A(n13547), .Y(n13548) );
  sky130_fd_sc_hd__nor2_1 U18784 ( .A(n17969), .B(n18091), .Y(n18153) );
  sky130_fd_sc_hd__nand4_1 U18785 ( .A(n18182), .B(n13549), .C(n13548), .D(
        n18153), .Y(n13563) );
  sky130_fd_sc_hd__nor4_1 U18786 ( .A(n13568), .B(n13551), .C(n17975), .D(
        n13550), .Y(n18152) );
  sky130_fd_sc_hd__nor4_1 U18787 ( .A(n18124), .B(n17963), .C(n18114), .D(
        n17957), .Y(n13552) );
  sky130_fd_sc_hd__a21oi_1 U18788 ( .A1(n18152), .A2(n13552), .B1(n18183), .Y(
        n13562) );
  sky130_fd_sc_hd__nor2_1 U18789 ( .A(n13554), .B(n13553), .Y(n13580) );
  sky130_fd_sc_hd__nand2_1 U18790 ( .A(n18095), .B(n18118), .Y(n18042) );
  sky130_fd_sc_hd__nand2_1 U18791 ( .A(n18086), .B(n13555), .Y(n13556) );
  sky130_fd_sc_hd__nor4bb_1 U18792 ( .C_N(n13580), .D_N(n13605), .A(n18042), 
        .B(n13556), .Y(n13560) );
  sky130_fd_sc_hd__nand2_1 U18793 ( .A(n18144), .B(n18035), .Y(n18016) );
  sky130_fd_sc_hd__nand2_1 U18794 ( .A(n18037), .B(n18086), .Y(n13558) );
  sky130_fd_sc_hd__nor4_1 U18795 ( .A(n18043), .B(n18016), .C(n13558), .D(
        n13557), .Y(n13559) );
  sky130_fd_sc_hd__o22ai_1 U18796 ( .A1(n13560), .A2(n18047), .B1(n13559), 
        .B2(n18172), .Y(n13561) );
  sky130_fd_sc_hd__a211oi_1 U18797 ( .A1(n18178), .A2(n13563), .B1(n13562), 
        .C1(n13561), .Y(n13577) );
  sky130_fd_sc_hd__nand2_1 U18798 ( .A(n13605), .B(n18086), .Y(n18097) );
  sky130_fd_sc_hd__nor2_1 U18799 ( .A(n18031), .B(n18097), .Y(n13612) );
  sky130_fd_sc_hd__a31oi_1 U18800 ( .A1(n13564), .A2(n13612), .A3(n13583), 
        .B1(n18183), .Y(n13575) );
  sky130_fd_sc_hd__nor2_1 U18801 ( .A(n18031), .B(n13568), .Y(n18083) );
  sky130_fd_sc_hd__nand2_1 U18802 ( .A(n18083), .B(n13571), .Y(n17974) );
  sky130_fd_sc_hd__nor4b_1 U18803 ( .D_N(n18153), .A(n18100), .B(n18005), .C(
        n17974), .Y(n13565) );
  sky130_fd_sc_hd__a31oi_1 U18804 ( .A1(n13565), .A2(n18173), .A3(n13587), 
        .B1(n18172), .Y(n13574) );
  sky130_fd_sc_hd__nand2_1 U18805 ( .A(n13600), .B(n18143), .Y(n18106) );
  sky130_fd_sc_hd__nor2_1 U18806 ( .A(n18026), .B(n18106), .Y(n18149) );
  sky130_fd_sc_hd__a31oi_1 U18807 ( .A1(n18149), .A2(n13566), .A3(n18180), 
        .B1(n18147), .Y(n13573) );
  sky130_fd_sc_hd__nor2_1 U18808 ( .A(n13567), .B(n18091), .Y(n18120) );
  sky130_fd_sc_hd__nor2_1 U18809 ( .A(n13568), .B(n17975), .Y(n18127) );
  sky130_fd_sc_hd__nand3b_1 U18810 ( .A_N(n17960), .B(n18120), .C(n18127), .Y(
        n18111) );
  sky130_fd_sc_hd__nor2_1 U18811 ( .A(n13569), .B(n18111), .Y(n13570) );
  sky130_fd_sc_hd__a31oi_1 U18812 ( .A1(n13571), .A2(n17981), .A3(n13570), 
        .B1(n18047), .Y(n13572) );
  sky130_fd_sc_hd__nor4_1 U18813 ( .A(n13575), .B(n13574), .C(n13573), .D(
        n13572), .Y(n13576) );
  sky130_fd_sc_hd__o22ai_1 U18814 ( .A1(n13577), .A2(n18107), .B1(n13576), 
        .B2(n18190), .Y(n13621) );
  sky130_fd_sc_hd__nor2_1 U18815 ( .A(n18031), .B(n13578), .Y(n18159) );
  sky130_fd_sc_hd__nor4_1 U18816 ( .A(n18041), .B(n13586), .C(n18100), .D(
        n17962), .Y(n13579) );
  sky130_fd_sc_hd__a31oi_1 U18817 ( .A1(n13580), .A2(n18159), .A3(n13579), 
        .B1(n18183), .Y(n13594) );
  sky130_fd_sc_hd__nand2_1 U18818 ( .A(n13581), .B(n18102), .Y(n13603) );
  sky130_fd_sc_hd__nor2_1 U18819 ( .A(n17984), .B(n13603), .Y(n18028) );
  sky130_fd_sc_hd__nor4_1 U18820 ( .A(n18045), .B(n18085), .C(n17996), .D(
        n18084), .Y(n13582) );
  sky130_fd_sc_hd__a31oi_1 U18821 ( .A1(n18028), .A2(n18135), .A3(n13582), 
        .B1(n18172), .Y(n13593) );
  sky130_fd_sc_hd__nand2_1 U18822 ( .A(n18173), .B(n13583), .Y(n18013) );
  sky130_fd_sc_hd__nor4_1 U18823 ( .A(n18101), .B(n18043), .C(n13584), .D(
        n18013), .Y(n13591) );
  sky130_fd_sc_hd__nor2_1 U18824 ( .A(n13586), .B(n13585), .Y(n17998) );
  sky130_fd_sc_hd__nand3_1 U18825 ( .A(n17998), .B(n18093), .C(n13587), .Y(
        n13588) );
  sky130_fd_sc_hd__nor4_1 U18826 ( .A(n13589), .B(n17960), .C(n17974), .D(
        n13588), .Y(n13590) );
  sky130_fd_sc_hd__o22ai_1 U18827 ( .A1(n13591), .A2(n18147), .B1(n13590), 
        .B2(n18047), .Y(n13592) );
  sky130_fd_sc_hd__nor3_1 U18828 ( .A(n13594), .B(n13593), .C(n13592), .Y(
        n13619) );
  sky130_fd_sc_hd__nor4_1 U18829 ( .A(n13595), .B(n18005), .C(n18100), .D(
        n13603), .Y(n13599) );
  sky130_fd_sc_hd__nand2_1 U18830 ( .A(n13598), .B(n13597), .Y(n13609) );
  sky130_fd_sc_hd__a21oi_1 U18831 ( .A1(n13599), .A2(n13609), .B1(n18047), .Y(
        n13617) );
  sky130_fd_sc_hd__nor2_1 U18832 ( .A(n18085), .B(n13607), .Y(n18018) );
  sky130_fd_sc_hd__nor4_1 U18833 ( .A(n18015), .B(n13603), .C(n13602), .D(
        n13601), .Y(n13604) );
  sky130_fd_sc_hd__a31oi_1 U18834 ( .A1(n13605), .A2(n18018), .A3(n13604), 
        .B1(n18147), .Y(n13616) );
  sky130_fd_sc_hd__nand4_1 U18835 ( .A(n18083), .B(n17993), .C(n18118), .D(
        n18133), .Y(n13606) );
  sky130_fd_sc_hd__nor4_1 U18836 ( .A(n13608), .B(n13607), .C(n18113), .D(
        n13606), .Y(n13614) );
  sky130_fd_sc_hd__nand3b_1 U18837 ( .A_N(n17996), .B(n13610), .C(n13609), .Y(
        n18014) );
  sky130_fd_sc_hd__nor3b_1 U18838 ( .C_N(n13612), .A(n18014), .B(n13611), .Y(
        n13613) );
  sky130_fd_sc_hd__o22ai_1 U18839 ( .A1(n13614), .A2(n18172), .B1(n13613), 
        .B2(n18183), .Y(n13615) );
  sky130_fd_sc_hd__nor3_1 U18840 ( .A(n13617), .B(n13616), .C(n13615), .Y(
        n13618) );
  sky130_fd_sc_hd__o22ai_1 U18841 ( .A1(n13619), .A2(n18164), .B1(n13618), 
        .B2(n18139), .Y(n13620) );
  sky130_fd_sc_hd__a22oi_1 U18843 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[274]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[50]), .Y(n13635) );
  sky130_fd_sc_hd__a22o_1 U18844 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[306]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[338]), .X(n13622) );
  sky130_fd_sc_hd__a21oi_1 U18845 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[370]), .B1(n13622), .Y(n13634) );
  sky130_fd_sc_hd__nand2_1 U18846 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[242]), .Y(n13626) );
  sky130_fd_sc_hd__a21oi_1 U18847 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[466]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n13625) );
  sky130_fd_sc_hd__nand2_1 U18848 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[402]), .Y(n13624) );
  sky130_fd_sc_hd__nand2_1 U18849 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[434]), .Y(n13623) );
  sky130_fd_sc_hd__nand4_1 U18850 ( .A(n13626), .B(n13625), .C(n13624), .D(
        n13623), .Y(n13627) );
  sky130_fd_sc_hd__a21oi_1 U18851 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[210]), .B1(n13627), .Y(n13633) );
  sky130_fd_sc_hd__a22o_1 U18852 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[18]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[82]), .X(n13628) );
  sky130_fd_sc_hd__a21oi_1 U18853 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[114]), .B1(n13628), .Y(n13630) );
  sky130_fd_sc_hd__a22oi_1 U18854 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[178]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[146]), .Y(n13629) );
  sky130_fd_sc_hd__nand2_1 U18855 ( .A(n13630), .B(n13629), .Y(n13631) );
  sky130_fd_sc_hd__nand2_1 U18856 ( .A(n13631), .B(n17639), .Y(n13632) );
  sky130_fd_sc_hd__nand4_1 U18857 ( .A(n13635), .B(n13634), .C(n13633), .D(
        n13632), .Y(n13643) );
  sky130_fd_sc_hd__nor2_1 U18858 ( .A(j202_soc_core_memory0_ram_dout0[498]), 
        .B(n18758), .Y(n13636) );
  sky130_fd_sc_hd__nor2_1 U18859 ( .A(n13636), .B(n18761), .Y(n13642) );
  sky130_fd_sc_hd__a22oi_1 U18860 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[18]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[50]), .Y(n13640) );
  sky130_fd_sc_hd__nand2_1 U18861 ( .A(n18727), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[82]), .Y(n13639) );
  sky130_fd_sc_hd__nand2_1 U18862 ( .A(n18379), .B(j202_soc_core_uart_div1[2]), 
        .Y(n13638) );
  sky130_fd_sc_hd__nand2_1 U18863 ( .A(n18629), .B(
        j202_soc_core_bldc_core_00_pwm_duty[6]), .Y(n13637) );
  sky130_fd_sc_hd__nand4_1 U18864 ( .A(n13640), .B(n13639), .C(n13638), .D(
        n13637), .Y(n13641) );
  sky130_fd_sc_hd__a21oi_1 U18865 ( .A1(n13643), .A2(n13642), .B1(n13641), .Y(
        n13644) );
  sky130_fd_sc_hd__nand2_1 U18866 ( .A(n13645), .B(n13644), .Y(n22523) );
  sky130_fd_sc_hd__nand2_1 U18867 ( .A(n22523), .B(n19737), .Y(n13647) );
  sky130_fd_sc_hd__a22oi_1 U18868 ( .A1(n19657), .A2(n21775), .B1(n19736), 
        .B2(n23304), .Y(n13646) );
  sky130_fd_sc_hd__nand2_1 U18869 ( .A(n13647), .B(n13646), .Y(n13648) );
  sky130_fd_sc_hd__a21oi_1 U18870 ( .A1(n21789), .A2(n19661), .B1(n13648), .Y(
        n13649) );
  sky130_fd_sc_hd__nand2_1 U18871 ( .A(n13650), .B(n13649), .Y(n25251) );
  sky130_fd_sc_hd__nand2_1 U18872 ( .A(j202_soc_core_j22_cpu_memop_MEM__1_), 
        .B(j202_soc_core_j22_cpu_memop_MEM__2_), .Y(n13651) );
  sky130_fd_sc_hd__nor2_1 U18873 ( .A(j202_soc_core_j22_cpu_memop_MEM__3_), 
        .B(n13651), .Y(n13656) );
  sky130_fd_sc_hd__nand3_1 U18874 ( .A(n23242), .B(n23240), .C(
        j202_soc_core_j22_cpu_memop_MEM__3_), .Y(n16686) );
  sky130_fd_sc_hd__clkinv_1 U18875 ( .A(n16686), .Y(n13655) );
  sky130_fd_sc_hd__nor2_1 U18876 ( .A(j202_soc_core_j22_cpu_memop_MEM__0_), 
        .B(n23245), .Y(n16689) );
  sky130_fd_sc_hd__nand2_1 U18877 ( .A(n21212), .B(n19917), .Y(n19500) );
  sky130_fd_sc_hd__o31ai_1 U18878 ( .A1(n13656), .A2(n13655), .A3(n19500), 
        .B1(n23239), .Y(n22821) );
  sky130_fd_sc_hd__nand2_1 U18879 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[350]), .Y(n13660) );
  sky130_fd_sc_hd__nand2_1 U18880 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[222]), .Y(n13659) );
  sky130_fd_sc_hd__nand2_1 U18881 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[414]), .Y(n13658) );
  sky130_fd_sc_hd__nand2_1 U18882 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[62]), .Y(n13657) );
  sky130_fd_sc_hd__nand4_1 U18883 ( .A(n13660), .B(n13659), .C(n13658), .D(
        n13657), .Y(n13666) );
  sky130_fd_sc_hd__nand2_1 U18884 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[382]), .Y(n13664) );
  sky130_fd_sc_hd__nand2_1 U18885 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[190]), .Y(n13663) );
  sky130_fd_sc_hd__nand2_1 U18886 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[446]), .Y(n13662) );
  sky130_fd_sc_hd__nand2_1 U18887 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[478]), .Y(n13661) );
  sky130_fd_sc_hd__nand4_1 U18888 ( .A(n13664), .B(n13663), .C(n13662), .D(
        n13661), .Y(n13665) );
  sky130_fd_sc_hd__nor2_1 U18889 ( .A(n13666), .B(n13665), .Y(n13680) );
  sky130_fd_sc_hd__nand2_1 U18890 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[318]), .Y(n13670) );
  sky130_fd_sc_hd__nand2_1 U18891 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[158]), .Y(n13669) );
  sky130_fd_sc_hd__nand2_1 U18892 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[126]), .Y(n13668) );
  sky130_fd_sc_hd__nand2_1 U18893 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[286]), .Y(n13667) );
  sky130_fd_sc_hd__and4_1 U18894 ( .A(n13670), .B(n13669), .C(n13668), .D(
        n13667), .X(n13679) );
  sky130_fd_sc_hd__nor2_1 U18895 ( .A(n13671), .B(n13919), .Y(n13677) );
  sky130_fd_sc_hd__a21oi_1 U18896 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[30]), .B1(n13920), .Y(n13675) );
  sky130_fd_sc_hd__nand2_1 U18897 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[510]), .Y(n13674) );
  sky130_fd_sc_hd__nand2_1 U18898 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[254]), .Y(n13673) );
  sky130_fd_sc_hd__nand2_1 U18899 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[94]), .Y(n13672) );
  sky130_fd_sc_hd__nand4_1 U18900 ( .A(n13675), .B(n13674), .C(n13673), .D(
        n13672), .Y(n13676) );
  sky130_fd_sc_hd__nor2_1 U18901 ( .A(n13677), .B(n13676), .Y(n13678) );
  sky130_fd_sc_hd__nand3_1 U18902 ( .A(n13680), .B(n13679), .C(n13678), .Y(
        n22579) );
  sky130_fd_sc_hd__nand2_1 U18903 ( .A(n22579), .B(n13681), .Y(n13708) );
  sky130_fd_sc_hd__nand2_1 U18904 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[191]), .Y(n13685) );
  sky130_fd_sc_hd__nand2_1 U18905 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[287]), .Y(n13684) );
  sky130_fd_sc_hd__nand2_1 U18906 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[415]), .Y(n13683) );
  sky130_fd_sc_hd__nand2_1 U18907 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[479]), .Y(n13682) );
  sky130_fd_sc_hd__nand4_1 U18908 ( .A(n13685), .B(n13684), .C(n13683), .D(
        n13682), .Y(n13691) );
  sky130_fd_sc_hd__nand2_1 U18909 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[351]), .Y(n13689) );
  sky130_fd_sc_hd__nand2_1 U18910 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[383]), .Y(n13688) );
  sky130_fd_sc_hd__nand2_1 U18911 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[511]), .Y(n13687) );
  sky130_fd_sc_hd__nand2_1 U18912 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[95]), .Y(n13686) );
  sky130_fd_sc_hd__nand4_1 U18913 ( .A(n13689), .B(n13688), .C(n13687), .D(
        n13686), .Y(n13690) );
  sky130_fd_sc_hd__nor2_1 U18914 ( .A(n13691), .B(n13690), .Y(n13705) );
  sky130_fd_sc_hd__nand2_1 U18915 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[223]), .Y(n13695) );
  sky130_fd_sc_hd__nand2_1 U18916 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[319]), .Y(n13694) );
  sky130_fd_sc_hd__nand2_1 U18917 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[127]), .Y(n13693) );
  sky130_fd_sc_hd__nand2_1 U18918 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[447]), .Y(n13692) );
  sky130_fd_sc_hd__and4_1 U18919 ( .A(n13695), .B(n13694), .C(n13693), .D(
        n13692), .X(n13704) );
  sky130_fd_sc_hd__nor2_1 U18920 ( .A(n13696), .B(n13919), .Y(n13702) );
  sky130_fd_sc_hd__a21oi_1 U18921 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[31]), .B1(n13920), .Y(n13700) );
  sky130_fd_sc_hd__nand2_1 U18922 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[63]), .Y(n13699) );
  sky130_fd_sc_hd__nand2_1 U18923 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[255]), .Y(n13698) );
  sky130_fd_sc_hd__nand2_1 U18924 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[159]), .Y(n13697) );
  sky130_fd_sc_hd__nand4_1 U18925 ( .A(n13700), .B(n13699), .C(n13698), .D(
        n13697), .Y(n13701) );
  sky130_fd_sc_hd__nor2_1 U18926 ( .A(n13702), .B(n13701), .Y(n13703) );
  sky130_fd_sc_hd__nand3_1 U18927 ( .A(n13705), .B(n13704), .C(n13703), .Y(
        n22591) );
  sky130_fd_sc_hd__nand2_1 U18928 ( .A(n22591), .B(n13706), .Y(n13707) );
  sky130_fd_sc_hd__nand2_1 U18929 ( .A(n13708), .B(n13707), .Y(n22424) );
  sky130_fd_sc_hd__nand2_1 U18930 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[191]), .Y(n13712) );
  sky130_fd_sc_hd__nand2_1 U18931 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[255]), .Y(n13711) );
  sky130_fd_sc_hd__nand2_1 U18932 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[511]), .Y(n13710) );
  sky130_fd_sc_hd__nand2_1 U18933 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[447]), .Y(n13709) );
  sky130_fd_sc_hd__nand4_1 U18934 ( .A(n13712), .B(n13711), .C(n13710), .D(
        n13709), .Y(n13718) );
  sky130_fd_sc_hd__nand2_1 U18935 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[415]), .Y(n13716) );
  sky130_fd_sc_hd__nand2_1 U18936 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[31]), .Y(n13715) );
  sky130_fd_sc_hd__nand2_1 U18937 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[63]), .Y(n13714) );
  sky130_fd_sc_hd__nand2_1 U18938 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[479]), .Y(n13713) );
  sky130_fd_sc_hd__nand4_1 U18939 ( .A(n13716), .B(n13715), .C(n13714), .D(
        n13713), .Y(n13717) );
  sky130_fd_sc_hd__nor2_1 U18940 ( .A(n13718), .B(n13717), .Y(n13726) );
  sky130_fd_sc_hd__a22oi_1 U18941 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[319]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[223]), .Y(n13725) );
  sky130_fd_sc_hd__a22oi_1 U18942 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[383]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[351]), .Y(n13724) );
  sky130_fd_sc_hd__nand2_1 U18943 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[159]), .Y(n13722) );
  sky130_fd_sc_hd__nand2_1 U18944 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[95]), .Y(n13721) );
  sky130_fd_sc_hd__nand2_1 U18945 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[127]), .Y(n13720) );
  sky130_fd_sc_hd__nand2_1 U18946 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[287]), .Y(n13719) );
  sky130_fd_sc_hd__and4_1 U18947 ( .A(n13722), .B(n13721), .C(n13720), .D(
        n13719), .X(n13723) );
  sky130_fd_sc_hd__nand4_1 U18948 ( .A(n13726), .B(n13725), .C(n13724), .D(
        n13723), .Y(n19647) );
  sky130_fd_sc_hd__nand2_1 U18949 ( .A(n19647), .B(n14086), .Y(n13736) );
  sky130_fd_sc_hd__nand2_1 U18950 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[31]), .Y(n13729) );
  sky130_fd_sc_hd__nand2_1 U18951 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[31]), .Y(n13728) );
  sky130_fd_sc_hd__nand2_1 U18952 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[511]), .Y(n13727) );
  sky130_fd_sc_hd__and4_1 U18953 ( .A(n13729), .B(n13728), .C(n14022), .D(
        n13727), .X(n13735) );
  sky130_fd_sc_hd__nand2_1 U18954 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[31]), .Y(n13733) );
  sky130_fd_sc_hd__nand2_1 U18955 ( .A(n14025), .B(
        j202_soc_core_j22_cpu_pc[31]), .Y(n13732) );
  sky130_fd_sc_hd__nand2_1 U18956 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[31]), .Y(n13731) );
  sky130_fd_sc_hd__nand2_1 U18957 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[31]), .Y(n13730) );
  sky130_fd_sc_hd__and4_1 U18958 ( .A(n13733), .B(n13732), .C(n13731), .D(
        n13730), .X(n13734) );
  sky130_fd_sc_hd__nand3_1 U18959 ( .A(n13736), .B(n13735), .C(n13734), .Y(
        n23344) );
  sky130_fd_sc_hd__nand2_1 U18960 ( .A(n23344), .B(n14089), .Y(n13737) );
  sky130_fd_sc_hd__o21a_1 U18961 ( .A1(n23344), .A2(n14087), .B1(n13737), .X(
        n22423) );
  sky130_fd_sc_hd__nand2_1 U18962 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[61]), .Y(n13741) );
  sky130_fd_sc_hd__nand2_1 U18963 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[477]), .Y(n13740) );
  sky130_fd_sc_hd__nand2_1 U18964 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[509]), .Y(n13739) );
  sky130_fd_sc_hd__nand2_1 U18965 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[93]), .Y(n13738) );
  sky130_fd_sc_hd__nand4_1 U18966 ( .A(n13741), .B(n13740), .C(n13739), .D(
        n13738), .Y(n13747) );
  sky130_fd_sc_hd__nand2_1 U18967 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[221]), .Y(n13745) );
  sky130_fd_sc_hd__nand2_1 U18968 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[317]), .Y(n13744) );
  sky130_fd_sc_hd__nand2_1 U18969 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[445]), .Y(n13743) );
  sky130_fd_sc_hd__nand2_1 U18970 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[157]), .Y(n13742) );
  sky130_fd_sc_hd__nand4_1 U18971 ( .A(n13745), .B(n13744), .C(n13743), .D(
        n13742), .Y(n13746) );
  sky130_fd_sc_hd__nor2_1 U18972 ( .A(n13747), .B(n13746), .Y(n13760) );
  sky130_fd_sc_hd__nand2_1 U18973 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[189]), .Y(n13751) );
  sky130_fd_sc_hd__nand2_1 U18974 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[349]), .Y(n13750) );
  sky130_fd_sc_hd__nand2_1 U18975 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[125]), .Y(n13749) );
  sky130_fd_sc_hd__nand2_1 U18976 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[285]), .Y(n13748) );
  sky130_fd_sc_hd__and4_1 U18977 ( .A(n13751), .B(n13750), .C(n13749), .D(
        n13748), .X(n13759) );
  sky130_fd_sc_hd__nor2_1 U18978 ( .A(n14076), .B(n13919), .Y(n13757) );
  sky130_fd_sc_hd__a21oi_1 U18979 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[29]), .B1(n13920), .Y(n13755) );
  sky130_fd_sc_hd__nand2_1 U18980 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[381]), .Y(n13754) );
  sky130_fd_sc_hd__nand2_1 U18981 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[253]), .Y(n13753) );
  sky130_fd_sc_hd__nand2_1 U18982 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[413]), .Y(n13752) );
  sky130_fd_sc_hd__nand4_1 U18983 ( .A(n13755), .B(n13754), .C(n13753), .D(
        n13752), .Y(n13756) );
  sky130_fd_sc_hd__nor2_1 U18984 ( .A(n13757), .B(n13756), .Y(n13758) );
  sky130_fd_sc_hd__nand3_1 U18985 ( .A(n13760), .B(n13759), .C(n13758), .Y(
        n22575) );
  sky130_fd_sc_hd__o22ai_1 U18986 ( .A1(n14042), .A2(n21048), .B1(n22604), 
        .B2(n20677), .Y(n14677) );
  sky130_fd_sc_hd__nand2_1 U18987 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[190]), .Y(n13764) );
  sky130_fd_sc_hd__nand2_1 U18988 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[254]), .Y(n13763) );
  sky130_fd_sc_hd__nand2_1 U18989 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[510]), .Y(n13762) );
  sky130_fd_sc_hd__nand2_1 U18990 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[446]), .Y(n13761) );
  sky130_fd_sc_hd__nand4_1 U18991 ( .A(n13764), .B(n13763), .C(n13762), .D(
        n13761), .Y(n13770) );
  sky130_fd_sc_hd__nand2_1 U18992 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[414]), .Y(n13768) );
  sky130_fd_sc_hd__nand2_1 U18993 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[30]), .Y(n13767) );
  sky130_fd_sc_hd__nand2_1 U18994 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[62]), .Y(n13766) );
  sky130_fd_sc_hd__nand2_1 U18995 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[478]), .Y(n13765) );
  sky130_fd_sc_hd__nand4_1 U18996 ( .A(n13768), .B(n13767), .C(n13766), .D(
        n13765), .Y(n13769) );
  sky130_fd_sc_hd__nor2_1 U18997 ( .A(n13770), .B(n13769), .Y(n13778) );
  sky130_fd_sc_hd__a22oi_1 U18998 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[318]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[222]), .Y(n13777) );
  sky130_fd_sc_hd__a22oi_1 U18999 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[382]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[350]), .Y(n13776) );
  sky130_fd_sc_hd__nand2_1 U19000 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[158]), .Y(n13774) );
  sky130_fd_sc_hd__nand2_1 U19001 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[94]), .Y(n13773) );
  sky130_fd_sc_hd__nand2_1 U19002 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[126]), .Y(n13772) );
  sky130_fd_sc_hd__nand2_1 U19003 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[286]), .Y(n13771) );
  sky130_fd_sc_hd__and4_1 U19004 ( .A(n13774), .B(n13773), .C(n13772), .D(
        n13771), .X(n13775) );
  sky130_fd_sc_hd__nand4_1 U19005 ( .A(n13778), .B(n13777), .C(n13776), .D(
        n13775), .Y(n19762) );
  sky130_fd_sc_hd__nand2_1 U19006 ( .A(n19762), .B(n14086), .Y(n13788) );
  sky130_fd_sc_hd__nand2_1 U19007 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[30]), .Y(n13781) );
  sky130_fd_sc_hd__nand2_1 U19008 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[30]), .Y(n13780) );
  sky130_fd_sc_hd__nand2_1 U19009 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[510]), .Y(n13779) );
  sky130_fd_sc_hd__and4_1 U19010 ( .A(n13781), .B(n13780), .C(n14022), .D(
        n13779), .X(n13787) );
  sky130_fd_sc_hd__nand2_1 U19011 ( .A(n14025), .B(
        j202_soc_core_j22_cpu_pc[30]), .Y(n13785) );
  sky130_fd_sc_hd__nand2_1 U19012 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[30]), .Y(n13784) );
  sky130_fd_sc_hd__nand2_1 U19013 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[30]), .Y(n13783) );
  sky130_fd_sc_hd__nand2_1 U19014 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[30]), .Y(n13782) );
  sky130_fd_sc_hd__and4_1 U19015 ( .A(n13785), .B(n13784), .C(n13783), .D(
        n13782), .X(n13786) );
  sky130_fd_sc_hd__nand3_1 U19016 ( .A(n13788), .B(n13787), .C(n13786), .Y(
        n23340) );
  sky130_fd_sc_hd__nand2_1 U19017 ( .A(n22603), .B(n14087), .Y(n13789) );
  sky130_fd_sc_hd__nand2_1 U19019 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[220]), .Y(n13793) );
  sky130_fd_sc_hd__nand2_1 U19020 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[92]), .Y(n13792) );
  sky130_fd_sc_hd__nand2_1 U19021 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[412]), .Y(n13791) );
  sky130_fd_sc_hd__nand2_1 U19022 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[508]), .Y(n13790) );
  sky130_fd_sc_hd__nand4_1 U19023 ( .A(n13793), .B(n13792), .C(n13791), .D(
        n13790), .Y(n13799) );
  sky130_fd_sc_hd__nand2_1 U19024 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[188]), .Y(n13797) );
  sky130_fd_sc_hd__nand2_1 U19025 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[316]), .Y(n13796) );
  sky130_fd_sc_hd__nand2_1 U19026 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[156]), .Y(n13795) );
  sky130_fd_sc_hd__nand2_1 U19027 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[444]), .Y(n13794) );
  sky130_fd_sc_hd__nand4_1 U19028 ( .A(n13797), .B(n13796), .C(n13795), .D(
        n13794), .Y(n13798) );
  sky130_fd_sc_hd__nor2_1 U19029 ( .A(n13799), .B(n13798), .Y(n13812) );
  sky130_fd_sc_hd__nor2_1 U19030 ( .A(n13860), .B(n13919), .Y(n13805) );
  sky130_fd_sc_hd__a21oi_1 U19031 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[28]), .B1(n13920), .Y(n13803) );
  sky130_fd_sc_hd__nand2_1 U19032 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[60]), .Y(n13802) );
  sky130_fd_sc_hd__nand2_1 U19033 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[252]), .Y(n13801) );
  sky130_fd_sc_hd__nand2_1 U19034 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[380]), .Y(n13800) );
  sky130_fd_sc_hd__nand4_1 U19035 ( .A(n13803), .B(n13802), .C(n13801), .D(
        n13800), .Y(n13804) );
  sky130_fd_sc_hd__nor2_1 U19036 ( .A(n13805), .B(n13804), .Y(n13811) );
  sky130_fd_sc_hd__nand2_1 U19037 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[348]), .Y(n13809) );
  sky130_fd_sc_hd__nand2_1 U19038 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[476]), .Y(n13808) );
  sky130_fd_sc_hd__nand2_1 U19039 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[124]), .Y(n13807) );
  sky130_fd_sc_hd__nand2_1 U19040 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[284]), .Y(n13806) );
  sky130_fd_sc_hd__and4_1 U19041 ( .A(n13809), .B(n13808), .C(n13807), .D(
        n13806), .X(n13810) );
  sky130_fd_sc_hd__nand3_1 U19042 ( .A(n13812), .B(n13811), .C(n13810), .Y(
        n22631) );
  sky130_fd_sc_hd__nand2_1 U19043 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[59]), .Y(n13816) );
  sky130_fd_sc_hd__nand2_1 U19044 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[91]), .Y(n13815) );
  sky130_fd_sc_hd__nand2_1 U19045 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[123]), .Y(n13814) );
  sky130_fd_sc_hd__nand2_1 U19046 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[507]), .Y(n13813) );
  sky130_fd_sc_hd__nand4_1 U19047 ( .A(n13816), .B(n13815), .C(n13814), .D(
        n13813), .Y(n13822) );
  sky130_fd_sc_hd__nand2_1 U19048 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[219]), .Y(n13820) );
  sky130_fd_sc_hd__nand2_1 U19049 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[315]), .Y(n13819) );
  sky130_fd_sc_hd__nand2_1 U19050 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[443]), .Y(n13818) );
  sky130_fd_sc_hd__nand2_1 U19051 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[347]), .Y(n13817) );
  sky130_fd_sc_hd__nand4_1 U19052 ( .A(n13820), .B(n13819), .C(n13818), .D(
        n13817), .Y(n13821) );
  sky130_fd_sc_hd__nor2_1 U19053 ( .A(n13822), .B(n13821), .Y(n13836) );
  sky130_fd_sc_hd__nor2_1 U19054 ( .A(n13823), .B(n13919), .Y(n13829) );
  sky130_fd_sc_hd__a21oi_1 U19055 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[27]), .B1(n13920), .Y(n13827) );
  sky130_fd_sc_hd__nand2_1 U19056 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[379]), .Y(n13826) );
  sky130_fd_sc_hd__nand2_1 U19057 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[251]), .Y(n13825) );
  sky130_fd_sc_hd__nand2_1 U19058 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[411]), .Y(n13824) );
  sky130_fd_sc_hd__nand4_1 U19059 ( .A(n13827), .B(n13826), .C(n13825), .D(
        n13824), .Y(n13828) );
  sky130_fd_sc_hd__nor2_1 U19060 ( .A(n13829), .B(n13828), .Y(n13835) );
  sky130_fd_sc_hd__nand2_1 U19061 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[187]), .Y(n13833) );
  sky130_fd_sc_hd__nand2_1 U19062 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[155]), .Y(n13832) );
  sky130_fd_sc_hd__nand2_1 U19063 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[283]), .Y(n13831) );
  sky130_fd_sc_hd__nand2_1 U19064 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[475]), .Y(n13830) );
  sky130_fd_sc_hd__and4_1 U19065 ( .A(n13833), .B(n13832), .C(n13831), .D(
        n13830), .X(n13834) );
  sky130_fd_sc_hd__nand3_1 U19066 ( .A(n13836), .B(n13835), .C(n13834), .Y(
        n22576) );
  sky130_fd_sc_hd__o22ai_1 U19067 ( .A1(n20677), .A2(n20955), .B1(n22610), 
        .B2(n14042), .Y(n14040) );
  sky130_fd_sc_hd__nand2_1 U19068 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[188]), .Y(n13840) );
  sky130_fd_sc_hd__nand2_1 U19069 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[252]), .Y(n13839) );
  sky130_fd_sc_hd__nand2_1 U19070 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[508]), .Y(n13838) );
  sky130_fd_sc_hd__nand2_1 U19071 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[444]), .Y(n13837) );
  sky130_fd_sc_hd__nand4_1 U19072 ( .A(n13840), .B(n13839), .C(n13838), .D(
        n13837), .Y(n13846) );
  sky130_fd_sc_hd__nand2_1 U19073 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[412]), .Y(n13844) );
  sky130_fd_sc_hd__nand2_1 U19074 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[28]), .Y(n13843) );
  sky130_fd_sc_hd__nand2_1 U19075 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[60]), .Y(n13842) );
  sky130_fd_sc_hd__nand2_1 U19076 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[476]), .Y(n13841) );
  sky130_fd_sc_hd__nand4_1 U19077 ( .A(n13844), .B(n13843), .C(n13842), .D(
        n13841), .Y(n13845) );
  sky130_fd_sc_hd__nor2_1 U19078 ( .A(n13846), .B(n13845), .Y(n13857) );
  sky130_fd_sc_hd__nand2_1 U19079 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[348]), .Y(n13850) );
  sky130_fd_sc_hd__nand2_1 U19080 ( .A(n11191), .B(
        j202_soc_core_j22_cpu_rf_gpr[220]), .Y(n13849) );
  sky130_fd_sc_hd__nand2_1 U19081 ( .A(n20285), .B(
        j202_soc_core_j22_cpu_rf_gpr[316]), .Y(n13848) );
  sky130_fd_sc_hd__nand2_1 U19082 ( .A(n20282), .B(
        j202_soc_core_j22_cpu_rf_gpr[380]), .Y(n13847) );
  sky130_fd_sc_hd__and4_1 U19083 ( .A(n13850), .B(n13849), .C(n13848), .D(
        n13847), .X(n13856) );
  sky130_fd_sc_hd__nand2_1 U19084 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[156]), .Y(n13854) );
  sky130_fd_sc_hd__nand2_1 U19085 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[92]), .Y(n13853) );
  sky130_fd_sc_hd__nand2_1 U19086 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[124]), .Y(n13852) );
  sky130_fd_sc_hd__nand2_1 U19087 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[284]), .Y(n13851) );
  sky130_fd_sc_hd__and4_1 U19088 ( .A(n13854), .B(n13853), .C(n13852), .D(
        n13851), .X(n13855) );
  sky130_fd_sc_hd__nand3_1 U19089 ( .A(n13857), .B(n13856), .C(n13855), .Y(
        n19785) );
  sky130_fd_sc_hd__a21oi_1 U19090 ( .A1(n14069), .A2(
        j202_soc_core_j22_cpu_rf_vbr[28]), .B1(n14068), .Y(n13866) );
  sky130_fd_sc_hd__a2bb2oi_1 U19091 ( .B1(j202_soc_core_j22_cpu_rf_gpr[508]), 
        .B2(n14072), .A1_N(n14071), .A2_N(n13858), .Y(n13865) );
  sky130_fd_sc_hd__o22a_1 U19092 ( .A1(n13860), .A2(n14075), .B1(n13859), .B2(
        n14073), .X(n13864) );
  sky130_fd_sc_hd__o22a_1 U19093 ( .A1(n13862), .A2(n14079), .B1(n13861), .B2(
        n14077), .X(n13863) );
  sky130_fd_sc_hd__nand4_1 U19094 ( .A(n13866), .B(n13865), .C(n13864), .D(
        n13863), .Y(n13867) );
  sky130_fd_sc_hd__a21oi_1 U19095 ( .A1(n19785), .A2(n14086), .B1(n13867), .Y(
        n22074) );
  sky130_fd_sc_hd__nand2_1 U19096 ( .A(n22074), .B(n14087), .Y(n13868) );
  sky130_fd_sc_hd__nor2_1 U19098 ( .A(n14040), .B(n14041), .Y(n14802) );
  sky130_fd_sc_hd__nand2_1 U19099 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[217]), .Y(n13872) );
  sky130_fd_sc_hd__nand2_1 U19100 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[89]), .Y(n13871) );
  sky130_fd_sc_hd__nand2_1 U19101 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[409]), .Y(n13870) );
  sky130_fd_sc_hd__nand2_1 U19102 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[505]), .Y(n13869) );
  sky130_fd_sc_hd__nand4_1 U19103 ( .A(n13872), .B(n13871), .C(n13870), .D(
        n13869), .Y(n13878) );
  sky130_fd_sc_hd__nand2_1 U19104 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[185]), .Y(n13876) );
  sky130_fd_sc_hd__nand2_1 U19105 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[313]), .Y(n13875) );
  sky130_fd_sc_hd__nand2_1 U19106 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[153]), .Y(n13874) );
  sky130_fd_sc_hd__nand2_1 U19107 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[441]), .Y(n13873) );
  sky130_fd_sc_hd__nand4_1 U19108 ( .A(n13876), .B(n13875), .C(n13874), .D(
        n13873), .Y(n13877) );
  sky130_fd_sc_hd__nor2_1 U19109 ( .A(n13878), .B(n13877), .Y(n13892) );
  sky130_fd_sc_hd__nor2_1 U19110 ( .A(n13879), .B(n13919), .Y(n13885) );
  sky130_fd_sc_hd__a21oi_1 U19111 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[25]), .B1(n13920), .Y(n13883) );
  sky130_fd_sc_hd__nand2_1 U19112 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[57]), .Y(n13882) );
  sky130_fd_sc_hd__nand2_1 U19113 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[249]), .Y(n13881) );
  sky130_fd_sc_hd__nand2_1 U19114 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[377]), .Y(n13880) );
  sky130_fd_sc_hd__nand4_1 U19115 ( .A(n13883), .B(n13882), .C(n13881), .D(
        n13880), .Y(n13884) );
  sky130_fd_sc_hd__nor2_1 U19116 ( .A(n13885), .B(n13884), .Y(n13891) );
  sky130_fd_sc_hd__nand2_1 U19117 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[345]), .Y(n13889) );
  sky130_fd_sc_hd__nand2_1 U19118 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[473]), .Y(n13888) );
  sky130_fd_sc_hd__nand2_1 U19119 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[121]), .Y(n13887) );
  sky130_fd_sc_hd__nand2_1 U19120 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[281]), .Y(n13886) );
  sky130_fd_sc_hd__and4_1 U19121 ( .A(n13889), .B(n13888), .C(n13887), .D(
        n13886), .X(n13890) );
  sky130_fd_sc_hd__nand3_1 U19122 ( .A(n13892), .B(n13891), .C(n13890), .Y(
        n22574) );
  sky130_fd_sc_hd__nand2_1 U19123 ( .A(n13893), .B(
        j202_soc_core_j22_cpu_rf_gpr[250]), .Y(n13900) );
  sky130_fd_sc_hd__nand2_1 U19124 ( .A(n13894), .B(
        j202_soc_core_j22_cpu_rf_gpr[58]), .Y(n13899) );
  sky130_fd_sc_hd__nand2_1 U19125 ( .A(n13895), .B(
        j202_soc_core_j22_cpu_rf_gpr[122]), .Y(n13898) );
  sky130_fd_sc_hd__nand2_1 U19126 ( .A(n13896), .B(
        j202_soc_core_j22_cpu_rf_gpr[90]), .Y(n13897) );
  sky130_fd_sc_hd__nand4_1 U19127 ( .A(n13900), .B(n13899), .C(n13898), .D(
        n13897), .Y(n13910) );
  sky130_fd_sc_hd__nand2_1 U19128 ( .A(n13901), .B(
        j202_soc_core_j22_cpu_rf_gpr[218]), .Y(n13908) );
  sky130_fd_sc_hd__nand2_1 U19129 ( .A(n13902), .B(
        j202_soc_core_j22_cpu_rf_gpr[346]), .Y(n13907) );
  sky130_fd_sc_hd__nand2_1 U19130 ( .A(n13903), .B(
        j202_soc_core_j22_cpu_rf_gpr[474]), .Y(n13906) );
  sky130_fd_sc_hd__nand2_1 U19131 ( .A(n13904), .B(
        j202_soc_core_j22_cpu_rf_gpr[282]), .Y(n13905) );
  sky130_fd_sc_hd__nand4_1 U19132 ( .A(n13908), .B(n13907), .C(n13906), .D(
        n13905), .Y(n13909) );
  sky130_fd_sc_hd__nor2_1 U19133 ( .A(n13910), .B(n13909), .Y(n13932) );
  sky130_fd_sc_hd__nand2_1 U19134 ( .A(n13911), .B(
        j202_soc_core_j22_cpu_rf_gpr[314]), .Y(n13918) );
  sky130_fd_sc_hd__nand2_1 U19135 ( .A(n13912), .B(
        j202_soc_core_j22_cpu_rf_gpr[154]), .Y(n13917) );
  sky130_fd_sc_hd__nand2_1 U19136 ( .A(n13913), .B(
        j202_soc_core_j22_cpu_rf_gpr[410]), .Y(n13916) );
  sky130_fd_sc_hd__nand2_1 U19137 ( .A(n13914), .B(
        j202_soc_core_j22_cpu_rf_gpr[442]), .Y(n13915) );
  sky130_fd_sc_hd__and4_1 U19138 ( .A(n13918), .B(n13917), .C(n13916), .D(
        n13915), .X(n13931) );
  sky130_fd_sc_hd__nor2_1 U19139 ( .A(n13956), .B(n13919), .Y(n13929) );
  sky130_fd_sc_hd__a21oi_1 U19140 ( .A1(n11184), .A2(
        j202_soc_core_j22_cpu_rf_tmp[26]), .B1(n13920), .Y(n13927) );
  sky130_fd_sc_hd__nand2_1 U19141 ( .A(n13921), .B(
        j202_soc_core_j22_cpu_rf_gpr[186]), .Y(n13926) );
  sky130_fd_sc_hd__nand2_1 U19142 ( .A(n13922), .B(
        j202_soc_core_j22_cpu_rf_gpr[378]), .Y(n13925) );
  sky130_fd_sc_hd__nand2_1 U19143 ( .A(n13923), .B(
        j202_soc_core_j22_cpu_rf_gpr[506]), .Y(n13924) );
  sky130_fd_sc_hd__nand4_1 U19144 ( .A(n13927), .B(n13926), .C(n13925), .D(
        n13924), .Y(n13928) );
  sky130_fd_sc_hd__nor2_1 U19145 ( .A(n13929), .B(n13928), .Y(n13930) );
  sky130_fd_sc_hd__nand3_1 U19146 ( .A(n13932), .B(n13931), .C(n13930), .Y(
        n22573) );
  sky130_fd_sc_hd__o22ai_1 U19147 ( .A1(n14042), .A2(n22606), .B1(n22601), 
        .B2(n20677), .Y(n14000) );
  sky130_fd_sc_hd__nand2_1 U19148 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[186]), .Y(n13936) );
  sky130_fd_sc_hd__nand2_1 U19149 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[250]), .Y(n13935) );
  sky130_fd_sc_hd__nand2_1 U19150 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[506]), .Y(n13934) );
  sky130_fd_sc_hd__nand2_1 U19151 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[442]), .Y(n13933) );
  sky130_fd_sc_hd__nand4_1 U19152 ( .A(n13936), .B(n13935), .C(n13934), .D(
        n13933), .Y(n13942) );
  sky130_fd_sc_hd__nand2_1 U19153 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[410]), .Y(n13940) );
  sky130_fd_sc_hd__nand2_1 U19154 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[26]), .Y(n13939) );
  sky130_fd_sc_hd__nand2_1 U19155 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[58]), .Y(n13938) );
  sky130_fd_sc_hd__nand2_1 U19156 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[474]), .Y(n13937) );
  sky130_fd_sc_hd__nand4_1 U19157 ( .A(n13940), .B(n13939), .C(n13938), .D(
        n13937), .Y(n13941) );
  sky130_fd_sc_hd__nor2_1 U19158 ( .A(n13942), .B(n13941), .Y(n13953) );
  sky130_fd_sc_hd__nand2_1 U19159 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[346]), .Y(n13946) );
  sky130_fd_sc_hd__nand2_1 U19160 ( .A(n11191), .B(
        j202_soc_core_j22_cpu_rf_gpr[218]), .Y(n13945) );
  sky130_fd_sc_hd__nand2_1 U19161 ( .A(n20285), .B(
        j202_soc_core_j22_cpu_rf_gpr[314]), .Y(n13944) );
  sky130_fd_sc_hd__nand2_1 U19162 ( .A(n20282), .B(
        j202_soc_core_j22_cpu_rf_gpr[378]), .Y(n13943) );
  sky130_fd_sc_hd__and4_1 U19163 ( .A(n13946), .B(n13945), .C(n13944), .D(
        n13943), .X(n13952) );
  sky130_fd_sc_hd__nand2_1 U19164 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[154]), .Y(n13950) );
  sky130_fd_sc_hd__nand2_1 U19165 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[90]), .Y(n13949) );
  sky130_fd_sc_hd__nand2_1 U19166 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[122]), .Y(n13948) );
  sky130_fd_sc_hd__nand2_1 U19167 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[282]), .Y(n13947) );
  sky130_fd_sc_hd__and4_1 U19168 ( .A(n13950), .B(n13949), .C(n13948), .D(
        n13947), .X(n13951) );
  sky130_fd_sc_hd__nand3_1 U19169 ( .A(n13953), .B(n13952), .C(n13951), .Y(
        n19575) );
  sky130_fd_sc_hd__a21oi_1 U19170 ( .A1(n14069), .A2(
        j202_soc_core_j22_cpu_rf_vbr[26]), .B1(n14068), .Y(n13962) );
  sky130_fd_sc_hd__a2bb2oi_1 U19171 ( .B1(j202_soc_core_j22_cpu_rf_gpr[506]), 
        .B2(n14072), .A1_N(n14071), .A2_N(n13954), .Y(n13961) );
  sky130_fd_sc_hd__o22a_1 U19172 ( .A1(n13956), .A2(n14075), .B1(n13955), .B2(
        n14073), .X(n13960) );
  sky130_fd_sc_hd__o22a_1 U19173 ( .A1(n13958), .A2(n14079), .B1(n13957), .B2(
        n14077), .X(n13959) );
  sky130_fd_sc_hd__nand4_1 U19174 ( .A(n13962), .B(n13961), .C(n13960), .D(
        n13959), .Y(n13963) );
  sky130_fd_sc_hd__a21oi_1 U19175 ( .A1(n19575), .A2(n14086), .B1(n13963), .Y(
        n22602) );
  sky130_fd_sc_hd__nand2_1 U19176 ( .A(n22602), .B(n14087), .Y(n13964) );
  sky130_fd_sc_hd__nor2_1 U19178 ( .A(n14000), .B(n14001), .Y(n14531) );
  sky130_fd_sc_hd__o21ai_1 U19179 ( .A1(n13967), .A2(n13966), .B1(n13965), .Y(
        n14274) );
  sky130_fd_sc_hd__o22ai_1 U19180 ( .A1(n20677), .A2(n22606), .B1(n22568), 
        .B2(n14042), .Y(n13997) );
  sky130_fd_sc_hd__nand2_1 U19181 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[185]), .Y(n13971) );
  sky130_fd_sc_hd__nand2_1 U19182 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[249]), .Y(n13970) );
  sky130_fd_sc_hd__nand2_1 U19183 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[505]), .Y(n13969) );
  sky130_fd_sc_hd__nand2_1 U19184 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[441]), .Y(n13968) );
  sky130_fd_sc_hd__nand4_1 U19185 ( .A(n13971), .B(n13970), .C(n13969), .D(
        n13968), .Y(n13977) );
  sky130_fd_sc_hd__nand2_1 U19186 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[409]), .Y(n13975) );
  sky130_fd_sc_hd__nand2_1 U19187 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[25]), .Y(n13974) );
  sky130_fd_sc_hd__nand2_1 U19188 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[57]), .Y(n13973) );
  sky130_fd_sc_hd__nand2_1 U19189 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[473]), .Y(n13972) );
  sky130_fd_sc_hd__nand4_1 U19190 ( .A(n13975), .B(n13974), .C(n13973), .D(
        n13972), .Y(n13976) );
  sky130_fd_sc_hd__nor2_1 U19191 ( .A(n13977), .B(n13976), .Y(n13985) );
  sky130_fd_sc_hd__a22oi_1 U19192 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[313]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[217]), .Y(n13984) );
  sky130_fd_sc_hd__a22oi_1 U19193 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[377]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[345]), .Y(n13983) );
  sky130_fd_sc_hd__nand2_1 U19194 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[153]), .Y(n13981) );
  sky130_fd_sc_hd__nand2_1 U19195 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[89]), .Y(n13980) );
  sky130_fd_sc_hd__nand2_1 U19196 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[121]), .Y(n13979) );
  sky130_fd_sc_hd__nand2_1 U19197 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[281]), .Y(n13978) );
  sky130_fd_sc_hd__and4_1 U19198 ( .A(n13981), .B(n13980), .C(n13979), .D(
        n13978), .X(n13982) );
  sky130_fd_sc_hd__nand4_1 U19199 ( .A(n13985), .B(n13984), .C(n13983), .D(
        n13982), .Y(n19997) );
  sky130_fd_sc_hd__nand2_1 U19200 ( .A(n19997), .B(n14086), .Y(n13995) );
  sky130_fd_sc_hd__nand2_1 U19201 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[25]), .Y(n13988) );
  sky130_fd_sc_hd__nand2_1 U19202 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[25]), .Y(n13987) );
  sky130_fd_sc_hd__nand2_1 U19203 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[505]), .Y(n13986) );
  sky130_fd_sc_hd__and4_1 U19204 ( .A(n13988), .B(n13987), .C(n14022), .D(
        n13986), .X(n13994) );
  sky130_fd_sc_hd__nand2_1 U19205 ( .A(n14025), .B(
        j202_soc_core_j22_cpu_pc[25]), .Y(n13992) );
  sky130_fd_sc_hd__nand2_1 U19206 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[25]), .Y(n13991) );
  sky130_fd_sc_hd__nand2_1 U19207 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[25]), .Y(n13990) );
  sky130_fd_sc_hd__nand2_1 U19208 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[25]), .Y(n13989) );
  sky130_fd_sc_hd__and4_1 U19209 ( .A(n13992), .B(n13991), .C(n13990), .D(
        n13989), .X(n13993) );
  sky130_fd_sc_hd__nand3_1 U19210 ( .A(n13995), .B(n13994), .C(n13993), .Y(
        n23324) );
  sky130_fd_sc_hd__nand2_1 U19211 ( .A(n22605), .B(n14087), .Y(n13996) );
  sky130_fd_sc_hd__o21ai_1 U19212 ( .A1(n14089), .A2(n22605), .B1(n13996), .Y(
        n13998) );
  sky130_fd_sc_hd__nand2_1 U19213 ( .A(n13998), .B(n13997), .Y(n14273) );
  sky130_fd_sc_hd__a21oi_1 U19214 ( .A1(n14274), .A2(n11189), .B1(n13999), .Y(
        n14535) );
  sky130_fd_sc_hd__nand2_1 U19215 ( .A(n14001), .B(n14000), .Y(n14532) );
  sky130_fd_sc_hd__o21ai_1 U19216 ( .A1(n14531), .A2(n14535), .B1(n14532), .Y(
        n14181) );
  sky130_fd_sc_hd__o22ai_1 U19217 ( .A1(n20677), .A2(n22610), .B1(n22601), 
        .B2(n14042), .Y(n14037) );
  sky130_fd_sc_hd__nand2_1 U19218 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[187]), .Y(n14005) );
  sky130_fd_sc_hd__nand2_1 U19219 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[251]), .Y(n14004) );
  sky130_fd_sc_hd__nand2_1 U19220 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[507]), .Y(n14003) );
  sky130_fd_sc_hd__nand2_1 U19221 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[443]), .Y(n14002) );
  sky130_fd_sc_hd__nand4_1 U19222 ( .A(n14005), .B(n14004), .C(n14003), .D(
        n14002), .Y(n14011) );
  sky130_fd_sc_hd__nand2_1 U19223 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[411]), .Y(n14009) );
  sky130_fd_sc_hd__nand2_1 U19224 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[27]), .Y(n14008) );
  sky130_fd_sc_hd__nand2_1 U19225 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[59]), .Y(n14007) );
  sky130_fd_sc_hd__nand2_1 U19226 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[475]), .Y(n14006) );
  sky130_fd_sc_hd__nand4_1 U19227 ( .A(n14009), .B(n14008), .C(n14007), .D(
        n14006), .Y(n14010) );
  sky130_fd_sc_hd__nor2_1 U19228 ( .A(n14011), .B(n14010), .Y(n14019) );
  sky130_fd_sc_hd__a22oi_1 U19229 ( .A1(n20285), .A2(
        j202_soc_core_j22_cpu_rf_gpr[315]), .B1(n11191), .B2(
        j202_soc_core_j22_cpu_rf_gpr[219]), .Y(n14018) );
  sky130_fd_sc_hd__a22oi_1 U19230 ( .A1(n20282), .A2(
        j202_soc_core_j22_cpu_rf_gpr[379]), .B1(n11193), .B2(
        j202_soc_core_j22_cpu_rf_gpr[347]), .Y(n14017) );
  sky130_fd_sc_hd__nand2_1 U19231 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[155]), .Y(n14015) );
  sky130_fd_sc_hd__nand2_1 U19232 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[91]), .Y(n14014) );
  sky130_fd_sc_hd__nand2_1 U19233 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[123]), .Y(n14013) );
  sky130_fd_sc_hd__nand2_1 U19234 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[283]), .Y(n14012) );
  sky130_fd_sc_hd__and4_1 U19235 ( .A(n14015), .B(n14014), .C(n14013), .D(
        n14012), .X(n14016) );
  sky130_fd_sc_hd__nand4_1 U19236 ( .A(n14019), .B(n14018), .C(n14017), .D(
        n14016), .Y(n19822) );
  sky130_fd_sc_hd__nand2_1 U19237 ( .A(n19822), .B(n14086), .Y(n14035) );
  sky130_fd_sc_hd__nand2_1 U19238 ( .A(n14069), .B(
        j202_soc_core_j22_cpu_rf_vbr[27]), .Y(n14024) );
  sky130_fd_sc_hd__nand2_1 U19239 ( .A(n14020), .B(
        j202_soc_core_j22_cpu_rf_tmp[27]), .Y(n14023) );
  sky130_fd_sc_hd__nand2_1 U19240 ( .A(n14072), .B(
        j202_soc_core_j22_cpu_rf_gpr[507]), .Y(n14021) );
  sky130_fd_sc_hd__and4_1 U19241 ( .A(n14024), .B(n14023), .C(n14022), .D(
        n14021), .X(n14034) );
  sky130_fd_sc_hd__nand2_1 U19242 ( .A(n14025), .B(
        j202_soc_core_j22_cpu_pc[27]), .Y(n14032) );
  sky130_fd_sc_hd__nand2_1 U19243 ( .A(n14026), .B(
        j202_soc_core_j22_cpu_rf_gpr[27]), .Y(n14031) );
  sky130_fd_sc_hd__nand2_1 U19244 ( .A(n14027), .B(
        j202_soc_core_j22_cpu_rf_pr[27]), .Y(n14030) );
  sky130_fd_sc_hd__nand2_1 U19245 ( .A(n14028), .B(
        j202_soc_core_j22_cpu_rf_gbr[27]), .Y(n14029) );
  sky130_fd_sc_hd__and4_1 U19246 ( .A(n14032), .B(n14031), .C(n14030), .D(
        n14029), .X(n14033) );
  sky130_fd_sc_hd__nand3_1 U19247 ( .A(n14035), .B(n14034), .C(n14033), .Y(
        n23330) );
  sky130_fd_sc_hd__nand2_1 U19248 ( .A(n22609), .B(n14087), .Y(n14036) );
  sky130_fd_sc_hd__nand2_1 U19250 ( .A(n14038), .B(n14037), .Y(n14180) );
  sky130_fd_sc_hd__a21oi_1 U19251 ( .A1(n14181), .A2(n11185), .B1(n14039), .Y(
        n14806) );
  sky130_fd_sc_hd__nand2_1 U19252 ( .A(n14041), .B(n14040), .Y(n14803) );
  sky130_fd_sc_hd__o21ai_1 U19253 ( .A1(n14802), .A2(n14806), .B1(n14803), .Y(
        n14396) );
  sky130_fd_sc_hd__o22ai_1 U19254 ( .A1(n14042), .A2(n20955), .B1(n21048), 
        .B2(n20677), .Y(n14090) );
  sky130_fd_sc_hd__nand2_1 U19255 ( .A(n20304), .B(
        j202_soc_core_j22_cpu_rf_gpr[189]), .Y(n14046) );
  sky130_fd_sc_hd__nand2_1 U19256 ( .A(n20301), .B(
        j202_soc_core_j22_cpu_rf_gpr[253]), .Y(n14045) );
  sky130_fd_sc_hd__nand2_1 U19257 ( .A(n20238), .B(
        j202_soc_core_j22_cpu_rf_gpr[509]), .Y(n14044) );
  sky130_fd_sc_hd__nand2_1 U19258 ( .A(n20288), .B(
        j202_soc_core_j22_cpu_rf_gpr[445]), .Y(n14043) );
  sky130_fd_sc_hd__nand4_1 U19259 ( .A(n14046), .B(n14045), .C(n14044), .D(
        n14043), .Y(n14053) );
  sky130_fd_sc_hd__nand2_1 U19260 ( .A(n14047), .B(
        j202_soc_core_j22_cpu_rf_gpr[413]), .Y(n14051) );
  sky130_fd_sc_hd__nand2_1 U19261 ( .A(n20250), .B(
        j202_soc_core_j22_cpu_rf_gpr[29]), .Y(n14050) );
  sky130_fd_sc_hd__nand2_1 U19262 ( .A(n20293), .B(
        j202_soc_core_j22_cpu_rf_gpr[61]), .Y(n14049) );
  sky130_fd_sc_hd__nand2_1 U19263 ( .A(n11183), .B(
        j202_soc_core_j22_cpu_rf_gpr[477]), .Y(n14048) );
  sky130_fd_sc_hd__nand4_1 U19264 ( .A(n14051), .B(n14050), .C(n14049), .D(
        n14048), .Y(n14052) );
  sky130_fd_sc_hd__nor2_1 U19265 ( .A(n14053), .B(n14052), .Y(n14067) );
  sky130_fd_sc_hd__nand2_1 U19266 ( .A(n11193), .B(
        j202_soc_core_j22_cpu_rf_gpr[349]), .Y(n14057) );
  sky130_fd_sc_hd__nand2_1 U19267 ( .A(n11191), .B(
        j202_soc_core_j22_cpu_rf_gpr[221]), .Y(n14056) );
  sky130_fd_sc_hd__nand2_1 U19268 ( .A(n20285), .B(
        j202_soc_core_j22_cpu_rf_gpr[317]), .Y(n14055) );
  sky130_fd_sc_hd__nand2_1 U19269 ( .A(n20282), .B(
        j202_soc_core_j22_cpu_rf_gpr[381]), .Y(n14054) );
  sky130_fd_sc_hd__and4_1 U19270 ( .A(n14057), .B(n14056), .C(n14055), .D(
        n14054), .X(n14066) );
  sky130_fd_sc_hd__nand2_1 U19271 ( .A(n14058), .B(
        j202_soc_core_j22_cpu_rf_gpr[157]), .Y(n14064) );
  sky130_fd_sc_hd__nand2_1 U19272 ( .A(n14059), .B(
        j202_soc_core_j22_cpu_rf_gpr[93]), .Y(n14063) );
  sky130_fd_sc_hd__nand2_1 U19273 ( .A(n20296), .B(
        j202_soc_core_j22_cpu_rf_gpr[125]), .Y(n14062) );
  sky130_fd_sc_hd__nand2_1 U19274 ( .A(n14060), .B(
        j202_soc_core_j22_cpu_rf_gpr[285]), .Y(n14061) );
  sky130_fd_sc_hd__and4_1 U19275 ( .A(n14064), .B(n14063), .C(n14062), .D(
        n14061), .X(n14065) );
  sky130_fd_sc_hd__nand3_1 U19276 ( .A(n14067), .B(n14066), .C(n14065), .Y(
        n19610) );
  sky130_fd_sc_hd__a21oi_1 U19277 ( .A1(n14069), .A2(
        j202_soc_core_j22_cpu_rf_vbr[29]), .B1(n14068), .Y(n14084) );
  sky130_fd_sc_hd__a2bb2oi_1 U19278 ( .B1(j202_soc_core_j22_cpu_rf_gpr[509]), 
        .B2(n14072), .A1_N(n14071), .A2_N(n14070), .Y(n14083) );
  sky130_fd_sc_hd__o22a_1 U19279 ( .A1(n14076), .A2(n14075), .B1(n14074), .B2(
        n14073), .X(n14082) );
  sky130_fd_sc_hd__o22a_1 U19280 ( .A1(n14080), .A2(n14079), .B1(n14078), .B2(
        n14077), .X(n14081) );
  sky130_fd_sc_hd__nand4_1 U19281 ( .A(n14084), .B(n14083), .C(n14082), .D(
        n14081), .Y(n14085) );
  sky130_fd_sc_hd__a21oi_1 U19282 ( .A1(n19610), .A2(n14086), .B1(n14085), .Y(
        n21985) );
  sky130_fd_sc_hd__nand2_1 U19283 ( .A(n21985), .B(n14087), .Y(n14088) );
  sky130_fd_sc_hd__o21ai_1 U19284 ( .A1(n14089), .A2(n21985), .B1(n14088), .Y(
        n14091) );
  sky130_fd_sc_hd__nand2_1 U19285 ( .A(n14091), .B(n14090), .Y(n14395) );
  sky130_fd_sc_hd__nand2_1 U19286 ( .A(n22426), .B(n19729), .Y(n14179) );
  sky130_fd_sc_hd__nor2_1 U19287 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(n14094), .Y(n14841) );
  sky130_fd_sc_hd__nand2_1 U19288 ( .A(n14096), .B(n14095), .Y(n14702) );
  sky130_fd_sc_hd__nor2_1 U19289 ( .A(n14099), .B(n14702), .Y(n14162) );
  sky130_fd_sc_hd__nor2_1 U19290 ( .A(n14412), .B(n14575), .Y(n14147) );
  sky130_fd_sc_hd__nor2_1 U19291 ( .A(n14162), .B(n14147), .Y(n14158) );
  sky130_fd_sc_hd__nand2_1 U19292 ( .A(n17533), .B(n14723), .Y(n14705) );
  sky130_fd_sc_hd__nand2_1 U19293 ( .A(n14158), .B(n14705), .Y(n14406) );
  sky130_fd_sc_hd__nand2_1 U19294 ( .A(n15016), .B(n14100), .Y(n14118) );
  sky130_fd_sc_hd__nor2_1 U19295 ( .A(n14097), .B(n14118), .Y(n14154) );
  sky130_fd_sc_hd__nor2_1 U19296 ( .A(j202_soc_core_bootrom_00_address_w[4]), 
        .B(n14702), .Y(n14738) );
  sky130_fd_sc_hd__nand2_1 U19297 ( .A(n14738), .B(
        j202_soc_core_bootrom_00_address_w[2]), .Y(n14446) );
  sky130_fd_sc_hd__nor2_1 U19298 ( .A(n14154), .B(n14401), .Y(n14488) );
  sky130_fd_sc_hd__nand2_1 U19299 ( .A(n17533), .B(n14404), .Y(n14678) );
  sky130_fd_sc_hd__nand2_1 U19300 ( .A(n18248), .B(n14999), .Y(n14838) );
  sky130_fd_sc_hd__nand2b_1 U19301 ( .A_N(n17970), .B(
        j202_soc_core_bootrom_00_address_w[3]), .Y(n14854) );
  sky130_fd_sc_hd__nor2b_1 U19302 ( .B_N(n14838), .A(n14861), .Y(n14774) );
  sky130_fd_sc_hd__nand2_1 U19303 ( .A(n14678), .B(n14774), .Y(n14727) );
  sky130_fd_sc_hd__nand3_1 U19304 ( .A(n14473), .B(n14098), .C(n15016), .Y(
        n14876) );
  sky130_fd_sc_hd__nor2_1 U19305 ( .A(n14100), .B(n14099), .Y(n14112) );
  sky130_fd_sc_hd__nor2b_1 U19306 ( .B_N(n14112), .A(n14120), .Y(n14822) );
  sky130_fd_sc_hd__nor2_1 U19307 ( .A(n14490), .B(n14822), .Y(n14773) );
  sky130_fd_sc_hd__nor2_1 U19308 ( .A(n14101), .B(n14702), .Y(n14157) );
  sky130_fd_sc_hd__nand2_1 U19309 ( .A(n14977), .B(n14102), .Y(n14837) );
  sky130_fd_sc_hd__nor2_1 U19310 ( .A(n14157), .B(n14117), .Y(n14711) );
  sky130_fd_sc_hd__nor2_1 U19311 ( .A(n14103), .B(n15009), .Y(n14881) );
  sky130_fd_sc_hd__nand3_1 U19312 ( .A(n14773), .B(n14711), .C(n14782), .Y(
        n14105) );
  sky130_fd_sc_hd__nor2_1 U19313 ( .A(n14727), .B(n14105), .Y(n14483) );
  sky130_fd_sc_hd__nor2_1 U19314 ( .A(j202_soc_core_bootrom_00_address_w[3]), 
        .B(n14155), .Y(n14448) );
  sky130_fd_sc_hd__nand4b_1 U19315 ( .A_N(n14406), .B(n14488), .C(n14483), .D(
        n14416), .Y(n14107) );
  sky130_fd_sc_hd__nor2_1 U19316 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(j202_soc_core_bootrom_00_address_w[5]), .Y(n14720) );
  sky130_fd_sc_hd__nand2_1 U19317 ( .A(n14724), .B(n14404), .Y(n14875) );
  sky130_fd_sc_hd__nand2_1 U19318 ( .A(n14777), .B(n14875), .Y(n14455) );
  sky130_fd_sc_hd__nand2_1 U19319 ( .A(n17604), .B(
        j202_soc_core_bootrom_00_address_w[7]), .Y(n14839) );
  sky130_fd_sc_hd__nand2b_1 U19320 ( .A_N(n14455), .B(n14839), .Y(n14737) );
  sky130_fd_sc_hd__nand2_1 U19321 ( .A(n14447), .B(
        j202_soc_core_bootrom_00_address_w[3]), .Y(n14874) );
  sky130_fd_sc_hd__nand2_1 U19322 ( .A(n14811), .B(n14874), .Y(n14767) );
  sky130_fd_sc_hd__nor2_1 U19323 ( .A(n14113), .B(n14118), .Y(n14415) );
  sky130_fd_sc_hd__nand2_1 U19324 ( .A(n17777), .B(n14104), .Y(n14146) );
  sky130_fd_sc_hd__nor2_1 U19325 ( .A(n14415), .B(n14417), .Y(n14495) );
  sky130_fd_sc_hd__or4b_2 U19326 ( .A(n14737), .B(n14767), .C(n14105), .D_N(
        n14495), .X(n14106) );
  sky130_fd_sc_hd__a22oi_1 U19327 ( .A1(n14841), .A2(n14107), .B1(n14720), 
        .B2(n14106), .Y(n14116) );
  sky130_fd_sc_hd__nand2_1 U19328 ( .A(n14977), .B(n14571), .Y(n14810) );
  sky130_fd_sc_hd__o211ai_1 U19329 ( .A1(n14108), .A2(n17442), .B1(n14810), 
        .C1(n14146), .Y(n14695) );
  sky130_fd_sc_hd__nand2_1 U19330 ( .A(n14990), .B(n14723), .Y(n14464) );
  sky130_fd_sc_hd__nand2_1 U19331 ( .A(n14778), .B(n14464), .Y(n14478) );
  sky130_fd_sc_hd__nand2_1 U19332 ( .A(n14119), .B(n14851), .Y(n14808) );
  sky130_fd_sc_hd__nand3_1 U19333 ( .A(n14494), .B(n14808), .C(n14839), .Y(
        n14833) );
  sky130_fd_sc_hd__nor2_1 U19334 ( .A(n14833), .B(n14727), .Y(n14465) );
  sky130_fd_sc_hd__nor2_1 U19335 ( .A(n14117), .B(n14406), .Y(n14829) );
  sky130_fd_sc_hd__nor2_1 U19336 ( .A(n14981), .B(n14296), .Y(n14477) );
  sky130_fd_sc_hd__nand2_1 U19337 ( .A(n14112), .B(n14456), .Y(n14148) );
  sky130_fd_sc_hd__nor2_1 U19338 ( .A(j202_soc_core_bootrom_00_address_w[10]), 
        .B(n14148), .Y(n14696) );
  sky130_fd_sc_hd__nor2_1 U19339 ( .A(n14477), .B(n14696), .Y(n14684) );
  sky130_fd_sc_hd__nand4_1 U19340 ( .A(n14465), .B(n14829), .C(n14684), .D(
        n14446), .Y(n14109) );
  sky130_fd_sc_hd__nor2_1 U19341 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .B(n14998), .Y(n14866) );
  sky130_fd_sc_hd__o21ai_1 U19342 ( .A1(n14478), .A2(n14109), .B1(n14866), .Y(
        n14115) );
  sky130_fd_sc_hd__nor2_1 U19343 ( .A(n17442), .B(n14110), .Y(n14880) );
  sky130_fd_sc_hd__nor2_1 U19344 ( .A(j202_soc_core_bootrom_00_address_w[3]), 
        .B(n14111), .Y(n14852) );
  sky130_fd_sc_hd__nor2_1 U19345 ( .A(n14852), .B(n14112), .Y(n14459) );
  sky130_fd_sc_hd__nor2_1 U19346 ( .A(n14459), .B(n14113), .Y(n14408) );
  sky130_fd_sc_hd__a21oi_1 U19347 ( .A1(n14723), .A2(n14724), .B1(n14408), .Y(
        n14450) );
  sky130_fd_sc_hd__nand2_1 U19348 ( .A(n14990), .B(n14314), .Y(n14419) );
  sky130_fd_sc_hd__nor2_1 U19349 ( .A(n14822), .B(n14422), .Y(n14144) );
  sky130_fd_sc_hd__nand2b_1 U19350 ( .A_N(n14120), .B(n14852), .Y(n14475) );
  sky130_fd_sc_hd__nand3_1 U19351 ( .A(n14450), .B(n14144), .C(n14475), .Y(
        n14703) );
  sky130_fd_sc_hd__nand2_1 U19352 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .B(j202_soc_core_bootrom_00_address_w[6]), .Y(n14815) );
  sky130_fd_sc_hd__o21ai_1 U19353 ( .A1(n14880), .A2(n14703), .B1(n14888), .Y(
        n14114) );
  sky130_fd_sc_hd__a31oi_1 U19354 ( .A1(n14116), .A2(n14115), .A3(n14114), 
        .B1(n18720), .Y(n14173) );
  sky130_fd_sc_hd__nor2_1 U19355 ( .A(n14417), .B(n14117), .Y(n14706) );
  sky130_fd_sc_hd__nor2_1 U19356 ( .A(n14120), .B(n14118), .Y(n14142) );
  sky130_fd_sc_hd__nand2_1 U19357 ( .A(n14706), .B(n14679), .Y(n14156) );
  sky130_fd_sc_hd__a21oi_1 U19358 ( .A1(n17469), .A2(n14399), .B1(n14142), .Y(
        n14454) );
  sky130_fd_sc_hd__nand2_1 U19359 ( .A(n14119), .B(n14852), .Y(n14474) );
  sky130_fd_sc_hd__nor2b_1 U19360 ( .B_N(n14851), .A(n14120), .Y(n14860) );
  sky130_fd_sc_hd__nand2_1 U19361 ( .A(n14474), .B(n14433), .Y(n14693) );
  sky130_fd_sc_hd__nor2_1 U19362 ( .A(n14880), .B(n14415), .Y(n14864) );
  sky130_fd_sc_hd__nand2b_1 U19363 ( .A_N(n14693), .B(n14864), .Y(n14428) );
  sky130_fd_sc_hd__nand2_1 U19364 ( .A(n14808), .B(n14837), .Y(n14766) );
  sky130_fd_sc_hd__nor2_1 U19365 ( .A(n14428), .B(n14766), .Y(n14739) );
  sky130_fd_sc_hd__o22ai_1 U19366 ( .A1(n14454), .A2(n14815), .B1(n14739), 
        .B2(n14871), .Y(n14121) );
  sky130_fd_sc_hd__a21oi_1 U19367 ( .A1(n14866), .A2(n14156), .B1(n14121), .Y(
        n14123) );
  sky130_fd_sc_hd__nand2_1 U19368 ( .A(n14475), .B(n14837), .Y(n14780) );
  sky130_fd_sc_hd__nand2_1 U19369 ( .A(n14476), .B(n14781), .Y(n14687) );
  sky130_fd_sc_hd__o21ai_1 U19370 ( .A1(n14780), .A2(n14687), .B1(n14841), .Y(
        n14122) );
  sky130_fd_sc_hd__a21oi_1 U19371 ( .A1(n14123), .A2(n14122), .B1(n18666), .Y(
        n14172) );
  sky130_fd_sc_hd__a22oi_1 U19372 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[255]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[223]), .Y(n14127) );
  sky130_fd_sc_hd__a22oi_1 U19373 ( .A1(n18734), .A2(
        j202_soc_core_memory0_ram_dout0[159]), .B1(n18733), .B2(
        j202_soc_core_memory0_ram_dout0[127]), .Y(n14126) );
  sky130_fd_sc_hd__a22oi_1 U19374 ( .A1(n18361), .A2(
        j202_soc_core_memory0_ram_dout0[63]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[95]), .Y(n14125) );
  sky130_fd_sc_hd__nand2_1 U19375 ( .A(n18735), .B(
        j202_soc_core_memory0_ram_dout0[191]), .Y(n14124) );
  sky130_fd_sc_hd__nand4_1 U19376 ( .A(n14127), .B(n14126), .C(n14125), .D(
        n14124), .Y(n14128) );
  sky130_fd_sc_hd__a21oi_1 U19377 ( .A1(n18367), .A2(
        j202_soc_core_memory0_ram_dout0[31]), .B1(n14128), .Y(n14136) );
  sky130_fd_sc_hd__a22oi_1 U19378 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[319]), .B1(n18062), .B2(
        j202_soc_core_memory0_ram_dout0[287]), .Y(n14135) );
  sky130_fd_sc_hd__nand2_1 U19379 ( .A(n18743), .B(
        j202_soc_core_memory0_ram_dout0[383]), .Y(n14132) );
  sky130_fd_sc_hd__a21oi_1 U19380 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[479]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n14131) );
  sky130_fd_sc_hd__nand2_1 U19381 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[415]), .Y(n14130) );
  sky130_fd_sc_hd__nand2_1 U19382 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[447]), .Y(n14129) );
  sky130_fd_sc_hd__nand4_1 U19383 ( .A(n14132), .B(n14131), .C(n14130), .D(
        n14129), .Y(n14133) );
  sky130_fd_sc_hd__a21oi_1 U19384 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[351]), .B1(n14133), .Y(n14134) );
  sky130_fd_sc_hd__o211ai_1 U19385 ( .A1(n18736), .A2(n14136), .B1(n14135), 
        .C1(n14134), .Y(n14137) );
  sky130_fd_sc_hd__a22oi_1 U19387 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[31]), .B1(n18379), .B2(
        j202_soc_core_uart_div0[7]), .Y(n14139) );
  sky130_fd_sc_hd__a22oi_1 U19388 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[95]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[63]), .Y(n14138) );
  sky130_fd_sc_hd__o211ai_1 U19389 ( .A1(n18761), .A2(n14140), .B1(n14139), 
        .C1(n14138), .Y(n14171) );
  sky130_fd_sc_hd__nand2_1 U19390 ( .A(n14782), .B(n14419), .Y(n14485) );
  sky130_fd_sc_hd__nand2_1 U19391 ( .A(n17469), .B(n14141), .Y(n14414) );
  sky130_fd_sc_hd__nor2_1 U19392 ( .A(n14142), .B(n14784), .Y(n14482) );
  sky130_fd_sc_hd__nand3b_1 U19393 ( .A_N(n14780), .B(n14774), .C(n14482), .Y(
        n14143) );
  sky130_fd_sc_hd__nand2_1 U19395 ( .A(n14414), .B(n14874), .Y(n14486) );
  sky130_fd_sc_hd__nand3_1 U19396 ( .A(n14462), .B(n14144), .C(n14839), .Y(
        n14858) );
  sky130_fd_sc_hd__nor3_1 U19397 ( .A(n14772), .B(n14727), .C(n14858), .Y(
        n14690) );
  sky130_fd_sc_hd__a31oi_1 U19398 ( .A1(n14495), .A2(n14690), .A3(n14474), 
        .B1(n14882), .Y(n14153) );
  sky130_fd_sc_hd__nor2_1 U19399 ( .A(n14448), .B(n14477), .Y(n14403) );
  sky130_fd_sc_hd__a31oi_1 U19400 ( .A1(n14864), .A2(n14145), .A3(n14874), 
        .B1(n14815), .Y(n14152) );
  sky130_fd_sc_hd__nor3_1 U19401 ( .A(n14861), .B(n14822), .C(n14833), .Y(
        n14421) );
  sky130_fd_sc_hd__nand2b_1 U19402 ( .A_N(n14485), .B(n14421), .Y(n14430) );
  sky130_fd_sc_hd__nor4_1 U19403 ( .A(n14490), .B(n14447), .C(n14738), .D(
        n14430), .Y(n14150) );
  sky130_fd_sc_hd__nand2_1 U19404 ( .A(n14146), .B(n14705), .Y(n14429) );
  sky130_fd_sc_hd__nor2_1 U19405 ( .A(n14422), .B(n14147), .Y(n14484) );
  sky130_fd_sc_hd__nand2_1 U19406 ( .A(n14484), .B(n14494), .Y(n14434) );
  sky130_fd_sc_hd__nand4_1 U19407 ( .A(n14148), .B(n14838), .C(n14475), .D(
        n14403), .Y(n14849) );
  sky130_fd_sc_hd__nor4_1 U19408 ( .A(n14881), .B(n14429), .C(n14434), .D(
        n14849), .Y(n14149) );
  sky130_fd_sc_hd__o22ai_1 U19409 ( .A1(n14150), .A2(n14884), .B1(n14149), 
        .B2(n14871), .Y(n14151) );
  sky130_fd_sc_hd__nor4b_1 U19410 ( .D_N(n14689), .A(n14153), .B(n14152), .C(
        n14151), .Y(n14169) );
  sky130_fd_sc_hd__nor2_1 U19411 ( .A(n14880), .B(n14162), .Y(n14776) );
  sky130_fd_sc_hd__nand2_1 U19412 ( .A(n14776), .B(n14782), .Y(n14821) );
  sky130_fd_sc_hd__nor2_1 U19413 ( .A(n14821), .B(n14458), .Y(n14423) );
  sky130_fd_sc_hd__o31a_1 U19415 ( .A1(n14444), .A2(n14835), .A3(n14154), .B1(
        n14841), .X(n14167) );
  sky130_fd_sc_hd__nor2_1 U19416 ( .A(n14477), .B(n14860), .Y(n14717) );
  sky130_fd_sc_hd__a31oi_1 U19417 ( .A1(n14778), .A2(n14717), .A3(n14155), 
        .B1(n14882), .Y(n14166) );
  sky130_fd_sc_hd__nand2_1 U19418 ( .A(n14875), .B(n14808), .Y(n14445) );
  sky130_fd_sc_hd__nor2_1 U19419 ( .A(n14157), .B(n14861), .Y(n14402) );
  sky130_fd_sc_hd__nand2_1 U19420 ( .A(n14402), .B(n14416), .Y(n14843) );
  sky130_fd_sc_hd__nor4b_1 U19421 ( .D_N(n14158), .A(n14784), .B(n14445), .C(
        n14843), .Y(n14159) );
  sky130_fd_sc_hd__a21oi_1 U19422 ( .A1(n14160), .A2(n14159), .B1(n14815), .Y(
        n14165) );
  sky130_fd_sc_hd__nand2_1 U19423 ( .A(n17533), .B(n14982), .Y(n17912) );
  sky130_fd_sc_hd__nor2_1 U19424 ( .A(n17442), .B(n14161), .Y(n14809) );
  sky130_fd_sc_hd__nor2_1 U19425 ( .A(n14680), .B(n14809), .Y(n14431) );
  sky130_fd_sc_hd__nand3_1 U19426 ( .A(n14476), .B(n14414), .C(n14431), .Y(
        n14400) );
  sky130_fd_sc_hd__nor4_1 U19427 ( .A(n14162), .B(n14415), .C(n17498), .D(
        n14400), .Y(n14163) );
  sky130_fd_sc_hd__a21oi_1 U19428 ( .A1(n14451), .A2(n14163), .B1(n14871), .Y(
        n14164) );
  sky130_fd_sc_hd__nor4_1 U19429 ( .A(n14167), .B(n14166), .C(n14165), .D(
        n14164), .Y(n14168) );
  sky130_fd_sc_hd__o22ai_1 U19430 ( .A1(n14169), .A2(n18722), .B1(n14168), 
        .B2(n18552), .Y(n14170) );
  sky130_fd_sc_hd__a22oi_1 U19431 ( .A1(n19657), .A2(n22591), .B1(n19736), 
        .B2(n23344), .Y(n14174) );
  sky130_fd_sc_hd__o21a_1 U19432 ( .A1(n14919), .A2(n22542), .B1(n14174), .X(
        n14178) );
  sky130_fd_sc_hd__ha_1 U19433 ( .A(j202_soc_core_j22_cpu_pc[24]), .B(n14175), 
        .COUT(n14276), .SUM(n21842) );
  sky130_fd_sc_hd__xor2_1 U19434 ( .A(n14176), .B(j202_soc_core_j22_cpu_pc[31]), .X(n22362) );
  sky130_fd_sc_hd__nand2_1 U19435 ( .A(n22362), .B(n19661), .Y(n14177) );
  sky130_fd_sc_hd__nand3_1 U19436 ( .A(n14179), .B(n14178), .C(n14177), .Y(
        n14965) );
  sky130_fd_sc_hd__nand2_1 U19437 ( .A(n11185), .B(n14180), .Y(n14182) );
  sky130_fd_sc_hd__xnor2_1 U19438 ( .A(n14182), .B(n14181), .Y(n21952) );
  sky130_fd_sc_hd__nand2_1 U19439 ( .A(n21952), .B(n19729), .Y(n14272) );
  sky130_fd_sc_hd__ha_1 U19440 ( .A(j202_soc_core_j22_cpu_pc[27]), .B(n14183), 
        .COUT(n14807), .SUM(n21954) );
  sky130_fd_sc_hd__nand4_1 U19441 ( .A(n14187), .B(n14288), .C(n14567), .D(
        n14186), .Y(n14192) );
  sky130_fd_sc_hd__a32oi_1 U19442 ( .A1(n14286), .A2(n14190), .A3(n14189), 
        .B1(n14639), .B2(n14190), .Y(n14191) );
  sky130_fd_sc_hd__a21oi_1 U19443 ( .A1(n14348), .A2(n14192), .B1(n14191), .Y(
        n14193) );
  sky130_fd_sc_hd__nand2b_1 U19444 ( .A_N(n14193), .B(n14308), .Y(n14248) );
  sky130_fd_sc_hd__nor4_1 U19445 ( .A(n14196), .B(n14195), .C(n14204), .D(
        n14194), .Y(n14197) );
  sky130_fd_sc_hd__a21oi_1 U19446 ( .A1(n14198), .A2(n14197), .B1(n15149), .Y(
        n14216) );
  sky130_fd_sc_hd__nor4b_1 U19447 ( .D_N(n14200), .A(n14538), .B(n14598), .C(
        n14199), .Y(n14355) );
  sky130_fd_sc_hd__a21oi_1 U19448 ( .A1(n14201), .A2(n14314), .B1(n14311), .Y(
        n14203) );
  sky130_fd_sc_hd__a31oi_1 U19449 ( .A1(n14355), .A2(n14203), .A3(n14202), 
        .B1(n14639), .Y(n14215) );
  sky130_fd_sc_hd__nor3_1 U19450 ( .A(n14232), .B(n14204), .C(n14354), .Y(
        n14213) );
  sky130_fd_sc_hd__nor2_1 U19451 ( .A(n14999), .B(n14205), .Y(n14238) );
  sky130_fd_sc_hd__nor3_1 U19452 ( .A(n14207), .B(n14206), .C(n14343), .Y(
        n14595) );
  sky130_fd_sc_hd__nand4b_1 U19453 ( .A_N(n14238), .B(n14209), .C(n14208), .D(
        n14595), .Y(n14210) );
  sky130_fd_sc_hd__nor3_1 U19454 ( .A(n14211), .B(n14325), .C(n14210), .Y(
        n14212) );
  sky130_fd_sc_hd__o22ai_1 U19455 ( .A1(n14213), .A2(n14619), .B1(n14212), 
        .B2(n14631), .Y(n14214) );
  sky130_fd_sc_hd__nor3_1 U19456 ( .A(n14216), .B(n14215), .C(n14214), .Y(
        n14226) );
  sky130_fd_sc_hd__a31oi_1 U19457 ( .A1(n14218), .A2(n14574), .A3(n14334), 
        .B1(n14631), .Y(n14224) );
  sky130_fd_sc_hd__a31oi_1 U19458 ( .A1(n14287), .A2(n14279), .A3(n14219), 
        .B1(n15149), .Y(n14223) );
  sky130_fd_sc_hd__a21oi_1 U19459 ( .A1(n14627), .A2(n14288), .B1(n14619), .Y(
        n14222) );
  sky130_fd_sc_hd__nor4_1 U19461 ( .A(n14224), .B(n14223), .C(n14222), .D(
        n14221), .Y(n14225) );
  sky130_fd_sc_hd__o22a_1 U19462 ( .A1(n14562), .A2(n14226), .B1(n14339), .B2(
        n14225), .X(n14247) );
  sky130_fd_sc_hd__a31oi_1 U19463 ( .A1(n14228), .A2(n14227), .A3(n14592), 
        .B1(n14639), .Y(n14243) );
  sky130_fd_sc_hd__nor2_1 U19464 ( .A(n14229), .B(n14238), .Y(n14318) );
  sky130_fd_sc_hd__nor4_1 U19465 ( .A(n14232), .B(n14325), .C(n14231), .D(
        n14230), .Y(n14233) );
  sky130_fd_sc_hd__a21oi_1 U19466 ( .A1(n14318), .A2(n14233), .B1(n15149), .Y(
        n14242) );
  sky130_fd_sc_hd__a21oi_1 U19467 ( .A1(n14236), .A2(n14235), .B1(n14234), .Y(
        n14237) );
  sky130_fd_sc_hd__a21oi_1 U19468 ( .A1(n14345), .A2(n14237), .B1(n14631), .Y(
        n14241) );
  sky130_fd_sc_hd__nor2_1 U19469 ( .A(n14310), .B(n14293), .Y(n14628) );
  sky130_fd_sc_hd__nor4_1 U19470 ( .A(n14598), .B(n14597), .C(n14238), .D(
        n14628), .Y(n14239) );
  sky130_fd_sc_hd__a21oi_1 U19471 ( .A1(n14596), .A2(n14239), .B1(n14619), .Y(
        n14240) );
  sky130_fd_sc_hd__nor4_1 U19472 ( .A(n14243), .B(n14242), .C(n14241), .D(
        n14240), .Y(n14245) );
  sky130_fd_sc_hd__nand2b_1 U19473 ( .A_N(n14245), .B(n14244), .Y(n14246) );
  sky130_fd_sc_hd__nand3_1 U19474 ( .A(n14248), .B(n14247), .C(n14246), .Y(
        n14267) );
  sky130_fd_sc_hd__a22oi_1 U19475 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[251]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[219]), .Y(n14252) );
  sky130_fd_sc_hd__a22oi_1 U19476 ( .A1(n18734), .A2(
        j202_soc_core_memory0_ram_dout0[155]), .B1(n18733), .B2(
        j202_soc_core_memory0_ram_dout0[123]), .Y(n14251) );
  sky130_fd_sc_hd__a22oi_1 U19477 ( .A1(n18361), .A2(
        j202_soc_core_memory0_ram_dout0[59]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[91]), .Y(n14250) );
  sky130_fd_sc_hd__nand2_1 U19478 ( .A(n18735), .B(
        j202_soc_core_memory0_ram_dout0[187]), .Y(n14249) );
  sky130_fd_sc_hd__nand4_1 U19479 ( .A(n14252), .B(n14251), .C(n14250), .D(
        n14249), .Y(n14253) );
  sky130_fd_sc_hd__a32oi_1 U19480 ( .A1(n18367), .A2(n17639), .A3(
        j202_soc_core_memory0_ram_dout0[27]), .B1(n14253), .B2(n17639), .Y(
        n14261) );
  sky130_fd_sc_hd__a22oi_1 U19481 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[315]), .B1(n18062), .B2(
        j202_soc_core_memory0_ram_dout0[283]), .Y(n14260) );
  sky130_fd_sc_hd__nand2_1 U19482 ( .A(n18743), .B(
        j202_soc_core_memory0_ram_dout0[379]), .Y(n14257) );
  sky130_fd_sc_hd__a21oi_1 U19483 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[475]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n14256) );
  sky130_fd_sc_hd__nand2_1 U19484 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[411]), .Y(n14255) );
  sky130_fd_sc_hd__nand2_1 U19485 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[443]), .Y(n14254) );
  sky130_fd_sc_hd__nand4_1 U19486 ( .A(n14257), .B(n14256), .C(n14255), .D(
        n14254), .Y(n14258) );
  sky130_fd_sc_hd__a21oi_1 U19487 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[347]), .B1(n14258), .Y(n14259) );
  sky130_fd_sc_hd__nand3_1 U19488 ( .A(n14261), .B(n14260), .C(n14259), .Y(
        n14262) );
  sky130_fd_sc_hd__o211ai_1 U19489 ( .A1(j202_soc_core_memory0_ram_dout0[507]), 
        .A2(n18758), .B1(n14906), .C1(n14262), .Y(n14265) );
  sky130_fd_sc_hd__a22oi_1 U19490 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[27]), .B1(n18727), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[91]), .Y(n14264) );
  sky130_fd_sc_hd__a22oi_1 U19491 ( .A1(n18726), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[59]), .B1(n18379), .B2(
        j202_soc_core_uart_div0[3]), .Y(n14263) );
  sky130_fd_sc_hd__nand3_1 U19492 ( .A(n14265), .B(n14264), .C(n14263), .Y(
        n14266) );
  sky130_fd_sc_hd__a21oi_1 U19493 ( .A1(n14267), .A2(n14668), .B1(n14266), .Y(
        n22538) );
  sky130_fd_sc_hd__a22oi_1 U19494 ( .A1(n19657), .A2(n22576), .B1(n19736), 
        .B2(n23330), .Y(n14269) );
  sky130_fd_sc_hd__nand2_1 U19495 ( .A(n21954), .B(n19517), .Y(n14268) );
  sky130_fd_sc_hd__o211ai_1 U19496 ( .A1(n22538), .A2(n14919), .B1(n14269), 
        .C1(n14268), .Y(n14270) );
  sky130_fd_sc_hd__a21oi_1 U19497 ( .A1(n19732), .A2(n21954), .B1(n14270), .Y(
        n14271) );
  sky130_fd_sc_hd__nand2_1 U19498 ( .A(n14272), .B(n14271), .Y(n14961) );
  sky130_fd_sc_hd__nand4_1 U19499 ( .A(n25257), .B(n25280), .C(n25252), .D(
        n25277), .Y(n14393) );
  sky130_fd_sc_hd__nand2_1 U19500 ( .A(n11189), .B(n14273), .Y(n14275) );
  sky130_fd_sc_hd__xnor2_1 U19501 ( .A(n14275), .B(n14274), .Y(n21765) );
  sky130_fd_sc_hd__ha_1 U19502 ( .A(j202_soc_core_j22_cpu_pc[25]), .B(n14276), 
        .COUT(n14536), .SUM(n21767) );
  sky130_fd_sc_hd__nand2_1 U19503 ( .A(n21767), .B(n19732), .Y(n14391) );
  sky130_fd_sc_hd__nand2_1 U19504 ( .A(n21767), .B(n19517), .Y(n14390) );
  sky130_fd_sc_hd__a22oi_1 U19505 ( .A1(n19657), .A2(n22574), .B1(n19736), 
        .B2(n23324), .Y(n14389) );
  sky130_fd_sc_hd__nor3b_1 U19506 ( .C_N(n14279), .A(n14278), .B(n14277), .Y(
        n14281) );
  sky130_fd_sc_hd__a21oi_1 U19507 ( .A1(n14281), .A2(n14280), .B1(n14619), .Y(
        n14306) );
  sky130_fd_sc_hd__nor3_1 U19508 ( .A(n14284), .B(n14283), .C(n14282), .Y(
        n14285) );
  sky130_fd_sc_hd__a21oi_1 U19509 ( .A1(n14286), .A2(n14285), .B1(n14631), .Y(
        n14305) );
  sky130_fd_sc_hd__nand3_1 U19510 ( .A(n14289), .B(n14288), .C(n14287), .Y(
        n14290) );
  sky130_fd_sc_hd__nor2_1 U19511 ( .A(n14291), .B(n14290), .Y(n14303) );
  sky130_fd_sc_hd__nor2_1 U19512 ( .A(n14294), .B(n14293), .Y(n14299) );
  sky130_fd_sc_hd__nor4_1 U19514 ( .A(n14300), .B(n14299), .C(n14298), .D(
        n14297), .Y(n14582) );
  sky130_fd_sc_hd__nor2_1 U19515 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(n17778), .Y(n17532) );
  sky130_fd_sc_hd__nand2_1 U19516 ( .A(n17532), .B(
        j202_soc_core_bootrom_00_address_w[9]), .Y(n14301) );
  sky130_fd_sc_hd__and3_1 U19517 ( .A(n14582), .B(n14567), .C(n14301), .X(
        n14302) );
  sky130_fd_sc_hd__o22ai_1 U19518 ( .A1(n14303), .A2(n15149), .B1(n14302), 
        .B2(n14639), .Y(n14304) );
  sky130_fd_sc_hd__nor4_1 U19519 ( .A(n14307), .B(n14306), .C(n14305), .D(
        n14304), .Y(n14366) );
  sky130_fd_sc_hd__nor2_1 U19520 ( .A(n14310), .B(n14309), .Y(n14312) );
  sky130_fd_sc_hd__nor3_1 U19521 ( .A(n14312), .B(n14598), .C(n14311), .Y(
        n14323) );
  sky130_fd_sc_hd__nand2_1 U19522 ( .A(n14314), .B(n14313), .Y(n14316) );
  sky130_fd_sc_hd__nand4_1 U19523 ( .A(n14317), .B(n14323), .C(n14316), .D(
        n14315), .Y(n14321) );
  sky130_fd_sc_hd__a31oi_1 U19524 ( .A1(n14319), .A2(n14593), .A3(n14318), 
        .B1(n15149), .Y(n14320) );
  sky130_fd_sc_hd__a21oi_1 U19525 ( .A1(n14348), .A2(n14321), .B1(n14320), .Y(
        n14329) );
  sky130_fd_sc_hd__o21ai_1 U19526 ( .A1(n14539), .A2(n14322), .B1(n14613), .Y(
        n14328) );
  sky130_fd_sc_hd__o31ai_1 U19527 ( .A1(n14326), .A2(n14325), .A3(n14324), 
        .B1(n14352), .Y(n14327) );
  sky130_fd_sc_hd__a31oi_1 U19528 ( .A1(n14329), .A2(n14328), .A3(n14327), 
        .B1(n14615), .Y(n14364) );
  sky130_fd_sc_hd__nand4_1 U19529 ( .A(n14331), .B(n14627), .C(n14330), .D(
        n14332), .Y(n14336) );
  sky130_fd_sc_hd__a31oi_1 U19530 ( .A1(n14334), .A2(n14333), .A3(n14332), 
        .B1(n14631), .Y(n14335) );
  sky130_fd_sc_hd__a211oi_1 U19531 ( .A1(n14352), .A2(n14336), .B1(n14335), 
        .C1(n14638), .Y(n14341) );
  sky130_fd_sc_hd__o21ai_1 U19532 ( .A1(n14338), .A2(n14623), .B1(n15093), .Y(
        n14340) );
  sky130_fd_sc_hd__a21oi_1 U19533 ( .A1(n14341), .A2(n14340), .B1(n14339), .Y(
        n14363) );
  sky130_fd_sc_hd__nand4b_1 U19534 ( .A_N(n14343), .B(n14351), .C(n14350), .D(
        n14342), .Y(n14347) );
  sky130_fd_sc_hd__a31oi_1 U19535 ( .A1(n14345), .A2(n14344), .A3(n14592), 
        .B1(n15149), .Y(n14346) );
  sky130_fd_sc_hd__a21oi_1 U19536 ( .A1(n14348), .A2(n14347), .B1(n14346), .Y(
        n14361) );
  sky130_fd_sc_hd__nor3b_1 U19537 ( .C_N(n14349), .A(n14539), .B(n14598), .Y(
        n14547) );
  sky130_fd_sc_hd__nand4_1 U19538 ( .A(n14351), .B(n14552), .C(n14547), .D(
        n14350), .Y(n14353) );
  sky130_fd_sc_hd__o31ai_1 U19540 ( .A1(n14358), .A2(n14357), .A3(n14356), 
        .B1(n14613), .Y(n14359) );
  sky130_fd_sc_hd__a31oi_1 U19541 ( .A1(n14361), .A2(n14360), .A3(n14359), 
        .B1(n14562), .Y(n14362) );
  sky130_fd_sc_hd__nor3_1 U19542 ( .A(n14364), .B(n14363), .C(n14362), .Y(
        n14365) );
  sky130_fd_sc_hd__nand2_1 U19544 ( .A(n14367), .B(n14668), .Y(n14387) );
  sky130_fd_sc_hd__a22oi_1 U19545 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[89]), .B1(n18725), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[25]), .Y(n14369) );
  sky130_fd_sc_hd__a22oi_1 U19546 ( .A1(n18726), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[57]), .B1(n18379), .B2(
        j202_soc_core_uart_div0[1]), .Y(n14368) );
  sky130_fd_sc_hd__and2_0 U19547 ( .A(n14369), .B(n14368), .X(n14386) );
  sky130_fd_sc_hd__a22oi_1 U19548 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[281]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[57]), .Y(n14383) );
  sky130_fd_sc_hd__a22o_1 U19549 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[313]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[345]), .X(n14370) );
  sky130_fd_sc_hd__a21oi_1 U19550 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[377]), .B1(n14370), .Y(n14382) );
  sky130_fd_sc_hd__nand2_1 U19551 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[249]), .Y(n14374) );
  sky130_fd_sc_hd__a21oi_1 U19552 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[473]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n14373) );
  sky130_fd_sc_hd__nand2_1 U19553 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[409]), .Y(n14372) );
  sky130_fd_sc_hd__nand2_1 U19554 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[441]), .Y(n14371) );
  sky130_fd_sc_hd__nand4_1 U19555 ( .A(n14374), .B(n14373), .C(n14372), .D(
        n14371), .Y(n14375) );
  sky130_fd_sc_hd__a21oi_1 U19556 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[217]), .B1(n14375), .Y(n14381) );
  sky130_fd_sc_hd__a22o_1 U19557 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[25]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[89]), .X(n14376) );
  sky130_fd_sc_hd__a21oi_1 U19558 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[121]), .B1(n14376), .Y(n14378) );
  sky130_fd_sc_hd__a22oi_1 U19559 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[185]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[153]), .Y(n14377) );
  sky130_fd_sc_hd__nand2_1 U19560 ( .A(n14378), .B(n14377), .Y(n14379) );
  sky130_fd_sc_hd__nand2_1 U19561 ( .A(n14379), .B(n17639), .Y(n14380) );
  sky130_fd_sc_hd__nand4_1 U19562 ( .A(n14383), .B(n14382), .C(n14381), .D(
        n14380), .Y(n14384) );
  sky130_fd_sc_hd__o211ai_1 U19563 ( .A1(j202_soc_core_memory0_ram_dout0[505]), 
        .A2(n18758), .B1(n14906), .C1(n14384), .Y(n14385) );
  sky130_fd_sc_hd__nand3_1 U19564 ( .A(n14387), .B(n14386), .C(n14385), .Y(
        n22541) );
  sky130_fd_sc_hd__nand2_1 U19565 ( .A(n22541), .B(n19737), .Y(n14388) );
  sky130_fd_sc_hd__nand4_1 U19566 ( .A(n14391), .B(n14390), .C(n14389), .D(
        n14388), .Y(n14392) );
  sky130_fd_sc_hd__a21oi_1 U19567 ( .A1(n21765), .A2(n19729), .B1(n14392), .Y(
        n14963) );
  sky130_fd_sc_hd__nor2_1 U19568 ( .A(n14393), .B(n14963), .Y(n14394) );
  sky130_fd_sc_hd__nand2_1 U19569 ( .A(n11194), .B(n14395), .Y(n14397) );
  sky130_fd_sc_hd__xnor2_1 U19570 ( .A(n14397), .B(n14396), .Y(n21984) );
  sky130_fd_sc_hd__nand2_1 U19571 ( .A(n21984), .B(n19729), .Y(n14529) );
  sky130_fd_sc_hd__ha_1 U19572 ( .A(j202_soc_core_j22_cpu_pc[29]), .B(n14398), 
        .COUT(n14795), .SUM(n21987) );
  sky130_fd_sc_hd__o22a_1 U19573 ( .A1(n21985), .A2(n18948), .B1(n21048), .B2(
        n19731), .X(n14525) );
  sky130_fd_sc_hd__nand2_1 U19574 ( .A(n14977), .B(n14399), .Y(n14685) );
  sky130_fd_sc_hd__nor3b_1 U19575 ( .C_N(n14685), .A(n14400), .B(n14737), .Y(
        n14731) );
  sky130_fd_sc_hd__nand2_1 U19576 ( .A(n14874), .B(n14838), .Y(n14452) );
  sky130_fd_sc_hd__nor2_1 U19577 ( .A(n14401), .B(n14452), .Y(n14817) );
  sky130_fd_sc_hd__nand4_1 U19578 ( .A(n14731), .B(n14403), .C(n14402), .D(
        n14817), .Y(n14411) );
  sky130_fd_sc_hd__nand2_1 U19579 ( .A(n14481), .B(n14810), .Y(n14405) );
  sky130_fd_sc_hd__nand2_1 U19580 ( .A(n14990), .B(n14404), .Y(n14862) );
  sky130_fd_sc_hd__nand2_1 U19581 ( .A(n14872), .B(n14862), .Y(n14812) );
  sky130_fd_sc_hd__nor2_1 U19582 ( .A(n14405), .B(n14812), .Y(n14691) );
  sky130_fd_sc_hd__nand2_1 U19583 ( .A(n14464), .B(n14495), .Y(n14487) );
  sky130_fd_sc_hd__nor2_1 U19584 ( .A(n14406), .B(n14487), .Y(n14407) );
  sky130_fd_sc_hd__nand4_1 U19585 ( .A(n14691), .B(n14421), .C(n14407), .D(
        n14433), .Y(n14715) );
  sky130_fd_sc_hd__nand2_1 U19586 ( .A(n14678), .B(n14475), .Y(n14832) );
  sky130_fd_sc_hd__nor2_1 U19587 ( .A(n14408), .B(n14832), .Y(n14770) );
  sky130_fd_sc_hd__nand2_1 U19588 ( .A(n14876), .B(n14679), .Y(n14479) );
  sky130_fd_sc_hd__nor2b_1 U19589 ( .B_N(n14488), .A(n14479), .Y(n14840) );
  sky130_fd_sc_hd__a31oi_1 U19590 ( .A1(n14409), .A2(n14770), .A3(n14840), 
        .B1(n14871), .Y(n14410) );
  sky130_fd_sc_hd__a21oi_1 U19591 ( .A1(n14841), .A2(n14411), .B1(n14410), .Y(
        n14427) );
  sky130_fd_sc_hd__nand4_1 U19592 ( .A(n14782), .B(n14702), .C(n14839), .D(
        n14464), .Y(n14887) );
  sky130_fd_sc_hd__nor2_1 U19593 ( .A(n14413), .B(n14412), .Y(n14865) );
  sky130_fd_sc_hd__nand2_1 U19594 ( .A(n14414), .B(n14810), .Y(n14453) );
  sky130_fd_sc_hd__nor2_1 U19595 ( .A(n14415), .B(n14490), .Y(n14692) );
  sky130_fd_sc_hd__nand3_1 U19596 ( .A(n14692), .B(n14416), .C(n14476), .Y(
        n14694) );
  sky130_fd_sc_hd__nor4_1 U19597 ( .A(n14417), .B(n14865), .C(n14453), .D(
        n14694), .Y(n14418) );
  sky130_fd_sc_hd__nand2b_1 U19598 ( .A_N(n14696), .B(n14418), .Y(n14730) );
  sky130_fd_sc_hd__nand4b_1 U19599 ( .A_N(n14730), .B(n14419), .C(n14838), .D(
        n14678), .Y(n14420) );
  sky130_fd_sc_hd__o21ai_1 U19600 ( .A1(n14887), .A2(n14420), .B1(n14888), .Y(
        n14426) );
  sky130_fd_sc_hd__nand2_1 U19601 ( .A(n14462), .B(n14421), .Y(n14721) );
  sky130_fd_sc_hd__nor2_1 U19602 ( .A(n14455), .B(n14479), .Y(n14718) );
  sky130_fd_sc_hd__nor2b_1 U19603 ( .B_N(n14718), .A(n14694), .Y(n14432) );
  sky130_fd_sc_hd__nor2_1 U19604 ( .A(n14422), .B(n14738), .Y(n14885) );
  sky130_fd_sc_hd__nand4_1 U19605 ( .A(n14432), .B(n14423), .C(n14885), .D(
        n14872), .Y(n14424) );
  sky130_fd_sc_hd__nand3_1 U19607 ( .A(n14427), .B(n14426), .C(n14425), .Y(
        n14443) );
  sky130_fd_sc_hd__nor4_1 U19608 ( .A(n14477), .B(n14430), .C(n14429), .D(
        n14428), .Y(n14441) );
  sky130_fd_sc_hd__nand2_1 U19609 ( .A(n14808), .B(n14838), .Y(n14859) );
  sky130_fd_sc_hd__nor4b_1 U19610 ( .D_N(n14431), .A(n14444), .B(n14737), .C(
        n14859), .Y(n14439) );
  sky130_fd_sc_hd__nand3_1 U19611 ( .A(n14432), .B(n14431), .C(n14854), .Y(
        n14437) );
  sky130_fd_sc_hd__nand2_1 U19612 ( .A(n14839), .B(n14433), .Y(n14728) );
  sky130_fd_sc_hd__nor3_1 U19613 ( .A(n14478), .B(n14728), .C(n14434), .Y(
        n14435) );
  sky130_fd_sc_hd__nand3_1 U19614 ( .A(n14435), .B(n14692), .C(n14874), .Y(
        n14436) );
  sky130_fd_sc_hd__a22oi_1 U19615 ( .A1(n14437), .A2(n14841), .B1(n14436), 
        .B2(n14720), .Y(n14438) );
  sky130_fd_sc_hd__o21a_1 U19616 ( .A1(n14815), .A2(n14439), .B1(n14438), .X(
        n14440) );
  sky130_fd_sc_hd__a22oi_1 U19618 ( .A1(n14443), .A2(n18610), .B1(n14442), 
        .B2(n17609), .Y(n14523) );
  sky130_fd_sc_hd__nor2_1 U19619 ( .A(n14809), .B(n14860), .Y(n14830) );
  sky130_fd_sc_hd__or4b_2 U19620 ( .A(n14445), .B(n14444), .C(n14479), .D_N(
        n14830), .X(n14470) );
  sky130_fd_sc_hd__nand2_1 U19621 ( .A(n14839), .B(n14446), .Y(n14879) );
  sky130_fd_sc_hd__nand2b_1 U19622 ( .A_N(n14879), .B(n14862), .Y(n14771) );
  sky130_fd_sc_hd__nor4_1 U19623 ( .A(n14448), .B(n14447), .C(n14822), .D(
        n14771), .Y(n14449) );
  sky130_fd_sc_hd__a31oi_1 U19624 ( .A1(n14451), .A2(n14450), .A3(n14449), 
        .B1(n14815), .Y(n14469) );
  sky130_fd_sc_hd__nand2_1 U19625 ( .A(n14811), .B(n14464), .Y(n14719) );
  sky130_fd_sc_hd__nor3_1 U19626 ( .A(n14453), .B(n14452), .C(n14719), .Y(
        n14707) );
  sky130_fd_sc_hd__nand2_1 U19627 ( .A(n14488), .B(n14454), .Y(n14736) );
  sky130_fd_sc_hd__nor4b_1 U19628 ( .D_N(n14707), .A(n14455), .B(n14693), .C(
        n14736), .Y(n14467) );
  sky130_fd_sc_hd__a211oi_1 U19629 ( .A1(n14850), .A2(n15016), .B1(n14458), 
        .C1(n14457), .Y(n14682) );
  sky130_fd_sc_hd__a21oi_1 U19630 ( .A1(n14850), .A2(n14460), .B1(n17785), .Y(
        n14461) );
  sky130_fd_sc_hd__nand4_1 U19631 ( .A(n14462), .B(n14682), .C(n14461), .D(
        n14476), .Y(n14463) );
  sky130_fd_sc_hd__and4b_1 U19632 ( .B(n14465), .C(n14484), .D(n14464), .A_N(
        n14463), .X(n14466) );
  sky130_fd_sc_hd__o22ai_1 U19633 ( .A1(n14467), .A2(n14884), .B1(n14466), 
        .B2(n14871), .Y(n14468) );
  sky130_fd_sc_hd__a211oi_1 U19634 ( .A1(n14866), .A2(n14470), .B1(n14469), 
        .C1(n14468), .Y(n14471) );
  sky130_fd_sc_hd__nand2b_1 U19635 ( .A_N(n14471), .B(n18605), .Y(n14522) );
  sky130_fd_sc_hd__nand3_1 U19636 ( .A(n14473), .B(
        j202_soc_core_bootrom_00_address_w[10]), .C(n14472), .Y(n17672) );
  sky130_fd_sc_hd__nand2_1 U19637 ( .A(n14474), .B(n17672), .Y(n14489) );
  sky130_fd_sc_hd__nor2_1 U19638 ( .A(n14696), .B(n14489), .Y(n14824) );
  sky130_fd_sc_hd__nand4_1 U19639 ( .A(n14824), .B(n14476), .C(n14875), .D(
        n14475), .Y(n14497) );
  sky130_fd_sc_hd__or4_1 U19640 ( .A(n14479), .B(n14478), .C(n14858), .D(
        n14477), .X(n14480) );
  sky130_fd_sc_hd__o21ai_1 U19641 ( .A1(n14497), .A2(n14480), .B1(n14841), .Y(
        n14500) );
  sky130_fd_sc_hd__nand4_1 U19642 ( .A(n14484), .B(n14483), .C(n14482), .D(
        n14481), .Y(n14493) );
  sky130_fd_sc_hd__nor2_1 U19643 ( .A(n14486), .B(n14485), .Y(n14742) );
  sky130_fd_sc_hd__nor2_1 U19644 ( .A(n14487), .B(n14812), .Y(n14836) );
  sky130_fd_sc_hd__nand2_1 U19645 ( .A(n14488), .B(n14836), .Y(n14783) );
  sky130_fd_sc_hd__nor4_1 U19646 ( .A(n14490), .B(n14814), .C(n14489), .D(
        n14783), .Y(n14491) );
  sky130_fd_sc_hd__a21oi_1 U19647 ( .A1(n14742), .A2(n14491), .B1(n14871), .Y(
        n14492) );
  sky130_fd_sc_hd__a21oi_1 U19648 ( .A1(n14866), .A2(n14493), .B1(n14492), .Y(
        n14499) );
  sky130_fd_sc_hd__nor2_1 U19649 ( .A(n14881), .B(n14768), .Y(n14726) );
  sky130_fd_sc_hd__nand4_1 U19650 ( .A(n14495), .B(n14707), .C(n14726), .D(
        n14494), .Y(n14496) );
  sky130_fd_sc_hd__nand3_1 U19652 ( .A(n14500), .B(n14499), .C(n14498), .Y(
        n14520) );
  sky130_fd_sc_hd__a22oi_1 U19653 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[29]), .B1(n18379), .B2(
        j202_soc_core_uart_div0[5]), .Y(n14502) );
  sky130_fd_sc_hd__a22oi_1 U19654 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[93]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[61]), .Y(n14501) );
  sky130_fd_sc_hd__nand2_1 U19655 ( .A(n14502), .B(n14501), .Y(n14518) );
  sky130_fd_sc_hd__a22oi_1 U19656 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[253]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[221]), .Y(n14506) );
  sky130_fd_sc_hd__a22oi_1 U19657 ( .A1(n18734), .A2(
        j202_soc_core_memory0_ram_dout0[157]), .B1(n18733), .B2(
        j202_soc_core_memory0_ram_dout0[125]), .Y(n14505) );
  sky130_fd_sc_hd__a22oi_1 U19658 ( .A1(n18361), .A2(
        j202_soc_core_memory0_ram_dout0[61]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[93]), .Y(n14504) );
  sky130_fd_sc_hd__nand2_1 U19659 ( .A(n18735), .B(
        j202_soc_core_memory0_ram_dout0[189]), .Y(n14503) );
  sky130_fd_sc_hd__nand4_1 U19660 ( .A(n14506), .B(n14505), .C(n14504), .D(
        n14503), .Y(n14507) );
  sky130_fd_sc_hd__a21oi_1 U19661 ( .A1(n18367), .A2(
        j202_soc_core_memory0_ram_dout0[29]), .B1(n14507), .Y(n14515) );
  sky130_fd_sc_hd__a22oi_1 U19662 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[317]), .B1(n18062), .B2(
        j202_soc_core_memory0_ram_dout0[285]), .Y(n14514) );
  sky130_fd_sc_hd__nand2_1 U19663 ( .A(n18743), .B(
        j202_soc_core_memory0_ram_dout0[381]), .Y(n14511) );
  sky130_fd_sc_hd__a21oi_1 U19664 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[477]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n14510) );
  sky130_fd_sc_hd__nand2_1 U19665 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[413]), .Y(n14509) );
  sky130_fd_sc_hd__nand2_1 U19666 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[445]), .Y(n14508) );
  sky130_fd_sc_hd__nand4_1 U19667 ( .A(n14511), .B(n14510), .C(n14509), .D(
        n14508), .Y(n14512) );
  sky130_fd_sc_hd__a21oi_1 U19668 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[349]), .B1(n14512), .Y(n14513) );
  sky130_fd_sc_hd__o211ai_1 U19669 ( .A1(n18736), .A2(n14515), .B1(n14514), 
        .C1(n14513), .Y(n14516) );
  sky130_fd_sc_hd__o211ai_1 U19670 ( .A1(j202_soc_core_memory0_ram_dout0[509]), 
        .A2(n18758), .B1(n14906), .C1(n14516), .Y(n14517) );
  sky130_fd_sc_hd__nand2b_1 U19671 ( .A_N(n14518), .B(n14517), .Y(n14519) );
  sky130_fd_sc_hd__a21oi_1 U19672 ( .A1(n14520), .A2(n18798), .B1(n14519), .Y(
        n14521) );
  sky130_fd_sc_hd__nand3_1 U19673 ( .A(n14523), .B(n14522), .C(n14521), .Y(
        n20546) );
  sky130_fd_sc_hd__nand2_1 U19674 ( .A(n20546), .B(n19737), .Y(n14524) );
  sky130_fd_sc_hd__o211ai_1 U19675 ( .A1(n21985), .A2(n19083), .B1(n14525), 
        .C1(n14524), .Y(n14526) );
  sky130_fd_sc_hd__a21oi_1 U19676 ( .A1(n21987), .A2(n19517), .B1(n14526), .Y(
        n14528) );
  sky130_fd_sc_hd__nand2_1 U19677 ( .A(n21987), .B(n19732), .Y(n14527) );
  sky130_fd_sc_hd__nand3_1 U19678 ( .A(n14529), .B(n14528), .C(n14527), .Y(
        n18472) );
  sky130_fd_sc_hd__nand3_1 U19679 ( .A(n14965), .B(n14530), .C(n18472), .Y(
        n18509) );
  sky130_fd_sc_hd__nand2_1 U19680 ( .A(n14533), .B(n14532), .Y(n14534) );
  sky130_fd_sc_hd__xor2_1 U19681 ( .A(n14535), .B(n14534), .X(n22252) );
  sky130_fd_sc_hd__nand2_1 U19682 ( .A(n22252), .B(n19729), .Y(n14675) );
  sky130_fd_sc_hd__ha_1 U19683 ( .A(j202_soc_core_j22_cpu_pc[26]), .B(n14536), 
        .COUT(n14183), .SUM(n22254) );
  sky130_fd_sc_hd__o22a_1 U19684 ( .A1(n22602), .A2(n18948), .B1(n22601), .B2(
        n19731), .X(n14671) );
  sky130_fd_sc_hd__nor4_1 U19685 ( .A(n14539), .B(n14538), .C(n14537), .D(
        n14600), .Y(n14541) );
  sky130_fd_sc_hd__a31oi_1 U19686 ( .A1(n14542), .A2(n14541), .A3(n14540), 
        .B1(n14639), .Y(n14561) );
  sky130_fd_sc_hd__nor2_1 U19687 ( .A(n14544), .B(n14543), .Y(n14545) );
  sky130_fd_sc_hd__a31oi_1 U19688 ( .A1(n14547), .A2(n14546), .A3(n14545), 
        .B1(n14631), .Y(n14560) );
  sky130_fd_sc_hd__a21oi_1 U19689 ( .A1(n14549), .A2(n14548), .B1(n14597), .Y(
        n14551) );
  sky130_fd_sc_hd__a31oi_1 U19690 ( .A1(n14552), .A2(n14551), .A3(n14550), 
        .B1(n15149), .Y(n14559) );
  sky130_fd_sc_hd__nor2_1 U19691 ( .A(n14554), .B(n14553), .Y(n14556) );
  sky130_fd_sc_hd__a31oi_1 U19692 ( .A1(n14557), .A2(n14556), .A3(n14555), 
        .B1(n14619), .Y(n14558) );
  sky130_fd_sc_hd__nor4_1 U19693 ( .A(n14561), .B(n14560), .C(n14559), .D(
        n14558), .Y(n14564) );
  sky130_fd_sc_hd__nand2b_1 U19694 ( .A_N(n14564), .B(n14563), .Y(n14649) );
  sky130_fd_sc_hd__a21oi_1 U19695 ( .A1(n14571), .A2(n14572), .B1(n14565), .Y(
        n14568) );
  sky130_fd_sc_hd__nand4_1 U19696 ( .A(n14569), .B(n14568), .C(n14567), .D(
        n14566), .Y(n14590) );
  sky130_fd_sc_hd__nand2_1 U19697 ( .A(n14572), .B(n14571), .Y(n14573) );
  sky130_fd_sc_hd__a31oi_1 U19698 ( .A1(n14574), .A2(n14581), .A3(n14573), 
        .B1(n14619), .Y(n14589) );
  sky130_fd_sc_hd__nor2_1 U19699 ( .A(n14576), .B(n14575), .Y(n14629) );
  sky130_fd_sc_hd__nor4_1 U19700 ( .A(n14579), .B(n14578), .C(n14629), .D(
        n14577), .Y(n14587) );
  sky130_fd_sc_hd__nand4_1 U19701 ( .A(n14583), .B(n14582), .C(n14581), .D(
        n14580), .Y(n14584) );
  sky130_fd_sc_hd__a211oi_1 U19704 ( .A1(n15093), .A2(n14590), .B1(n14589), 
        .C1(n14588), .Y(n14616) );
  sky130_fd_sc_hd__nand4_1 U19705 ( .A(n14594), .B(n14593), .C(n14592), .D(
        n14591), .Y(n14612) );
  sky130_fd_sc_hd__a21oi_1 U19706 ( .A1(n14596), .A2(n14595), .B1(n14619), .Y(
        n14611) );
  sky130_fd_sc_hd__nor4_1 U19707 ( .A(n14602), .B(n14601), .C(n14600), .D(
        n14599), .Y(n14609) );
  sky130_fd_sc_hd__nor2_1 U19709 ( .A(n14607), .B(n14606), .Y(n14608) );
  sky130_fd_sc_hd__o22ai_1 U19710 ( .A1(n14631), .A2(n14609), .B1(n14608), 
        .B2(n15149), .Y(n14610) );
  sky130_fd_sc_hd__a211oi_1 U19711 ( .A1(n14613), .A2(n14612), .B1(n14611), 
        .C1(n14610), .Y(n14614) );
  sky130_fd_sc_hd__o22a_1 U19712 ( .A1(n14617), .A2(n14616), .B1(n14615), .B2(
        n14614), .X(n14648) );
  sky130_fd_sc_hd__a31oi_1 U19713 ( .A1(n14622), .A2(n14621), .A3(n14620), 
        .B1(n14619), .Y(n14644) );
  sky130_fd_sc_hd__nor3_1 U19714 ( .A(n14624), .B(n14630), .C(n14623), .Y(
        n14626) );
  sky130_fd_sc_hd__a31oi_1 U19715 ( .A1(n14626), .A2(n14637), .A3(n14625), 
        .B1(n15149), .Y(n14643) );
  sky130_fd_sc_hd__or3b_2 U19716 ( .A(n14629), .B(n14628), .C_N(n14627), .X(
        n14635) );
  sky130_fd_sc_hd__nor2_1 U19717 ( .A(n14630), .B(n14635), .Y(n14633) );
  sky130_fd_sc_hd__a31oi_1 U19718 ( .A1(n14634), .A2(n14633), .A3(n14632), 
        .B1(n14631), .Y(n14642) );
  sky130_fd_sc_hd__nor3b_1 U19719 ( .C_N(n14637), .A(n14636), .B(n14635), .Y(
        n14640) );
  sky130_fd_sc_hd__o21bai_1 U19720 ( .A1(n14640), .A2(n14639), .B1_N(n14638), 
        .Y(n14641) );
  sky130_fd_sc_hd__nor4_1 U19721 ( .A(n14644), .B(n14643), .C(n14642), .D(
        n14641), .Y(n14646) );
  sky130_fd_sc_hd__nand2b_1 U19722 ( .A_N(n14646), .B(n14645), .Y(n14647) );
  sky130_fd_sc_hd__nand3_1 U19723 ( .A(n14649), .B(n14648), .C(n14647), .Y(
        n14669) );
  sky130_fd_sc_hd__a22oi_1 U19724 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[250]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[218]), .Y(n14653) );
  sky130_fd_sc_hd__a22oi_1 U19725 ( .A1(n18734), .A2(
        j202_soc_core_memory0_ram_dout0[154]), .B1(n18733), .B2(
        j202_soc_core_memory0_ram_dout0[122]), .Y(n14652) );
  sky130_fd_sc_hd__a22oi_1 U19726 ( .A1(n18361), .A2(
        j202_soc_core_memory0_ram_dout0[58]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[90]), .Y(n14651) );
  sky130_fd_sc_hd__nand2_1 U19727 ( .A(n18735), .B(
        j202_soc_core_memory0_ram_dout0[186]), .Y(n14650) );
  sky130_fd_sc_hd__nand4_1 U19728 ( .A(n14653), .B(n14652), .C(n14651), .D(
        n14650), .Y(n14654) );
  sky130_fd_sc_hd__a32oi_1 U19729 ( .A1(n18367), .A2(n17639), .A3(
        j202_soc_core_memory0_ram_dout0[26]), .B1(n14654), .B2(n17639), .Y(
        n14662) );
  sky130_fd_sc_hd__a22oi_1 U19730 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[314]), .B1(n18062), .B2(
        j202_soc_core_memory0_ram_dout0[282]), .Y(n14661) );
  sky130_fd_sc_hd__nand2_1 U19731 ( .A(n18743), .B(
        j202_soc_core_memory0_ram_dout0[378]), .Y(n14658) );
  sky130_fd_sc_hd__a21oi_1 U19732 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[474]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n14657) );
  sky130_fd_sc_hd__nand2_1 U19733 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[410]), .Y(n14656) );
  sky130_fd_sc_hd__nand2_1 U19734 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[442]), .Y(n14655) );
  sky130_fd_sc_hd__nand4_1 U19735 ( .A(n14658), .B(n14657), .C(n14656), .D(
        n14655), .Y(n14659) );
  sky130_fd_sc_hd__a21oi_1 U19736 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[346]), .B1(n14659), .Y(n14660) );
  sky130_fd_sc_hd__nand3_1 U19737 ( .A(n14662), .B(n14661), .C(n14660), .Y(
        n14663) );
  sky130_fd_sc_hd__o211ai_1 U19738 ( .A1(j202_soc_core_memory0_ram_dout0[506]), 
        .A2(n18758), .B1(n14906), .C1(n14663), .Y(n14666) );
  sky130_fd_sc_hd__a22oi_1 U19739 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[26]), .B1(n18727), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[90]), .Y(n14665) );
  sky130_fd_sc_hd__a22oi_1 U19740 ( .A1(n18726), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[58]), .B1(n18379), .B2(
        j202_soc_core_uart_div0[2]), .Y(n14664) );
  sky130_fd_sc_hd__nand3_1 U19741 ( .A(n14666), .B(n14665), .C(n14664), .Y(
        n14667) );
  sky130_fd_sc_hd__a21o_1 U19742 ( .A1(n14669), .A2(n14668), .B1(n14667), .X(
        n20825) );
  sky130_fd_sc_hd__nand2_1 U19743 ( .A(n20825), .B(n19737), .Y(n14670) );
  sky130_fd_sc_hd__o211ai_1 U19744 ( .A1(n22602), .A2(n19083), .B1(n14671), 
        .C1(n14670), .Y(n14672) );
  sky130_fd_sc_hd__a21oi_1 U19745 ( .A1(n22254), .A2(n19517), .B1(n14672), .Y(
        n14674) );
  sky130_fd_sc_hd__nand2_1 U19746 ( .A(n22254), .B(n19732), .Y(n14673) );
  sky130_fd_sc_hd__nand3_1 U19747 ( .A(n14675), .B(n14674), .C(n14673), .Y(
        n18506) );
  sky130_fd_sc_hd__nand3_1 U19748 ( .A(n18506), .B(n25281), .C(n25250), .Y(
        n14799) );
  sky130_fd_sc_hd__nand2_1 U19749 ( .A(n14679), .B(n14678), .Y(n14819) );
  sky130_fd_sc_hd__nor4_1 U19750 ( .A(n14680), .B(n14879), .C(n14849), .D(
        n14819), .Y(n14681) );
  sky130_fd_sc_hd__a21oi_1 U19751 ( .A1(n14682), .A2(n14681), .B1(n14871), .Y(
        n14701) );
  sky130_fd_sc_hd__nor4b_1 U19752 ( .D_N(n14684), .A(n14683), .B(n14809), .C(
        n14821), .Y(n14686) );
  sky130_fd_sc_hd__a21oi_1 U19753 ( .A1(n14686), .A2(n14685), .B1(n14884), .Y(
        n14700) );
  sky130_fd_sc_hd__nand4b_1 U19754 ( .A_N(n14687), .B(n14774), .C(n14839), .D(
        n14705), .Y(n14688) );
  sky130_fd_sc_hd__nand2_1 U19755 ( .A(n14841), .B(n14688), .Y(n14790) );
  sky130_fd_sc_hd__nand2_1 U19756 ( .A(n14689), .B(n14790), .Y(n14856) );
  sky130_fd_sc_hd__and4_1 U19757 ( .A(n14692), .B(n14691), .C(n14690), .D(
        n14877), .X(n14698) );
  sky130_fd_sc_hd__nor4b_1 U19758 ( .D_N(n14875), .A(n14696), .B(n14695), .C(
        n14712), .Y(n14697) );
  sky130_fd_sc_hd__o22ai_1 U19759 ( .A1(n14698), .A2(n14882), .B1(n14697), 
        .B2(n14815), .Y(n14699) );
  sky130_fd_sc_hd__nor4_1 U19760 ( .A(n14701), .B(n14700), .C(n14856), .D(
        n14699), .Y(n14794) );
  sky130_fd_sc_hd__nand4_1 U19761 ( .A(n14702), .B(n14810), .C(n14838), .D(
        n14862), .Y(n14704) );
  sky130_fd_sc_hd__nor3_1 U19762 ( .A(n14704), .B(n14728), .C(n14703), .Y(
        n14710) );
  sky130_fd_sc_hd__nand4_1 U19763 ( .A(n14885), .B(n14707), .C(n14706), .D(
        n14705), .Y(n14708) );
  sky130_fd_sc_hd__o21ai_1 U19764 ( .A1(n14833), .A2(n14708), .B1(n14720), .Y(
        n14709) );
  sky130_fd_sc_hd__nand2b_1 U19766 ( .A_N(n14771), .B(n14711), .Y(n14820) );
  sky130_fd_sc_hd__o31a_1 U19767 ( .A1(n14820), .A2(n14727), .A3(n14712), .B1(
        n14841), .X(n14713) );
  sky130_fd_sc_hd__a211oi_1 U19768 ( .A1(n14866), .A2(n14715), .B1(n14714), 
        .C1(n14713), .Y(n14716) );
  sky130_fd_sc_hd__nor2_1 U19769 ( .A(n18720), .B(n14716), .Y(n14765) );
  sky130_fd_sc_hd__o21ai_1 U19770 ( .A1(n14722), .A2(n14721), .B1(n14720), .Y(
        n14735) );
  sky130_fd_sc_hd__nand2_1 U19771 ( .A(n14724), .B(n14723), .Y(n14725) );
  sky130_fd_sc_hd__nand2_1 U19773 ( .A(n14732), .B(n14841), .Y(n14733) );
  sky130_fd_sc_hd__nand3_1 U19774 ( .A(n14735), .B(n14734), .C(n14733), .Y(
        n14744) );
  sky130_fd_sc_hd__nor4b_1 U19775 ( .D_N(n14739), .A(n14738), .B(n14737), .C(
        n14843), .Y(n14740) );
  sky130_fd_sc_hd__a31oi_1 U19776 ( .A1(n14742), .A2(n14741), .A3(n14740), 
        .B1(n14882), .Y(n14743) );
  sky130_fd_sc_hd__a22oi_1 U19778 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[30]), .B1(n18727), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[94]), .Y(n14762) );
  sky130_fd_sc_hd__a22oi_1 U19779 ( .A1(n18726), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[62]), .B1(n18379), .B2(
        j202_soc_core_uart_div0[6]), .Y(n14761) );
  sky130_fd_sc_hd__a22oi_1 U19780 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[254]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[222]), .Y(n14748) );
  sky130_fd_sc_hd__a22oi_1 U19781 ( .A1(n18734), .A2(
        j202_soc_core_memory0_ram_dout0[158]), .B1(n18733), .B2(
        j202_soc_core_memory0_ram_dout0[126]), .Y(n14747) );
  sky130_fd_sc_hd__a22oi_1 U19782 ( .A1(n18361), .A2(
        j202_soc_core_memory0_ram_dout0[62]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[94]), .Y(n14746) );
  sky130_fd_sc_hd__nand2_1 U19783 ( .A(n18735), .B(
        j202_soc_core_memory0_ram_dout0[190]), .Y(n14745) );
  sky130_fd_sc_hd__nand4_1 U19784 ( .A(n14748), .B(n14747), .C(n14746), .D(
        n14745), .Y(n14749) );
  sky130_fd_sc_hd__a21oi_1 U19785 ( .A1(n18367), .A2(
        j202_soc_core_memory0_ram_dout0[30]), .B1(n14749), .Y(n14750) );
  sky130_fd_sc_hd__nand2b_1 U19786 ( .A_N(n14750), .B(n17639), .Y(n14758) );
  sky130_fd_sc_hd__a22oi_1 U19787 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[318]), .B1(n18062), .B2(
        j202_soc_core_memory0_ram_dout0[286]), .Y(n14757) );
  sky130_fd_sc_hd__nand2_1 U19788 ( .A(n18743), .B(
        j202_soc_core_memory0_ram_dout0[382]), .Y(n14754) );
  sky130_fd_sc_hd__a21oi_1 U19789 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[478]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n14753) );
  sky130_fd_sc_hd__nand2_1 U19790 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[414]), .Y(n14752) );
  sky130_fd_sc_hd__nand2_1 U19791 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[446]), .Y(n14751) );
  sky130_fd_sc_hd__nand4_1 U19792 ( .A(n14754), .B(n14753), .C(n14752), .D(
        n14751), .Y(n14755) );
  sky130_fd_sc_hd__a21oi_1 U19793 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[350]), .B1(n14755), .Y(n14756) );
  sky130_fd_sc_hd__nand3_1 U19794 ( .A(n14758), .B(n14757), .C(n14756), .Y(
        n14759) );
  sky130_fd_sc_hd__o211ai_1 U19795 ( .A1(j202_soc_core_memory0_ram_dout0[510]), 
        .A2(n18758), .B1(n14906), .C1(n14759), .Y(n14760) );
  sky130_fd_sc_hd__nand4_1 U19796 ( .A(n14763), .B(n14762), .C(n14761), .D(
        n14760), .Y(n14764) );
  sky130_fd_sc_hd__nor2_1 U19797 ( .A(n14765), .B(n14764), .Y(n14793) );
  sky130_fd_sc_hd__nor3_1 U19798 ( .A(n14768), .B(n14767), .C(n14766), .Y(
        n14769) );
  sky130_fd_sc_hd__a31oi_1 U19799 ( .A1(n14836), .A2(n14770), .A3(n14769), 
        .B1(n14884), .Y(n14789) );
  sky130_fd_sc_hd__nor2_1 U19800 ( .A(n14772), .B(n14771), .Y(n14873) );
  sky130_fd_sc_hd__a31oi_1 U19801 ( .A1(n14776), .A2(n14873), .A3(n14775), 
        .B1(n14882), .Y(n14788) );
  sky130_fd_sc_hd__nand4b_1 U19802 ( .A_N(n14858), .B(n14778), .C(n14777), .D(
        n17970), .Y(n14779) );
  sky130_fd_sc_hd__nor4_1 U19803 ( .A(n14881), .B(n14814), .C(n14780), .D(
        n14779), .Y(n14786) );
  sky130_fd_sc_hd__nand2_1 U19804 ( .A(n14782), .B(n14781), .Y(n14831) );
  sky130_fd_sc_hd__nor4_1 U19805 ( .A(n14880), .B(n14784), .C(n14783), .D(
        n14831), .Y(n14785) );
  sky130_fd_sc_hd__o22ai_1 U19806 ( .A1(n14786), .A2(n14815), .B1(n14785), 
        .B2(n14871), .Y(n14787) );
  sky130_fd_sc_hd__nor4b_1 U19807 ( .D_N(n14790), .A(n14789), .B(n14788), .C(
        n14787), .Y(n14791) );
  sky130_fd_sc_hd__nand2b_1 U19808 ( .A_N(n14791), .B(n18798), .Y(n14792) );
  sky130_fd_sc_hd__o211a_2 U19809 ( .A1(n18722), .A2(n14794), .B1(n14793), 
        .C1(n14792), .X(n21045) );
  sky130_fd_sc_hd__a22oi_1 U19810 ( .A1(n19657), .A2(n22579), .B1(n19736), 
        .B2(n23340), .Y(n14797) );
  sky130_fd_sc_hd__ha_1 U19811 ( .A(j202_soc_core_j22_cpu_pc[30]), .B(n14795), 
        .COUT(n14176), .SUM(n21894) );
  sky130_fd_sc_hd__nand2_1 U19812 ( .A(n21894), .B(n19661), .Y(n14796) );
  sky130_fd_sc_hd__o211ai_1 U19813 ( .A1(n21045), .A2(n14919), .B1(n14797), 
        .C1(n14796), .Y(n14798) );
  sky130_fd_sc_hd__a21oi_1 U19814 ( .A1(n21892), .A2(n19729), .B1(n14798), .Y(
        n18508) );
  sky130_fd_sc_hd__nor2_1 U19815 ( .A(n14799), .B(n18508), .Y(n14800) );
  sky130_fd_sc_hd__nand2b_1 U19816 ( .A_N(n18509), .B(n14800), .Y(n14956) );
  sky130_fd_sc_hd__nand2_1 U19817 ( .A(n14801), .B(io_in[14]), .Y(n14972) );
  sky130_fd_sc_hd__nand2_1 U19818 ( .A(n14956), .B(n14972), .Y(n14955) );
  sky130_fd_sc_hd__nand2_1 U19819 ( .A(n14804), .B(n14803), .Y(n14805) );
  sky130_fd_sc_hd__xor2_1 U19820 ( .A(n14806), .B(n14805), .X(n22073) );
  sky130_fd_sc_hd__nand2_1 U19821 ( .A(n22073), .B(n19729), .Y(n14923) );
  sky130_fd_sc_hd__ha_1 U19822 ( .A(j202_soc_core_j22_cpu_pc[28]), .B(n14807), 
        .COUT(n14398), .SUM(n22080) );
  sky130_fd_sc_hd__nand2_1 U19823 ( .A(n14808), .B(n14839), .Y(n14813) );
  sky130_fd_sc_hd__nor2b_1 U19824 ( .B_N(n14810), .A(n14809), .Y(n14816) );
  sky130_fd_sc_hd__nand2_1 U19825 ( .A(n14816), .B(n14811), .Y(n14834) );
  sky130_fd_sc_hd__o31a_1 U19826 ( .A1(n14813), .A2(n14812), .A3(n14834), .B1(
        n14841), .X(n14827) );
  sky130_fd_sc_hd__nor2_1 U19827 ( .A(n14881), .B(n14814), .Y(n14818) );
  sky130_fd_sc_hd__a31oi_1 U19828 ( .A1(n14818), .A2(n14817), .A3(n14816), 
        .B1(n14815), .Y(n14826) );
  sky130_fd_sc_hd__nor4_1 U19829 ( .A(n14822), .B(n14821), .C(n14820), .D(
        n14819), .Y(n14823) );
  sky130_fd_sc_hd__o22ai_1 U19830 ( .A1(n14824), .A2(n14871), .B1(n14823), 
        .B2(n14882), .Y(n14825) );
  sky130_fd_sc_hd__nor3_1 U19831 ( .A(n14827), .B(n14826), .C(n14825), .Y(
        n14916) );
  sky130_fd_sc_hd__a31oi_1 U19832 ( .A1(n14830), .A2(n14829), .A3(n14828), 
        .B1(n14871), .Y(n14848) );
  sky130_fd_sc_hd__o31a_1 U19833 ( .A1(n14833), .A2(n14832), .A3(n14831), .B1(
        n14888), .X(n14847) );
  sky130_fd_sc_hd__nor4b_1 U19834 ( .D_N(n14836), .A(n14861), .B(n14835), .C(
        n14834), .Y(n14845) );
  sky130_fd_sc_hd__nand4_1 U19835 ( .A(n14840), .B(n14839), .C(n14838), .D(
        n14837), .Y(n14842) );
  sky130_fd_sc_hd__nor3_1 U19838 ( .A(n14848), .B(n14847), .C(n14846), .Y(
        n14914) );
  sky130_fd_sc_hd__o21ai_1 U19839 ( .A1(n14852), .A2(n14851), .B1(n14850), .Y(
        n14853) );
  sky130_fd_sc_hd__a31oi_1 U19840 ( .A1(n14855), .A2(n14854), .A3(n14853), 
        .B1(n14871), .Y(n14857) );
  sky130_fd_sc_hd__nor2_1 U19841 ( .A(n14857), .B(n14856), .Y(n14869) );
  sky130_fd_sc_hd__nor4_1 U19842 ( .A(n14861), .B(n14860), .C(n14859), .D(
        n14858), .Y(n14863) );
  sky130_fd_sc_hd__nand4b_1 U19843 ( .A_N(n14865), .B(n14864), .C(n14863), .D(
        n14862), .Y(n14867) );
  sky130_fd_sc_hd__nand2_1 U19844 ( .A(n14867), .B(n14866), .Y(n14868) );
  sky130_fd_sc_hd__nand2_1 U19845 ( .A(n14869), .B(n14868), .Y(n14870) );
  sky130_fd_sc_hd__nand2_1 U19846 ( .A(n14870), .B(n18605), .Y(n14913) );
  sky130_fd_sc_hd__a21oi_1 U19847 ( .A1(n14873), .A2(n14872), .B1(n14871), .Y(
        n14890) );
  sky130_fd_sc_hd__nand4_1 U19848 ( .A(n14877), .B(n14876), .C(n14875), .D(
        n14874), .Y(n14878) );
  sky130_fd_sc_hd__nor4_1 U19849 ( .A(n14881), .B(n14880), .C(n14879), .D(
        n14878), .Y(n14883) );
  sky130_fd_sc_hd__o22ai_1 U19850 ( .A1(n14885), .A2(n14884), .B1(n14883), 
        .B2(n14882), .Y(n14886) );
  sky130_fd_sc_hd__a21oi_1 U19851 ( .A1(n14888), .A2(n14887), .B1(n14886), .Y(
        n14889) );
  sky130_fd_sc_hd__nand2b_1 U19852 ( .A_N(n14890), .B(n14889), .Y(n14911) );
  sky130_fd_sc_hd__a22oi_1 U19853 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[252]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[220]), .Y(n14894) );
  sky130_fd_sc_hd__a22oi_1 U19854 ( .A1(n18734), .A2(
        j202_soc_core_memory0_ram_dout0[156]), .B1(n18733), .B2(
        j202_soc_core_memory0_ram_dout0[124]), .Y(n14893) );
  sky130_fd_sc_hd__a22oi_1 U19855 ( .A1(n18361), .A2(
        j202_soc_core_memory0_ram_dout0[60]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[92]), .Y(n14892) );
  sky130_fd_sc_hd__nand2_1 U19856 ( .A(n18735), .B(
        j202_soc_core_memory0_ram_dout0[188]), .Y(n14891) );
  sky130_fd_sc_hd__nand4_1 U19857 ( .A(n14894), .B(n14893), .C(n14892), .D(
        n14891), .Y(n14895) );
  sky130_fd_sc_hd__a21oi_1 U19858 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[28]), .B1(n14895), .Y(n14896) );
  sky130_fd_sc_hd__nand2b_1 U19859 ( .A_N(n14896), .B(n17639), .Y(n14904) );
  sky130_fd_sc_hd__a22oi_1 U19860 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[316]), .B1(n18062), .B2(
        j202_soc_core_memory0_ram_dout0[284]), .Y(n14903) );
  sky130_fd_sc_hd__nand2_1 U19861 ( .A(n18743), .B(
        j202_soc_core_memory0_ram_dout0[380]), .Y(n14900) );
  sky130_fd_sc_hd__a21oi_1 U19862 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[476]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n14899) );
  sky130_fd_sc_hd__nand2_1 U19863 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[412]), .Y(n14898) );
  sky130_fd_sc_hd__nand2_1 U19864 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[444]), .Y(n14897) );
  sky130_fd_sc_hd__nand4_1 U19865 ( .A(n14900), .B(n14899), .C(n14898), .D(
        n14897), .Y(n14901) );
  sky130_fd_sc_hd__a21oi_1 U19866 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[348]), .B1(n14901), .Y(n14902) );
  sky130_fd_sc_hd__nand3_1 U19867 ( .A(n14904), .B(n14903), .C(n14902), .Y(
        n14905) );
  sky130_fd_sc_hd__o211ai_1 U19868 ( .A1(j202_soc_core_memory0_ram_dout0[508]), 
        .A2(n18758), .B1(n14906), .C1(n14905), .Y(n14909) );
  sky130_fd_sc_hd__a22oi_1 U19869 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[28]), .B1(n18727), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[92]), .Y(n14908) );
  sky130_fd_sc_hd__a22oi_1 U19870 ( .A1(n18726), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[60]), .B1(n18379), .B2(
        j202_soc_core_uart_div0[4]), .Y(n14907) );
  sky130_fd_sc_hd__nand3_1 U19871 ( .A(n14909), .B(n14908), .C(n14907), .Y(
        n14910) );
  sky130_fd_sc_hd__a21oi_1 U19872 ( .A1(n14911), .A2(n18610), .B1(n14910), .Y(
        n14912) );
  sky130_fd_sc_hd__o211a_2 U19873 ( .A1(n18720), .A2(n14914), .B1(n14913), 
        .C1(n14912), .X(n14915) );
  sky130_fd_sc_hd__o21a_1 U19874 ( .A1(n14916), .A2(n18552), .B1(n14915), .X(
        n22525) );
  sky130_fd_sc_hd__o22a_1 U19875 ( .A1(n22074), .A2(n18948), .B1(n20955), .B2(
        n19731), .X(n14917) );
  sky130_fd_sc_hd__o21a_1 U19876 ( .A1(n22074), .A2(n19083), .B1(n14917), .X(
        n14918) );
  sky130_fd_sc_hd__o21ai_1 U19877 ( .A1(n14919), .A2(n22525), .B1(n14918), .Y(
        n14920) );
  sky130_fd_sc_hd__a21oi_1 U19878 ( .A1(n22080), .A2(n19517), .B1(n14920), .Y(
        n14922) );
  sky130_fd_sc_hd__nand2_1 U19879 ( .A(n22080), .B(n19732), .Y(n14921) );
  sky130_fd_sc_hd__nand3_1 U19880 ( .A(n14923), .B(n14922), .C(n14921), .Y(
        n21074) );
  sky130_fd_sc_hd__nor2_1 U19881 ( .A(n11182), .B(n25299), .Y(n14938) );
  sky130_fd_sc_hd__nor3_1 U19882 ( .A(j202_soc_core_j22_cpu_id_op2_v_), .B(
        j202_soc_core_j22_cpu_id_opn_v_), .C(n23235), .Y(n14924) );
  sky130_fd_sc_hd__a31oi_1 U19883 ( .A1(n23239), .A2(n14938), .A3(n14943), 
        .B1(n14924), .Y(n14936) );
  sky130_fd_sc_hd__nand2_1 U19884 ( .A(n20488), .B(n22807), .Y(n22799) );
  sky130_fd_sc_hd__a22oi_1 U19885 ( .A1(n14926), .A2(
        j202_soc_core_j22_cpu_rfuo_sr__i__3_), .B1(
        j202_soc_core_j22_cpu_rfuo_sr__i__2_), .B2(n14925), .Y(n14933) );
  sky130_fd_sc_hd__nand2_1 U19886 ( .A(j202_soc_core_j22_cpu_rfuo_sr__i__1_), 
        .B(n14927), .Y(n14928) );
  sky130_fd_sc_hd__nand3_1 U19887 ( .A(n14928), .B(n17064), .C(
        j202_soc_core_intr_level__0_), .Y(n14931) );
  sky130_fd_sc_hd__nand2_1 U19888 ( .A(n19052), .B(
        j202_soc_core_intr_level__2_), .Y(n14930) );
  sky130_fd_sc_hd__nand2_1 U19889 ( .A(n19180), .B(
        j202_soc_core_intr_level__1_), .Y(n14929) );
  sky130_fd_sc_hd__nand3_1 U19890 ( .A(n14931), .B(n14930), .C(n14929), .Y(
        n14932) );
  sky130_fd_sc_hd__nand2_1 U19891 ( .A(n14933), .B(n14932), .Y(n14935) );
  sky130_fd_sc_hd__a21oi_1 U19892 ( .A1(n16692), .A2(
        j202_soc_core_intr_level__3_), .B1(j202_soc_core_intr_level__4_), .Y(
        n14934) );
  sky130_fd_sc_hd__a21oi_1 U19893 ( .A1(n14935), .A2(n14934), .B1(n21399), .Y(
        n22792) );
  sky130_fd_sc_hd__nand2_1 U19894 ( .A(n23239), .B(n22792), .Y(n22802) );
  sky130_fd_sc_hd__nand4_1 U19895 ( .A(n14936), .B(n22799), .C(n25731), .D(
        n22802), .Y(n22798) );
  sky130_fd_sc_hd__o21ai_1 U19896 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        n24894), .B1(j202_soc_core_j22_cpu_id_opn_v_), .Y(n14937) );
  sky130_fd_sc_hd__nand2_1 U19897 ( .A(n14938), .B(n14937), .Y(n14941) );
  sky130_fd_sc_hd__o211ai_1 U19898 ( .A1(n14939), .A2(n22789), .B1(n25543), 
        .C1(n21338), .Y(n14940) );
  sky130_fd_sc_hd__a21oi_1 U19899 ( .A1(n14941), .A2(n22789), .B1(n14940), .Y(
        n14942) );
  sky130_fd_sc_hd__nand2b_1 U19900 ( .A_N(n22798), .B(n14942), .Y(n23241) );
  sky130_fd_sc_hd__nand2_1 U19901 ( .A(n23241), .B(n14944), .Y(n14959) );
  sky130_fd_sc_hd__nor2_1 U19902 ( .A(n14945), .B(n25251), .Y(n14946) );
  sky130_fd_sc_hd__o21a_1 U19903 ( .A1(n14962), .A2(n21074), .B1(n14946), .X(
        n14954) );
  sky130_fd_sc_hd__nor2_1 U19904 ( .A(n25277), .B(n25280), .Y(n14968) );
  sky130_fd_sc_hd__nor3_1 U19905 ( .A(n25252), .B(n25250), .C(n25281), .Y(
        n14947) );
  sky130_fd_sc_hd__nand4_1 U19906 ( .A(n14963), .B(n14948), .C(n14968), .D(
        n14947), .Y(n14949) );
  sky130_fd_sc_hd__nor3_1 U19907 ( .A(n14961), .B(n14949), .C(n21074), .Y(
        n14950) );
  sky130_fd_sc_hd__nand4b_1 U19908 ( .A_N(n14965), .B(n21075), .C(n18508), .D(
        n14950), .Y(n14952) );
  sky130_fd_sc_hd__nand2_1 U19909 ( .A(n14952), .B(n14951), .Y(n14953) );
  sky130_fd_sc_hd__and3_1 U19910 ( .A(n11036), .B(n25488), .C(n22403), .X(
        n25248) );
  sky130_fd_sc_hd__nand2_1 U19911 ( .A(n22403), .B(n14959), .Y(n22381) );
  sky130_fd_sc_hd__nand2_1 U19912 ( .A(n21253), .B(
        j202_soc_core_ahbcs_6__HREADY_), .Y(n14960) );
  sky130_fd_sc_hd__nand4_1 U19913 ( .A(n18508), .B(n14964), .C(n14963), .D(
        n14962), .Y(n14966) );
  sky130_fd_sc_hd__nor2_1 U19914 ( .A(n14966), .B(n14965), .Y(n18476) );
  sky130_fd_sc_hd__nor3_1 U19915 ( .A(n25252), .B(n25251), .C(n25250), .Y(
        n14967) );
  sky130_fd_sc_hd__nand3_1 U19916 ( .A(n14968), .B(n18504), .C(n14967), .Y(
        n14969) );
  sky130_fd_sc_hd__nor2_1 U19917 ( .A(n25257), .B(n14969), .Y(n14970) );
  sky130_fd_sc_hd__nand3_1 U19918 ( .A(n22099), .B(n18476), .C(n14970), .Y(
        n21076) );
  sky130_fd_sc_hd__nand2_1 U19919 ( .A(n14971), .B(io_in[15]), .Y(n18473) );
  sky130_fd_sc_hd__nand2_1 U19920 ( .A(n14972), .B(n18473), .Y(n14973) );
  sky130_fd_sc_hd__mux2i_1 U19921 ( .A0(n18472), .A1(n18475), .S(n14973), .Y(
        n14975) );
  sky130_fd_sc_hd__nand2_1 U19922 ( .A(n21075), .B(n21074), .Y(n14974) );
  sky130_fd_sc_hd__nor2_1 U19923 ( .A(j202_soc_core_bootrom_00_address_w[5]), 
        .B(n14999), .Y(n17543) );
  sky130_fd_sc_hd__nor2_1 U19924 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(n17799), .Y(n17662) );
  sky130_fd_sc_hd__nand2_1 U19925 ( .A(n14980), .B(
        j202_soc_core_bootrom_00_address_w[6]), .Y(n16740) );
  sky130_fd_sc_hd__nand2_1 U19926 ( .A(n14977), .B(n14997), .Y(n17875) );
  sky130_fd_sc_hd__nor2_1 U19927 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(n14978), .Y(n16744) );
  sky130_fd_sc_hd__nor2_1 U19928 ( .A(n15009), .B(n14979), .Y(n17945) );
  sky130_fd_sc_hd__nor2_1 U19929 ( .A(n14998), .B(n18519), .Y(n18392) );
  sky130_fd_sc_hd__nand2_1 U19930 ( .A(n14980), .B(n14998), .Y(n17441) );
  sky130_fd_sc_hd__nor2_1 U19931 ( .A(n14981), .B(n17441), .Y(n18435) );
  sky130_fd_sc_hd__nand2_1 U19932 ( .A(n17757), .B(n17771), .Y(n17867) );
  sky130_fd_sc_hd__nor2_1 U19933 ( .A(n17945), .B(n17867), .Y(n17599) );
  sky130_fd_sc_hd__nand2_1 U19934 ( .A(n14982), .B(
        j202_soc_core_bootrom_00_address_w[6]), .Y(n14992) );
  sky130_fd_sc_hd__nor2_1 U19935 ( .A(n14992), .B(n17731), .Y(n18397) );
  sky130_fd_sc_hd__nand2_1 U19936 ( .A(n17599), .B(n17617), .Y(n17806) );
  sky130_fd_sc_hd__nor3_1 U19937 ( .A(n17662), .B(n17746), .C(n17806), .Y(
        n17418) );
  sky130_fd_sc_hd__nand2_1 U19938 ( .A(n14983), .B(n14998), .Y(n14984) );
  sky130_fd_sc_hd__nor2_1 U19939 ( .A(n14984), .B(n18296), .Y(n18398) );
  sky130_fd_sc_hd__nand2_1 U19940 ( .A(n18398), .B(n14985), .Y(n17478) );
  sky130_fd_sc_hd__nand2_1 U19941 ( .A(n14986), .B(
        j202_soc_core_bootrom_00_address_w[6]), .Y(n14993) );
  sky130_fd_sc_hd__nor2_1 U19942 ( .A(n14993), .B(n17442), .Y(n17509) );
  sky130_fd_sc_hd__nor2_1 U19943 ( .A(n18418), .B(n17509), .Y(n17470) );
  sky130_fd_sc_hd__nor2_1 U19944 ( .A(n14998), .B(n17778), .Y(n15018) );
  sky130_fd_sc_hd__nand2_1 U19945 ( .A(n17777), .B(n15018), .Y(n17548) );
  sky130_fd_sc_hd__nor2_1 U19946 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(n17672), .Y(n17915) );
  sky130_fd_sc_hd__nand2_1 U19947 ( .A(n15016), .B(n15017), .Y(n14987) );
  sky130_fd_sc_hd__nor2_1 U19948 ( .A(n14987), .B(n16740), .Y(n17624) );
  sky130_fd_sc_hd__nor2_1 U19949 ( .A(n17915), .B(n17624), .Y(n17557) );
  sky130_fd_sc_hd__nor2_1 U19950 ( .A(n17621), .B(n17744), .Y(n16739) );
  sky130_fd_sc_hd__nor2_1 U19951 ( .A(n14987), .B(n17441), .Y(n17737) );
  sky130_fd_sc_hd__nor2_1 U19952 ( .A(n14989), .B(n14988), .Y(n17508) );
  sky130_fd_sc_hd__nand2_1 U19953 ( .A(n17508), .B(n14998), .Y(n18446) );
  sky130_fd_sc_hd__nor2_1 U19954 ( .A(n17737), .B(n17944), .Y(n17908) );
  sky130_fd_sc_hd__nand4_1 U19955 ( .A(n17418), .B(n17528), .C(n16739), .D(
        n17908), .Y(n14996) );
  sky130_fd_sc_hd__nand2_1 U19956 ( .A(n17469), .B(n17532), .Y(n17911) );
  sky130_fd_sc_hd__nand2_1 U19957 ( .A(n16737), .B(n17911), .Y(n17943) );
  sky130_fd_sc_hd__nand2_1 U19958 ( .A(n17469), .B(n15018), .Y(n18399) );
  sky130_fd_sc_hd__nand2_1 U19959 ( .A(n17620), .B(n18399), .Y(n17530) );
  sky130_fd_sc_hd__nor2_1 U19960 ( .A(n18392), .B(n17530), .Y(n17750) );
  sky130_fd_sc_hd__nand2_1 U19961 ( .A(n17469), .B(n14997), .Y(n18346) );
  sky130_fd_sc_hd__nor2_1 U19962 ( .A(n14998), .B(n17912), .Y(n17784) );
  sky130_fd_sc_hd__nand2_1 U19963 ( .A(n16744), .B(n14990), .Y(n16736) );
  sky130_fd_sc_hd__nor2_1 U19964 ( .A(n17784), .B(n18354), .Y(n17623) );
  sky130_fd_sc_hd__nand2_1 U19965 ( .A(n17508), .B(
        j202_soc_core_bootrom_00_address_w[6]), .Y(n18341) );
  sky130_fd_sc_hd__nand2_1 U19966 ( .A(n17623), .B(n18341), .Y(n17669) );
  sky130_fd_sc_hd__nor2_1 U19967 ( .A(n17752), .B(n17669), .Y(n17417) );
  sky130_fd_sc_hd__nor2_1 U19968 ( .A(n14998), .B(n17672), .Y(n17842) );
  sky130_fd_sc_hd__nor2_1 U19969 ( .A(n17624), .B(n17842), .Y(n18402) );
  sky130_fd_sc_hd__nand2_1 U19970 ( .A(n17533), .B(n16744), .Y(n17923) );
  sky130_fd_sc_hd__nand3_1 U19971 ( .A(n18402), .B(n17923), .C(n17771), .Y(
        n17482) );
  sky130_fd_sc_hd__nor2_1 U19972 ( .A(j202_soc_core_bootrom_00_address_w[6]), 
        .B(n14991), .Y(n17910) );
  sky130_fd_sc_hd__nor2_1 U19973 ( .A(n14992), .B(n15009), .Y(n17866) );
  sky130_fd_sc_hd__nand2_1 U19974 ( .A(n17779), .B(n18347), .Y(n17526) );
  sky130_fd_sc_hd__nor2_1 U19975 ( .A(n15009), .B(n14993), .Y(n17774) );
  sky130_fd_sc_hd__nand2_1 U19976 ( .A(n17777), .B(n17532), .Y(n17791) );
  sky130_fd_sc_hd__nand2_1 U19977 ( .A(n17596), .B(n17791), .Y(n18390) );
  sky130_fd_sc_hd__nor3_1 U19978 ( .A(n17482), .B(n17526), .C(n18390), .Y(
        n14994) );
  sky130_fd_sc_hd__a31oi_1 U19979 ( .A1(n17750), .A2(n17417), .A3(n14994), 
        .B1(n18423), .Y(n14995) );
  sky130_fd_sc_hd__a21oi_1 U19980 ( .A1(n17543), .A2(n14996), .B1(n14995), .Y(
        n15004) );
  sky130_fd_sc_hd__nor2_1 U19981 ( .A(j202_soc_core_bootrom_00_address_w[7]), 
        .B(j202_soc_core_bootrom_00_address_w[5]), .Y(n17812) );
  sky130_fd_sc_hd__nand2_1 U19982 ( .A(n17596), .B(n16736), .Y(n15036) );
  sky130_fd_sc_hd__nand2_1 U19983 ( .A(n17923), .B(n17478), .Y(n16767) );
  sky130_fd_sc_hd__nor2_1 U19984 ( .A(n17866), .B(n16767), .Y(n16714) );
  sky130_fd_sc_hd__nor2_1 U19985 ( .A(n14998), .B(n17768), .Y(n17916) );
  sky130_fd_sc_hd__nand2_1 U19986 ( .A(n17604), .B(
        j202_soc_core_bootrom_00_address_w[6]), .Y(n17863) );
  sky130_fd_sc_hd__nand2_1 U19987 ( .A(n17868), .B(n17863), .Y(n17928) );
  sky130_fd_sc_hd__nand2_1 U19988 ( .A(n17678), .B(n18346), .Y(n17865) );
  sky130_fd_sc_hd__nand2_1 U19989 ( .A(n17845), .B(n18341), .Y(n15007) );
  sky130_fd_sc_hd__nor2_1 U19990 ( .A(n17928), .B(n15007), .Y(n16747) );
  sky130_fd_sc_hd__nand2_1 U19991 ( .A(n17469), .B(n17930), .Y(n17756) );
  sky130_fd_sc_hd__nand2_1 U19992 ( .A(n17593), .B(n14998), .Y(n17676) );
  sky130_fd_sc_hd__nand2_1 U19993 ( .A(n17756), .B(n17676), .Y(n17870) );
  sky130_fd_sc_hd__nor2_1 U19994 ( .A(n17727), .B(n17870), .Y(n17525) );
  sky130_fd_sc_hd__nand4_1 U19995 ( .A(n15011), .B(n16714), .C(n16747), .D(
        n17525), .Y(n15002) );
  sky130_fd_sc_hd__nor3_1 U19996 ( .A(n17774), .B(n17662), .C(n17727), .Y(
        n16765) );
  sky130_fd_sc_hd__nand2_1 U19997 ( .A(n17757), .B(n17923), .Y(n17670) );
  sky130_fd_sc_hd__nand2_1 U19998 ( .A(n18398), .B(
        j202_soc_core_bootrom_00_address_w[4]), .Y(n17618) );
  sky130_fd_sc_hd__nor2_1 U19999 ( .A(n18436), .B(n17866), .Y(n17739) );
  sky130_fd_sc_hd__nand2_1 U20000 ( .A(n17777), .B(n14997), .Y(n17675) );
  sky130_fd_sc_hd__nand2_1 U20001 ( .A(n17739), .B(n17675), .Y(n17751) );
  sky130_fd_sc_hd__nand3_1 U20002 ( .A(n17676), .B(n17617), .C(n18399), .Y(
        n17759) );
  sky130_fd_sc_hd__nand2_1 U20003 ( .A(n17604), .B(n14998), .Y(n17554) );
  sky130_fd_sc_hd__nand2_1 U20004 ( .A(n17554), .B(n18346), .Y(n16769) );
  sky130_fd_sc_hd__nor4_1 U20005 ( .A(n17915), .B(n17751), .C(n17759), .D(
        n16769), .Y(n15000) );
  sky130_fd_sc_hd__nand2_1 U20006 ( .A(n14999), .B(
        j202_soc_core_bootrom_00_address_w[5]), .Y(n18439) );
  sky130_fd_sc_hd__a31oi_1 U20007 ( .A1(n16765), .A2(n17876), .A3(n15000), 
        .B1(n18439), .Y(n15001) );
  sky130_fd_sc_hd__a21oi_1 U20008 ( .A1(n17812), .A2(n15002), .B1(n15001), .Y(
        n15003) );
  sky130_fd_sc_hd__a21oi_1 U20009 ( .A1(n15004), .A2(n15003), .B1(n18666), .Y(
        n15062) );
  sky130_fd_sc_hd__nand2_1 U20010 ( .A(n17478), .B(n17676), .Y(n17773) );
  sky130_fd_sc_hd__nand2_1 U20011 ( .A(n17653), .B(n17615), .Y(n17536) );
  sky130_fd_sc_hd__nor2_1 U20012 ( .A(n18248), .B(n17536), .Y(n15005) );
  sky130_fd_sc_hd__nand2_1 U20013 ( .A(n17923), .B(n18346), .Y(n17661) );
  sky130_fd_sc_hd__nor2_1 U20014 ( .A(n17915), .B(n17661), .Y(n17614) );
  sky130_fd_sc_hd__a31oi_1 U20015 ( .A1(n15005), .A2(n17614), .A3(n16737), 
        .B1(n18437), .Y(n15015) );
  sky130_fd_sc_hd__nor2_1 U20016 ( .A(n17842), .B(n17795), .Y(n17849) );
  sky130_fd_sc_hd__nand2_1 U20017 ( .A(n17756), .B(n17548), .Y(n17495) );
  sky130_fd_sc_hd__nand4_1 U20018 ( .A(n17912), .B(n17771), .C(n18399), .D(
        n18430), .Y(n17552) );
  sky130_fd_sc_hd__nor3_1 U20019 ( .A(n17916), .B(n17943), .C(n17552), .Y(
        n15006) );
  sky130_fd_sc_hd__a31oi_1 U20020 ( .A1(n17849), .A2(n17845), .A3(n15006), 
        .B1(n18439), .Y(n15014) );
  sky130_fd_sc_hd__nor2_1 U20021 ( .A(n17774), .B(n17866), .Y(n17591) );
  sky130_fd_sc_hd__nor2_1 U20022 ( .A(n17592), .B(n18397), .Y(n17848) );
  sky130_fd_sc_hd__nor4b_1 U20023 ( .D_N(n17848), .A(n17498), .B(n17795), .C(
        n15007), .Y(n17440) );
  sky130_fd_sc_hd__nor2_1 U20024 ( .A(n17624), .B(n17795), .Y(n17735) );
  sky130_fd_sc_hd__nand2_1 U20025 ( .A(n17502), .B(n17618), .Y(n17517) );
  sky130_fd_sc_hd__a21oi_1 U20026 ( .A1(n15010), .A2(n15009), .B1(n15008), .Y(
        n17616) );
  sky130_fd_sc_hd__a21oi_1 U20027 ( .A1(n17930), .A2(n17931), .B1(n17616), .Y(
        n16746) );
  sky130_fd_sc_hd__nand2_1 U20028 ( .A(n16746), .B(n15011), .Y(n17443) );
  sky130_fd_sc_hd__nor4b_1 U20029 ( .D_N(n17735), .A(n17517), .B(n17495), .C(
        n17443), .Y(n15012) );
  sky130_fd_sc_hd__o22ai_1 U20030 ( .A1(n17440), .A2(n18423), .B1(n15012), 
        .B2(n18445), .Y(n15013) );
  sky130_fd_sc_hd__nor3_1 U20031 ( .A(n15015), .B(n15014), .C(n15013), .Y(
        n15029) );
  sky130_fd_sc_hd__nand3_1 U20032 ( .A(n15019), .B(n15018), .C(n15017), .Y(
        n15020) );
  sky130_fd_sc_hd__nand2_1 U20033 ( .A(n17779), .B(n17771), .Y(n17529) );
  sky130_fd_sc_hd__nand2_1 U20034 ( .A(n17757), .B(n17791), .Y(n17420) );
  sky130_fd_sc_hd__nor3_1 U20035 ( .A(n17529), .B(n17420), .C(n17556), .Y(
        n15021) );
  sky130_fd_sc_hd__a21oi_1 U20036 ( .A1(n15022), .A2(n15021), .B1(n18445), .Y(
        n15027) );
  sky130_fd_sc_hd__nor2_1 U20037 ( .A(n18418), .B(n17842), .Y(n17724) );
  sky130_fd_sc_hd__nand2_1 U20038 ( .A(n17875), .B(n18345), .Y(n17725) );
  sky130_fd_sc_hd__nor2_1 U20039 ( .A(n17725), .B(n15036), .Y(n17524) );
  sky130_fd_sc_hd__a31oi_1 U20040 ( .A1(n17724), .A2(n17524), .A3(n17534), 
        .B1(n18423), .Y(n15026) );
  sky130_fd_sc_hd__o31a_1 U20041 ( .A1(n17759), .A2(n17928), .A3(n18435), .B1(
        n17543), .X(n15025) );
  sky130_fd_sc_hd__nand3_1 U20042 ( .A(n17653), .B(n17923), .C(n17618), .Y(
        n17783) );
  sky130_fd_sc_hd__nand2_1 U20043 ( .A(n17591), .B(n17623), .Y(n17516) );
  sky130_fd_sc_hd__nor2_1 U20044 ( .A(n17783), .B(n17516), .Y(n17445) );
  sky130_fd_sc_hd__nand2_1 U20045 ( .A(n17478), .B(n17617), .Y(n17864) );
  sky130_fd_sc_hd__nor4_1 U20046 ( .A(n17604), .B(n17593), .C(n17624), .D(
        n17864), .Y(n15023) );
  sky130_fd_sc_hd__a21oi_1 U20047 ( .A1(n17445), .A2(n15023), .B1(n18439), .Y(
        n15024) );
  sky130_fd_sc_hd__nor4_1 U20048 ( .A(n15027), .B(n15026), .C(n15025), .D(
        n15024), .Y(n15028) );
  sky130_fd_sc_hd__o22ai_1 U20049 ( .A1(n15029), .A2(n18722), .B1(n15028), 
        .B2(n18552), .Y(n15061) );
  sky130_fd_sc_hd__nand2_1 U20050 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[66]), .B(n18727), .Y(
        n15035) );
  sky130_fd_sc_hd__a22oi_1 U20051 ( .A1(n18724), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[98]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[34]), .Y(n15034) );
  sky130_fd_sc_hd__a22oi_1 U20052 ( .A1(n18242), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[10]), .B1(n18243), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[2]), .Y(n15031) );
  sky130_fd_sc_hd__a22oi_1 U20053 ( .A1(n18244), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[18]), .B1(n18241), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[26]), .Y(n15030) );
  sky130_fd_sc_hd__a21oi_1 U20054 ( .A1(n15031), .A2(n15030), .B1(n18245), .Y(
        n15032) );
  sky130_fd_sc_hd__a21oi_1 U20055 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[2]), .B1(n15032), .Y(
        n15033) );
  sky130_fd_sc_hd__nand3_1 U20056 ( .A(n15035), .B(n15034), .C(n15033), .Y(
        n15060) );
  sky130_fd_sc_hd__nor2_1 U20057 ( .A(n17537), .B(n17552), .Y(n17479) );
  sky130_fd_sc_hd__a21oi_1 U20058 ( .A1(n18402), .A2(n17479), .B1(n18437), .Y(
        n15042) );
  sky130_fd_sc_hd__nor2_1 U20059 ( .A(n18436), .B(n17624), .Y(n15037) );
  sky130_fd_sc_hd__nor3_1 U20060 ( .A(n17600), .B(n17943), .C(n15036), .Y(
        n17514) );
  sky130_fd_sc_hd__a31oi_1 U20061 ( .A1(n15037), .A2(n17514), .A3(n17768), 
        .B1(n18439), .Y(n15041) );
  sky130_fd_sc_hd__nor2_1 U20062 ( .A(n17752), .B(n17944), .Y(n17622) );
  sky130_fd_sc_hd__nand2_1 U20063 ( .A(n17534), .B(n17791), .Y(n17942) );
  sky130_fd_sc_hd__nand2_1 U20064 ( .A(n17622), .B(n17656), .Y(n17555) );
  sky130_fd_sc_hd__nor4b_1 U20065 ( .D_N(n15037), .A(n17529), .B(n17870), .C(
        n17555), .Y(n15039) );
  sky130_fd_sc_hd__nor2_1 U20066 ( .A(n17941), .B(n17725), .Y(n18428) );
  sky130_fd_sc_hd__nand2_1 U20067 ( .A(n18428), .B(n18399), .Y(n17444) );
  sky130_fd_sc_hd__nor2_1 U20068 ( .A(n17444), .B(n17942), .Y(n15038) );
  sky130_fd_sc_hd__o22ai_1 U20069 ( .A1(n15039), .A2(n18445), .B1(n15038), 
        .B2(n18423), .Y(n15040) );
  sky130_fd_sc_hd__nor3_1 U20070 ( .A(n15042), .B(n15041), .C(n15040), .Y(
        n15058) );
  sky130_fd_sc_hd__a22o_1 U20071 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[2]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[66]), .X(n15043) );
  sky130_fd_sc_hd__a21oi_1 U20072 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[98]), .B1(n15043), .Y(n15045) );
  sky130_fd_sc_hd__a22oi_1 U20073 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[162]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[130]), .Y(n15044) );
  sky130_fd_sc_hd__a21oi_1 U20074 ( .A1(n15045), .A2(n15044), .B1(n18736), .Y(
        n15056) );
  sky130_fd_sc_hd__a22oi_1 U20075 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[258]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[34]), .Y(n15054) );
  sky130_fd_sc_hd__a22o_1 U20076 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[290]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[322]), .X(n15046) );
  sky130_fd_sc_hd__a21oi_1 U20077 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[354]), .B1(n15046), .Y(n15053) );
  sky130_fd_sc_hd__nand2_1 U20078 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[226]), .Y(n15050) );
  sky130_fd_sc_hd__a21oi_1 U20079 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[450]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n15049) );
  sky130_fd_sc_hd__nand2_1 U20080 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[386]), .Y(n15048) );
  sky130_fd_sc_hd__nand2_1 U20081 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[418]), .Y(n15047) );
  sky130_fd_sc_hd__nand4_1 U20082 ( .A(n15050), .B(n15049), .C(n15048), .D(
        n15047), .Y(n15051) );
  sky130_fd_sc_hd__a21oi_1 U20083 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[194]), .B1(n15051), .Y(n15052) );
  sky130_fd_sc_hd__nand3_1 U20084 ( .A(n15054), .B(n15053), .C(n15052), .Y(
        n15055) );
  sky130_fd_sc_hd__o22ai_1 U20085 ( .A1(j202_soc_core_memory0_ram_dout0[482]), 
        .A2(n18758), .B1(n15056), .B2(n15055), .Y(n15057) );
  sky130_fd_sc_hd__o22ai_1 U20086 ( .A1(n15058), .A2(n18720), .B1(n18761), 
        .B2(n15057), .Y(n15059) );
  sky130_fd_sc_hd__nor4_1 U20087 ( .A(n15062), .B(n15061), .C(n15060), .D(
        n15059), .Y(n15072) );
  sky130_fd_sc_hd__nor2_1 U20088 ( .A(n15065), .B(n19742), .Y(n25159) );
  sky130_fd_sc_hd__nor2_1 U20089 ( .A(n15064), .B(n15063), .Y(n17711) );
  sky130_fd_sc_hd__nand2_1 U20090 ( .A(n17427), .B(
        j202_soc_core_bldc_core_00_comm[2]), .Y(n15068) );
  sky130_fd_sc_hd__nand2_1 U20091 ( .A(n17716), .B(j202_soc_core_aquc_ADR__3_), 
        .Y(n15066) );
  sky130_fd_sc_hd__nor2_1 U20092 ( .A(n15066), .B(n15065), .Y(n17715) );
  sky130_fd_sc_hd__nand2_1 U20093 ( .A(n17715), .B(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[2]), .Y(n15067) );
  sky130_fd_sc_hd__nand2_1 U20094 ( .A(n15068), .B(n15067), .Y(n15070) );
  sky130_fd_sc_hd__a22oi_1 U20095 ( .A1(n18629), .A2(
        j202_soc_core_bldc_core_00_pwm_period[2]), .B1(n15070), .B2(n15069), 
        .Y(n15071) );
  sky130_fd_sc_hd__nand2_1 U20096 ( .A(n15072), .B(n15071), .Y(n25246) );
  sky130_fd_sc_hd__nand2_1 U20097 ( .A(n15075), .B(n15074), .Y(n15078) );
  sky130_fd_sc_hd__o21ai_1 U20098 ( .A1(n17824), .A2(n17828), .B1(n17825), .Y(
        n15077) );
  sky130_fd_sc_hd__xnor2_1 U20099 ( .A(n15078), .B(n15077), .Y(n22262) );
  sky130_fd_sc_hd__nand2_1 U20100 ( .A(n22262), .B(n19729), .Y(n15084) );
  sky130_fd_sc_hd__ha_1 U20101 ( .A(j202_soc_core_j22_cpu_pc[2]), .B(
        j202_soc_core_j22_cpu_pc[1]), .COUT(n17836), .SUM(n22259) );
  sky130_fd_sc_hd__o22ai_1 U20102 ( .A1(n22267), .A2(n19078), .B1(n22487), 
        .B2(n19731), .Y(n15079) );
  sky130_fd_sc_hd__a21oi_1 U20103 ( .A1(n19080), .A2(n22181), .B1(n15079), .Y(
        n15081) );
  sky130_fd_sc_hd__nand2_1 U20104 ( .A(n19517), .B(n22259), .Y(n15080) );
  sky130_fd_sc_hd__o211ai_1 U20105 ( .A1(n22264), .A2(n19083), .B1(n15081), 
        .C1(n15080), .Y(n15082) );
  sky130_fd_sc_hd__a21oi_1 U20106 ( .A1(n25246), .A2(n19737), .B1(n15082), .Y(
        n15083) );
  sky130_fd_sc_hd__nand2_1 U20107 ( .A(n15084), .B(n15083), .Y(n25333) );
  sky130_fd_sc_hd__nor2_1 U20108 ( .A(n18512), .B(n18597), .Y(n16889) );
  sky130_fd_sc_hd__nand2_1 U20109 ( .A(n16889), .B(n18713), .Y(n18678) );
  sky130_fd_sc_hd__nor4_1 U20110 ( .A(n16987), .B(n16924), .C(n18678), .D(
        n15085), .Y(n15086) );
  sky130_fd_sc_hd__nand3_1 U20111 ( .A(n18574), .B(n15086), .C(n18662), .Y(
        n18601) );
  sky130_fd_sc_hd__nand2_1 U20112 ( .A(n18522), .B(n15087), .Y(n18790) );
  sky130_fd_sc_hd__nand2_1 U20113 ( .A(n18681), .B(n18588), .Y(n18685) );
  sky130_fd_sc_hd__nor4_1 U20114 ( .A(n18645), .B(n18512), .C(n18584), .D(
        n18685), .Y(n15088) );
  sky130_fd_sc_hd__o22ai_1 U20115 ( .A1(n18589), .A2(n18783), .B1(n15088), 
        .B2(n18792), .Y(n15089) );
  sky130_fd_sc_hd__a21oi_1 U20116 ( .A1(n18655), .A2(n18601), .B1(n15089), .Y(
        n15092) );
  sky130_fd_sc_hd__nor2_1 U20117 ( .A(n16741), .B(n15090), .Y(n16896) );
  sky130_fd_sc_hd__o21ai_1 U20118 ( .A1(n15186), .A2(n16896), .B1(n18664), .Y(
        n15091) );
  sky130_fd_sc_hd__a21oi_1 U20119 ( .A1(n15092), .A2(n15091), .B1(n18666), .Y(
        n15135) );
  sky130_fd_sc_hd__nand2_1 U20120 ( .A(n18555), .B(n18680), .Y(n18672) );
  sky130_fd_sc_hd__nor2_1 U20121 ( .A(n18770), .B(n18672), .Y(n18544) );
  sky130_fd_sc_hd__a21oi_1 U20122 ( .A1(n15093), .A2(n18534), .B1(n16987), .Y(
        n18538) );
  sky130_fd_sc_hd__nand3_1 U20123 ( .A(n18544), .B(n18538), .C(n16901), .Y(
        n18778) );
  sky130_fd_sc_hd__nor3_1 U20124 ( .A(n18645), .B(n18702), .C(n18769), .Y(
        n18604) );
  sky130_fd_sc_hd__nand2_1 U20125 ( .A(n18559), .B(n18698), .Y(n18511) );
  sky130_fd_sc_hd__nor2_1 U20126 ( .A(n18703), .B(n18511), .Y(n18781) );
  sky130_fd_sc_hd__nand2_1 U20127 ( .A(n18593), .B(n18675), .Y(n18602) );
  sky130_fd_sc_hd__nand2b_1 U20128 ( .A_N(n18602), .B(n16916), .Y(n15094) );
  sky130_fd_sc_hd__nor4_1 U20129 ( .A(n18687), .B(n18250), .C(n16924), .D(
        n15094), .Y(n15095) );
  sky130_fd_sc_hd__a31oi_1 U20130 ( .A1(n18604), .A2(n18781), .A3(n15095), 
        .B1(n18771), .Y(n15100) );
  sky130_fd_sc_hd__nand2_1 U20131 ( .A(n18559), .B(n18662), .Y(n18322) );
  sky130_fd_sc_hd__nand4_1 U20132 ( .A(n18291), .B(n18675), .C(n15122), .D(
        n18588), .Y(n18697) );
  sky130_fd_sc_hd__nor3_1 U20133 ( .A(n18790), .B(n18322), .C(n18697), .Y(
        n15098) );
  sky130_fd_sc_hd__nor3_1 U20134 ( .A(n18557), .B(n15186), .C(n18644), .Y(
        n15136) );
  sky130_fd_sc_hd__nor2_1 U20135 ( .A(n18564), .B(n18540), .Y(n18648) );
  sky130_fd_sc_hd__and4b_1 U20136 ( .B(n15136), .C(n18648), .D(n18558), .A_N(
        n15096), .X(n15097) );
  sky130_fd_sc_hd__o22ai_1 U20137 ( .A1(n15098), .A2(n18779), .B1(n15097), 
        .B2(n18783), .Y(n15099) );
  sky130_fd_sc_hd__a211oi_1 U20138 ( .A1(n18651), .A2(n18778), .B1(n15100), 
        .C1(n15099), .Y(n15116) );
  sky130_fd_sc_hd__a22oi_1 U20139 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[239]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[207]), .Y(n15104) );
  sky130_fd_sc_hd__a22oi_1 U20140 ( .A1(n18734), .A2(
        j202_soc_core_memory0_ram_dout0[143]), .B1(n18733), .B2(
        j202_soc_core_memory0_ram_dout0[111]), .Y(n15103) );
  sky130_fd_sc_hd__a22oi_1 U20141 ( .A1(n18361), .A2(
        j202_soc_core_memory0_ram_dout0[47]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[79]), .Y(n15102) );
  sky130_fd_sc_hd__nand2_1 U20142 ( .A(n18735), .B(
        j202_soc_core_memory0_ram_dout0[175]), .Y(n15101) );
  sky130_fd_sc_hd__nand4_1 U20143 ( .A(n15104), .B(n15103), .C(n15102), .D(
        n15101), .Y(n15105) );
  sky130_fd_sc_hd__a21oi_1 U20144 ( .A1(n18367), .A2(
        j202_soc_core_memory0_ram_dout0[15]), .B1(n15105), .Y(n15113) );
  sky130_fd_sc_hd__a22oi_1 U20145 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[303]), .B1(n18062), .B2(
        j202_soc_core_memory0_ram_dout0[271]), .Y(n15112) );
  sky130_fd_sc_hd__nand2_1 U20146 ( .A(n18743), .B(
        j202_soc_core_memory0_ram_dout0[367]), .Y(n15109) );
  sky130_fd_sc_hd__a21oi_1 U20147 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[463]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n15108) );
  sky130_fd_sc_hd__nand2_1 U20148 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[399]), .Y(n15107) );
  sky130_fd_sc_hd__nand2_1 U20149 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[431]), .Y(n15106) );
  sky130_fd_sc_hd__nand4_1 U20150 ( .A(n15109), .B(n15108), .C(n15107), .D(
        n15106), .Y(n15110) );
  sky130_fd_sc_hd__a21oi_1 U20151 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[335]), .B1(n15110), .Y(n15111) );
  sky130_fd_sc_hd__o211ai_1 U20152 ( .A1(n18736), .A2(n15113), .B1(n15112), 
        .C1(n15111), .Y(n15114) );
  sky130_fd_sc_hd__o22ai_1 U20154 ( .A1(n15116), .A2(n18720), .B1(n18761), 
        .B2(n15115), .Y(n15134) );
  sky130_fd_sc_hd__nand2_1 U20155 ( .A(n18698), .B(n18675), .Y(n18323) );
  sky130_fd_sc_hd__nand3_1 U20156 ( .A(n18514), .B(n16977), .C(n15184), .Y(
        n15198) );
  sky130_fd_sc_hd__nor4_1 U20157 ( .A(n18323), .B(n16976), .C(n15117), .D(
        n15198), .Y(n15120) );
  sky130_fd_sc_hd__nand2_1 U20158 ( .A(n16974), .B(n18291), .Y(n18562) );
  sky130_fd_sc_hd__nor2_1 U20159 ( .A(n18770), .B(n18527), .Y(n18520) );
  sky130_fd_sc_hd__nand2_1 U20160 ( .A(n18520), .B(n18593), .Y(n16930) );
  sky130_fd_sc_hd__nor4_1 U20161 ( .A(n18766), .B(n15118), .C(n18562), .D(
        n16930), .Y(n15119) );
  sky130_fd_sc_hd__o22ai_1 U20162 ( .A1(n15120), .A2(n18792), .B1(n15119), 
        .B2(n18779), .Y(n15128) );
  sky130_fd_sc_hd__nor2_1 U20163 ( .A(n18250), .B(n15121), .Y(n18573) );
  sky130_fd_sc_hd__and4_1 U20164 ( .A(n18661), .B(n15189), .C(n18514), .D(
        n16901), .X(n18566) );
  sky130_fd_sc_hd__nand2_1 U20165 ( .A(n18566), .B(n18592), .Y(n18583) );
  sky130_fd_sc_hd__nor3b_1 U20166 ( .C_N(n18573), .A(n18685), .B(n18583), .Y(
        n15126) );
  sky130_fd_sc_hd__nand2_1 U20167 ( .A(n15122), .B(n18588), .Y(n15124) );
  sky130_fd_sc_hd__nand2_1 U20168 ( .A(n18559), .B(n18289), .Y(n15123) );
  sky130_fd_sc_hd__nor4_1 U20169 ( .A(n18641), .B(n18672), .C(n15124), .D(
        n15123), .Y(n15125) );
  sky130_fd_sc_hd__o22ai_1 U20170 ( .A1(n15126), .A2(n18783), .B1(n15125), 
        .B2(n18771), .Y(n15127) );
  sky130_fd_sc_hd__nor2_1 U20171 ( .A(n15128), .B(n15127), .Y(n15129) );
  sky130_fd_sc_hd__o22ai_1 U20172 ( .A1(n15129), .A2(n18552), .B1(n18759), 
        .B2(n25188), .Y(n15133) );
  sky130_fd_sc_hd__a22oi_1 U20173 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[15]), .B1(n18724), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[111]), .Y(n15131) );
  sky130_fd_sc_hd__a22oi_1 U20174 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[79]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[47]), .Y(n15130) );
  sky130_fd_sc_hd__nand2_1 U20175 ( .A(n15131), .B(n15130), .Y(n15132) );
  sky130_fd_sc_hd__nor4_1 U20176 ( .A(n15135), .B(n15134), .C(n15133), .D(
        n15132), .Y(n15148) );
  sky130_fd_sc_hd__nor3_1 U20177 ( .A(n18253), .B(n18673), .C(n18702), .Y(
        n18537) );
  sky130_fd_sc_hd__nand4_1 U20178 ( .A(n18537), .B(n18267), .C(n18573), .D(
        n15136), .Y(n15139) );
  sky130_fd_sc_hd__nor4_1 U20179 ( .A(n18703), .B(n18585), .C(n18512), .D(
        n18775), .Y(n15137) );
  sky130_fd_sc_hd__a31oi_1 U20180 ( .A1(n18292), .A2(n15137), .A3(n18661), 
        .B1(n18783), .Y(n15138) );
  sky130_fd_sc_hd__a21o_1 U20181 ( .A1(n18651), .A2(n15139), .B1(n15138), .X(
        n15146) );
  sky130_fd_sc_hd__nand4_1 U20182 ( .A(n18292), .B(n18574), .C(n18588), .D(
        n18522), .Y(n16989) );
  sky130_fd_sc_hd__nand2_1 U20183 ( .A(n16974), .B(n18681), .Y(n18670) );
  sky130_fd_sc_hd__nor3_1 U20184 ( .A(n18709), .B(n16989), .C(n18670), .Y(
        n15144) );
  sky130_fd_sc_hd__nand3_1 U20185 ( .A(n16916), .B(n18554), .C(n18713), .Y(
        n15141) );
  sky130_fd_sc_hd__nor3_1 U20186 ( .A(n18557), .B(n16924), .C(n15182), .Y(
        n18659) );
  sky130_fd_sc_hd__nand2_1 U20187 ( .A(n18659), .B(n18698), .Y(n18686) );
  sky130_fd_sc_hd__nor4_1 U20188 ( .A(n15142), .B(n18641), .C(n15141), .D(
        n18686), .Y(n15143) );
  sky130_fd_sc_hd__o22ai_1 U20189 ( .A1(n15144), .A2(n18771), .B1(n15143), 
        .B2(n18779), .Y(n15145) );
  sky130_fd_sc_hd__nand2_1 U20191 ( .A(n15148), .B(n15147), .Y(n25388) );
  sky130_fd_sc_hd__nor2_1 U20192 ( .A(n16924), .B(n15182), .Y(n18270) );
  sky130_fd_sc_hd__nor2b_1 U20193 ( .B_N(n18534), .A(n15149), .Y(n16897) );
  sky130_fd_sc_hd__nor2_1 U20194 ( .A(n18766), .B(n16897), .Y(n16915) );
  sky130_fd_sc_hd__nor2_1 U20195 ( .A(n16898), .B(n18674), .Y(n15150) );
  sky130_fd_sc_hd__nand4_1 U20196 ( .A(n18270), .B(n16915), .C(n15150), .D(
        n18698), .Y(n15157) );
  sky130_fd_sc_hd__a31oi_1 U20197 ( .A1(n15152), .A2(n15151), .A3(n16901), 
        .B1(n18771), .Y(n15156) );
  sky130_fd_sc_hd__nor4_1 U20198 ( .A(n16898), .B(n15153), .C(n16983), .D(
        n16896), .Y(n15155) );
  sky130_fd_sc_hd__a211oi_1 U20201 ( .A1(n18651), .A2(n15157), .B1(n15156), 
        .C1(n16891), .Y(n15158) );
  sky130_fd_sc_hd__o22ai_1 U20202 ( .A1(n15158), .A2(n18722), .B1(n18759), 
        .B2(n25180), .Y(n15180) );
  sky130_fd_sc_hd__a22o_1 U20203 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[7]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[71]), .X(n15159) );
  sky130_fd_sc_hd__a21oi_1 U20204 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[103]), .B1(n15159), .Y(n15161) );
  sky130_fd_sc_hd__a22oi_1 U20205 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[167]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[135]), .Y(n15160) );
  sky130_fd_sc_hd__a21oi_1 U20206 ( .A1(n15161), .A2(n15160), .B1(n18736), .Y(
        n15172) );
  sky130_fd_sc_hd__a22oi_1 U20207 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[263]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[39]), .Y(n15170) );
  sky130_fd_sc_hd__a22o_1 U20208 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[295]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[327]), .X(n15162) );
  sky130_fd_sc_hd__a21oi_1 U20209 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[359]), .B1(n15162), .Y(n15169) );
  sky130_fd_sc_hd__nand2_1 U20210 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[231]), .Y(n15166) );
  sky130_fd_sc_hd__a21oi_1 U20211 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[455]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n15165) );
  sky130_fd_sc_hd__nand2_1 U20212 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[391]), .Y(n15164) );
  sky130_fd_sc_hd__nand2_1 U20213 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[423]), .Y(n15163) );
  sky130_fd_sc_hd__nand4_1 U20214 ( .A(n15166), .B(n15165), .C(n15164), .D(
        n15163), .Y(n15167) );
  sky130_fd_sc_hd__a21oi_1 U20215 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[199]), .B1(n15167), .Y(n15168) );
  sky130_fd_sc_hd__nand3_1 U20216 ( .A(n15170), .B(n15169), .C(n15168), .Y(
        n15171) );
  sky130_fd_sc_hd__o22ai_1 U20217 ( .A1(j202_soc_core_memory0_ram_dout0[487]), 
        .A2(n18758), .B1(n15172), .B2(n15171), .Y(n15178) );
  sky130_fd_sc_hd__a22oi_1 U20218 ( .A1(n18242), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[15]), .B1(n18244), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[23]), .Y(n15174) );
  sky130_fd_sc_hd__a22oi_1 U20219 ( .A1(n18241), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[31]), .B1(n18243), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[7]), .Y(n15173) );
  sky130_fd_sc_hd__a21oi_1 U20220 ( .A1(n15174), .A2(n15173), .B1(n18245), .Y(
        n15175) );
  sky130_fd_sc_hd__a21oi_1 U20221 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[7]), .B1(n15175), .Y(
        n15177) );
  sky130_fd_sc_hd__a22oi_1 U20222 ( .A1(n18724), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[103]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[39]), .Y(n15176) );
  sky130_fd_sc_hd__o211ai_1 U20223 ( .A1(n18761), .A2(n15178), .B1(n15177), 
        .C1(n15176), .Y(n15179) );
  sky130_fd_sc_hd__a211oi_1 U20224 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[71]), .B1(n15180), .C1(
        n15179), .Y(n15211) );
  sky130_fd_sc_hd__nor2_1 U20225 ( .A(n18256), .B(n18770), .Y(n16988) );
  sky130_fd_sc_hd__nor4_1 U20226 ( .A(n18709), .B(n15182), .C(n17001), .D(
        n15181), .Y(n15188) );
  sky130_fd_sc_hd__nand2_1 U20227 ( .A(n18642), .B(n18680), .Y(n18767) );
  sky130_fd_sc_hd__nor2_1 U20228 ( .A(n18767), .B(n18777), .Y(n15183) );
  sky130_fd_sc_hd__nand3_1 U20229 ( .A(n15183), .B(n18514), .C(n18639), .Y(
        n18315) );
  sky130_fd_sc_hd__nand2b_1 U20230 ( .A_N(n18315), .B(n15184), .Y(n15185) );
  sky130_fd_sc_hd__nor4_1 U20231 ( .A(n15186), .B(n18512), .C(n18568), .D(
        n15185), .Y(n15187) );
  sky130_fd_sc_hd__o22ai_1 U20232 ( .A1(n15188), .A2(n18771), .B1(n15187), 
        .B2(n18779), .Y(n15193) );
  sky130_fd_sc_hd__nand2_1 U20233 ( .A(n15189), .B(n18680), .Y(n18299) );
  sky130_fd_sc_hd__nor3_1 U20234 ( .A(n18250), .B(n18299), .C(n18273), .Y(
        n15190) );
  sky130_fd_sc_hd__o22ai_1 U20235 ( .A1(n15191), .A2(n18783), .B1(n15190), 
        .B2(n18792), .Y(n15192) );
  sky130_fd_sc_hd__o21ai_1 U20236 ( .A1(n15193), .A2(n15192), .B1(n18798), .Y(
        n15210) );
  sky130_fd_sc_hd__nor2_1 U20237 ( .A(n18644), .B(n16924), .Y(n18321) );
  sky130_fd_sc_hd__a21oi_1 U20238 ( .A1(n18321), .A2(n18291), .B1(n18771), .Y(
        n15203) );
  sky130_fd_sc_hd__nor2_1 U20239 ( .A(n18645), .B(n16896), .Y(n18652) );
  sky130_fd_sc_hd__and3_1 U20240 ( .A(n18652), .B(n18698), .C(n16977), .X(
        n15205) );
  sky130_fd_sc_hd__nand2_1 U20241 ( .A(n18784), .B(n18660), .Y(n18776) );
  sky130_fd_sc_hd__nor3_1 U20242 ( .A(n18673), .B(n18568), .C(n18776), .Y(
        n15195) );
  sky130_fd_sc_hd__a31oi_1 U20243 ( .A1(n15205), .A2(n18520), .A3(n15195), 
        .B1(n18792), .Y(n15202) );
  sky130_fd_sc_hd__nand2_1 U20244 ( .A(n16990), .B(n18698), .Y(n15196) );
  sky130_fd_sc_hd__nor4_1 U20245 ( .A(n18670), .B(n15198), .C(n15197), .D(
        n15196), .Y(n15200) );
  sky130_fd_sc_hd__o22ai_1 U20246 ( .A1(n15200), .A2(n18779), .B1(n18783), 
        .B2(n15199), .Y(n15201) );
  sky130_fd_sc_hd__o31ai_1 U20247 ( .A1(n15203), .A2(n15202), .A3(n15201), 
        .B1(n17609), .Y(n15209) );
  sky130_fd_sc_hd__o22ai_1 U20248 ( .A1(n15205), .A2(n18783), .B1(n15204), 
        .B2(n18792), .Y(n16921) );
  sky130_fd_sc_hd__o21ai_1 U20250 ( .A1(n18252), .A2(n18779), .B1(n15206), .Y(
        n15207) );
  sky130_fd_sc_hd__nand4_1 U20252 ( .A(n15211), .B(n15210), .C(n15209), .D(
        n15208), .Y(n25247) );
  sky130_fd_sc_hd__nor2_1 U20253 ( .A(n23240), .B(n19917), .Y(n21222) );
  sky130_fd_sc_hd__nor2_1 U20254 ( .A(n21222), .B(n19379), .Y(n19317) );
  sky130_fd_sc_hd__nand2_1 U20255 ( .A(n15216), .B(n15212), .Y(n19977) );
  sky130_fd_sc_hd__clkinv_1 U20256 ( .A(n19977), .Y(n16812) );
  sky130_fd_sc_hd__nor2_1 U20257 ( .A(n15214), .B(n15213), .Y(n19985) );
  sky130_fd_sc_hd__a22oi_1 U20258 ( .A1(n16812), .A2(
        j202_soc_core_j22_cpu_pc[15]), .B1(n19985), .B2(
        j202_soc_core_j22_cpu_rf_vbr[15]), .Y(n15226) );
  sky130_fd_sc_hd__nand2_1 U20259 ( .A(n15216), .B(n15215), .Y(n19975) );
  sky130_fd_sc_hd__o22a_1 U20260 ( .A1(n15218), .A2(n19971), .B1(n15217), .B2(
        n19975), .X(n15225) );
  sky130_fd_sc_hd__nand2_1 U20261 ( .A(n15219), .B(n15220), .Y(n19981) );
  sky130_fd_sc_hd__nand2b_1 U20262 ( .A_N(n15221), .B(n15220), .Y(n19986) );
  sky130_fd_sc_hd__a2bb2oi_1 U20263 ( .B1(j202_soc_core_j22_cpu_rf_tmp[15]), 
        .B2(n19843), .A1_N(n15222), .A2_N(n19986), .Y(n15224) );
  sky130_fd_sc_hd__nand2_1 U20264 ( .A(n19842), .B(
        j202_soc_core_j22_cpu_rf_gpr[15]), .Y(n15223) );
  sky130_fd_sc_hd__nand4_1 U20265 ( .A(n15226), .B(n15225), .C(n15224), .D(
        n15223), .Y(n15227) );
  sky130_fd_sc_hd__a21oi_1 U20266 ( .A1(n15228), .A2(n19969), .B1(n15227), .Y(
        n19649) );
  sky130_fd_sc_hd__xnor2_1 U20267 ( .A(j202_soc_core_j22_cpu_ml_bufa[27]), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .Y(n15402) );
  sky130_fd_sc_hd__xor2_1 U20268 ( .A(j202_soc_core_j22_cpu_ml_bufa[28]), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n15403) );
  sky130_fd_sc_hd__nand2b_1 U20269 ( .A_N(n15402), .B(n15403), .Y(n16551) );
  sky130_fd_sc_hd__nand2_1 U20270 ( .A(j202_soc_core_j22_cpu_ml_bufb[0]), .B(
        j202_soc_core_j22_cpu_ml_bufb[1]), .Y(n15370) );
  sky130_fd_sc_hd__nand2_1 U20271 ( .A(n15229), .B(n15370), .Y(n16164) );
  sky130_fd_sc_hd__nor2_1 U20272 ( .A(n15402), .B(n15403), .Y(n16549) );
  sky130_fd_sc_hd__xnor2_1 U20273 ( .A(j202_soc_core_j22_cpu_ml_bufa[28]), .B(
        j202_soc_core_j22_cpu_ml_bufa[27]), .Y(n15401) );
  sky130_fd_sc_hd__nor2b_1 U20274 ( .B_N(n15402), .A(n15401), .Y(n16548) );
  sky130_fd_sc_hd__a22oi_1 U20275 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15230) );
  sky130_fd_sc_hd__o21ai_1 U20276 ( .A1(n16551), .A2(n16164), .B1(n15230), .Y(
        n15231) );
  sky130_fd_sc_hd__xor2_1 U20277 ( .A(n15231), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16195) );
  sky130_fd_sc_hd__nand2b_1 U20278 ( .A_N(n15233), .B(n15235), .Y(n16599) );
  sky130_fd_sc_hd__nand2b_1 U20279 ( .A_N(n21723), .B(n15234), .Y(n16592) );
  sky130_fd_sc_hd__nor2_1 U20280 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[4]), .B(n15235), .Y(n15238) );
  sky130_fd_sc_hd__nand2_1 U20282 ( .A(n15240), .B(n15239), .Y(n15243) );
  sky130_fd_sc_hd__nand2_1 U20283 ( .A(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[0]), .Y(n21724) );
  sky130_fd_sc_hd__o21ai_1 U20284 ( .A1(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .A2(n21724), .B1(n15241), 
        .Y(n15242) );
  sky130_fd_sc_hd__nand2_1 U20285 ( .A(n15243), .B(n15242), .Y(n16593) );
  sky130_fd_sc_hd__nor2_1 U20286 ( .A(j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]), .B(j202_soc_core_j22_cpu_ml_X_macop_MAC_[4]), .Y(n16590) );
  sky130_fd_sc_hd__o22ai_1 U20287 ( .A1(n16191), .A2(n17039), .B1(n15804), 
        .B2(n16189), .Y(n15407) );
  sky130_fd_sc_hd__xnor2_1 U20288 ( .A(j202_soc_core_j22_cpu_ml_bufa[24]), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .Y(n15249) );
  sky130_fd_sc_hd__xor2_1 U20289 ( .A(j202_soc_core_j22_cpu_ml_bufa[25]), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n15250) );
  sky130_fd_sc_hd__nand2b_1 U20290 ( .A_N(n15249), .B(n15250), .Y(n16373) );
  sky130_fd_sc_hd__nor2_1 U20291 ( .A(j202_soc_core_j22_cpu_ml_bufb[4]), .B(
        j202_soc_core_j22_cpu_ml_bufb[3]), .Y(n15268) );
  sky130_fd_sc_hd__nand2_1 U20292 ( .A(j202_soc_core_j22_cpu_ml_bufb[3]), .B(
        j202_soc_core_j22_cpu_ml_bufb[4]), .Y(n15344) );
  sky130_fd_sc_hd__nand2_1 U20293 ( .A(n15346), .B(n15344), .Y(n15247) );
  sky130_fd_sc_hd__nand2_1 U20294 ( .A(j202_soc_core_j22_cpu_ml_bufb[2]), .B(
        j202_soc_core_j22_cpu_ml_bufb[3]), .Y(n15263) );
  sky130_fd_sc_hd__nand2_1 U20295 ( .A(j202_soc_core_j22_cpu_ml_bufb[2]), .B(
        j202_soc_core_j22_cpu_ml_bufb[1]), .Y(n15369) );
  sky130_fd_sc_hd__nand2_1 U20296 ( .A(n15263), .B(n15369), .Y(n15245) );
  sky130_fd_sc_hd__a21oi_1 U20297 ( .A1(n11196), .A2(n15246), .B1(n15245), .Y(
        n15272) );
  sky130_fd_sc_hd__xor2_1 U20298 ( .A(n15247), .B(n15347), .X(n16193) );
  sky130_fd_sc_hd__nor2_1 U20299 ( .A(n15249), .B(n15250), .Y(n16371) );
  sky130_fd_sc_hd__xnor2_1 U20300 ( .A(j202_soc_core_j22_cpu_ml_bufa[25]), .B(
        j202_soc_core_j22_cpu_ml_bufa[24]), .Y(n15248) );
  sky130_fd_sc_hd__nor2b_1 U20301 ( .B_N(n15249), .A(n15248), .Y(n16370) );
  sky130_fd_sc_hd__and3_1 U20302 ( .A(n15250), .B(n15249), .C(n15248), .X(
        n16369) );
  sky130_fd_sc_hd__a222oi_1 U20303 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .Y(n15251) );
  sky130_fd_sc_hd__o21ai_1 U20304 ( .A1(n16373), .A2(n16193), .B1(n15251), .Y(
        n15252) );
  sky130_fd_sc_hd__xor2_1 U20305 ( .A(n15252), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n15406) );
  sky130_fd_sc_hd__nand2_1 U20306 ( .A(n16549), .B(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15253) );
  sky130_fd_sc_hd__o21ai_1 U20307 ( .A1(n15962), .A2(n16551), .B1(n15253), .Y(
        n15254) );
  sky130_fd_sc_hd__xor2_1 U20308 ( .A(n15254), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n15360) );
  sky130_fd_sc_hd__a22oi_1 U20309 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15255) );
  sky130_fd_sc_hd__o21ai_1 U20310 ( .A1(n16373), .A2(n16164), .B1(n15255), .Y(
        n15256) );
  sky130_fd_sc_hd__xor2_1 U20311 ( .A(n15256), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n15368) );
  sky130_fd_sc_hd__xnor2_1 U20312 ( .A(j202_soc_core_j22_cpu_ml_bufa[9]), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .Y(n15258) );
  sky130_fd_sc_hd__xor2_1 U20313 ( .A(j202_soc_core_j22_cpu_ml_bufa[10]), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15259) );
  sky130_fd_sc_hd__nand2b_1 U20314 ( .A_N(n15258), .B(n15259), .Y(n16046) );
  sky130_fd_sc_hd__nor2_1 U20315 ( .A(n15258), .B(n15259), .Y(n16044) );
  sky130_fd_sc_hd__xnor2_1 U20316 ( .A(j202_soc_core_j22_cpu_ml_bufa[10]), .B(
        j202_soc_core_j22_cpu_ml_bufa[9]), .Y(n15257) );
  sky130_fd_sc_hd__nor2b_1 U20317 ( .B_N(n15258), .A(n15257), .Y(n16043) );
  sky130_fd_sc_hd__and3_1 U20318 ( .A(n15259), .B(n15258), .C(n15257), .X(
        n16042) );
  sky130_fd_sc_hd__a222oi_1 U20319 ( .A1(n16044), .A2(n11170), .B1(n16043), 
        .B2(n11170), .C1(n16042), .C2(n11170), .Y(n15260) );
  sky130_fd_sc_hd__o21ai_1 U20320 ( .A1(n11169), .A2(n16046), .B1(n15260), .Y(
        n15261) );
  sky130_fd_sc_hd__xnor2_1 U20321 ( .A(j202_soc_core_j22_cpu_ml_bufa[11]), .B(
        n15261), .Y(n15442) );
  sky130_fd_sc_hd__o22ai_1 U20322 ( .A1(n16191), .A2(n15262), .B1(n15853), 
        .B2(n16189), .Y(n15441) );
  sky130_fd_sc_hd__nand2_1 U20323 ( .A(n11196), .B(n15263), .Y(n15265) );
  sky130_fd_sc_hd__nand2_1 U20324 ( .A(n15369), .B(n15370), .Y(n15264) );
  sky130_fd_sc_hd__xor2_1 U20325 ( .A(n15265), .B(n15264), .X(n16159) );
  sky130_fd_sc_hd__a222oi_1 U20326 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .Y(n15266) );
  sky130_fd_sc_hd__o21ai_1 U20327 ( .A1(n16373), .A2(n16159), .B1(n15266), .Y(
        n15267) );
  sky130_fd_sc_hd__xor2_1 U20328 ( .A(n15267), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n15440) );
  sky130_fd_sc_hd__xnor2_1 U20329 ( .A(j202_soc_core_j22_cpu_ml_bufa[18]), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .Y(n15280) );
  sky130_fd_sc_hd__xor2_1 U20330 ( .A(j202_soc_core_j22_cpu_ml_bufa[19]), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n15278) );
  sky130_fd_sc_hd__nand2b_1 U20331 ( .A_N(n15280), .B(n15278), .Y(n16265) );
  sky130_fd_sc_hd__nor2_1 U20332 ( .A(j202_soc_core_j22_cpu_ml_bufb[10]), .B(
        j202_soc_core_j22_cpu_ml_bufb[9]), .Y(n15284) );
  sky130_fd_sc_hd__nand2_1 U20333 ( .A(j202_soc_core_j22_cpu_ml_bufb[9]), .B(
        j202_soc_core_j22_cpu_ml_bufb[10]), .Y(n15391) );
  sky130_fd_sc_hd__nand2_1 U20334 ( .A(n15393), .B(n15391), .Y(n15277) );
  sky130_fd_sc_hd__nor2_1 U20335 ( .A(j202_soc_core_j22_cpu_ml_bufb[9]), .B(
        j202_soc_core_j22_cpu_ml_bufb[8]), .Y(n15430) );
  sky130_fd_sc_hd__nor2_1 U20336 ( .A(j202_soc_core_j22_cpu_ml_bufb[7]), .B(
        j202_soc_core_j22_cpu_ml_bufb[8]), .Y(n15435) );
  sky130_fd_sc_hd__nor2_1 U20337 ( .A(n15430), .B(n15435), .Y(n15390) );
  sky130_fd_sc_hd__nor2_1 U20338 ( .A(j202_soc_core_j22_cpu_ml_bufb[4]), .B(
        j202_soc_core_j22_cpu_ml_bufb[5]), .Y(n15348) );
  sky130_fd_sc_hd__nor2_1 U20339 ( .A(n15268), .B(n15348), .Y(n15301) );
  sky130_fd_sc_hd__nor2_1 U20340 ( .A(j202_soc_core_j22_cpu_ml_bufb[7]), .B(
        j202_soc_core_j22_cpu_ml_bufb[6]), .Y(n15297) );
  sky130_fd_sc_hd__nor2_1 U20341 ( .A(j202_soc_core_j22_cpu_ml_bufb[6]), .B(
        j202_soc_core_j22_cpu_ml_bufb[5]), .Y(n15361) );
  sky130_fd_sc_hd__nor2_1 U20342 ( .A(n15297), .B(n15361), .Y(n15270) );
  sky130_fd_sc_hd__nand2_1 U20343 ( .A(n15301), .B(n15270), .Y(n15273) );
  sky130_fd_sc_hd__nand2_1 U20344 ( .A(j202_soc_core_j22_cpu_ml_bufb[5]), .B(
        j202_soc_core_j22_cpu_ml_bufb[4]), .Y(n15349) );
  sky130_fd_sc_hd__nand2_1 U20345 ( .A(n15349), .B(n15344), .Y(n15300) );
  sky130_fd_sc_hd__nand2_1 U20346 ( .A(j202_soc_core_j22_cpu_ml_bufb[6]), .B(
        j202_soc_core_j22_cpu_ml_bufb[7]), .Y(n15298) );
  sky130_fd_sc_hd__nand2_1 U20347 ( .A(j202_soc_core_j22_cpu_ml_bufb[5]), .B(
        j202_soc_core_j22_cpu_ml_bufb[6]), .Y(n15362) );
  sky130_fd_sc_hd__nand2_1 U20348 ( .A(n15298), .B(n15362), .Y(n15269) );
  sky130_fd_sc_hd__a21oi_1 U20349 ( .A1(n15300), .A2(n15270), .B1(n15269), .Y(
        n15271) );
  sky130_fd_sc_hd__nand2_1 U20351 ( .A(j202_soc_core_j22_cpu_ml_bufb[8]), .B(
        j202_soc_core_j22_cpu_ml_bufb[9]), .Y(n15431) );
  sky130_fd_sc_hd__nand2_1 U20352 ( .A(j202_soc_core_j22_cpu_ml_bufb[8]), .B(
        j202_soc_core_j22_cpu_ml_bufb[7]), .Y(n15433) );
  sky130_fd_sc_hd__nand2_1 U20353 ( .A(n15431), .B(n15433), .Y(n15394) );
  sky130_fd_sc_hd__o21ai_1 U20354 ( .A1(n15275), .A2(n15434), .B1(n15274), .Y(
        n15276) );
  sky130_fd_sc_hd__xor2_1 U20355 ( .A(n15277), .B(n15276), .X(n16354) );
  sky130_fd_sc_hd__nor2_1 U20356 ( .A(n15278), .B(n15280), .Y(n16263) );
  sky130_fd_sc_hd__xnor2_1 U20357 ( .A(j202_soc_core_j22_cpu_ml_bufa[19]), .B(
        j202_soc_core_j22_cpu_ml_bufa[18]), .Y(n15279) );
  sky130_fd_sc_hd__nor2b_1 U20358 ( .B_N(n15280), .A(n15279), .Y(n16262) );
  sky130_fd_sc_hd__and3_1 U20359 ( .A(n15280), .B(n15279), .C(n15278), .X(
        n16261) );
  sky130_fd_sc_hd__a222oi_1 U20360 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .Y(n15281) );
  sky130_fd_sc_hd__o21ai_1 U20361 ( .A1(n16265), .A2(n16354), .B1(n15281), .Y(
        n15282) );
  sky130_fd_sc_hd__xor2_1 U20362 ( .A(n15282), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n15326) );
  sky130_fd_sc_hd__xnor2_1 U20363 ( .A(j202_soc_core_j22_cpu_ml_bufa[15]), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .Y(n15293) );
  sky130_fd_sc_hd__xor2_1 U20364 ( .A(j202_soc_core_j22_cpu_ml_bufa[16]), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n15294) );
  sky130_fd_sc_hd__nand2b_1 U20365 ( .A_N(n15293), .B(n15294), .Y(n16227) );
  sky130_fd_sc_hd__nor2_1 U20366 ( .A(j202_soc_core_j22_cpu_ml_bufb[13]), .B(
        j202_soc_core_j22_cpu_ml_bufb[12]), .Y(n15310) );
  sky130_fd_sc_hd__nand2_1 U20367 ( .A(j202_soc_core_j22_cpu_ml_bufb[12]), .B(
        j202_soc_core_j22_cpu_ml_bufb[13]), .Y(n15311) );
  sky130_fd_sc_hd__nand2_1 U20368 ( .A(n15283), .B(n15311), .Y(n15291) );
  sky130_fd_sc_hd__nor2_1 U20369 ( .A(j202_soc_core_j22_cpu_ml_bufb[10]), .B(
        j202_soc_core_j22_cpu_ml_bufb[11]), .Y(n15387) );
  sky130_fd_sc_hd__nor2_1 U20370 ( .A(n15284), .B(n15387), .Y(n15286) );
  sky130_fd_sc_hd__nand2_1 U20371 ( .A(n15390), .B(n15286), .Y(n15335) );
  sky130_fd_sc_hd__nor2_1 U20372 ( .A(j202_soc_core_j22_cpu_ml_bufb[12]), .B(
        j202_soc_core_j22_cpu_ml_bufb[11]), .Y(n15309) );
  sky130_fd_sc_hd__nand2_1 U20373 ( .A(n15416), .B(n15333), .Y(n15289) );
  sky130_fd_sc_hd__nand2_1 U20374 ( .A(j202_soc_core_j22_cpu_ml_bufb[11]), .B(
        j202_soc_core_j22_cpu_ml_bufb[10]), .Y(n15388) );
  sky130_fd_sc_hd__nand2_1 U20375 ( .A(n15388), .B(n15391), .Y(n15285) );
  sky130_fd_sc_hd__a21oi_1 U20376 ( .A1(n15394), .A2(n15286), .B1(n15285), .Y(
        n15334) );
  sky130_fd_sc_hd__nand2_1 U20377 ( .A(j202_soc_core_j22_cpu_ml_bufb[11]), .B(
        j202_soc_core_j22_cpu_ml_bufb[12]), .Y(n15332) );
  sky130_fd_sc_hd__a21oi_1 U20378 ( .A1(n15423), .A2(n15333), .B1(n15287), .Y(
        n15288) );
  sky130_fd_sc_hd__o21ai_1 U20379 ( .A1(n15289), .A2(n15434), .B1(n15288), .Y(
        n15290) );
  sky130_fd_sc_hd__xor2_1 U20380 ( .A(n15291), .B(n15290), .X(n16402) );
  sky130_fd_sc_hd__nor2_1 U20381 ( .A(n15293), .B(n15294), .Y(n16225) );
  sky130_fd_sc_hd__xnor2_1 U20382 ( .A(j202_soc_core_j22_cpu_ml_bufa[16]), .B(
        j202_soc_core_j22_cpu_ml_bufa[15]), .Y(n15292) );
  sky130_fd_sc_hd__nor2b_1 U20383 ( .B_N(n15293), .A(n15292), .Y(n16224) );
  sky130_fd_sc_hd__and3_1 U20384 ( .A(n15294), .B(n15293), .C(n15292), .X(
        n16223) );
  sky130_fd_sc_hd__a222oi_1 U20385 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .Y(n15295) );
  sky130_fd_sc_hd__o21ai_1 U20386 ( .A1(n16227), .A2(n16402), .B1(n15295), .Y(
        n15296) );
  sky130_fd_sc_hd__xor2_1 U20387 ( .A(n15296), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n15331) );
  sky130_fd_sc_hd__xnor2_1 U20388 ( .A(j202_soc_core_j22_cpu_ml_bufa[20]), .B(
        j202_soc_core_j22_cpu_ml_bufa[21]), .Y(n15304) );
  sky130_fd_sc_hd__xor2_1 U20389 ( .A(j202_soc_core_j22_cpu_ml_bufa[22]), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n15306) );
  sky130_fd_sc_hd__nand2b_1 U20390 ( .A_N(n15304), .B(n15306), .Y(n16327) );
  sky130_fd_sc_hd__nand2_1 U20391 ( .A(n15299), .B(n15298), .Y(n15303) );
  sky130_fd_sc_hd__a21oi_1 U20392 ( .A1(n15347), .A2(n15301), .B1(n15300), .Y(
        n15365) );
  sky130_fd_sc_hd__xor2_1 U20394 ( .A(n15303), .B(n15302), .X(n16305) );
  sky130_fd_sc_hd__nor2_1 U20395 ( .A(n15304), .B(n15306), .Y(n16325) );
  sky130_fd_sc_hd__xnor2_1 U20396 ( .A(j202_soc_core_j22_cpu_ml_bufa[22]), .B(
        j202_soc_core_j22_cpu_ml_bufa[21]), .Y(n15305) );
  sky130_fd_sc_hd__nor2b_1 U20397 ( .B_N(n15304), .A(n15305), .Y(n16324) );
  sky130_fd_sc_hd__and3_1 U20398 ( .A(n15306), .B(n15305), .C(n15304), .X(
        n16323) );
  sky130_fd_sc_hd__a222oi_1 U20399 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .Y(n15307) );
  sky130_fd_sc_hd__o21ai_1 U20400 ( .A1(n16327), .A2(n16305), .B1(n15307), .Y(
        n15308) );
  sky130_fd_sc_hd__xor2_1 U20401 ( .A(n15308), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n15330) );
  sky130_fd_sc_hd__xnor2_1 U20402 ( .A(j202_soc_core_j22_cpu_ml_bufa[12]), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .Y(n15322) );
  sky130_fd_sc_hd__xor2_1 U20403 ( .A(j202_soc_core_j22_cpu_ml_bufa[13]), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15323) );
  sky130_fd_sc_hd__nand2b_1 U20404 ( .A_N(n15322), .B(n15323), .Y(n16052) );
  sky130_fd_sc_hd__nor2_1 U20405 ( .A(j202_soc_core_j22_cpu_ml_bufb[15]), .B(
        j202_soc_core_j22_cpu_ml_bufb[14]), .Y(n15411) );
  sky130_fd_sc_hd__nor2_1 U20406 ( .A(j202_soc_core_j22_cpu_ml_bufb[13]), .B(
        j202_soc_core_j22_cpu_ml_bufb[14]), .Y(n15420) );
  sky130_fd_sc_hd__nor2_1 U20407 ( .A(n15411), .B(n15420), .Y(n15313) );
  sky130_fd_sc_hd__nor2_1 U20408 ( .A(n15310), .B(n15309), .Y(n15414) );
  sky130_fd_sc_hd__nand2_1 U20409 ( .A(n15313), .B(n15414), .Y(n15315) );
  sky130_fd_sc_hd__nor2_1 U20410 ( .A(n15315), .B(n15335), .Y(n15317) );
  sky130_fd_sc_hd__nand2_1 U20411 ( .A(n15311), .B(n15332), .Y(n15417) );
  sky130_fd_sc_hd__nand2_1 U20412 ( .A(j202_soc_core_j22_cpu_ml_bufb[14]), .B(
        j202_soc_core_j22_cpu_ml_bufb[15]), .Y(n15412) );
  sky130_fd_sc_hd__nand2_1 U20413 ( .A(j202_soc_core_j22_cpu_ml_bufb[14]), .B(
        j202_soc_core_j22_cpu_ml_bufb[13]), .Y(n15418) );
  sky130_fd_sc_hd__nand2_1 U20414 ( .A(n15412), .B(n15418), .Y(n15312) );
  sky130_fd_sc_hd__a21oi_1 U20415 ( .A1(n15313), .A2(n15417), .B1(n15312), .Y(
        n15314) );
  sky130_fd_sc_hd__o21ai_1 U20416 ( .A1(n15315), .A2(n15334), .B1(n15314), .Y(
        n15316) );
  sky130_fd_sc_hd__a21oi_1 U20417 ( .A1(n15318), .A2(n15317), .B1(n15316), .Y(
        n15356) );
  sky130_fd_sc_hd__nor2_1 U20418 ( .A(j202_soc_core_j22_cpu_ml_bufb[15]), .B(
        n11170), .Y(n15357) );
  sky130_fd_sc_hd__nand2_1 U20419 ( .A(n11170), .B(
        j202_soc_core_j22_cpu_ml_bufb[15]), .Y(n15355) );
  sky130_fd_sc_hd__nand2_1 U20420 ( .A(n15319), .B(n15355), .Y(n15320) );
  sky130_fd_sc_hd__xnor2_1 U20421 ( .A(n15356), .B(n15320), .Y(n16537) );
  sky130_fd_sc_hd__nor2_1 U20422 ( .A(n15322), .B(n15323), .Y(n16050) );
  sky130_fd_sc_hd__xnor2_1 U20423 ( .A(j202_soc_core_j22_cpu_ml_bufa[13]), .B(
        j202_soc_core_j22_cpu_ml_bufa[12]), .Y(n15321) );
  sky130_fd_sc_hd__nor2b_1 U20424 ( .B_N(n15322), .A(n15321), .Y(n16049) );
  sky130_fd_sc_hd__and3_1 U20425 ( .A(n15323), .B(n15322), .C(n15321), .X(
        n16048) );
  sky130_fd_sc_hd__a222oi_1 U20426 ( .A1(n16050), .A2(n11170), .B1(n16049), 
        .B2(j202_soc_core_j22_cpu_ml_bufb[15]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .Y(n15324) );
  sky130_fd_sc_hd__xor2_1 U20428 ( .A(n15325), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15329) );
  sky130_fd_sc_hd__fa_1 U20429 ( .A(n15328), .B(n15327), .CIN(n15326), .COUT(
        n15471), .SUM(n15508) );
  sky130_fd_sc_hd__fa_1 U20430 ( .A(n15331), .B(n15330), .CIN(n15329), .COUT(
        n15470), .SUM(n15507) );
  sky130_fd_sc_hd__nand2_1 U20431 ( .A(n15333), .B(n15332), .Y(n15337) );
  sky130_fd_sc_hd__xor2_1 U20433 ( .A(n15337), .B(n15336), .X(n16367) );
  sky130_fd_sc_hd__a222oi_1 U20434 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .Y(n15338) );
  sky130_fd_sc_hd__xor2_1 U20436 ( .A(n15339), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n15514) );
  sky130_fd_sc_hd__nand2_1 U20437 ( .A(n15340), .B(n15433), .Y(n15341) );
  sky130_fd_sc_hd__xnor2_1 U20438 ( .A(n15434), .B(n15341), .Y(n16311) );
  sky130_fd_sc_hd__a222oi_1 U20439 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .Y(n15342) );
  sky130_fd_sc_hd__o21ai_1 U20440 ( .A1(n16265), .A2(n16311), .B1(n15342), .Y(
        n15343) );
  sky130_fd_sc_hd__xor2_1 U20441 ( .A(n15343), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n15517) );
  sky130_fd_sc_hd__a21oi_1 U20442 ( .A1(n15347), .A2(n15346), .B1(n15345), .Y(
        n15352) );
  sky130_fd_sc_hd__nand2_1 U20443 ( .A(n15350), .B(n15349), .Y(n15351) );
  sky130_fd_sc_hd__xnor2_1 U20444 ( .A(n15352), .B(n15351), .Y(n16247) );
  sky130_fd_sc_hd__a222oi_1 U20445 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .Y(n15353) );
  sky130_fd_sc_hd__o21ai_1 U20446 ( .A1(n16327), .A2(n16247), .B1(n15353), .Y(
        n15354) );
  sky130_fd_sc_hd__xor2_1 U20447 ( .A(n15354), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n15516) );
  sky130_fd_sc_hd__o21a_1 U20448 ( .A1(n15357), .A2(n15356), .B1(n15355), .X(
        n16584) );
  sky130_fd_sc_hd__a222oi_1 U20449 ( .A1(n16044), .A2(n11170), .B1(n16043), 
        .B2(n11170), .C1(n16042), .C2(j202_soc_core_j22_cpu_ml_bufb[15]), .Y(
        n15358) );
  sky130_fd_sc_hd__xor2_1 U20451 ( .A(n15359), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15515) );
  sky130_fd_sc_hd__fa_1 U20452 ( .A(j202_soc_core_j22_cpu_ml_bufa[29]), .B(
        n15360), .CIN(n15368), .COUT(n15328), .SUM(n15410) );
  sky130_fd_sc_hd__nand2_1 U20453 ( .A(n15363), .B(n15362), .Y(n15364) );
  sky130_fd_sc_hd__xnor2_1 U20454 ( .A(n15365), .B(n15364), .Y(n16278) );
  sky130_fd_sc_hd__a222oi_1 U20455 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .Y(n15366) );
  sky130_fd_sc_hd__o21ai_1 U20456 ( .A1(n16327), .A2(n16278), .B1(n15366), .Y(
        n15367) );
  sky130_fd_sc_hd__xor2_1 U20457 ( .A(n15367), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n15409) );
  sky130_fd_sc_hd__nand2_1 U20458 ( .A(n11198), .B(n15369), .Y(n15371) );
  sky130_fd_sc_hd__xnor2_1 U20459 ( .A(n15371), .B(n15370), .Y(n16168) );
  sky130_fd_sc_hd__a222oi_1 U20460 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15372) );
  sky130_fd_sc_hd__xor2_1 U20462 ( .A(n15373), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n15481) );
  sky130_fd_sc_hd__o22ai_1 U20463 ( .A1(n16191), .A2(n16798), .B1(n15841), 
        .B2(n16189), .Y(n15480) );
  sky130_fd_sc_hd__a222oi_1 U20464 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .Y(n15374) );
  sky130_fd_sc_hd__o21ai_1 U20465 ( .A1(n16327), .A2(n16311), .B1(n15374), .Y(
        n15375) );
  sky130_fd_sc_hd__xor2_1 U20466 ( .A(n15375), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n15447) );
  sky130_fd_sc_hd__a222oi_1 U20467 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .Y(n15376) );
  sky130_fd_sc_hd__o21ai_1 U20468 ( .A1(n16373), .A2(n16247), .B1(n15376), .Y(
        n15377) );
  sky130_fd_sc_hd__xor2_1 U20469 ( .A(n15377), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n15446) );
  sky130_fd_sc_hd__a222oi_1 U20470 ( .A1(n16050), .A2(n11170), .B1(n16049), 
        .B2(n11170), .C1(n16048), .C2(j202_soc_core_j22_cpu_ml_bufb[15]), .Y(
        n15378) );
  sky130_fd_sc_hd__o21ai_1 U20471 ( .A1(n16052), .A2(n16584), .B1(n15378), .Y(
        n15379) );
  sky130_fd_sc_hd__xor2_1 U20472 ( .A(n15379), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15445) );
  sky130_fd_sc_hd__nand2_1 U20473 ( .A(n15380), .B(n15418), .Y(n15384) );
  sky130_fd_sc_hd__nand2_1 U20474 ( .A(n15416), .B(n15414), .Y(n15382) );
  sky130_fd_sc_hd__a21oi_1 U20475 ( .A1(n15423), .A2(n15414), .B1(n15417), .Y(
        n15381) );
  sky130_fd_sc_hd__o21ai_1 U20476 ( .A1(n15382), .A2(n15434), .B1(n15381), .Y(
        n15383) );
  sky130_fd_sc_hd__xor2_1 U20477 ( .A(n15384), .B(n15383), .X(n16557) );
  sky130_fd_sc_hd__a222oi_1 U20478 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .Y(n15385) );
  sky130_fd_sc_hd__o21ai_1 U20479 ( .A1(n16227), .A2(n16557), .B1(n15385), .Y(
        n15386) );
  sky130_fd_sc_hd__xor2_1 U20480 ( .A(n15386), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n15460) );
  sky130_fd_sc_hd__nand2_1 U20481 ( .A(n15389), .B(n15388), .Y(n15398) );
  sky130_fd_sc_hd__nand2_1 U20482 ( .A(n15390), .B(n15393), .Y(n15396) );
  sky130_fd_sc_hd__a21oi_1 U20483 ( .A1(n15394), .A2(n15393), .B1(n15392), .Y(
        n15395) );
  sky130_fd_sc_hd__o21ai_1 U20484 ( .A1(n15396), .A2(n15434), .B1(n15395), .Y(
        n15397) );
  sky130_fd_sc_hd__xor2_1 U20485 ( .A(n15398), .B(n15397), .X(n16379) );
  sky130_fd_sc_hd__a222oi_1 U20486 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .Y(n15399) );
  sky130_fd_sc_hd__o21ai_1 U20487 ( .A1(n16265), .A2(n16379), .B1(n15399), .Y(
        n15400) );
  sky130_fd_sc_hd__xor2_1 U20488 ( .A(n15400), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n15459) );
  sky130_fd_sc_hd__and3_1 U20489 ( .A(n15403), .B(n15402), .C(n15401), .X(
        n16547) );
  sky130_fd_sc_hd__a222oi_1 U20490 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15404) );
  sky130_fd_sc_hd__xor2_1 U20492 ( .A(n15405), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n15453) );
  sky130_fd_sc_hd__o22ai_1 U20493 ( .A1(n16191), .A2(n19104), .B1(n15796), 
        .B2(n16189), .Y(n15452) );
  sky130_fd_sc_hd__fa_1 U20494 ( .A(n15454), .B(n15407), .CIN(n15406), .COUT(
        n15472), .SUM(n15475) );
  sky130_fd_sc_hd__fa_1 U20495 ( .A(n15410), .B(n15409), .CIN(n15408), .COUT(
        n15474), .SUM(n15512) );
  sky130_fd_sc_hd__nand2_1 U20496 ( .A(n15413), .B(n15412), .Y(n15427) );
  sky130_fd_sc_hd__nor2_1 U20497 ( .A(n15420), .B(n15415), .Y(n15422) );
  sky130_fd_sc_hd__nand2_1 U20498 ( .A(n15422), .B(n15416), .Y(n15425) );
  sky130_fd_sc_hd__a21oi_1 U20500 ( .A1(n15423), .A2(n15422), .B1(n15421), .Y(
        n15424) );
  sky130_fd_sc_hd__xor2_1 U20502 ( .A(n15427), .B(n15426), .X(n16540) );
  sky130_fd_sc_hd__a222oi_1 U20503 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[15]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .Y(n15428) );
  sky130_fd_sc_hd__o21ai_1 U20504 ( .A1(n16052), .A2(n16540), .B1(n15428), .Y(
        n15429) );
  sky130_fd_sc_hd__xor2_1 U20505 ( .A(n15429), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15484) );
  sky130_fd_sc_hd__nand2_1 U20506 ( .A(n15432), .B(n15431), .Y(n15437) );
  sky130_fd_sc_hd__o21ai_1 U20507 ( .A1(n15435), .A2(n15434), .B1(n15433), .Y(
        n15436) );
  sky130_fd_sc_hd__xor2_1 U20508 ( .A(n15437), .B(n15436), .X(n16319) );
  sky130_fd_sc_hd__a222oi_1 U20509 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .Y(n15438) );
  sky130_fd_sc_hd__o21ai_1 U20510 ( .A1(n16265), .A2(n16319), .B1(n15438), .Y(
        n15439) );
  sky130_fd_sc_hd__xor2_1 U20511 ( .A(n15439), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n15483) );
  sky130_fd_sc_hd__fa_1 U20512 ( .A(n15442), .B(n15441), .CIN(n15440), .COUT(
        n15327), .SUM(n15482) );
  sky130_fd_sc_hd__a222oi_1 U20513 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .Y(n15443) );
  sky130_fd_sc_hd__xor2_1 U20515 ( .A(n15444), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n16454) );
  sky130_fd_sc_hd__fa_1 U20516 ( .A(n15447), .B(n15446), .CIN(n15445), .COUT(
        n16453), .SUM(n15457) );
  sky130_fd_sc_hd__xnor2_1 U20517 ( .A(j202_soc_core_j22_cpu_ml_bufa[30]), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .Y(n16157) );
  sky130_fd_sc_hd__xor2_1 U20518 ( .A(j202_soc_core_j22_cpu_ml_bufa[31]), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16155) );
  sky130_fd_sc_hd__nor2_1 U20519 ( .A(n16155), .B(n16157), .Y(n19334) );
  sky130_fd_sc_hd__nand2_1 U20520 ( .A(n19334), .B(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15448) );
  sky130_fd_sc_hd__o21ai_1 U20521 ( .A1(n15962), .A2(n19336), .B1(n15448), .Y(
        n15449) );
  sky130_fd_sc_hd__xor2_1 U20522 ( .A(n15449), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16196) );
  sky130_fd_sc_hd__a222oi_1 U20523 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .Y(n15450) );
  sky130_fd_sc_hd__o21ai_1 U20524 ( .A1(n16373), .A2(n16278), .B1(n15450), .Y(
        n15451) );
  sky130_fd_sc_hd__xor2_1 U20525 ( .A(n15451), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n16438) );
  sky130_fd_sc_hd__fa_1 U20526 ( .A(n15454), .B(n15453), .CIN(n15452), .COUT(
        n16437), .SUM(n15458) );
  sky130_fd_sc_hd__fa_1 U20527 ( .A(n15457), .B(n15456), .CIN(n15455), .COUT(
        n16432), .SUM(n15509) );
  sky130_fd_sc_hd__fa_1 U20528 ( .A(n15460), .B(n15459), .CIN(n15458), .COUT(
        n16445), .SUM(n15456) );
  sky130_fd_sc_hd__a222oi_1 U20529 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[15]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .Y(n15461) );
  sky130_fd_sc_hd__o21ai_1 U20530 ( .A1(n16227), .A2(n16540), .B1(n15461), .Y(
        n15462) );
  sky130_fd_sc_hd__xor2_1 U20531 ( .A(n15462), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n16442) );
  sky130_fd_sc_hd__a222oi_1 U20532 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .Y(n15463) );
  sky130_fd_sc_hd__o21ai_1 U20533 ( .A1(n16327), .A2(n16319), .B1(n15463), .Y(
        n15464) );
  sky130_fd_sc_hd__xor2_1 U20534 ( .A(n15464), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n16441) );
  sky130_fd_sc_hd__a222oi_1 U20535 ( .A1(n16050), .A2(n11170), .B1(n16049), 
        .B2(n11170), .C1(n16048), .C2(n11170), .Y(n15465) );
  sky130_fd_sc_hd__o21ai_1 U20536 ( .A1(n11169), .A2(n16052), .B1(n15465), .Y(
        n15466) );
  sky130_fd_sc_hd__xnor2_1 U20537 ( .A(j202_soc_core_j22_cpu_ml_bufa[14]), .B(
        n15466), .Y(n16199) );
  sky130_fd_sc_hd__o22ai_1 U20538 ( .A1(n16191), .A2(n15467), .B1(n15709), 
        .B2(n16189), .Y(n16198) );
  sky130_fd_sc_hd__a222oi_1 U20539 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .Y(n15468) );
  sky130_fd_sc_hd__xor2_1 U20541 ( .A(n15469), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16197) );
  sky130_fd_sc_hd__fa_1 U20542 ( .A(n15472), .B(n15471), .CIN(n15470), .COUT(
        n16443), .SUM(n15511) );
  sky130_fd_sc_hd__nor2_1 U20543 ( .A(n16145), .B(n16146), .Y(n18979) );
  sky130_fd_sc_hd__fa_1 U20544 ( .A(n15475), .B(n15474), .CIN(n15473), .COUT(
        n15455), .SUM(n15542) );
  sky130_fd_sc_hd__a222oi_1 U20545 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .Y(n15476) );
  sky130_fd_sc_hd__o21ai_1 U20546 ( .A1(n16052), .A2(n16557), .B1(n15476), .Y(
        n15477) );
  sky130_fd_sc_hd__xor2_1 U20547 ( .A(n15477), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15520) );
  sky130_fd_sc_hd__a222oi_1 U20548 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .Y(n15478) );
  sky130_fd_sc_hd__xor2_1 U20550 ( .A(n15479), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n15519) );
  sky130_fd_sc_hd__fa_1 U20551 ( .A(n15523), .B(n15481), .CIN(n15480), .COUT(
        n15408), .SUM(n15518) );
  sky130_fd_sc_hd__fa_1 U20552 ( .A(n15484), .B(n15483), .CIN(n15482), .COUT(
        n15473), .SUM(n15538) );
  sky130_fd_sc_hd__o22ai_1 U20553 ( .A1(n16191), .A2(n20006), .B1(n15894), 
        .B2(n16189), .Y(n15522) );
  sky130_fd_sc_hd__a222oi_1 U20554 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .Y(n15485) );
  sky130_fd_sc_hd__o21ai_1 U20555 ( .A1(n16327), .A2(n16193), .B1(n15485), .Y(
        n15486) );
  sky130_fd_sc_hd__xor2_1 U20556 ( .A(n15486), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n15521) );
  sky130_fd_sc_hd__nand2_1 U20557 ( .A(n16371), .B(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15487) );
  sky130_fd_sc_hd__xor2_1 U20559 ( .A(n15488), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n15524) );
  sky130_fd_sc_hd__a22oi_1 U20560 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15489) );
  sky130_fd_sc_hd__xor2_1 U20562 ( .A(n15490), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n15527) );
  sky130_fd_sc_hd__xnor2_1 U20563 ( .A(j202_soc_core_j22_cpu_ml_bufa[6]), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .Y(n15492) );
  sky130_fd_sc_hd__xor2_1 U20564 ( .A(j202_soc_core_j22_cpu_ml_bufa[7]), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15493) );
  sky130_fd_sc_hd__nand2b_1 U20565 ( .A_N(n15492), .B(n15493), .Y(n16067) );
  sky130_fd_sc_hd__nor2_1 U20566 ( .A(n15492), .B(n15493), .Y(n16065) );
  sky130_fd_sc_hd__xnor2_1 U20567 ( .A(j202_soc_core_j22_cpu_ml_bufa[7]), .B(
        j202_soc_core_j22_cpu_ml_bufa[6]), .Y(n15491) );
  sky130_fd_sc_hd__nor2b_1 U20568 ( .B_N(n15492), .A(n15491), .Y(n16064) );
  sky130_fd_sc_hd__and3_1 U20569 ( .A(n15493), .B(n15492), .C(n15491), .X(
        n16063) );
  sky130_fd_sc_hd__a222oi_1 U20570 ( .A1(n16065), .A2(n11170), .B1(n16064), 
        .B2(n11170), .C1(n16063), .C2(n11170), .Y(n15494) );
  sky130_fd_sc_hd__o21ai_1 U20571 ( .A1(n11169), .A2(n16067), .B1(n15494), .Y(
        n15495) );
  sky130_fd_sc_hd__xnor2_1 U20572 ( .A(j202_soc_core_j22_cpu_ml_bufa[8]), .B(
        n15495), .Y(n15536) );
  sky130_fd_sc_hd__o22ai_1 U20573 ( .A1(n16191), .A2(n19303), .B1(n15880), 
        .B2(n16189), .Y(n15535) );
  sky130_fd_sc_hd__a222oi_1 U20574 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .Y(n15496) );
  sky130_fd_sc_hd__xor2_1 U20576 ( .A(n15497), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n15534) );
  sky130_fd_sc_hd__a222oi_1 U20577 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .Y(n15498) );
  sky130_fd_sc_hd__o21ai_1 U20578 ( .A1(n16227), .A2(n16354), .B1(n15498), .Y(
        n15499) );
  sky130_fd_sc_hd__xor2_1 U20579 ( .A(n15499), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n15546) );
  sky130_fd_sc_hd__a222oi_1 U20580 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .Y(n15500) );
  sky130_fd_sc_hd__o21ai_1 U20581 ( .A1(n16052), .A2(n16402), .B1(n15500), .Y(
        n15501) );
  sky130_fd_sc_hd__xor2_1 U20582 ( .A(n15501), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15551) );
  sky130_fd_sc_hd__a222oi_1 U20583 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .Y(n15502) );
  sky130_fd_sc_hd__o21ai_1 U20584 ( .A1(n16265), .A2(n16305), .B1(n15502), .Y(
        n15503) );
  sky130_fd_sc_hd__xor2_1 U20585 ( .A(n15503), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n15550) );
  sky130_fd_sc_hd__a222oi_1 U20586 ( .A1(n16044), .A2(n11170), .B1(n16043), 
        .B2(j202_soc_core_j22_cpu_ml_bufb[15]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .Y(n15504) );
  sky130_fd_sc_hd__xor2_1 U20588 ( .A(n15505), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15549) );
  sky130_fd_sc_hd__fa_1 U20589 ( .A(n15508), .B(n15507), .CIN(n15506), .COUT(
        n15510), .SUM(n15540) );
  sky130_fd_sc_hd__fa_1 U20590 ( .A(n15511), .B(n15510), .CIN(n15509), .COUT(
        n16145), .SUM(n16144) );
  sky130_fd_sc_hd__nor2_1 U20591 ( .A(n16143), .B(n16144), .Y(n18977) );
  sky130_fd_sc_hd__nor2_1 U20592 ( .A(n18979), .B(n18977), .Y(n16148) );
  sky130_fd_sc_hd__fa_1 U20593 ( .A(n15514), .B(n15513), .CIN(n15512), .COUT(
        n15506), .SUM(n15568) );
  sky130_fd_sc_hd__fa_1 U20594 ( .A(n15517), .B(n15516), .CIN(n15515), .COUT(
        n15513), .SUM(n15565) );
  sky130_fd_sc_hd__fa_1 U20595 ( .A(n15520), .B(n15519), .CIN(n15518), .COUT(
        n15539), .SUM(n15564) );
  sky130_fd_sc_hd__fa_1 U20596 ( .A(n15523), .B(n15522), .CIN(n15521), .COUT(
        n15545), .SUM(n15685) );
  sky130_fd_sc_hd__fa_1 U20597 ( .A(j202_soc_core_j22_cpu_ml_bufa[26]), .B(
        n15524), .CIN(n15527), .COUT(n15548), .SUM(n15562) );
  sky130_fd_sc_hd__a222oi_1 U20598 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .Y(n15525) );
  sky130_fd_sc_hd__o21ai_1 U20599 ( .A1(n16265), .A2(n16278), .B1(n15525), .Y(
        n15526) );
  sky130_fd_sc_hd__xor2_1 U20600 ( .A(n15526), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n15561) );
  sky130_fd_sc_hd__a222oi_1 U20601 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15528) );
  sky130_fd_sc_hd__o21ai_1 U20602 ( .A1(n16327), .A2(n16168), .B1(n15528), .Y(
        n15529) );
  sky130_fd_sc_hd__xor2_1 U20603 ( .A(n15529), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n15616) );
  sky130_fd_sc_hd__o22ai_1 U20604 ( .A1(n16191), .A2(n16628), .B1(n15875), 
        .B2(n16189), .Y(n15615) );
  sky130_fd_sc_hd__a222oi_1 U20605 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[15]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .Y(n15530) );
  sky130_fd_sc_hd__o21ai_1 U20606 ( .A1(n16046), .A2(n16540), .B1(n15530), .Y(
        n15531) );
  sky130_fd_sc_hd__xor2_1 U20607 ( .A(n15531), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15643) );
  sky130_fd_sc_hd__a222oi_1 U20608 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .Y(n15532) );
  sky130_fd_sc_hd__o21ai_1 U20609 ( .A1(n16227), .A2(n16319), .B1(n15532), .Y(
        n15533) );
  sky130_fd_sc_hd__xor2_1 U20610 ( .A(n15533), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n15642) );
  sky130_fd_sc_hd__fa_1 U20611 ( .A(n15536), .B(n15535), .CIN(n15534), .COUT(
        n15547), .SUM(n15641) );
  sky130_fd_sc_hd__fa_1 U20612 ( .A(n15539), .B(n15538), .CIN(n15537), .COUT(
        n15541), .SUM(n15566) );
  sky130_fd_sc_hd__fa_1 U20613 ( .A(n15542), .B(n15541), .CIN(n15540), .COUT(
        n16143), .SUM(n16142) );
  sky130_fd_sc_hd__nor2_1 U20614 ( .A(n16141), .B(n16142), .Y(n17034) );
  sky130_fd_sc_hd__fa_1 U20615 ( .A(n15545), .B(n15544), .CIN(n15543), .COUT(
        n15537), .SUM(n15697) );
  sky130_fd_sc_hd__fa_1 U20616 ( .A(n15548), .B(n15547), .CIN(n15546), .COUT(
        n15544), .SUM(n15691) );
  sky130_fd_sc_hd__fa_1 U20617 ( .A(n15551), .B(n15550), .CIN(n15549), .COUT(
        n15543), .SUM(n15690) );
  sky130_fd_sc_hd__a222oi_1 U20618 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .Y(n15552) );
  sky130_fd_sc_hd__xor2_1 U20620 ( .A(n15553), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15634) );
  sky130_fd_sc_hd__a222oi_1 U20621 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .Y(n15554) );
  sky130_fd_sc_hd__o21ai_1 U20622 ( .A1(n16227), .A2(n16311), .B1(n15554), .Y(
        n15555) );
  sky130_fd_sc_hd__xor2_1 U20623 ( .A(n15555), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n15612) );
  sky130_fd_sc_hd__a222oi_1 U20624 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .Y(n15556) );
  sky130_fd_sc_hd__o21ai_1 U20625 ( .A1(n16265), .A2(n16247), .B1(n15556), .Y(
        n15557) );
  sky130_fd_sc_hd__xor2_1 U20626 ( .A(n15557), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n15611) );
  sky130_fd_sc_hd__a222oi_1 U20627 ( .A1(n16065), .A2(n11170), .B1(n16064), 
        .B2(n11170), .C1(n16063), .C2(j202_soc_core_j22_cpu_ml_bufb[15]), .Y(
        n15558) );
  sky130_fd_sc_hd__o21ai_1 U20628 ( .A1(n16067), .A2(n16584), .B1(n15558), .Y(
        n15559) );
  sky130_fd_sc_hd__xor2_1 U20629 ( .A(n15559), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15610) );
  sky130_fd_sc_hd__fa_1 U20630 ( .A(n15562), .B(n15561), .CIN(n15560), .COUT(
        n15684), .SUM(n15632) );
  sky130_fd_sc_hd__fa_1 U20631 ( .A(n15565), .B(n15564), .CIN(n15563), .COUT(
        n15567), .SUM(n15695) );
  sky130_fd_sc_hd__fa_1 U20632 ( .A(n15568), .B(n15567), .CIN(n15566), .COUT(
        n16141), .SUM(n16140) );
  sky130_fd_sc_hd__nor2_1 U20633 ( .A(n16139), .B(n16140), .Y(n17032) );
  sky130_fd_sc_hd__nor2_1 U20634 ( .A(n17034), .B(n17032), .Y(n18972) );
  sky130_fd_sc_hd__nand2_1 U20635 ( .A(n16148), .B(n18972), .Y(n16150) );
  sky130_fd_sc_hd__a222oi_1 U20636 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .Y(n15569) );
  sky130_fd_sc_hd__xor2_1 U20638 ( .A(n15570), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15646) );
  sky130_fd_sc_hd__a222oi_1 U20639 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .Y(n15571) );
  sky130_fd_sc_hd__o21ai_1 U20640 ( .A1(n16265), .A2(n16193), .B1(n15571), .Y(
        n15572) );
  sky130_fd_sc_hd__xor2_1 U20641 ( .A(n15572), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n15590) );
  sky130_fd_sc_hd__xnor2_1 U20642 ( .A(j202_soc_core_j22_cpu_ml_bufa[3]), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .Y(n15575) );
  sky130_fd_sc_hd__xor2_1 U20643 ( .A(j202_soc_core_j22_cpu_ml_bufa[5]), .B(
        j202_soc_core_j22_cpu_ml_bufa[4]), .X(n15574) );
  sky130_fd_sc_hd__nand2b_1 U20644 ( .A_N(n15575), .B(n15574), .Y(n16058) );
  sky130_fd_sc_hd__nor2_1 U20645 ( .A(n15574), .B(n15575), .Y(n16056) );
  sky130_fd_sc_hd__xnor2_1 U20646 ( .A(j202_soc_core_j22_cpu_ml_bufa[4]), .B(
        j202_soc_core_j22_cpu_ml_bufa[3]), .Y(n15573) );
  sky130_fd_sc_hd__nor2b_1 U20647 ( .B_N(n15575), .A(n15573), .Y(n16055) );
  sky130_fd_sc_hd__and3_1 U20648 ( .A(n15575), .B(n15574), .C(n15573), .X(
        n16054) );
  sky130_fd_sc_hd__a222oi_1 U20649 ( .A1(n16056), .A2(n11170), .B1(n16055), 
        .B2(n11170), .C1(n16054), .C2(n11170), .Y(n15576) );
  sky130_fd_sc_hd__o21ai_1 U20650 ( .A1(n11169), .A2(n16058), .B1(n15576), .Y(
        n15577) );
  sky130_fd_sc_hd__xnor2_1 U20651 ( .A(j202_soc_core_j22_cpu_ml_bufa[5]), .B(
        n15577), .Y(n15631) );
  sky130_fd_sc_hd__o22ai_1 U20652 ( .A1(n16191), .A2(n19136), .B1(n15925), 
        .B2(n16189), .Y(n15630) );
  sky130_fd_sc_hd__a222oi_1 U20653 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .Y(n15578) );
  sky130_fd_sc_hd__o21ai_1 U20654 ( .A1(n16265), .A2(n16159), .B1(n15578), .Y(
        n15579) );
  sky130_fd_sc_hd__xor2_1 U20655 ( .A(n15579), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n15629) );
  sky130_fd_sc_hd__a222oi_1 U20656 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .Y(n15580) );
  sky130_fd_sc_hd__o21ai_1 U20657 ( .A1(n16052), .A2(n16354), .B1(n15580), .Y(
        n15581) );
  sky130_fd_sc_hd__xor2_1 U20658 ( .A(n15581), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15588) );
  sky130_fd_sc_hd__a222oi_1 U20659 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .Y(n15582) );
  sky130_fd_sc_hd__xor2_1 U20661 ( .A(n15583), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15593) );
  sky130_fd_sc_hd__a222oi_1 U20662 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .Y(n15584) );
  sky130_fd_sc_hd__o21ai_1 U20663 ( .A1(n16227), .A2(n16305), .B1(n15584), .Y(
        n15585) );
  sky130_fd_sc_hd__xor2_1 U20664 ( .A(n15585), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n15592) );
  sky130_fd_sc_hd__a222oi_1 U20665 ( .A1(n16065), .A2(n11170), .B1(n16064), 
        .B2(j202_soc_core_j22_cpu_ml_bufb[15]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .Y(n15586) );
  sky130_fd_sc_hd__o21ai_1 U20666 ( .A1(n16067), .A2(n16537), .B1(n15586), .Y(
        n15587) );
  sky130_fd_sc_hd__xor2_1 U20667 ( .A(n15587), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15591) );
  sky130_fd_sc_hd__fa_1 U20668 ( .A(n15590), .B(n15589), .CIN(n15588), .COUT(
        n15645), .SUM(n15676) );
  sky130_fd_sc_hd__fa_1 U20669 ( .A(n15593), .B(n15592), .CIN(n15591), .COUT(
        n15644), .SUM(n15675) );
  sky130_fd_sc_hd__a222oi_1 U20670 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .Y(n15594) );
  sky130_fd_sc_hd__o21ai_1 U20671 ( .A1(n16046), .A2(n16367), .B1(n15594), .Y(
        n15595) );
  sky130_fd_sc_hd__xor2_1 U20672 ( .A(n15595), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n16041) );
  sky130_fd_sc_hd__a222oi_1 U20673 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .Y(n15596) );
  sky130_fd_sc_hd__o21ai_1 U20674 ( .A1(n16052), .A2(n16311), .B1(n15596), .Y(
        n15597) );
  sky130_fd_sc_hd__xor2_1 U20675 ( .A(n15597), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15673) );
  sky130_fd_sc_hd__a222oi_1 U20676 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .Y(n15598) );
  sky130_fd_sc_hd__o21ai_1 U20677 ( .A1(n16227), .A2(n16247), .B1(n15598), .Y(
        n15599) );
  sky130_fd_sc_hd__xor2_1 U20678 ( .A(n15599), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n15672) );
  sky130_fd_sc_hd__a22oi_1 U20679 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15600) );
  sky130_fd_sc_hd__o21ai_1 U20680 ( .A1(n16265), .A2(n16164), .B1(n15600), .Y(
        n15601) );
  sky130_fd_sc_hd__xor2_1 U20681 ( .A(n15601), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n15670) );
  sky130_fd_sc_hd__o22ai_1 U20682 ( .A1(n16191), .A2(n15602), .B1(n20037), 
        .B2(n16189), .Y(n15669) );
  sky130_fd_sc_hd__nand2_1 U20683 ( .A(n16325), .B(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15603) );
  sky130_fd_sc_hd__o21ai_1 U20684 ( .A1(n16327), .A2(n15962), .B1(n15603), .Y(
        n15604) );
  sky130_fd_sc_hd__xor2_1 U20685 ( .A(n15604), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n15618) );
  sky130_fd_sc_hd__a222oi_1 U20686 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .Y(n15605) );
  sky130_fd_sc_hd__xor2_1 U20688 ( .A(n15606), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n15623) );
  sky130_fd_sc_hd__a222oi_1 U20689 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15607) );
  sky130_fd_sc_hd__xor2_1 U20691 ( .A(n15608), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n15655) );
  sky130_fd_sc_hd__o22ai_1 U20692 ( .A1(n16191), .A2(n17092), .B1(n15609), 
        .B2(n16189), .Y(n15654) );
  sky130_fd_sc_hd__fa_1 U20693 ( .A(n15612), .B(n15611), .CIN(n15610), .COUT(
        n15633), .SUM(n15637) );
  sky130_fd_sc_hd__a222oi_1 U20694 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .Y(n15613) );
  sky130_fd_sc_hd__o21ai_1 U20695 ( .A1(n16046), .A2(n16557), .B1(n15613), .Y(
        n15614) );
  sky130_fd_sc_hd__xor2_1 U20696 ( .A(n15614), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15640) );
  sky130_fd_sc_hd__fa_1 U20697 ( .A(n15621), .B(n15616), .CIN(n15615), .COUT(
        n15560), .SUM(n15639) );
  sky130_fd_sc_hd__o22ai_1 U20698 ( .A1(n16191), .A2(n15617), .B1(n19533), 
        .B2(n16189), .Y(n15620) );
  sky130_fd_sc_hd__fa_1 U20699 ( .A(j202_soc_core_j22_cpu_ml_bufa[20]), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .CIN(n15618), .COUT(n15619), .SUM(
        n15624) );
  sky130_fd_sc_hd__fa_1 U20700 ( .A(n15621), .B(n15620), .CIN(n15619), .COUT(
        n15638), .SUM(n15649) );
  sky130_fd_sc_hd__fa_1 U20701 ( .A(n15624), .B(n15623), .CIN(n15622), .COUT(
        n15648), .SUM(n16039) );
  sky130_fd_sc_hd__a222oi_1 U20702 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[15]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .Y(n15625) );
  sky130_fd_sc_hd__o21ai_1 U20703 ( .A1(n16067), .A2(n16540), .B1(n15625), .Y(
        n15626) );
  sky130_fd_sc_hd__xor2_1 U20704 ( .A(n15626), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15658) );
  sky130_fd_sc_hd__a222oi_1 U20705 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .Y(n15627) );
  sky130_fd_sc_hd__o21ai_1 U20706 ( .A1(n16052), .A2(n16319), .B1(n15627), .Y(
        n15628) );
  sky130_fd_sc_hd__xor2_1 U20707 ( .A(n15628), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15657) );
  sky130_fd_sc_hd__fa_1 U20708 ( .A(n15631), .B(n15630), .CIN(n15629), .COUT(
        n15589), .SUM(n15656) );
  sky130_fd_sc_hd__fa_1 U20709 ( .A(n15634), .B(n15633), .CIN(n15632), .COUT(
        n15689), .SUM(n15682) );
  sky130_fd_sc_hd__fa_1 U20710 ( .A(n15637), .B(n15636), .CIN(n15635), .COUT(
        n15681), .SUM(n15677) );
  sky130_fd_sc_hd__fa_1 U20711 ( .A(n15640), .B(n15639), .CIN(n15638), .COUT(
        n15688), .SUM(n15636) );
  sky130_fd_sc_hd__fa_1 U20712 ( .A(n15643), .B(n15642), .CIN(n15641), .COUT(
        n15683), .SUM(n15687) );
  sky130_fd_sc_hd__fa_1 U20713 ( .A(n15646), .B(n15645), .CIN(n15644), .COUT(
        n15686), .SUM(n15679) );
  sky130_fd_sc_hd__nor2_1 U20714 ( .A(n16131), .B(n16132), .Y(n19295) );
  sky130_fd_sc_hd__fa_1 U20715 ( .A(n15649), .B(n15648), .CIN(n15647), .COUT(
        n15635), .SUM(n16080) );
  sky130_fd_sc_hd__a222oi_1 U20716 ( .A1(n16056), .A2(n11170), .B1(n16055), 
        .B2(n11170), .C1(n16054), .C2(j202_soc_core_j22_cpu_ml_bufb[15]), .Y(
        n15650) );
  sky130_fd_sc_hd__o21ai_1 U20717 ( .A1(n16058), .A2(n16584), .B1(n15650), .Y(
        n15651) );
  sky130_fd_sc_hd__xor2_1 U20718 ( .A(n15651), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n16062) );
  sky130_fd_sc_hd__a222oi_1 U20719 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .Y(n15652) );
  sky130_fd_sc_hd__o21ai_1 U20720 ( .A1(n16046), .A2(n16379), .B1(n15652), .Y(
        n15653) );
  sky130_fd_sc_hd__xor2_1 U20721 ( .A(n15653), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n16061) );
  sky130_fd_sc_hd__fa_1 U20722 ( .A(n15783), .B(n15655), .CIN(n15654), .COUT(
        n15622), .SUM(n16060) );
  sky130_fd_sc_hd__fa_1 U20723 ( .A(n15658), .B(n15657), .CIN(n15656), .COUT(
        n15647), .SUM(n16076) );
  sky130_fd_sc_hd__a222oi_1 U20724 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .Y(n15659) );
  sky130_fd_sc_hd__xor2_1 U20726 ( .A(n15660), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n16083) );
  sky130_fd_sc_hd__a222oi_1 U20727 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .Y(n15661) );
  sky130_fd_sc_hd__o21ai_1 U20728 ( .A1(n16227), .A2(n16193), .B1(n15661), .Y(
        n15662) );
  sky130_fd_sc_hd__xor2_1 U20729 ( .A(n15662), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n16086) );
  sky130_fd_sc_hd__nand2_1 U20730 ( .A(n16263), .B(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15663) );
  sky130_fd_sc_hd__o21ai_1 U20731 ( .A1(n15962), .A2(n16265), .B1(n15663), .Y(
        n15664) );
  sky130_fd_sc_hd__xor2_1 U20732 ( .A(n15664), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n15782) );
  sky130_fd_sc_hd__xor2_1 U20733 ( .A(j202_soc_core_j22_cpu_ml_bufa[1]), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15665) );
  sky130_fd_sc_hd__nand2b_1 U20734 ( .A_N(n22247), .B(n15665), .Y(n15959) );
  sky130_fd_sc_hd__nor2_1 U20735 ( .A(n22247), .B(n15665), .Y(n15957) );
  sky130_fd_sc_hd__nor2b_1 U20736 ( .B_N(n22247), .A(n15666), .Y(n15956) );
  sky130_fd_sc_hd__and3_1 U20737 ( .A(n15666), .B(n15665), .C(n22247), .X(
        n15955) );
  sky130_fd_sc_hd__a222oi_1 U20738 ( .A1(n15957), .A2(n11170), .B1(n15956), 
        .B2(n11170), .C1(n15955), .C2(n11170), .Y(n15667) );
  sky130_fd_sc_hd__xnor2_1 U20740 ( .A(j202_soc_core_j22_cpu_ml_bufa[2]), .B(
        n15668), .Y(n15781) );
  sky130_fd_sc_hd__fa_1 U20741 ( .A(n15783), .B(n15670), .CIN(n15669), .COUT(
        n15671), .SUM(n16084) );
  sky130_fd_sc_hd__fa_1 U20742 ( .A(n15673), .B(n15672), .CIN(n15671), .COUT(
        n16040), .SUM(n16081) );
  sky130_fd_sc_hd__fa_1 U20743 ( .A(n15676), .B(n15675), .CIN(n15674), .COUT(
        n15678), .SUM(n16078) );
  sky130_fd_sc_hd__fa_1 U20744 ( .A(n15679), .B(n15678), .CIN(n15677), .COUT(
        n16131), .SUM(n16130) );
  sky130_fd_sc_hd__nor2_1 U20745 ( .A(n16129), .B(n16130), .Y(n19300) );
  sky130_fd_sc_hd__nor2_1 U20746 ( .A(n19295), .B(n19300), .Y(n16787) );
  sky130_fd_sc_hd__fa_1 U20747 ( .A(n15682), .B(n15681), .CIN(n15680), .COUT(
        n16133), .SUM(n16132) );
  sky130_fd_sc_hd__fa_1 U20748 ( .A(n15685), .B(n15684), .CIN(n15683), .COUT(
        n15563), .SUM(n15694) );
  sky130_fd_sc_hd__fa_1 U20749 ( .A(n15688), .B(n15687), .CIN(n15686), .COUT(
        n15693), .SUM(n15680) );
  sky130_fd_sc_hd__fa_1 U20750 ( .A(n15691), .B(n15690), .CIN(n15689), .COUT(
        n15696), .SUM(n15692) );
  sky130_fd_sc_hd__nor2_1 U20751 ( .A(n16133), .B(n16134), .Y(n16791) );
  sky130_fd_sc_hd__fa_1 U20752 ( .A(n15694), .B(n15693), .CIN(n15692), .COUT(
        n16135), .SUM(n16134) );
  sky130_fd_sc_hd__fa_1 U20753 ( .A(n15697), .B(n15696), .CIN(n15695), .COUT(
        n16139), .SUM(n16136) );
  sky130_fd_sc_hd__nor2_1 U20754 ( .A(n16135), .B(n16136), .Y(n16793) );
  sky130_fd_sc_hd__nor2_1 U20755 ( .A(n16791), .B(n16793), .Y(n16138) );
  sky130_fd_sc_hd__nand2_1 U20756 ( .A(n16787), .B(n16138), .Y(n17031) );
  sky130_fd_sc_hd__nor2_1 U20757 ( .A(n16150), .B(n17031), .Y(n16152) );
  sky130_fd_sc_hd__a222oi_1 U20758 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .Y(n15698) );
  sky130_fd_sc_hd__o21ai_1 U20759 ( .A1(n16046), .A2(n16305), .B1(n15698), .Y(
        n15699) );
  sky130_fd_sc_hd__xor2_1 U20760 ( .A(n15699), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15762) );
  sky130_fd_sc_hd__a222oi_1 U20761 ( .A1(n15957), .A2(n11170), .B1(n15956), 
        .B2(j202_soc_core_j22_cpu_ml_bufb[15]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .Y(n15700) );
  sky130_fd_sc_hd__o21ai_1 U20762 ( .A1(n15959), .A2(n16537), .B1(n15700), .Y(
        n15701) );
  sky130_fd_sc_hd__xor2_1 U20763 ( .A(n15701), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15761) );
  sky130_fd_sc_hd__a22oi_1 U20764 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15702) );
  sky130_fd_sc_hd__o21ai_1 U20765 ( .A1(n16227), .A2(n16164), .B1(n15702), .Y(
        n15703) );
  sky130_fd_sc_hd__xor2_1 U20766 ( .A(n15703), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n15743) );
  sky130_fd_sc_hd__o22ai_1 U20767 ( .A1(n16191), .A2(n15704), .B1(n15942), 
        .B2(n16189), .Y(n15742) );
  sky130_fd_sc_hd__a222oi_1 U20768 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .Y(n15705) );
  sky130_fd_sc_hd__xor2_1 U20770 ( .A(n15706), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15741) );
  sky130_fd_sc_hd__a222oi_1 U20771 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15707) );
  sky130_fd_sc_hd__xor2_1 U20773 ( .A(n15708), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15801) );
  sky130_fd_sc_hd__o22ai_1 U20774 ( .A1(n20036), .A2(n15709), .B1(n18992), 
        .B2(n16189), .Y(n15800) );
  sky130_fd_sc_hd__a222oi_1 U20775 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .Y(n15710) );
  sky130_fd_sc_hd__o21ai_1 U20776 ( .A1(n16067), .A2(n16311), .B1(n15710), .Y(
        n15711) );
  sky130_fd_sc_hd__xor2_1 U20777 ( .A(n15711), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15799) );
  sky130_fd_sc_hd__a222oi_1 U20778 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .Y(n15712) );
  sky130_fd_sc_hd__o21ai_1 U20779 ( .A1(n16046), .A2(n16247), .B1(n15712), .Y(
        n15713) );
  sky130_fd_sc_hd__xor2_1 U20780 ( .A(n15713), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15817) );
  sky130_fd_sc_hd__a222oi_1 U20781 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .Y(n15714) );
  sky130_fd_sc_hd__o21ai_1 U20782 ( .A1(n15959), .A2(n16557), .B1(n15714), .Y(
        n15715) );
  sky130_fd_sc_hd__xor2_1 U20783 ( .A(n15715), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15816) );
  sky130_fd_sc_hd__a222oi_1 U20784 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .Y(n15716) );
  sky130_fd_sc_hd__o21ai_1 U20785 ( .A1(n16058), .A2(n16379), .B1(n15716), .Y(
        n15717) );
  sky130_fd_sc_hd__xor2_1 U20786 ( .A(n15717), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15815) );
  sky130_fd_sc_hd__a222oi_1 U20787 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .Y(n15718) );
  sky130_fd_sc_hd__o21ai_1 U20788 ( .A1(n16052), .A2(n16159), .B1(n15718), .Y(
        n15719) );
  sky130_fd_sc_hd__xor2_1 U20789 ( .A(n15719), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15726) );
  sky130_fd_sc_hd__a222oi_1 U20790 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .Y(n15720) );
  sky130_fd_sc_hd__o21ai_1 U20791 ( .A1(n16046), .A2(n16278), .B1(n15720), .Y(
        n15721) );
  sky130_fd_sc_hd__xor2_1 U20792 ( .A(n15721), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15725) );
  sky130_fd_sc_hd__nand2_1 U20793 ( .A(n16225), .B(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15722) );
  sky130_fd_sc_hd__xor2_1 U20795 ( .A(n15723), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n15734) );
  sky130_fd_sc_hd__o22ai_1 U20796 ( .A1(n20036), .A2(n16190), .B1(n16608), 
        .B2(n16189), .Y(n15733) );
  sky130_fd_sc_hd__fa_1 U20797 ( .A(n15726), .B(n15725), .CIN(n15724), .COUT(
        n15750), .SUM(n15809) );
  sky130_fd_sc_hd__a222oi_1 U20798 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[15]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .Y(n15727) );
  sky130_fd_sc_hd__o21ai_1 U20799 ( .A1(n15959), .A2(n16540), .B1(n15727), .Y(
        n15728) );
  sky130_fd_sc_hd__xor2_1 U20800 ( .A(n15728), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15793) );
  sky130_fd_sc_hd__a222oi_1 U20801 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .Y(n15729) );
  sky130_fd_sc_hd__o21ai_1 U20802 ( .A1(n16067), .A2(n16319), .B1(n15729), .Y(
        n15730) );
  sky130_fd_sc_hd__xor2_1 U20803 ( .A(n15730), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15792) );
  sky130_fd_sc_hd__a222oi_1 U20804 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .Y(n15731) );
  sky130_fd_sc_hd__o21ai_1 U20805 ( .A1(n16058), .A2(n16367), .B1(n15731), .Y(
        n15732) );
  sky130_fd_sc_hd__xor2_1 U20806 ( .A(n15732), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15791) );
  sky130_fd_sc_hd__fa_1 U20807 ( .A(j202_soc_core_j22_cpu_ml_bufa[17]), .B(
        n15734), .CIN(n15733), .COUT(n15753), .SUM(n15724) );
  sky130_fd_sc_hd__a222oi_1 U20808 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .Y(n15735) );
  sky130_fd_sc_hd__xor2_1 U20810 ( .A(n15736), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15752) );
  sky130_fd_sc_hd__a222oi_1 U20811 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .Y(n15737) );
  sky130_fd_sc_hd__o21ai_1 U20812 ( .A1(n16058), .A2(n16402), .B1(n15737), .Y(
        n15738) );
  sky130_fd_sc_hd__xor2_1 U20813 ( .A(n15738), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15751) );
  sky130_fd_sc_hd__a222oi_1 U20814 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .Y(n15739) );
  sky130_fd_sc_hd__xor2_1 U20816 ( .A(n15740), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15790) );
  sky130_fd_sc_hd__fa_1 U20817 ( .A(n15743), .B(n15742), .CIN(n15741), .COUT(
        n15789), .SUM(n15760) );
  sky130_fd_sc_hd__a222oi_1 U20818 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15744) );
  sky130_fd_sc_hd__o21ai_1 U20819 ( .A1(n16227), .A2(n16168), .B1(n15744), .Y(
        n15745) );
  sky130_fd_sc_hd__xor2_1 U20820 ( .A(n15745), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n15770) );
  sky130_fd_sc_hd__o22ai_1 U20821 ( .A1(n16191), .A2(n19860), .B1(n15941), 
        .B2(n16189), .Y(n15769) );
  sky130_fd_sc_hd__a222oi_1 U20822 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .Y(n15746) );
  sky130_fd_sc_hd__o21ai_1 U20823 ( .A1(n16046), .A2(n16311), .B1(n15746), .Y(
        n15747) );
  sky130_fd_sc_hd__xor2_1 U20824 ( .A(n15747), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15768) );
  sky130_fd_sc_hd__fa_1 U20825 ( .A(n15750), .B(n15749), .CIN(n15748), .COUT(
        n15764), .SUM(n15812) );
  sky130_fd_sc_hd__fa_1 U20826 ( .A(n15753), .B(n15752), .CIN(n15751), .COUT(
        n15777), .SUM(n15748) );
  sky130_fd_sc_hd__a222oi_1 U20827 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .Y(n15754) );
  sky130_fd_sc_hd__o21ai_1 U20828 ( .A1(n16052), .A2(n16247), .B1(n15754), .Y(
        n15755) );
  sky130_fd_sc_hd__xor2_1 U20829 ( .A(n15755), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15780) );
  sky130_fd_sc_hd__a222oi_1 U20830 ( .A1(n15957), .A2(n11170), .B1(n15956), 
        .B2(n11170), .C1(n15955), .C2(j202_soc_core_j22_cpu_ml_bufb[15]), .Y(
        n15756) );
  sky130_fd_sc_hd__o21ai_1 U20831 ( .A1(n15959), .A2(n16584), .B1(n15756), .Y(
        n15757) );
  sky130_fd_sc_hd__xor2_1 U20832 ( .A(n15757), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15779) );
  sky130_fd_sc_hd__a222oi_1 U20833 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .Y(n15758) );
  sky130_fd_sc_hd__o21ai_1 U20834 ( .A1(n16058), .A2(n16557), .B1(n15758), .Y(
        n15759) );
  sky130_fd_sc_hd__xor2_1 U20835 ( .A(n15759), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15778) );
  sky130_fd_sc_hd__fa_1 U20836 ( .A(n15762), .B(n15761), .CIN(n15760), .COUT(
        n15775), .SUM(n15814) );
  sky130_fd_sc_hd__nor2_1 U20837 ( .A(n16033), .B(n16034), .Y(n19855) );
  sky130_fd_sc_hd__fa_1 U20838 ( .A(n15765), .B(n15764), .CIN(n15763), .COUT(
        n16035), .SUM(n16034) );
  sky130_fd_sc_hd__a222oi_1 U20839 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .Y(n15766) );
  sky130_fd_sc_hd__xor2_1 U20841 ( .A(n15767), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n16092) );
  sky130_fd_sc_hd__fa_1 U20842 ( .A(n15770), .B(n15769), .CIN(n15768), .COUT(
        n16091), .SUM(n15788) );
  sky130_fd_sc_hd__o22ai_1 U20843 ( .A1(n16191), .A2(n16835), .B1(n15951), 
        .B2(n16189), .Y(n16071) );
  sky130_fd_sc_hd__a222oi_1 U20844 ( .A1(n16225), .A2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .B1(n16224), .B2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .Y(n15771) );
  sky130_fd_sc_hd__o21ai_1 U20845 ( .A1(n16227), .A2(n16159), .B1(n15771), .Y(
        n15772) );
  sky130_fd_sc_hd__xor2_1 U20846 ( .A(n15772), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n16070) );
  sky130_fd_sc_hd__a222oi_1 U20847 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .Y(n15773) );
  sky130_fd_sc_hd__o21ai_1 U20848 ( .A1(n16052), .A2(n16278), .B1(n15773), .Y(
        n15774) );
  sky130_fd_sc_hd__xor2_1 U20849 ( .A(n15774), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n16069) );
  sky130_fd_sc_hd__fa_1 U20850 ( .A(n15777), .B(n15776), .CIN(n15775), .COUT(
        n16100), .SUM(n15763) );
  sky130_fd_sc_hd__fa_1 U20851 ( .A(n15780), .B(n15779), .CIN(n15778), .COUT(
        n16107), .SUM(n15776) );
  sky130_fd_sc_hd__fa_1 U20852 ( .A(n15783), .B(n15782), .CIN(n15781), .COUT(
        n16085), .SUM(n16074) );
  sky130_fd_sc_hd__a222oi_1 U20853 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[15]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .Y(n15784) );
  sky130_fd_sc_hd__o21ai_1 U20854 ( .A1(n16058), .A2(n16540), .B1(n15784), .Y(
        n15785) );
  sky130_fd_sc_hd__xor2_1 U20855 ( .A(n15785), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n16073) );
  sky130_fd_sc_hd__a222oi_1 U20856 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .Y(n15786) );
  sky130_fd_sc_hd__o21ai_1 U20857 ( .A1(n16046), .A2(n16319), .B1(n15786), .Y(
        n15787) );
  sky130_fd_sc_hd__xor2_1 U20858 ( .A(n15787), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n16072) );
  sky130_fd_sc_hd__fa_1 U20859 ( .A(n15790), .B(n15789), .CIN(n15788), .COUT(
        n16105), .SUM(n15765) );
  sky130_fd_sc_hd__nor2_1 U20860 ( .A(n16035), .B(n16036), .Y(n16829) );
  sky130_fd_sc_hd__nor2_1 U20861 ( .A(n19855), .B(n16829), .Y(n16038) );
  sky130_fd_sc_hd__fa_1 U20862 ( .A(n15793), .B(n15792), .CIN(n15791), .COUT(
        n15749), .SUM(n15834) );
  sky130_fd_sc_hd__a22oi_1 U20863 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15794) );
  sky130_fd_sc_hd__o21ai_1 U20864 ( .A1(n16052), .A2(n16164), .B1(n15794), .Y(
        n15795) );
  sky130_fd_sc_hd__xor2_1 U20865 ( .A(n15795), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15822) );
  sky130_fd_sc_hd__o22ai_1 U20866 ( .A1(n20036), .A2(n15796), .B1(n19112), 
        .B2(n16189), .Y(n15821) );
  sky130_fd_sc_hd__a222oi_1 U20867 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .Y(n15797) );
  sky130_fd_sc_hd__xor2_1 U20869 ( .A(n15798), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15820) );
  sky130_fd_sc_hd__fa_1 U20870 ( .A(n15801), .B(n15800), .CIN(n15799), .COUT(
        n15811), .SUM(n15830) );
  sky130_fd_sc_hd__nand2_1 U20871 ( .A(n16050), .B(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15802) );
  sky130_fd_sc_hd__o21ai_1 U20872 ( .A1(n15962), .A2(n16052), .B1(n15802), .Y(
        n15803) );
  sky130_fd_sc_hd__xor2_1 U20873 ( .A(n15803), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n15828) );
  sky130_fd_sc_hd__o22ai_1 U20874 ( .A1(n20036), .A2(n15804), .B1(n17048), 
        .B2(n16189), .Y(n15827) );
  sky130_fd_sc_hd__a222oi_1 U20875 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .Y(n15805) );
  sky130_fd_sc_hd__o21ai_1 U20876 ( .A1(n15959), .A2(n16402), .B1(n15805), .Y(
        n15806) );
  sky130_fd_sc_hd__xor2_1 U20877 ( .A(n15806), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15857) );
  sky130_fd_sc_hd__a222oi_1 U20878 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .Y(n15807) );
  sky130_fd_sc_hd__xor2_1 U20880 ( .A(n15808), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15856) );
  sky130_fd_sc_hd__fa_1 U20881 ( .A(n15811), .B(n15810), .CIN(n15809), .COUT(
        n15813), .SUM(n15832) );
  sky130_fd_sc_hd__fa_1 U20882 ( .A(n15814), .B(n15813), .CIN(n15812), .COUT(
        n16033), .SUM(n16029) );
  sky130_fd_sc_hd__fa_1 U20883 ( .A(n15817), .B(n15816), .CIN(n15815), .COUT(
        n15810), .SUM(n15870) );
  sky130_fd_sc_hd__a222oi_1 U20884 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .Y(n15818) );
  sky130_fd_sc_hd__o21ai_1 U20885 ( .A1(n16067), .A2(n16305), .B1(n15818), .Y(
        n15819) );
  sky130_fd_sc_hd__xor2_1 U20886 ( .A(n15819), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15864) );
  sky130_fd_sc_hd__fa_1 U20887 ( .A(n15822), .B(n15821), .CIN(n15820), .COUT(
        n15831), .SUM(n15863) );
  sky130_fd_sc_hd__a222oi_1 U20888 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .Y(n15823) );
  sky130_fd_sc_hd__o21ai_1 U20889 ( .A1(n16046), .A2(n16159), .B1(n15823), .Y(
        n15824) );
  sky130_fd_sc_hd__xor2_1 U20890 ( .A(n15824), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15846) );
  sky130_fd_sc_hd__a222oi_1 U20891 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .Y(n15825) );
  sky130_fd_sc_hd__xor2_1 U20893 ( .A(n15826), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15845) );
  sky130_fd_sc_hd__fa_1 U20894 ( .A(j202_soc_core_j22_cpu_ml_bufa[14]), .B(
        n15828), .CIN(n15827), .COUT(n15858), .SUM(n15844) );
  sky130_fd_sc_hd__fa_1 U20895 ( .A(n15831), .B(n15830), .CIN(n15829), .COUT(
        n15833), .SUM(n15868) );
  sky130_fd_sc_hd__fa_1 U20896 ( .A(n15834), .B(n15833), .CIN(n15832), .COUT(
        n16028), .SUM(n16027) );
  sky130_fd_sc_hd__nand2_1 U20897 ( .A(n19226), .B(n19223), .Y(n16032) );
  sky130_fd_sc_hd__a222oi_1 U20898 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .Y(n15835) );
  sky130_fd_sc_hd__o21ai_1 U20899 ( .A1(n16067), .A2(n16247), .B1(n15835), .Y(
        n15836) );
  sky130_fd_sc_hd__xor2_1 U20900 ( .A(n15836), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n16003) );
  sky130_fd_sc_hd__a222oi_1 U20901 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .Y(n15837) );
  sky130_fd_sc_hd__o21ai_1 U20902 ( .A1(n15959), .A2(n16379), .B1(n15837), .Y(
        n15838) );
  sky130_fd_sc_hd__xor2_1 U20903 ( .A(n15838), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n16002) );
  sky130_fd_sc_hd__a22oi_1 U20904 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15839) );
  sky130_fd_sc_hd__o21ai_1 U20905 ( .A1(n16046), .A2(n16164), .B1(n15839), .Y(
        n15840) );
  sky130_fd_sc_hd__xor2_1 U20906 ( .A(n15840), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15900) );
  sky130_fd_sc_hd__o22ai_1 U20907 ( .A1(n20036), .A2(n15841), .B1(n16808), 
        .B2(n16189), .Y(n15899) );
  sky130_fd_sc_hd__a222oi_1 U20908 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .Y(n15842) );
  sky130_fd_sc_hd__o21ai_1 U20909 ( .A1(n16067), .A2(n16193), .B1(n15842), .Y(
        n15843) );
  sky130_fd_sc_hd__xor2_1 U20910 ( .A(n15843), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15898) );
  sky130_fd_sc_hd__fa_1 U20911 ( .A(n15846), .B(n15845), .CIN(n15844), .COUT(
        n15862), .SUM(n16005) );
  sky130_fd_sc_hd__a222oi_1 U20912 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .Y(n15847) );
  sky130_fd_sc_hd__o21ai_1 U20913 ( .A1(n15959), .A2(n16367), .B1(n15847), .Y(
        n15848) );
  sky130_fd_sc_hd__xor2_1 U20914 ( .A(n15848), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15861) );
  sky130_fd_sc_hd__a222oi_1 U20915 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .Y(n15849) );
  sky130_fd_sc_hd__o21ai_1 U20916 ( .A1(n16058), .A2(n16319), .B1(n15849), .Y(
        n15850) );
  sky130_fd_sc_hd__xor2_1 U20917 ( .A(n15850), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15860) );
  sky130_fd_sc_hd__a222oi_1 U20918 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15851) );
  sky130_fd_sc_hd__xor2_1 U20920 ( .A(n15852), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15997) );
  sky130_fd_sc_hd__o22ai_1 U20921 ( .A1(n20036), .A2(n15853), .B1(n18869), 
        .B2(n16189), .Y(n15996) );
  sky130_fd_sc_hd__a222oi_1 U20922 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .Y(n15854) );
  sky130_fd_sc_hd__xor2_1 U20924 ( .A(n15855), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15995) );
  sky130_fd_sc_hd__fa_1 U20925 ( .A(n15858), .B(n15857), .CIN(n15856), .COUT(
        n15829), .SUM(n15867) );
  sky130_fd_sc_hd__fa_1 U20926 ( .A(n15861), .B(n15860), .CIN(n15859), .COUT(
        n15866), .SUM(n16004) );
  sky130_fd_sc_hd__fa_1 U20927 ( .A(n15864), .B(n15863), .CIN(n15862), .COUT(
        n15869), .SUM(n15865) );
  sky130_fd_sc_hd__nor2_1 U20928 ( .A(n16020), .B(n16021), .Y(n19107) );
  sky130_fd_sc_hd__fa_1 U20929 ( .A(n15867), .B(n15866), .CIN(n15865), .COUT(
        n16022), .SUM(n16021) );
  sky130_fd_sc_hd__fa_1 U20930 ( .A(n15870), .B(n15869), .CIN(n15868), .COUT(
        n16026), .SUM(n16023) );
  sky130_fd_sc_hd__nor2_1 U20931 ( .A(n16022), .B(n16023), .Y(n18986) );
  sky130_fd_sc_hd__nor2_1 U20932 ( .A(n19107), .B(n18986), .Y(n16025) );
  sky130_fd_sc_hd__a222oi_1 U20933 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .Y(n15871) );
  sky130_fd_sc_hd__o21ai_1 U20934 ( .A1(n16058), .A2(n16247), .B1(n15871), .Y(
        n15872) );
  sky130_fd_sc_hd__xor2_1 U20935 ( .A(n15872), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15986) );
  sky130_fd_sc_hd__a22oi_1 U20936 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15873) );
  sky130_fd_sc_hd__o21ai_1 U20937 ( .A1(n16067), .A2(n16164), .B1(n15873), .Y(
        n15874) );
  sky130_fd_sc_hd__xor2_1 U20938 ( .A(n15874), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15922) );
  sky130_fd_sc_hd__o22ai_1 U20939 ( .A1(n20036), .A2(n15875), .B1(n16636), 
        .B2(n16189), .Y(n15921) );
  sky130_fd_sc_hd__a222oi_1 U20940 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .Y(n15876) );
  sky130_fd_sc_hd__xor2_1 U20942 ( .A(n15877), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15920) );
  sky130_fd_sc_hd__a222oi_1 U20943 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15878) );
  sky130_fd_sc_hd__o21ai_1 U20944 ( .A1(n16067), .A2(n16168), .B1(n15878), .Y(
        n15879) );
  sky130_fd_sc_hd__xor2_1 U20945 ( .A(n15879), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15887) );
  sky130_fd_sc_hd__o22ai_1 U20946 ( .A1(n20036), .A2(n15880), .B1(n19312), 
        .B2(n16189), .Y(n15886) );
  sky130_fd_sc_hd__a222oi_1 U20947 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .Y(n15881) );
  sky130_fd_sc_hd__o21ai_1 U20948 ( .A1(n15959), .A2(n16311), .B1(n15881), .Y(
        n15882) );
  sky130_fd_sc_hd__xor2_1 U20949 ( .A(n15882), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15885) );
  sky130_fd_sc_hd__a222oi_1 U20950 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .Y(n15883) );
  sky130_fd_sc_hd__xor2_1 U20952 ( .A(n15884), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15897) );
  sky130_fd_sc_hd__fa_1 U20953 ( .A(n15887), .B(n15886), .CIN(n15885), .COUT(
        n15896), .SUM(n15984) );
  sky130_fd_sc_hd__a222oi_1 U20954 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .Y(n15888) );
  sky130_fd_sc_hd__o21ai_1 U20955 ( .A1(n16067), .A2(n16159), .B1(n15888), .Y(
        n15889) );
  sky130_fd_sc_hd__xor2_1 U20956 ( .A(n15889), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15903) );
  sky130_fd_sc_hd__a222oi_1 U20957 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .Y(n15890) );
  sky130_fd_sc_hd__xor2_1 U20959 ( .A(n15891), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15902) );
  sky130_fd_sc_hd__nand2_1 U20960 ( .A(n16044), .B(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15892) );
  sky130_fd_sc_hd__xor2_1 U20962 ( .A(n15893), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n15905) );
  sky130_fd_sc_hd__o22ai_1 U20963 ( .A1(n20036), .A2(n15894), .B1(n20013), 
        .B2(n16189), .Y(n15904) );
  sky130_fd_sc_hd__nor2_1 U20964 ( .A(n15989), .B(n15990), .Y(n19954) );
  sky130_fd_sc_hd__fa_1 U20965 ( .A(n15897), .B(n15896), .CIN(n15895), .COUT(
        n15991), .SUM(n15990) );
  sky130_fd_sc_hd__fa_1 U20966 ( .A(n15900), .B(n15899), .CIN(n15898), .COUT(
        n16001), .SUM(n16009) );
  sky130_fd_sc_hd__fa_1 U20967 ( .A(n15903), .B(n15902), .CIN(n15901), .COUT(
        n16008), .SUM(n15895) );
  sky130_fd_sc_hd__fa_1 U20968 ( .A(j202_soc_core_j22_cpu_ml_bufa[11]), .B(
        n15905), .CIN(n15904), .COUT(n16000), .SUM(n15901) );
  sky130_fd_sc_hd__a222oi_1 U20969 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .Y(n15906) );
  sky130_fd_sc_hd__o21ai_1 U20970 ( .A1(n15959), .A2(n16354), .B1(n15906), .Y(
        n15907) );
  sky130_fd_sc_hd__xor2_1 U20971 ( .A(n15907), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15999) );
  sky130_fd_sc_hd__a222oi_1 U20972 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .Y(n15908) );
  sky130_fd_sc_hd__xor2_1 U20974 ( .A(n15909), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15998) );
  sky130_fd_sc_hd__nor2_1 U20975 ( .A(n15991), .B(n15992), .Y(n16802) );
  sky130_fd_sc_hd__nor2_1 U20976 ( .A(n19954), .B(n16802), .Y(n15994) );
  sky130_fd_sc_hd__a222oi_1 U20977 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .Y(n15910) );
  sky130_fd_sc_hd__o21ai_1 U20978 ( .A1(n16058), .A2(n16159), .B1(n15910), .Y(
        n15911) );
  sky130_fd_sc_hd__xor2_1 U20979 ( .A(n15911), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15930) );
  sky130_fd_sc_hd__a222oi_1 U20980 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .Y(n15912) );
  sky130_fd_sc_hd__o21ai_1 U20981 ( .A1(n15959), .A2(n16278), .B1(n15912), .Y(
        n15913) );
  sky130_fd_sc_hd__xor2_1 U20982 ( .A(n15913), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15929) );
  sky130_fd_sc_hd__nand2_1 U20983 ( .A(n16065), .B(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15914) );
  sky130_fd_sc_hd__xor2_1 U20985 ( .A(n15915), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n15917) );
  sky130_fd_sc_hd__o22ai_1 U20986 ( .A1(n20036), .A2(n19533), .B1(n19017), 
        .B2(n16189), .Y(n15916) );
  sky130_fd_sc_hd__fa_1 U20987 ( .A(j202_soc_core_j22_cpu_ml_bufa[8]), .B(
        n15917), .CIN(n15916), .COUT(n15983), .SUM(n15928) );
  sky130_fd_sc_hd__a222oi_1 U20988 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .Y(n15918) );
  sky130_fd_sc_hd__o21ai_1 U20989 ( .A1(n15959), .A2(n16305), .B1(n15918), .Y(
        n15919) );
  sky130_fd_sc_hd__xor2_1 U20990 ( .A(n15919), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15982) );
  sky130_fd_sc_hd__fa_1 U20991 ( .A(n15922), .B(n15921), .CIN(n15920), .COUT(
        n15985), .SUM(n15981) );
  sky130_fd_sc_hd__a222oi_1 U20992 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15923) );
  sky130_fd_sc_hd__o21ai_1 U20993 ( .A1(n16058), .A2(n16168), .B1(n15923), .Y(
        n15924) );
  sky130_fd_sc_hd__xor2_1 U20994 ( .A(n15924), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15938) );
  sky130_fd_sc_hd__o22ai_1 U20995 ( .A1(n20036), .A2(n15925), .B1(n19144), 
        .B2(n16189), .Y(n15937) );
  sky130_fd_sc_hd__a222oi_1 U20996 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .Y(n15926) );
  sky130_fd_sc_hd__o21ai_1 U20997 ( .A1(n15959), .A2(n16247), .B1(n15926), .Y(
        n15927) );
  sky130_fd_sc_hd__xor2_1 U20998 ( .A(n15927), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15936) );
  sky130_fd_sc_hd__fa_1 U20999 ( .A(n15930), .B(n15929), .CIN(n15928), .COUT(
        n15978), .SUM(n15977) );
  sky130_fd_sc_hd__nor2_1 U21000 ( .A(n15976), .B(n15977), .Y(n19012) );
  sky130_fd_sc_hd__a22oi_1 U21001 ( .A1(n16056), .A2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .B1(n16055), .B2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15931) );
  sky130_fd_sc_hd__xor2_1 U21003 ( .A(n15932), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15970) );
  sky130_fd_sc_hd__a22o_1 U21004 ( .A1(j202_soc_core_j22_cpu_ml_macl[20]), 
        .A2(n19959), .B1(n15933), .B2(j202_soc_core_j22_cpu_ml_macl[4]), .X(
        n15969) );
  sky130_fd_sc_hd__a222oi_1 U21005 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .Y(n15934) );
  sky130_fd_sc_hd__o21ai_1 U21006 ( .A1(n15959), .A2(n16193), .B1(n15934), .Y(
        n15935) );
  sky130_fd_sc_hd__xor2_1 U21007 ( .A(n15935), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15968) );
  sky130_fd_sc_hd__fa_1 U21008 ( .A(n15938), .B(n15937), .CIN(n15936), .COUT(
        n15976), .SUM(n15974) );
  sky130_fd_sc_hd__a22oi_1 U21009 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15939) );
  sky130_fd_sc_hd__o21ai_1 U21010 ( .A1(n15959), .A2(n16164), .B1(n15939), .Y(
        n15940) );
  sky130_fd_sc_hd__xor2_1 U21011 ( .A(n15940), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15947) );
  sky130_fd_sc_hd__o22ai_1 U21012 ( .A1(n20036), .A2(n15941), .B1(n19869), 
        .B2(n16189), .Y(n15948) );
  sky130_fd_sc_hd__nor2_1 U21013 ( .A(n15947), .B(n15948), .Y(n19864) );
  sky130_fd_sc_hd__o22ai_1 U21014 ( .A1(n20036), .A2(n15942), .B1(n19235), 
        .B2(n16189), .Y(n19234) );
  sky130_fd_sc_hd__nand2_1 U21015 ( .A(n15957), .B(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15943) );
  sky130_fd_sc_hd__xor2_1 U21017 ( .A(n19232), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15944) );
  sky130_fd_sc_hd__a21oi_1 U21018 ( .A1(n19234), .A2(n15946), .B1(n15945), .Y(
        n19867) );
  sky130_fd_sc_hd__nand2_1 U21019 ( .A(n15948), .B(n15947), .Y(n19865) );
  sky130_fd_sc_hd__a222oi_1 U21021 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15949) );
  sky130_fd_sc_hd__o21ai_1 U21022 ( .A1(n15959), .A2(n16168), .B1(n15949), .Y(
        n15950) );
  sky130_fd_sc_hd__xor2_1 U21023 ( .A(n15950), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15952) );
  sky130_fd_sc_hd__o22ai_1 U21024 ( .A1(n20036), .A2(n15951), .B1(n16843), 
        .B2(n16189), .Y(n15953) );
  sky130_fd_sc_hd__nand2_1 U21025 ( .A(n15953), .B(n15952), .Y(n16839) );
  sky130_fd_sc_hd__a21oi_1 U21026 ( .A1(n16841), .A2(n16840), .B1(n15954), .Y(
        n18886) );
  sky130_fd_sc_hd__a222oi_1 U21027 ( .A1(n15957), .A2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .B1(n15956), .B2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .C1(n15955), .C2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .Y(n15958) );
  sky130_fd_sc_hd__xor2_1 U21029 ( .A(n15960), .B(
        j202_soc_core_j22_cpu_ml_bufa[2]), .X(n15964) );
  sky130_fd_sc_hd__nand2_1 U21030 ( .A(n16056), .B(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n15961) );
  sky130_fd_sc_hd__xor2_1 U21032 ( .A(n15963), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n15967) );
  sky130_fd_sc_hd__o22ai_1 U21033 ( .A1(n20036), .A2(n20037), .B1(n18888), 
        .B2(n16189), .Y(n15966) );
  sky130_fd_sc_hd__nor2_1 U21034 ( .A(n15964), .B(n15965), .Y(n18883) );
  sky130_fd_sc_hd__nand2_1 U21035 ( .A(n15965), .B(n15964), .Y(n18884) );
  sky130_fd_sc_hd__o21a_1 U21036 ( .A1(n18886), .A2(n18883), .B1(n18884), .X(
        n17097) );
  sky130_fd_sc_hd__fa_1 U21037 ( .A(j202_soc_core_j22_cpu_ml_bufa[5]), .B(
        n15967), .CIN(n15966), .COUT(n15971), .SUM(n15965) );
  sky130_fd_sc_hd__fa_1 U21038 ( .A(n15970), .B(n15969), .CIN(n15968), .COUT(
        n15973), .SUM(n15972) );
  sky130_fd_sc_hd__nor2_1 U21039 ( .A(n15971), .B(n15972), .Y(n17094) );
  sky130_fd_sc_hd__nand2_1 U21040 ( .A(n15972), .B(n15971), .Y(n17095) );
  sky130_fd_sc_hd__nand2_1 U21042 ( .A(n15974), .B(n15973), .Y(n19140) );
  sky130_fd_sc_hd__a21oi_1 U21043 ( .A1(n19141), .A2(n19143), .B1(n15975), .Y(
        n19015) );
  sky130_fd_sc_hd__nand2_1 U21044 ( .A(n15977), .B(n15976), .Y(n19013) );
  sky130_fd_sc_hd__nand2_1 U21046 ( .A(n15979), .B(n15978), .Y(n16632) );
  sky130_fd_sc_hd__a21oi_1 U21047 ( .A1(n16633), .A2(n16635), .B1(n15980), .Y(
        n19310) );
  sky130_fd_sc_hd__fa_1 U21048 ( .A(n15983), .B(n15982), .CIN(n15981), .COUT(
        n15987), .SUM(n15979) );
  sky130_fd_sc_hd__fa_1 U21049 ( .A(n15986), .B(n15985), .CIN(n15984), .COUT(
        n15989), .SUM(n15988) );
  sky130_fd_sc_hd__nor2_1 U21050 ( .A(n15987), .B(n15988), .Y(n19307) );
  sky130_fd_sc_hd__nand2_1 U21051 ( .A(n15988), .B(n15987), .Y(n19308) );
  sky130_fd_sc_hd__nand2_1 U21053 ( .A(n15990), .B(n15989), .Y(n19955) );
  sky130_fd_sc_hd__nand2_1 U21054 ( .A(n15992), .B(n15991), .Y(n16803) );
  sky130_fd_sc_hd__o21ai_1 U21055 ( .A1(n19955), .A2(n16802), .B1(n16803), .Y(
        n15993) );
  sky130_fd_sc_hd__a21oi_1 U21056 ( .A1(n15994), .A2(n16805), .B1(n15993), .Y(
        n17042) );
  sky130_fd_sc_hd__fa_1 U21057 ( .A(n15997), .B(n15996), .CIN(n15995), .COUT(
        n15859), .SUM(n16012) );
  sky130_fd_sc_hd__fa_1 U21058 ( .A(n16000), .B(n15999), .CIN(n15998), .COUT(
        n16011), .SUM(n16007) );
  sky130_fd_sc_hd__fa_1 U21059 ( .A(n16003), .B(n16002), .CIN(n16001), .COUT(
        n16006), .SUM(n16010) );
  sky130_fd_sc_hd__fa_1 U21060 ( .A(n16006), .B(n16005), .CIN(n16004), .COUT(
        n16020), .SUM(n16016) );
  sky130_fd_sc_hd__fa_1 U21061 ( .A(n16009), .B(n16008), .CIN(n16007), .COUT(
        n16013), .SUM(n15992) );
  sky130_fd_sc_hd__fa_1 U21062 ( .A(n16012), .B(n16011), .CIN(n16010), .COUT(
        n16015), .SUM(n16014) );
  sky130_fd_sc_hd__nand2_1 U21063 ( .A(n17045), .B(n18866), .Y(n16019) );
  sky130_fd_sc_hd__nand2_1 U21064 ( .A(n16014), .B(n16013), .Y(n18865) );
  sky130_fd_sc_hd__nand2_1 U21065 ( .A(n16016), .B(n16015), .Y(n17044) );
  sky130_fd_sc_hd__a21oi_1 U21066 ( .A1(n17045), .A2(n17043), .B1(n16017), .Y(
        n16018) );
  sky130_fd_sc_hd__nand2_1 U21068 ( .A(n16021), .B(n16020), .Y(n19108) );
  sky130_fd_sc_hd__nand2_1 U21069 ( .A(n16023), .B(n16022), .Y(n18987) );
  sky130_fd_sc_hd__a21oi_1 U21071 ( .A1(n16025), .A2(n18989), .B1(n16024), .Y(
        n16605) );
  sky130_fd_sc_hd__nand2_1 U21072 ( .A(n16027), .B(n16026), .Y(n16604) );
  sky130_fd_sc_hd__nand2_1 U21073 ( .A(n16029), .B(n16028), .Y(n19225) );
  sky130_fd_sc_hd__a21oi_1 U21074 ( .A1(n19226), .A2(n19222), .B1(n16030), .Y(
        n16031) );
  sky130_fd_sc_hd__nand2_1 U21076 ( .A(n16034), .B(n16033), .Y(n19856) );
  sky130_fd_sc_hd__nand2_1 U21077 ( .A(n16036), .B(n16035), .Y(n16830) );
  sky130_fd_sc_hd__a21oi_1 U21079 ( .A1(n16038), .A2(n16832), .B1(n16037), .Y(
        n17082) );
  sky130_fd_sc_hd__fa_1 U21080 ( .A(n16041), .B(n16040), .CIN(n16039), .COUT(
        n15674), .SUM(n16098) );
  sky130_fd_sc_hd__a222oi_1 U21081 ( .A1(n16044), .A2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .B1(n16043), .B2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .C1(n16042), .C2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .Y(n16045) );
  sky130_fd_sc_hd__o21ai_1 U21082 ( .A1(n16046), .A2(n16354), .B1(n16045), .Y(
        n16047) );
  sky130_fd_sc_hd__xor2_1 U21083 ( .A(n16047), .B(
        j202_soc_core_j22_cpu_ml_bufa[11]), .X(n16089) );
  sky130_fd_sc_hd__a222oi_1 U21084 ( .A1(n16050), .A2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .B1(n16049), .B2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .C1(n16048), .C2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .Y(n16051) );
  sky130_fd_sc_hd__o21ai_1 U21085 ( .A1(n16052), .A2(n16305), .B1(n16051), .Y(
        n16053) );
  sky130_fd_sc_hd__xor2_1 U21086 ( .A(n16053), .B(
        j202_soc_core_j22_cpu_ml_bufa[14]), .X(n16088) );
  sky130_fd_sc_hd__a222oi_1 U21087 ( .A1(n16056), .A2(n11170), .B1(n16055), 
        .B2(j202_soc_core_j22_cpu_ml_bufb[15]), .C1(n16054), .C2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .Y(n16057) );
  sky130_fd_sc_hd__o21ai_1 U21088 ( .A1(n16058), .A2(n16537), .B1(n16057), .Y(
        n16059) );
  sky130_fd_sc_hd__xor2_1 U21089 ( .A(n16059), .B(
        j202_soc_core_j22_cpu_ml_bufa[5]), .X(n16087) );
  sky130_fd_sc_hd__fa_1 U21090 ( .A(n16062), .B(n16061), .CIN(n16060), .COUT(
        n16077), .SUM(n16094) );
  sky130_fd_sc_hd__a222oi_1 U21091 ( .A1(n16065), .A2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .B1(n16064), .B2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .C1(n16063), .C2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .Y(n16066) );
  sky130_fd_sc_hd__xor2_1 U21093 ( .A(n16068), .B(
        j202_soc_core_j22_cpu_ml_bufa[8]), .X(n16104) );
  sky130_fd_sc_hd__fa_1 U21094 ( .A(n16071), .B(n16070), .CIN(n16069), .COUT(
        n16103), .SUM(n16090) );
  sky130_fd_sc_hd__fa_1 U21095 ( .A(n16074), .B(n16073), .CIN(n16072), .COUT(
        n16102), .SUM(n16106) );
  sky130_fd_sc_hd__fa_1 U21096 ( .A(n16077), .B(n16076), .CIN(n16075), .COUT(
        n16079), .SUM(n16096) );
  sky130_fd_sc_hd__fa_1 U21097 ( .A(n16080), .B(n16079), .CIN(n16078), .COUT(
        n16129), .SUM(n16124) );
  sky130_fd_sc_hd__nor2_1 U21098 ( .A(n16123), .B(n16124), .Y(n19002) );
  sky130_fd_sc_hd__fa_1 U21099 ( .A(n16083), .B(n16082), .CIN(n16081), .COUT(
        n16075), .SUM(n16116) );
  sky130_fd_sc_hd__fa_1 U21100 ( .A(n16086), .B(n16085), .CIN(n16084), .COUT(
        n16082), .SUM(n16110) );
  sky130_fd_sc_hd__fa_1 U21101 ( .A(n16089), .B(n16088), .CIN(n16087), .COUT(
        n16095), .SUM(n16109) );
  sky130_fd_sc_hd__fa_1 U21102 ( .A(n16092), .B(n16091), .CIN(n16090), .COUT(
        n16108), .SUM(n16101) );
  sky130_fd_sc_hd__fa_1 U21103 ( .A(n16095), .B(n16094), .CIN(n16093), .COUT(
        n16097), .SUM(n16114) );
  sky130_fd_sc_hd__fa_1 U21104 ( .A(n16098), .B(n16097), .CIN(n16096), .COUT(
        n16123), .SUM(n16122) );
  sky130_fd_sc_hd__nor2_1 U21105 ( .A(n16121), .B(n16122), .Y(n19131) );
  sky130_fd_sc_hd__nor2_1 U21106 ( .A(n19002), .B(n19131), .Y(n16126) );
  sky130_fd_sc_hd__fa_1 U21107 ( .A(n16101), .B(n16100), .CIN(n16099), .COUT(
        n16117), .SUM(n16036) );
  sky130_fd_sc_hd__fa_1 U21108 ( .A(n16104), .B(n16103), .CIN(n16102), .COUT(
        n16093), .SUM(n16113) );
  sky130_fd_sc_hd__fa_1 U21109 ( .A(n16107), .B(n16106), .CIN(n16105), .COUT(
        n16112), .SUM(n16099) );
  sky130_fd_sc_hd__fa_1 U21110 ( .A(n16110), .B(n16109), .CIN(n16108), .COUT(
        n16115), .SUM(n16111) );
  sky130_fd_sc_hd__nor2_1 U21111 ( .A(n16117), .B(n16118), .Y(n17083) );
  sky130_fd_sc_hd__fa_1 U21112 ( .A(n16113), .B(n16112), .CIN(n16111), .COUT(
        n16119), .SUM(n16118) );
  sky130_fd_sc_hd__fa_1 U21113 ( .A(n16116), .B(n16115), .CIN(n16114), .COUT(
        n16121), .SUM(n16120) );
  sky130_fd_sc_hd__nor2_1 U21114 ( .A(n16119), .B(n16120), .Y(n17085) );
  sky130_fd_sc_hd__nor2_1 U21115 ( .A(n17083), .B(n17085), .Y(n19006) );
  sky130_fd_sc_hd__nand2_1 U21116 ( .A(n16126), .B(n19006), .Y(n16128) );
  sky130_fd_sc_hd__nand2_1 U21117 ( .A(n16118), .B(n16117), .Y(n18878) );
  sky130_fd_sc_hd__nand2_1 U21118 ( .A(n16120), .B(n16119), .Y(n17086) );
  sky130_fd_sc_hd__nand2_1 U21120 ( .A(n16122), .B(n16121), .Y(n19132) );
  sky130_fd_sc_hd__nand2_1 U21121 ( .A(n16124), .B(n16123), .Y(n19003) );
  sky130_fd_sc_hd__a21oi_1 U21123 ( .A1(n16126), .A2(n19005), .B1(n16125), .Y(
        n16127) );
  sky130_fd_sc_hd__nand2_1 U21125 ( .A(n16130), .B(n16129), .Y(n19298) );
  sky130_fd_sc_hd__nand2_1 U21126 ( .A(n16132), .B(n16131), .Y(n19296) );
  sky130_fd_sc_hd__o21ai_1 U21127 ( .A1(n19298), .A2(n19295), .B1(n19296), .Y(
        n16788) );
  sky130_fd_sc_hd__nand2_1 U21128 ( .A(n16134), .B(n16133), .Y(n19949) );
  sky130_fd_sc_hd__nand2_1 U21129 ( .A(n16136), .B(n16135), .Y(n16794) );
  sky130_fd_sc_hd__a21oi_1 U21131 ( .A1(n16788), .A2(n16138), .B1(n16137), .Y(
        n17030) );
  sky130_fd_sc_hd__nand2_1 U21132 ( .A(n16140), .B(n16139), .Y(n18860) );
  sky130_fd_sc_hd__nand2_1 U21133 ( .A(n16142), .B(n16141), .Y(n17035) );
  sky130_fd_sc_hd__nand2_1 U21135 ( .A(n16144), .B(n16143), .Y(n19100) );
  sky130_fd_sc_hd__nand2_1 U21136 ( .A(n16146), .B(n16145), .Y(n18980) );
  sky130_fd_sc_hd__o21ai_1 U21137 ( .A1(n19100), .A2(n18979), .B1(n18980), .Y(
        n16147) );
  sky130_fd_sc_hd__a21oi_1 U21138 ( .A1(n16148), .A2(n18973), .B1(n16147), .Y(
        n16149) );
  sky130_fd_sc_hd__a21oi_1 U21140 ( .A1(n16152), .A2(n16625), .B1(n16151), .Y(
        n19361) );
  sky130_fd_sc_hd__a222oi_1 U21141 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .Y(n16153) );
  sky130_fd_sc_hd__xor2_1 U21143 ( .A(n16154), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n16255) );
  sky130_fd_sc_hd__xnor2_1 U21144 ( .A(j202_soc_core_j22_cpu_ml_bufa[31]), .B(
        j202_soc_core_j22_cpu_ml_bufa[30]), .Y(n16156) );
  sky130_fd_sc_hd__nor2b_1 U21145 ( .B_N(n16157), .A(n16156), .Y(n19333) );
  sky130_fd_sc_hd__and3_1 U21146 ( .A(n16157), .B(n16156), .C(n16155), .X(
        n19332) );
  sky130_fd_sc_hd__a222oi_1 U21147 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .Y(n16158) );
  sky130_fd_sc_hd__o21ai_1 U21148 ( .A1(n19336), .A2(n16159), .B1(n16158), .Y(
        n16160) );
  sky130_fd_sc_hd__xor2_1 U21149 ( .A(n16160), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16231) );
  sky130_fd_sc_hd__a222oi_1 U21150 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .Y(n16161) );
  sky130_fd_sc_hd__xor2_1 U21152 ( .A(n16162), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16230) );
  sky130_fd_sc_hd__a22oi_1 U21153 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n16163) );
  sky130_fd_sc_hd__o21ai_1 U21154 ( .A1(n19336), .A2(n16164), .B1(n16163), .Y(
        n16165) );
  sky130_fd_sc_hd__xor2_1 U21155 ( .A(n16165), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16184) );
  sky130_fd_sc_hd__a22oi_1 U21156 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[16]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[0]), .Y(n16166) );
  sky130_fd_sc_hd__nand2_1 U21157 ( .A(n16546), .B(n16166), .Y(n16181) );
  sky130_fd_sc_hd__a222oi_1 U21158 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[1]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[0]), .Y(n16167) );
  sky130_fd_sc_hd__o21ai_1 U21159 ( .A1(n19336), .A2(n16168), .B1(n16167), .Y(
        n16169) );
  sky130_fd_sc_hd__xor2_1 U21160 ( .A(n16169), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16180) );
  sky130_fd_sc_hd__a22oi_1 U21161 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[18]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[2]), .Y(n16170) );
  sky130_fd_sc_hd__nand2_1 U21162 ( .A(n16546), .B(n16170), .Y(n16270) );
  sky130_fd_sc_hd__a222oi_1 U21163 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .Y(n16171) );
  sky130_fd_sc_hd__xor2_1 U21165 ( .A(n16172), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16235) );
  sky130_fd_sc_hd__a222oi_1 U21166 ( .A1(n16225), .A2(n11170), .B1(n16224), 
        .B2(n11170), .C1(n16223), .C2(n11170), .Y(n16173) );
  sky130_fd_sc_hd__o21ai_1 U21167 ( .A1(n11169), .A2(n16227), .B1(n16173), .Y(
        n16174) );
  sky130_fd_sc_hd__xnor2_1 U21168 ( .A(j202_soc_core_j22_cpu_ml_bufa[17]), .B(
        n16174), .Y(n16183) );
  sky130_fd_sc_hd__a22oi_1 U21169 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[17]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[1]), .Y(n16175) );
  sky130_fd_sc_hd__nand2_1 U21170 ( .A(n16546), .B(n16175), .Y(n16182) );
  sky130_fd_sc_hd__a222oi_1 U21171 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .Y(n16176) );
  sky130_fd_sc_hd__o21ai_1 U21172 ( .A1(n16265), .A2(n16557), .B1(n16176), .Y(
        n16177) );
  sky130_fd_sc_hd__xor2_1 U21173 ( .A(n16177), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n16469) );
  sky130_fd_sc_hd__a222oi_1 U21174 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .Y(n16178) );
  sky130_fd_sc_hd__o21ai_1 U21175 ( .A1(n16327), .A2(n16379), .B1(n16178), .Y(
        n16179) );
  sky130_fd_sc_hd__xor2_1 U21176 ( .A(n16179), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n16468) );
  sky130_fd_sc_hd__fa_1 U21177 ( .A(n16436), .B(n16181), .CIN(n16180), .COUT(
        n16229), .SUM(n16467) );
  sky130_fd_sc_hd__fa_1 U21178 ( .A(n16184), .B(n16183), .CIN(n16182), .COUT(
        n16234), .SUM(n16210) );
  sky130_fd_sc_hd__a222oi_1 U21179 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[15]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .Y(n16185) );
  sky130_fd_sc_hd__o21ai_1 U21180 ( .A1(n16265), .A2(n16540), .B1(n16185), .Y(
        n16186) );
  sky130_fd_sc_hd__xor2_1 U21181 ( .A(n16186), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n16209) );
  sky130_fd_sc_hd__a222oi_1 U21182 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .Y(n16187) );
  sky130_fd_sc_hd__o21ai_1 U21183 ( .A1(n16373), .A2(n16319), .B1(n16187), .Y(
        n16188) );
  sky130_fd_sc_hd__xor2_1 U21184 ( .A(n16188), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n16208) );
  sky130_fd_sc_hd__o22ai_1 U21185 ( .A1(n16191), .A2(n16582), .B1(n16190), 
        .B2(n16189), .Y(n16435) );
  sky130_fd_sc_hd__a222oi_1 U21186 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[2]), .Y(n16192) );
  sky130_fd_sc_hd__xor2_1 U21188 ( .A(n16194), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16434) );
  sky130_fd_sc_hd__fa_1 U21189 ( .A(j202_soc_core_j22_cpu_ml_bufa[32]), .B(
        n16196), .CIN(n16195), .COUT(n16448), .SUM(n16439) );
  sky130_fd_sc_hd__fa_1 U21190 ( .A(n16199), .B(n16198), .CIN(n16197), .COUT(
        n16447), .SUM(n16440) );
  sky130_fd_sc_hd__a222oi_1 U21191 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .Y(n16200) );
  sky130_fd_sc_hd__o21ai_1 U21192 ( .A1(n16327), .A2(n16354), .B1(n16200), .Y(
        n16201) );
  sky130_fd_sc_hd__xor2_1 U21193 ( .A(n16201), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n16446) );
  sky130_fd_sc_hd__a222oi_1 U21194 ( .A1(n16263), .A2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .B1(n16262), .B2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .Y(n16202) );
  sky130_fd_sc_hd__o21ai_1 U21195 ( .A1(n16265), .A2(n16402), .B1(n16202), .Y(
        n16203) );
  sky130_fd_sc_hd__xor2_1 U21196 ( .A(n16203), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n16451) );
  sky130_fd_sc_hd__a222oi_1 U21197 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .Y(n16204) );
  sky130_fd_sc_hd__o21ai_1 U21198 ( .A1(n16373), .A2(n16305), .B1(n16204), .Y(
        n16205) );
  sky130_fd_sc_hd__xor2_1 U21199 ( .A(n16205), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n16450) );
  sky130_fd_sc_hd__a222oi_1 U21200 ( .A1(n16225), .A2(n11170), .B1(n16224), 
        .B2(j202_soc_core_j22_cpu_ml_bufb[15]), .C1(n16223), .C2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .Y(n16206) );
  sky130_fd_sc_hd__xor2_1 U21202 ( .A(n16207), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n16449) );
  sky130_fd_sc_hd__fa_1 U21203 ( .A(n16210), .B(n16209), .CIN(n16208), .COUT(
        n16242), .SUM(n16480) );
  sky130_fd_sc_hd__a222oi_1 U21204 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .Y(n16211) );
  sky130_fd_sc_hd__o21ai_1 U21205 ( .A1(n16373), .A2(n16354), .B1(n16211), .Y(
        n16212) );
  sky130_fd_sc_hd__xor2_1 U21206 ( .A(n16212), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n16245) );
  sky130_fd_sc_hd__a222oi_1 U21207 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .Y(n16213) );
  sky130_fd_sc_hd__o21ai_1 U21208 ( .A1(n16551), .A2(n16305), .B1(n16213), .Y(
        n16214) );
  sky130_fd_sc_hd__xor2_1 U21209 ( .A(n16214), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16244) );
  sky130_fd_sc_hd__a222oi_1 U21210 ( .A1(n16263), .A2(n11170), .B1(n16262), 
        .B2(j202_soc_core_j22_cpu_ml_bufb[15]), .C1(n16261), .C2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .Y(n16215) );
  sky130_fd_sc_hd__o21ai_1 U21211 ( .A1(n16265), .A2(n16537), .B1(n16215), .Y(
        n16216) );
  sky130_fd_sc_hd__xor2_1 U21212 ( .A(n16216), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n16243) );
  sky130_fd_sc_hd__a222oi_1 U21213 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .Y(n16217) );
  sky130_fd_sc_hd__o21ai_1 U21214 ( .A1(n16327), .A2(n16367), .B1(n16217), .Y(
        n16218) );
  sky130_fd_sc_hd__xor2_1 U21215 ( .A(n16218), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n16475) );
  sky130_fd_sc_hd__a222oi_1 U21216 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .Y(n16219) );
  sky130_fd_sc_hd__o21ai_1 U21217 ( .A1(n16373), .A2(n16311), .B1(n16219), .Y(
        n16220) );
  sky130_fd_sc_hd__xor2_1 U21218 ( .A(n16220), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n16466) );
  sky130_fd_sc_hd__a222oi_1 U21219 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .Y(n16221) );
  sky130_fd_sc_hd__o21ai_1 U21220 ( .A1(n16551), .A2(n16247), .B1(n16221), .Y(
        n16222) );
  sky130_fd_sc_hd__xor2_1 U21221 ( .A(n16222), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16465) );
  sky130_fd_sc_hd__a222oi_1 U21222 ( .A1(n16225), .A2(n11170), .B1(n16224), 
        .B2(n11170), .C1(n16223), .C2(j202_soc_core_j22_cpu_ml_bufb[15]), .Y(
        n16226) );
  sky130_fd_sc_hd__xor2_1 U21224 ( .A(n16228), .B(
        j202_soc_core_j22_cpu_ml_bufa[17]), .X(n16464) );
  sky130_fd_sc_hd__fa_1 U21225 ( .A(n16231), .B(n16230), .CIN(n16229), .COUT(
        n16254), .SUM(n16473) );
  sky130_fd_sc_hd__a222oi_1 U21226 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .Y(n16232) );
  sky130_fd_sc_hd__o21ai_1 U21227 ( .A1(n16373), .A2(n16379), .B1(n16232), .Y(
        n16233) );
  sky130_fd_sc_hd__xor2_1 U21228 ( .A(n16233), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n16286) );
  sky130_fd_sc_hd__fa_1 U21229 ( .A(n16236), .B(n16235), .CIN(n16234), .COUT(
        n16285), .SUM(n16253) );
  sky130_fd_sc_hd__a22oi_1 U21230 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[19]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[3]), .Y(n16237) );
  sky130_fd_sc_hd__nand2_1 U21231 ( .A(n16546), .B(n16237), .Y(n16298) );
  sky130_fd_sc_hd__a222oi_1 U21232 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .Y(n16238) );
  sky130_fd_sc_hd__o21ai_1 U21233 ( .A1(n16551), .A2(n16311), .B1(n16238), .Y(
        n16239) );
  sky130_fd_sc_hd__xor2_1 U21234 ( .A(n16239), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16268) );
  sky130_fd_sc_hd__fa_1 U21235 ( .A(n16242), .B(n16241), .CIN(n16240), .COUT(
        n16257), .SUM(n16482) );
  sky130_fd_sc_hd__fa_1 U21236 ( .A(n16245), .B(n16244), .CIN(n16243), .COUT(
        n16273), .SUM(n16241) );
  sky130_fd_sc_hd__a222oi_1 U21237 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[3]), .Y(n16246) );
  sky130_fd_sc_hd__o21ai_1 U21238 ( .A1(n19336), .A2(n16247), .B1(n16246), .Y(
        n16248) );
  sky130_fd_sc_hd__xor2_1 U21239 ( .A(n16248), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16276) );
  sky130_fd_sc_hd__a222oi_1 U21240 ( .A1(n16263), .A2(n11170), .B1(n16262), 
        .B2(n11170), .C1(n16261), .C2(j202_soc_core_j22_cpu_ml_bufb[15]), .Y(
        n16249) );
  sky130_fd_sc_hd__o21ai_1 U21241 ( .A1(n16265), .A2(n16584), .B1(n16249), .Y(
        n16250) );
  sky130_fd_sc_hd__xor2_1 U21242 ( .A(n16250), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .X(n16275) );
  sky130_fd_sc_hd__a222oi_1 U21243 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .Y(n16251) );
  sky130_fd_sc_hd__o21ai_1 U21244 ( .A1(n16327), .A2(n16557), .B1(n16251), .Y(
        n16252) );
  sky130_fd_sc_hd__xor2_1 U21245 ( .A(n16252), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n16274) );
  sky130_fd_sc_hd__fa_1 U21246 ( .A(n16255), .B(n16254), .CIN(n16253), .COUT(
        n16271), .SUM(n16484) );
  sky130_fd_sc_hd__nor2_1 U21247 ( .A(n16501), .B(n16502), .Y(n18873) );
  sky130_fd_sc_hd__fa_1 U21248 ( .A(n16258), .B(n16257), .CIN(n16256), .COUT(
        n16503), .SUM(n16502) );
  sky130_fd_sc_hd__a222oi_1 U21249 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .Y(n16259) );
  sky130_fd_sc_hd__xor2_1 U21251 ( .A(n16260), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n16418) );
  sky130_fd_sc_hd__a222oi_1 U21252 ( .A1(n16263), .A2(n11170), .B1(n16262), 
        .B2(n11170), .C1(n16261), .C2(n11170), .Y(n16264) );
  sky130_fd_sc_hd__xnor2_1 U21254 ( .A(j202_soc_core_j22_cpu_ml_bufa[20]), .B(
        n16266), .Y(n16299) );
  sky130_fd_sc_hd__a22oi_1 U21255 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[20]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[4]), .Y(n16267) );
  sky130_fd_sc_hd__nand2_1 U21256 ( .A(n16546), .B(n16267), .Y(n16297) );
  sky130_fd_sc_hd__fa_1 U21257 ( .A(n16270), .B(n16269), .CIN(n16268), .COUT(
        n16416), .SUM(n16284) );
  sky130_fd_sc_hd__fa_1 U21258 ( .A(n16273), .B(n16272), .CIN(n16271), .COUT(
        n16414), .SUM(n16256) );
  sky130_fd_sc_hd__fa_1 U21259 ( .A(n16276), .B(n16275), .CIN(n16274), .COUT(
        n16424), .SUM(n16272) );
  sky130_fd_sc_hd__a222oi_1 U21260 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[4]), .Y(n16277) );
  sky130_fd_sc_hd__o21ai_1 U21261 ( .A1(n19336), .A2(n16278), .B1(n16277), .Y(
        n16279) );
  sky130_fd_sc_hd__xor2_1 U21262 ( .A(n16279), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16295) );
  sky130_fd_sc_hd__a222oi_1 U21263 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .Y(n16280) );
  sky130_fd_sc_hd__o21ai_1 U21264 ( .A1(n16551), .A2(n16319), .B1(n16280), .Y(
        n16281) );
  sky130_fd_sc_hd__xor2_1 U21265 ( .A(n16281), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16294) );
  sky130_fd_sc_hd__a222oi_1 U21266 ( .A1(n16325), .A2(
        j202_soc_core_j22_cpu_ml_bufb[15]), .B1(n16324), .B2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .Y(n16282) );
  sky130_fd_sc_hd__o21ai_1 U21267 ( .A1(n16327), .A2(n16540), .B1(n16282), .Y(
        n16283) );
  sky130_fd_sc_hd__xor2_1 U21268 ( .A(n16283), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n16293) );
  sky130_fd_sc_hd__fa_1 U21269 ( .A(n16286), .B(n16285), .CIN(n16284), .COUT(
        n16422), .SUM(n16258) );
  sky130_fd_sc_hd__nor2_1 U21270 ( .A(n16503), .B(n16504), .Y(n17076) );
  sky130_fd_sc_hd__nor2_1 U21271 ( .A(n18873), .B(n17076), .Y(n16619) );
  sky130_fd_sc_hd__a222oi_1 U21272 ( .A1(n16325), .A2(n11170), .B1(n16324), 
        .B2(n11170), .C1(n16323), .C2(j202_soc_core_j22_cpu_ml_bufb[15]), .Y(
        n16287) );
  sky130_fd_sc_hd__o21ai_1 U21273 ( .A1(n16327), .A2(n16584), .B1(n16287), .Y(
        n16288) );
  sky130_fd_sc_hd__xor2_1 U21274 ( .A(n16288), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n16340) );
  sky130_fd_sc_hd__a222oi_1 U21275 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .Y(n16289) );
  sky130_fd_sc_hd__o21ai_1 U21276 ( .A1(n16551), .A2(n16379), .B1(n16289), .Y(
        n16290) );
  sky130_fd_sc_hd__xor2_1 U21277 ( .A(n16290), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16339) );
  sky130_fd_sc_hd__a222oi_1 U21278 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .Y(n16291) );
  sky130_fd_sc_hd__xor2_1 U21280 ( .A(n16292), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n16338) );
  sky130_fd_sc_hd__fa_1 U21281 ( .A(n16295), .B(n16294), .CIN(n16293), .COUT(
        n16421), .SUM(n16423) );
  sky130_fd_sc_hd__a22oi_1 U21282 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[21]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[5]), .Y(n16296) );
  sky130_fd_sc_hd__nand2_1 U21283 ( .A(n16546), .B(n16296), .Y(n16346) );
  sky130_fd_sc_hd__fa_1 U21284 ( .A(n16299), .B(n16298), .CIN(n16297), .COUT(
        n16314), .SUM(n16417) );
  sky130_fd_sc_hd__a222oi_1 U21285 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .Y(n16300) );
  sky130_fd_sc_hd__o21ai_1 U21286 ( .A1(n16373), .A2(n16402), .B1(n16300), .Y(
        n16301) );
  sky130_fd_sc_hd__xor2_1 U21287 ( .A(n16301), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n16313) );
  sky130_fd_sc_hd__a222oi_1 U21288 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .Y(n16302) );
  sky130_fd_sc_hd__o21ai_1 U21289 ( .A1(n16551), .A2(n16354), .B1(n16302), .Y(
        n16303) );
  sky130_fd_sc_hd__xor2_1 U21290 ( .A(n16303), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16317) );
  sky130_fd_sc_hd__a222oi_1 U21291 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[5]), .Y(n16304) );
  sky130_fd_sc_hd__o21ai_1 U21292 ( .A1(n19336), .A2(n16305), .B1(n16304), .Y(
        n16306) );
  sky130_fd_sc_hd__xor2_1 U21293 ( .A(n16306), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16316) );
  sky130_fd_sc_hd__a222oi_1 U21294 ( .A1(n16325), .A2(n11170), .B1(n16324), 
        .B2(j202_soc_core_j22_cpu_ml_bufb[15]), .C1(n16323), .C2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .Y(n16307) );
  sky130_fd_sc_hd__xor2_1 U21296 ( .A(n16308), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .X(n16315) );
  sky130_fd_sc_hd__a22oi_1 U21297 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[22]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[6]), .Y(n16309) );
  sky130_fd_sc_hd__nand2_1 U21298 ( .A(n16546), .B(n16309), .Y(n16337) );
  sky130_fd_sc_hd__a222oi_1 U21299 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[6]), .Y(n16310) );
  sky130_fd_sc_hd__o21ai_1 U21300 ( .A1(n19336), .A2(n16311), .B1(n16310), .Y(
        n16312) );
  sky130_fd_sc_hd__xor2_1 U21301 ( .A(n16312), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16335) );
  sky130_fd_sc_hd__fa_1 U21302 ( .A(n16336), .B(n16314), .CIN(n16313), .COUT(
        n16331), .SUM(n16420) );
  sky130_fd_sc_hd__fa_1 U21303 ( .A(n16317), .B(n16316), .CIN(n16315), .COUT(
        n16330), .SUM(n16419) );
  sky130_fd_sc_hd__a222oi_1 U21304 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[7]), .Y(n16318) );
  sky130_fd_sc_hd__o21ai_1 U21305 ( .A1(n19336), .A2(n16319), .B1(n16318), .Y(
        n16320) );
  sky130_fd_sc_hd__xor2_1 U21306 ( .A(n16320), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16360) );
  sky130_fd_sc_hd__a222oi_1 U21307 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .Y(n16321) );
  sky130_fd_sc_hd__xor2_1 U21309 ( .A(n16322), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16359) );
  sky130_fd_sc_hd__a222oi_1 U21310 ( .A1(n16325), .A2(n11170), .B1(n16324), 
        .B2(n11170), .C1(n16323), .C2(n11170), .Y(n16326) );
  sky130_fd_sc_hd__o21ai_1 U21311 ( .A1(n11169), .A2(n16327), .B1(n16326), .Y(
        n16328) );
  sky130_fd_sc_hd__xnor2_1 U21312 ( .A(j202_soc_core_j22_cpu_ml_bufa[23]), .B(
        n16328), .Y(n16347) );
  sky130_fd_sc_hd__a22oi_1 U21313 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[23]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[7]), .Y(n16329) );
  sky130_fd_sc_hd__nand2_1 U21314 ( .A(n16546), .B(n16329), .Y(n16345) );
  sky130_fd_sc_hd__fa_1 U21315 ( .A(n16332), .B(n16331), .CIN(n16330), .COUT(
        n16342), .SUM(n16425) );
  sky130_fd_sc_hd__a222oi_1 U21316 ( .A1(n16371), .A2(
        j202_soc_core_j22_cpu_ml_bufb[15]), .B1(n16370), .B2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .Y(n16333) );
  sky130_fd_sc_hd__o21ai_1 U21317 ( .A1(n16373), .A2(n16540), .B1(n16333), .Y(
        n16334) );
  sky130_fd_sc_hd__xor2_1 U21318 ( .A(n16334), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n16352) );
  sky130_fd_sc_hd__fa_1 U21319 ( .A(n16337), .B(n16336), .CIN(n16335), .COUT(
        n16351), .SUM(n16332) );
  sky130_fd_sc_hd__fa_1 U21320 ( .A(n16340), .B(n16339), .CIN(n16338), .COUT(
        n16350), .SUM(n16427) );
  sky130_fd_sc_hd__nor2_1 U21321 ( .A(n16511), .B(n16512), .Y(n19292) );
  sky130_fd_sc_hd__fa_1 U21322 ( .A(n16343), .B(n16342), .CIN(n16341), .COUT(
        n16513), .SUM(n16512) );
  sky130_fd_sc_hd__a22oi_1 U21323 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[24]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[8]), .Y(n16344) );
  sky130_fd_sc_hd__nand2_1 U21324 ( .A(n16546), .B(n16344), .Y(n16399) );
  sky130_fd_sc_hd__fa_1 U21325 ( .A(n16347), .B(n16346), .CIN(n16345), .COUT(
        n16382), .SUM(n16358) );
  sky130_fd_sc_hd__a222oi_1 U21326 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .Y(n16348) );
  sky130_fd_sc_hd__xor2_1 U21328 ( .A(n16349), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16381) );
  sky130_fd_sc_hd__fa_1 U21329 ( .A(n16352), .B(n16351), .CIN(n16350), .COUT(
        n16408), .SUM(n16341) );
  sky130_fd_sc_hd__a222oi_1 U21330 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[8]), .Y(n16353) );
  sky130_fd_sc_hd__o21ai_1 U21331 ( .A1(n19336), .A2(n16354), .B1(n16353), .Y(
        n16355) );
  sky130_fd_sc_hd__xor2_1 U21332 ( .A(n16355), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16388) );
  sky130_fd_sc_hd__a222oi_1 U21333 ( .A1(n16371), .A2(n11170), .B1(n16370), 
        .B2(j202_soc_core_j22_cpu_ml_bufb[15]), .C1(n16369), .C2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .Y(n16356) );
  sky130_fd_sc_hd__o21ai_1 U21334 ( .A1(n16373), .A2(n16537), .B1(n16356), .Y(
        n16357) );
  sky130_fd_sc_hd__xor2_1 U21335 ( .A(n16357), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n16387) );
  sky130_fd_sc_hd__fa_1 U21336 ( .A(n16360), .B(n16359), .CIN(n16358), .COUT(
        n16386), .SUM(n16343) );
  sky130_fd_sc_hd__nor2_1 U21337 ( .A(n16513), .B(n16514), .Y(n19287) );
  sky130_fd_sc_hd__nor2_1 U21338 ( .A(n19292), .B(n19287), .Y(n16784) );
  sky130_fd_sc_hd__a22oi_1 U21339 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[25]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[9]), .Y(n16361) );
  sky130_fd_sc_hd__nand2_1 U21340 ( .A(n16546), .B(n16361), .Y(n16385) );
  sky130_fd_sc_hd__a222oi_1 U21341 ( .A1(n16371), .A2(n11170), .B1(n16370), 
        .B2(n11170), .C1(n16369), .C2(j202_soc_core_j22_cpu_ml_bufb[15]), .Y(
        n16362) );
  sky130_fd_sc_hd__o21ai_1 U21342 ( .A1(n16373), .A2(n16584), .B1(n16362), .Y(
        n16363) );
  sky130_fd_sc_hd__xor2_1 U21343 ( .A(n16363), .B(
        j202_soc_core_j22_cpu_ml_bufa[26]), .X(n16383) );
  sky130_fd_sc_hd__a222oi_1 U21344 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[15]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .Y(n16364) );
  sky130_fd_sc_hd__o21ai_1 U21345 ( .A1(n16551), .A2(n16540), .B1(n16364), .Y(
        n16365) );
  sky130_fd_sc_hd__xor2_1 U21346 ( .A(n16365), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16396) );
  sky130_fd_sc_hd__a222oi_1 U21347 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .Y(n16366) );
  sky130_fd_sc_hd__xor2_1 U21349 ( .A(n16368), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16395) );
  sky130_fd_sc_hd__a222oi_1 U21350 ( .A1(n16371), .A2(n11170), .B1(n16370), 
        .B2(n11170), .C1(n16369), .C2(n11170), .Y(n16372) );
  sky130_fd_sc_hd__o21ai_1 U21351 ( .A1(n11169), .A2(n16373), .B1(n16372), .Y(
        n16374) );
  sky130_fd_sc_hd__xnor2_1 U21352 ( .A(j202_soc_core_j22_cpu_ml_bufa[26]), .B(
        n16374), .Y(n16400) );
  sky130_fd_sc_hd__a22oi_1 U21353 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[26]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[10]), .Y(n16375) );
  sky130_fd_sc_hd__nand2_1 U21354 ( .A(n16546), .B(n16375), .Y(n16398) );
  sky130_fd_sc_hd__a222oi_1 U21355 ( .A1(n16549), .A2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .B1(n16548), .B2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .Y(n16376) );
  sky130_fd_sc_hd__o21ai_1 U21356 ( .A1(n16551), .A2(n16557), .B1(n16376), .Y(
        n16377) );
  sky130_fd_sc_hd__xor2_1 U21357 ( .A(n16377), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16391) );
  sky130_fd_sc_hd__a222oi_1 U21358 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[10]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[9]), .Y(n16378) );
  sky130_fd_sc_hd__o21ai_1 U21359 ( .A1(n19336), .A2(n16379), .B1(n16378), .Y(
        n16380) );
  sky130_fd_sc_hd__xor2_1 U21360 ( .A(n16380), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16390) );
  sky130_fd_sc_hd__fa_1 U21361 ( .A(n16384), .B(n16382), .CIN(n16381), .COUT(
        n16389), .SUM(n16409) );
  sky130_fd_sc_hd__fa_1 U21362 ( .A(n16385), .B(n16384), .CIN(n16383), .COUT(
        n16406), .SUM(n16412) );
  sky130_fd_sc_hd__fa_1 U21363 ( .A(n16388), .B(n16387), .CIN(n16386), .COUT(
        n16411), .SUM(n16407) );
  sky130_fd_sc_hd__fa_1 U21364 ( .A(n16391), .B(n16390), .CIN(n16389), .COUT(
        n16404), .SUM(n16410) );
  sky130_fd_sc_hd__a222oi_1 U21365 ( .A1(n16549), .A2(n11170), .B1(n16548), 
        .B2(j202_soc_core_j22_cpu_ml_bufb[15]), .C1(n16547), .C2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .Y(n16392) );
  sky130_fd_sc_hd__o21ai_1 U21366 ( .A1(n16551), .A2(n16537), .B1(n16392), .Y(
        n16393) );
  sky130_fd_sc_hd__xor2_1 U21367 ( .A(n16393), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16555) );
  sky130_fd_sc_hd__fa_1 U21368 ( .A(n16396), .B(n16395), .CIN(n16394), .COUT(
        n16554), .SUM(n16405) );
  sky130_fd_sc_hd__a22oi_1 U21369 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[27]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[11]), .Y(n16397) );
  sky130_fd_sc_hd__nand2_1 U21370 ( .A(n16546), .B(n16397), .Y(n16543) );
  sky130_fd_sc_hd__fa_1 U21371 ( .A(n16400), .B(n16399), .CIN(n16398), .COUT(
        n16560), .SUM(n16394) );
  sky130_fd_sc_hd__a222oi_1 U21372 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[11]), .Y(n16401) );
  sky130_fd_sc_hd__o21ai_1 U21373 ( .A1(n19336), .A2(n16402), .B1(n16401), .Y(
        n16403) );
  sky130_fd_sc_hd__xor2_1 U21374 ( .A(n16403), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16559) );
  sky130_fd_sc_hd__fa_1 U21375 ( .A(n16406), .B(n16405), .CIN(n16404), .COUT(
        n16520), .SUM(n16517) );
  sky130_fd_sc_hd__nand2_1 U21376 ( .A(n18853), .B(n18856), .Y(n16523) );
  sky130_fd_sc_hd__fa_1 U21377 ( .A(n16409), .B(n16408), .CIN(n16407), .COUT(
        n16515), .SUM(n16514) );
  sky130_fd_sc_hd__fa_1 U21378 ( .A(n16412), .B(n16411), .CIN(n16410), .COUT(
        n16518), .SUM(n16516) );
  sky130_fd_sc_hd__nor2_1 U21379 ( .A(n16515), .B(n16516), .Y(n19941) );
  sky130_fd_sc_hd__nor2_1 U21380 ( .A(n16523), .B(n19941), .Y(n16525) );
  sky130_fd_sc_hd__nand2_1 U21381 ( .A(n16784), .B(n16525), .Y(n16527) );
  sky130_fd_sc_hd__fa_1 U21382 ( .A(n16415), .B(n16414), .CIN(n16413), .COUT(
        n16505), .SUM(n16504) );
  sky130_fd_sc_hd__fa_1 U21383 ( .A(n16418), .B(n16417), .CIN(n16416), .COUT(
        n16430), .SUM(n16415) );
  sky130_fd_sc_hd__fa_1 U21384 ( .A(n16421), .B(n16420), .CIN(n16419), .COUT(
        n16426), .SUM(n16429) );
  sky130_fd_sc_hd__fa_1 U21385 ( .A(n16424), .B(n16423), .CIN(n16422), .COUT(
        n16428), .SUM(n16413) );
  sky130_fd_sc_hd__nor2_1 U21386 ( .A(n16505), .B(n16506), .Y(n18999) );
  sky130_fd_sc_hd__fa_1 U21387 ( .A(n16427), .B(n16426), .CIN(n16425), .COUT(
        n16511), .SUM(n16507) );
  sky130_fd_sc_hd__fa_1 U21388 ( .A(n16430), .B(n16429), .CIN(n16428), .COUT(
        n16508), .SUM(n16506) );
  sky130_fd_sc_hd__nand2_1 U21389 ( .A(n19128), .B(n18997), .Y(n16620) );
  sky130_fd_sc_hd__nor2_1 U21390 ( .A(n16527), .B(n16620), .Y(n16529) );
  sky130_fd_sc_hd__nand2_1 U21391 ( .A(n16619), .B(n16529), .Y(n16531) );
  sky130_fd_sc_hd__fa_1 U21392 ( .A(n16433), .B(n16432), .CIN(n16431), .COUT(
        n16491), .SUM(n16146) );
  sky130_fd_sc_hd__fa_1 U21393 ( .A(n16436), .B(n16435), .CIN(n16434), .COUT(
        n16460), .SUM(n16472) );
  sky130_fd_sc_hd__fa_1 U21394 ( .A(n16439), .B(n16438), .CIN(n16437), .COUT(
        n16471), .SUM(n16452) );
  sky130_fd_sc_hd__fa_1 U21395 ( .A(n16442), .B(n16441), .CIN(n16440), .COUT(
        n16470), .SUM(n16444) );
  sky130_fd_sc_hd__fa_1 U21396 ( .A(n16445), .B(n16444), .CIN(n16443), .COUT(
        n16456), .SUM(n16431) );
  sky130_fd_sc_hd__fa_1 U21397 ( .A(n16448), .B(n16447), .CIN(n16446), .COUT(
        n16459), .SUM(n16463) );
  sky130_fd_sc_hd__fa_1 U21398 ( .A(n16451), .B(n16450), .CIN(n16449), .COUT(
        n16458), .SUM(n16462) );
  sky130_fd_sc_hd__fa_1 U21399 ( .A(n16454), .B(n16453), .CIN(n16452), .COUT(
        n16461), .SUM(n16433) );
  sky130_fd_sc_hd__nor2_1 U21400 ( .A(n16491), .B(n16492), .Y(n16600) );
  sky130_fd_sc_hd__fa_1 U21401 ( .A(n16457), .B(n16456), .CIN(n16455), .COUT(
        n16493), .SUM(n16492) );
  sky130_fd_sc_hd__fa_1 U21402 ( .A(n16460), .B(n16459), .CIN(n16458), .COUT(
        n16479), .SUM(n16487) );
  sky130_fd_sc_hd__fa_1 U21403 ( .A(n16463), .B(n16462), .CIN(n16461), .COUT(
        n16486), .SUM(n16455) );
  sky130_fd_sc_hd__fa_1 U21404 ( .A(n16466), .B(n16465), .CIN(n16464), .COUT(
        n16474), .SUM(n16478) );
  sky130_fd_sc_hd__fa_1 U21405 ( .A(n16469), .B(n16468), .CIN(n16467), .COUT(
        n16481), .SUM(n16477) );
  sky130_fd_sc_hd__fa_1 U21406 ( .A(n16472), .B(n16471), .CIN(n16470), .COUT(
        n16476), .SUM(n16457) );
  sky130_fd_sc_hd__nor2_1 U21407 ( .A(n16493), .B(n16494), .Y(n19217) );
  sky130_fd_sc_hd__nor2_1 U21408 ( .A(n16600), .B(n19217), .Y(n16826) );
  sky130_fd_sc_hd__fa_1 U21409 ( .A(n16475), .B(n16474), .CIN(n16473), .COUT(
        n16240), .SUM(n16490) );
  sky130_fd_sc_hd__fa_1 U21410 ( .A(n16478), .B(n16477), .CIN(n16476), .COUT(
        n16489), .SUM(n16485) );
  sky130_fd_sc_hd__fa_1 U21411 ( .A(n16481), .B(n16480), .CIN(n16479), .COUT(
        n16483), .SUM(n16488) );
  sky130_fd_sc_hd__fa_1 U21412 ( .A(n16484), .B(n16483), .CIN(n16482), .COUT(
        n16501), .SUM(n16498) );
  sky130_fd_sc_hd__nor2_1 U21413 ( .A(n16497), .B(n16498), .Y(n16822) );
  sky130_fd_sc_hd__fa_1 U21414 ( .A(n16487), .B(n16486), .CIN(n16485), .COUT(
        n16495), .SUM(n16494) );
  sky130_fd_sc_hd__fa_1 U21415 ( .A(n16490), .B(n16489), .CIN(n16488), .COUT(
        n16497), .SUM(n16496) );
  sky130_fd_sc_hd__nor2_1 U21416 ( .A(n16495), .B(n16496), .Y(n19850) );
  sky130_fd_sc_hd__nor2_1 U21417 ( .A(n16822), .B(n19850), .Y(n16500) );
  sky130_fd_sc_hd__nand2_1 U21418 ( .A(n16826), .B(n16500), .Y(n16614) );
  sky130_fd_sc_hd__nor2_1 U21419 ( .A(n16531), .B(n16614), .Y(n19347) );
  sky130_fd_sc_hd__nand2_1 U21420 ( .A(n16492), .B(n16491), .Y(n19213) );
  sky130_fd_sc_hd__nand2_1 U21421 ( .A(n16494), .B(n16493), .Y(n19218) );
  sky130_fd_sc_hd__o21ai_1 U21422 ( .A1(n19213), .A2(n19217), .B1(n19218), .Y(
        n16825) );
  sky130_fd_sc_hd__nand2_1 U21423 ( .A(n16496), .B(n16495), .Y(n19851) );
  sky130_fd_sc_hd__nand2_1 U21424 ( .A(n16498), .B(n16497), .Y(n16823) );
  sky130_fd_sc_hd__o21ai_1 U21425 ( .A1(n19851), .A2(n16822), .B1(n16823), .Y(
        n16499) );
  sky130_fd_sc_hd__a21oi_1 U21426 ( .A1(n16825), .A2(n16500), .B1(n16499), .Y(
        n16615) );
  sky130_fd_sc_hd__nand2_1 U21427 ( .A(n16502), .B(n16501), .Y(n18874) );
  sky130_fd_sc_hd__nand2_1 U21428 ( .A(n16504), .B(n16503), .Y(n17077) );
  sky130_fd_sc_hd__nand2_1 U21430 ( .A(n16506), .B(n16505), .Y(n19127) );
  sky130_fd_sc_hd__nand2_1 U21431 ( .A(n16508), .B(n16507), .Y(n18996) );
  sky130_fd_sc_hd__a21oi_1 U21432 ( .A1(n16510), .A2(n18997), .B1(n16509), .Y(
        n16621) );
  sky130_fd_sc_hd__nand2_1 U21433 ( .A(n16512), .B(n16511), .Y(n19290) );
  sky130_fd_sc_hd__nand2_1 U21434 ( .A(n16514), .B(n16513), .Y(n19288) );
  sky130_fd_sc_hd__nand2_1 U21436 ( .A(n16516), .B(n16515), .Y(n19942) );
  sky130_fd_sc_hd__nand2_1 U21437 ( .A(n16518), .B(n16517), .Y(n16782) );
  sky130_fd_sc_hd__nand2_1 U21438 ( .A(n16520), .B(n16519), .Y(n18855) );
  sky130_fd_sc_hd__a21oi_1 U21439 ( .A1(n18852), .A2(n18856), .B1(n16521), .Y(
        n16522) );
  sky130_fd_sc_hd__a21oi_1 U21441 ( .A1(n16783), .A2(n16525), .B1(n16524), .Y(
        n16526) );
  sky130_fd_sc_hd__a21oi_1 U21443 ( .A1(n16618), .A2(n16529), .B1(n16528), .Y(
        n16530) );
  sky130_fd_sc_hd__a21oi_1 U21445 ( .A1(n19216), .A2(n19347), .B1(n19359), .Y(
        n19096) );
  sky130_fd_sc_hd__a22oi_1 U21446 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[30]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[14]), .Y(n16532) );
  sky130_fd_sc_hd__nand2_1 U21447 ( .A(n16546), .B(n16532), .Y(n19345) );
  sky130_fd_sc_hd__a222oi_1 U21448 ( .A1(n16549), .A2(n11170), .B1(n16548), 
        .B2(n11170), .C1(n16547), .C2(n11170), .Y(n16533) );
  sky130_fd_sc_hd__o21ai_1 U21449 ( .A1(n11169), .A2(n16551), .B1(n16533), .Y(
        n16534) );
  sky130_fd_sc_hd__xnor2_1 U21450 ( .A(j202_soc_core_j22_cpu_ml_bufa[29]), .B(
        n16534), .Y(n16544) );
  sky130_fd_sc_hd__a22oi_1 U21451 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[29]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[13]), .Y(n16535) );
  sky130_fd_sc_hd__nand2_1 U21452 ( .A(n16546), .B(n16535), .Y(n16542) );
  sky130_fd_sc_hd__a222oi_1 U21453 ( .A1(n19334), .A2(n11170), .B1(n19333), 
        .B2(j202_soc_core_j22_cpu_ml_bufb[15]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .Y(n16536) );
  sky130_fd_sc_hd__o21ai_1 U21454 ( .A1(n19336), .A2(n16537), .B1(n16536), .Y(
        n16538) );
  sky130_fd_sc_hd__xor2_1 U21455 ( .A(n16538), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16578) );
  sky130_fd_sc_hd__a222oi_1 U21456 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[15]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .Y(n16539) );
  sky130_fd_sc_hd__xor2_1 U21458 ( .A(n16541), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16569) );
  sky130_fd_sc_hd__fa_1 U21459 ( .A(n16544), .B(n16543), .CIN(n16542), .COUT(
        n16579), .SUM(n16568) );
  sky130_fd_sc_hd__a22oi_1 U21460 ( .A1(n20025), .A2(
        j202_soc_core_j22_cpu_ml_mach[28]), .B1(n16580), .B2(
        j202_soc_core_j22_cpu_ml_mach[12]), .Y(n16545) );
  sky130_fd_sc_hd__nand2_1 U21461 ( .A(n16546), .B(n16545), .Y(n16563) );
  sky130_fd_sc_hd__a222oi_1 U21462 ( .A1(n16549), .A2(n11170), .B1(n16548), 
        .B2(n11170), .C1(n16547), .C2(j202_soc_core_j22_cpu_ml_bufb[15]), .Y(
        n16550) );
  sky130_fd_sc_hd__o21ai_1 U21463 ( .A1(n16551), .A2(n16584), .B1(n16550), .Y(
        n16552) );
  sky130_fd_sc_hd__xor2_1 U21464 ( .A(n16552), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .X(n16561) );
  sky130_fd_sc_hd__nor2_1 U21465 ( .A(n16576), .B(n16577), .Y(n18967) );
  sky130_fd_sc_hd__fa_1 U21466 ( .A(n16555), .B(n16554), .CIN(n16553), .COUT(
        n16570), .SUM(n16519) );
  sky130_fd_sc_hd__a222oi_1 U21467 ( .A1(n19334), .A2(
        j202_soc_core_j22_cpu_ml_bufb[14]), .B1(n19333), .B2(
        j202_soc_core_j22_cpu_ml_bufb[13]), .C1(n19332), .C2(
        j202_soc_core_j22_cpu_ml_bufb[12]), .Y(n16556) );
  sky130_fd_sc_hd__o21ai_1 U21468 ( .A1(n19336), .A2(n16557), .B1(n16556), .Y(
        n16558) );
  sky130_fd_sc_hd__xor2_1 U21469 ( .A(n16558), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n16566) );
  sky130_fd_sc_hd__fa_1 U21470 ( .A(n16562), .B(n16560), .CIN(n16559), .COUT(
        n16565), .SUM(n16553) );
  sky130_fd_sc_hd__fa_1 U21471 ( .A(n16563), .B(n16562), .CIN(n16561), .COUT(
        n16567), .SUM(n16564) );
  sky130_fd_sc_hd__nor2_1 U21472 ( .A(n16570), .B(n16571), .Y(n19097) );
  sky130_fd_sc_hd__fa_1 U21473 ( .A(n16566), .B(n16565), .CIN(n16564), .COUT(
        n16572), .SUM(n16571) );
  sky130_fd_sc_hd__fa_1 U21474 ( .A(n16569), .B(n16568), .CIN(n16567), .COUT(
        n16577), .SUM(n16573) );
  sky130_fd_sc_hd__nand2_1 U21475 ( .A(n17028), .B(n19094), .Y(n18963) );
  sky130_fd_sc_hd__nor2_1 U21476 ( .A(n18967), .B(n18963), .Y(n19343) );
  sky130_fd_sc_hd__nand2_1 U21477 ( .A(n16571), .B(n16570), .Y(n19095) );
  sky130_fd_sc_hd__nand2_1 U21478 ( .A(n16573), .B(n16572), .Y(n19093) );
  sky130_fd_sc_hd__a21oi_1 U21479 ( .A1(n16575), .A2(n19094), .B1(n16574), .Y(
        n18964) );
  sky130_fd_sc_hd__nand2_1 U21480 ( .A(n16577), .B(n16576), .Y(n18968) );
  sky130_fd_sc_hd__a21oi_1 U21482 ( .A1(n19920), .A2(n19343), .B1(n19351), .Y(
        n16589) );
  sky130_fd_sc_hd__fa_1 U21483 ( .A(n19341), .B(n16579), .CIN(n16578), .COUT(
        n16586), .SUM(n16576) );
  sky130_fd_sc_hd__a21oi_1 U21484 ( .A1(j202_soc_core_j22_cpu_ml_mach[31]), 
        .A2(n20025), .B1(n16581), .Y(n19338) );
  sky130_fd_sc_hd__o21ai_1 U21485 ( .A1(n19623), .A2(n16582), .B1(n19338), .Y(
        n19342) );
  sky130_fd_sc_hd__a222oi_1 U21486 ( .A1(n19334), .A2(n11170), .B1(n19333), 
        .B2(n11170), .C1(n19332), .C2(j202_soc_core_j22_cpu_ml_bufb[15]), .Y(
        n16583) );
  sky130_fd_sc_hd__o21ai_1 U21487 ( .A1(n19336), .A2(n16584), .B1(n16583), .Y(
        n16585) );
  sky130_fd_sc_hd__xor2_1 U21488 ( .A(n16585), .B(
        j202_soc_core_j22_cpu_ml_bufa[32]), .X(n19340) );
  sky130_fd_sc_hd__nand2_1 U21489 ( .A(n16587), .B(n16586), .Y(n19348) );
  sky130_fd_sc_hd__nand2_1 U21490 ( .A(n19350), .B(n19348), .Y(n16588) );
  sky130_fd_sc_hd__xor2_1 U21491 ( .A(n16589), .B(n16588), .X(n21695) );
  sky130_fd_sc_hd__nand3_1 U21492 ( .A(n16593), .B(n16592), .C(n22246), .Y(
        n16598) );
  sky130_fd_sc_hd__o31ai_1 U21493 ( .A1(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .A2(n16597), .A3(n16596), 
        .B1(n16595), .Y(n16607) );
  sky130_fd_sc_hd__nand2_1 U21494 ( .A(n20005), .B(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[3]), .Y(n21663) );
  sky130_fd_sc_hd__nand2_1 U21495 ( .A(n21695), .B(n20030), .Y(n16603) );
  sky130_fd_sc_hd__nand2_1 U21496 ( .A(n19215), .B(n19213), .Y(n16601) );
  sky130_fd_sc_hd__xnor2_1 U21497 ( .A(n16601), .B(n19216), .Y(n21701) );
  sky130_fd_sc_hd__a22oi_1 U21498 ( .A1(j202_soc_core_j22_cpu_ml_mach[15]), 
        .A2(n20032), .B1(n21701), .B2(n20025), .Y(n16602) );
  sky130_fd_sc_hd__nand2_1 U21499 ( .A(n16603), .B(n16602), .Y(n22203) );
  sky130_fd_sc_hd__nand2_1 U21500 ( .A(n22203), .B(n22125), .Y(n16611) );
  sky130_fd_sc_hd__nand2_1 U21501 ( .A(n19223), .B(n16604), .Y(n16606) );
  sky130_fd_sc_hd__xnor2_1 U21502 ( .A(n16606), .B(n19224), .Y(n22227) );
  sky130_fd_sc_hd__nor2_1 U21503 ( .A(n16607), .B(n20030), .Y(n21795) );
  sky130_fd_sc_hd__nand2_1 U21504 ( .A(n22225), .B(
        j202_soc_core_j22_cpu_macop_MAC_[0]), .Y(n20014) );
  sky130_fd_sc_hd__nand2b_1 U21505 ( .A_N(n20007), .B(n22125), .Y(n19565) );
  sky130_fd_sc_hd__nand2_1 U21506 ( .A(n20014), .B(n19565), .Y(n19931) );
  sky130_fd_sc_hd__nand2_1 U21507 ( .A(n17099), .B(
        j202_soc_core_j22_cpu_macop_MAC_[0]), .Y(n20012) );
  sky130_fd_sc_hd__o22ai_1 U21508 ( .A1(n20043), .A2(n22229), .B1(n16608), 
        .B2(n20012), .Y(n16609) );
  sky130_fd_sc_hd__a21oi_1 U21509 ( .A1(n22227), .A2(n20016), .B1(n16609), .Y(
        n16610) );
  sky130_fd_sc_hd__nand2_1 U21510 ( .A(n16611), .B(n16610), .Y(n20640) );
  sky130_fd_sc_hd__nand3_1 U21511 ( .A(n23245), .B(
        j202_soc_core_j22_cpu_memop_MEM__0_), .C(
        j202_soc_core_j22_cpu_memop_MEM__2_), .Y(n21211) );
  sky130_fd_sc_hd__nand2_1 U21512 ( .A(n20640), .B(n20019), .Y(n16705) );
  sky130_fd_sc_hd__nand2_1 U21513 ( .A(n16613), .B(n19290), .Y(n16624) );
  sky130_fd_sc_hd__a21oi_1 U21514 ( .A1(n19216), .A2(n16617), .B1(n16616), .Y(
        n17079) );
  sky130_fd_sc_hd__a21oi_1 U21515 ( .A1(n18876), .A2(n16619), .B1(n16618), .Y(
        n18998) );
  sky130_fd_sc_hd__a21oi_1 U21516 ( .A1(n19129), .A2(n16623), .B1(n16622), .Y(
        n19291) );
  sky130_fd_sc_hd__xnor2_1 U21517 ( .A(n16624), .B(n16785), .Y(n21694) );
  sky130_fd_sc_hd__nand2_1 U21518 ( .A(n21694), .B(n20030), .Y(n16631) );
  sky130_fd_sc_hd__nand2_1 U21519 ( .A(n16626), .B(n19298), .Y(n16627) );
  sky130_fd_sc_hd__xor2_1 U21520 ( .A(n19299), .B(n16627), .X(n19376) );
  sky130_fd_sc_hd__o22ai_1 U21521 ( .A1(n20007), .A2(n22235), .B1(n16628), 
        .B2(n20005), .Y(n16629) );
  sky130_fd_sc_hd__a21oi_1 U21522 ( .A1(n19376), .A2(n20025), .B1(n16629), .Y(
        n16630) );
  sky130_fd_sc_hd__nand2_1 U21523 ( .A(n16631), .B(n16630), .Y(n22208) );
  sky130_fd_sc_hd__nand2_1 U21524 ( .A(n22208), .B(n22125), .Y(n16639) );
  sky130_fd_sc_hd__nand2_1 U21525 ( .A(n16633), .B(n16632), .Y(n16634) );
  sky130_fd_sc_hd__xnor2_1 U21526 ( .A(n16635), .B(n16634), .Y(n22233) );
  sky130_fd_sc_hd__o22ai_1 U21527 ( .A1(n20014), .A2(n22235), .B1(n16636), 
        .B2(n20012), .Y(n16637) );
  sky130_fd_sc_hd__a21oi_1 U21528 ( .A1(n22233), .A2(n20016), .B1(n16637), .Y(
        n16638) );
  sky130_fd_sc_hd__nand2_1 U21529 ( .A(n16639), .B(n16638), .Y(n19463) );
  sky130_fd_sc_hd__nand2_1 U21530 ( .A(n19463), .B(n21137), .Y(n16685) );
  sky130_fd_sc_hd__nand2b_1 U21531 ( .A_N(n22687), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n16642) );
  sky130_fd_sc_hd__a22oi_1 U21532 ( .A1(j202_soc_core_j22_cpu_exuop_EXU_[3]), 
        .A2(j202_soc_core_j22_cpu_exuop_EXU_[0]), .B1(n22697), .B2(
        j202_soc_core_j22_cpu_exuop_EXU_[4]), .Y(n16641) );
  sky130_fd_sc_hd__nand2_1 U21533 ( .A(n22790), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[5]), .Y(n16640) );
  sky130_fd_sc_hd__nand2_1 U21534 ( .A(n22510), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[5]), .Y(n21011) );
  sky130_fd_sc_hd__nand2_1 U21535 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[1]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[0]), .Y(n22693) );
  sky130_fd_sc_hd__nand3_1 U21536 ( .A(n22689), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .C(n22670), .Y(n20839) );
  sky130_fd_sc_hd__nand2_1 U21537 ( .A(n20839), .B(n22509), .Y(n21063) );
  sky130_fd_sc_hd__nand2_1 U21538 ( .A(n21139), .B(n21063), .Y(n21027) );
  sky130_fd_sc_hd__nor2_1 U21539 ( .A(j202_soc_core_j22_cpu_ma_M_address[0]), 
        .B(n16643), .Y(n16860) );
  sky130_fd_sc_hd__clkinv_1 U21540 ( .A(n16860), .Y(n16859) );
  sky130_fd_sc_hd__nand2_1 U21541 ( .A(n22542), .B(n16650), .Y(n16645) );
  sky130_fd_sc_hd__nand2b_1 U21542 ( .A_N(n25388), .B(
        j202_soc_core_j22_cpu_ma_M_address[1]), .Y(n16644) );
  sky130_fd_sc_hd__nand2_1 U21543 ( .A(n16645), .B(n16644), .Y(n20353) );
  sky130_fd_sc_hd__nand3_1 U21544 ( .A(j202_soc_core_j22_cpu_ma_M_address[0]), 
        .B(n16650), .C(j202_soc_core_j22_cpu_ma_M_MEM[1]), .Y(n16861) );
  sky130_fd_sc_hd__nand4_1 U21545 ( .A(j202_soc_core_j22_cpu_ma_M_MEM[1]), .B(
        j202_soc_core_j22_cpu_ma_M_address[1]), .C(
        j202_soc_core_j22_cpu_ma_M_address[0]), .D(n25247), .Y(n16646) );
  sky130_fd_sc_hd__nand2_1 U21546 ( .A(n20352), .B(
        j202_soc_core_j22_cpu_ma_M_address[1]), .Y(n16649) );
  sky130_fd_sc_hd__nand2_1 U21547 ( .A(n22551), .B(n16649), .Y(n20706) );
  sky130_fd_sc_hd__nand2_1 U21548 ( .A(n16650), .B(n20352), .Y(n20616) );
  sky130_fd_sc_hd__a22oi_1 U21549 ( .A1(n25247), .A2(n20706), .B1(n22531), 
        .B2(n20707), .Y(n22537) );
  sky130_fd_sc_hd__nand2_1 U21550 ( .A(n20708), .B(n22537), .Y(n22495) );
  sky130_fd_sc_hd__nand2_1 U21551 ( .A(n22715), .B(n22790), .Y(n16651) );
  sky130_fd_sc_hd__nand2_1 U21552 ( .A(n22670), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[3]), .Y(n22700) );
  sky130_fd_sc_hd__nor2_1 U21553 ( .A(n16651), .B(n22700), .Y(n20829) );
  sky130_fd_sc_hd__nand2_1 U21554 ( .A(n21139), .B(n20829), .Y(n21150) );
  sky130_fd_sc_hd__nor2_1 U21555 ( .A(n22691), .B(n20931), .Y(n21146) );
  sky130_fd_sc_hd__a21oi_1 U21556 ( .A1(n22704), .A2(n21089), .B1(n21146), .Y(
        n16655) );
  sky130_fd_sc_hd__nand2_1 U21557 ( .A(n22510), .B(n16652), .Y(n16653) );
  sky130_fd_sc_hd__nand2_1 U21558 ( .A(n22495), .B(n21170), .Y(n16654) );
  sky130_fd_sc_hd__o211ai_1 U21559 ( .A1(n21027), .A2(n22495), .B1(n16655), 
        .C1(n16654), .Y(n16678) );
  sky130_fd_sc_hd__nand3_1 U21561 ( .A(n22495), .B(n21063), .C(n16656), .Y(
        n16676) );
  sky130_fd_sc_hd__nor2_1 U21562 ( .A(n22711), .B(n22037), .Y(n20360) );
  sky130_fd_sc_hd__nand2_1 U21563 ( .A(n22185), .B(n22707), .Y(n19880) );
  sky130_fd_sc_hd__nand2_1 U21564 ( .A(n20360), .B(n16668), .Y(n19875) );
  sky130_fd_sc_hd__nor2_1 U21565 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[3]), 
        .B(n22715), .Y(n19172) );
  sky130_fd_sc_hd__nand2_1 U21566 ( .A(n21139), .B(n19172), .Y(n19028) );
  sky130_fd_sc_hd__nand2_1 U21567 ( .A(n19875), .B(n19028), .Y(n20711) );
  sky130_fd_sc_hd__nor2_1 U21568 ( .A(n21011), .B(n22185), .Y(n22592) );
  sky130_fd_sc_hd__nor2_1 U21569 ( .A(n22705), .B(n22176), .Y(n19152) );
  sky130_fd_sc_hd__nand2_1 U21570 ( .A(n19152), .B(n22179), .Y(n16662) );
  sky130_fd_sc_hd__a22oi_1 U21571 ( .A1(n20711), .A2(n21828), .B1(n21164), 
        .B2(n19173), .Y(n16675) );
  sky130_fd_sc_hd__nand2_1 U21572 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[5]), 
        .B(j202_soc_core_j22_cpu_exuop_EXU_[3]), .Y(n16658) );
  sky130_fd_sc_hd__nand2_1 U21573 ( .A(n22584), .B(n16657), .Y(n21018) );
  sky130_fd_sc_hd__nor2_1 U21574 ( .A(n22141), .B(n21019), .Y(n16659) );
  sky130_fd_sc_hd__nand2_1 U21575 ( .A(n20365), .B(n16659), .Y(n20364) );
  sky130_fd_sc_hd__nor2_1 U21576 ( .A(n20931), .B(n20364), .Y(n20716) );
  sky130_fd_sc_hd__nor2_1 U21577 ( .A(n16658), .B(n22584), .Y(n20649) );
  sky130_fd_sc_hd__nand2_1 U21578 ( .A(n20649), .B(n22487), .Y(n20371) );
  sky130_fd_sc_hd__nand2b_1 U21579 ( .A_N(n20371), .B(n21139), .Y(n20712) );
  sky130_fd_sc_hd__a2bb2oi_1 U21580 ( .B1(n23319), .B2(n20716), .A1_N(n22275), 
        .A2_N(n20712), .Y(n16674) );
  sky130_fd_sc_hd__nor2_1 U21581 ( .A(n16658), .B(n22487), .Y(n16661) );
  sky130_fd_sc_hd__nand2_1 U21582 ( .A(n20365), .B(n22581), .Y(n16660) );
  sky130_fd_sc_hd__nand2_1 U21583 ( .A(n16660), .B(n20370), .Y(n20524) );
  sky130_fd_sc_hd__o21a_1 U21584 ( .A1(n16661), .A2(n20524), .B1(n21139), .X(
        n19884) );
  sky130_fd_sc_hd__nand2b_1 U21585 ( .A_N(n16662), .B(n16668), .Y(n21163) );
  sky130_fd_sc_hd__nand2b_1 U21586 ( .A_N(n22711), .B(n22264), .Y(n16669) );
  sky130_fd_sc_hd__nand2_1 U21587 ( .A(n16669), .B(n22592), .Y(n21155) );
  sky130_fd_sc_hd__nand2_1 U21588 ( .A(n21139), .B(n16663), .Y(n21145) );
  sky130_fd_sc_hd__nand3_1 U21589 ( .A(n16664), .B(n22790), .C(
        j202_soc_core_j22_cpu_exuop_EXU_[2]), .Y(n17108) );
  sky130_fd_sc_hd__o21a_1 U21590 ( .A1(n21145), .A2(n22704), .B1(n21174), .X(
        n16667) );
  sky130_fd_sc_hd__xor2_1 U21591 ( .A(n22496), .B(n22704), .X(n22435) );
  sky130_fd_sc_hd__nor2_1 U21592 ( .A(n20835), .B(n20931), .Y(n21147) );
  sky130_fd_sc_hd__nand2_1 U21593 ( .A(n22435), .B(n21147), .Y(n16666) );
  sky130_fd_sc_hd__o211a_2 U21594 ( .A1(n22612), .A2(n21155), .B1(n16667), 
        .C1(n16666), .X(n16671) );
  sky130_fd_sc_hd__nor2_1 U21595 ( .A(n22646), .B(n19880), .Y(n21156) );
  sky130_fd_sc_hd__nand2_1 U21596 ( .A(n16669), .B(n16668), .Y(n21154) );
  sky130_fd_sc_hd__a2bb2oi_1 U21597 ( .B1(n21156), .B2(n22136), .A1_N(n22558), 
        .A2_N(n21154), .Y(n16670) );
  sky130_fd_sc_hd__o211ai_1 U21598 ( .A1(n22559), .A2(n21163), .B1(n16671), 
        .C1(n16670), .Y(n16672) );
  sky130_fd_sc_hd__a21oi_1 U21599 ( .A1(n19884), .A2(n22704), .B1(n16672), .Y(
        n16673) );
  sky130_fd_sc_hd__nand4_1 U21600 ( .A(n16676), .B(n16675), .C(n16674), .D(
        n16673), .Y(n16677) );
  sky130_fd_sc_hd__a21oi_1 U21601 ( .A1(n16678), .A2(n22496), .B1(n16677), .Y(
        n16684) );
  sky130_fd_sc_hd__nand2_1 U21602 ( .A(n16680), .B(n19724), .Y(n16681) );
  sky130_fd_sc_hd__xor2_1 U21603 ( .A(n19725), .B(n16681), .X(n22292) );
  sky130_fd_sc_hd__nand2_1 U21604 ( .A(n22292), .B(n21178), .Y(n16683) );
  sky130_fd_sc_hd__o21ai_0 U21605 ( .A1(j202_soc_core_j22_cpu_memop_MEM__2_), 
        .A2(n23240), .B1(n16686), .Y(n16688) );
  sky130_fd_sc_hd__nor2_1 U21606 ( .A(n23243), .B(n21220), .Y(n16687) );
  sky130_fd_sc_hd__nor2_1 U21607 ( .A(n16688), .B(n16687), .Y(n21237) );
  sky130_fd_sc_hd__nand2b_1 U21608 ( .A_N(n16689), .B(n23242), .Y(n21251) );
  sky130_fd_sc_hd__nand2_1 U21609 ( .A(n16690), .B(n21251), .Y(n21241) );
  sky130_fd_sc_hd__nand2_1 U21610 ( .A(n22286), .B(n19905), .Y(n19464) );
  sky130_fd_sc_hd__o22ai_1 U21611 ( .A1(n16692), .A2(n19973), .B1(n16691), 
        .B2(n19971), .Y(n16696) );
  sky130_fd_sc_hd__o22ai_1 U21612 ( .A1(n16694), .A2(n19977), .B1(n16693), 
        .B2(n19975), .Y(n16695) );
  sky130_fd_sc_hd__nor2_1 U21613 ( .A(n16696), .B(n16695), .Y(n16701) );
  sky130_fd_sc_hd__a2bb2oi_1 U21614 ( .B1(j202_soc_core_j22_cpu_rf_vbr[7]), 
        .B2(n19985), .A1_N(n16697), .A2_N(n19986), .Y(n16700) );
  sky130_fd_sc_hd__nand2_1 U21615 ( .A(n19842), .B(
        j202_soc_core_j22_cpu_rf_gpr[7]), .Y(n16699) );
  sky130_fd_sc_hd__nand2_1 U21616 ( .A(n19843), .B(
        j202_soc_core_j22_cpu_rf_tmp[7]), .Y(n16698) );
  sky130_fd_sc_hd__nand4_1 U21617 ( .A(n16701), .B(n16700), .C(n16699), .D(
        n16698), .Y(n16702) );
  sky130_fd_sc_hd__a21oi_1 U21618 ( .A1(n16703), .A2(n19969), .B1(n16702), .Y(
        n19466) );
  sky130_fd_sc_hd__nor2_1 U21619 ( .A(j202_soc_core_j22_cpu_memop_MEM__0_), 
        .B(n19917), .Y(n19285) );
  sky130_fd_sc_hd__nand2b_1 U21620 ( .A_N(n19466), .B(n19285), .Y(n16704) );
  sky130_fd_sc_hd__o211ai_1 U21621 ( .A1(n19317), .A2(n19649), .B1(n16705), 
        .C1(n19651), .Y(n25345) );
  sky130_fd_sc_hd__nand2_1 U21622 ( .A(n25731), .B(
        j202_soc_core_qspi_wb_wdat[15]), .Y(n24432) );
  sky130_fd_sc_hd__nand2_1 U21623 ( .A(n22292), .B(n19729), .Y(n16711) );
  sky130_fd_sc_hd__ha_1 U21624 ( .A(j202_soc_core_j22_cpu_pc[7]), .B(n16706), 
        .COUT(n19730), .SUM(n22289) );
  sky130_fd_sc_hd__nand2_1 U21625 ( .A(n19661), .B(n22289), .Y(n16708) );
  sky130_fd_sc_hd__nand2_1 U21626 ( .A(n19736), .B(n22704), .Y(n16707) );
  sky130_fd_sc_hd__o211ai_1 U21627 ( .A1(n22645), .A2(n19731), .B1(n16708), 
        .C1(n16707), .Y(n16709) );
  sky130_fd_sc_hd__a21oi_1 U21628 ( .A1(n25247), .A2(n19737), .B1(n16709), .Y(
        n16710) );
  sky130_fd_sc_hd__nand2_1 U21629 ( .A(n16711), .B(n16710), .Y(n25338) );
  sky130_fd_sc_hd__nand2_1 U21630 ( .A(n17868), .B(n17534), .Y(n18349) );
  sky130_fd_sc_hd__nor2_1 U21631 ( .A(n18390), .B(n18349), .Y(n18400) );
  sky130_fd_sc_hd__nand3_1 U21632 ( .A(n17653), .B(n17779), .C(n17675), .Y(
        n18395) );
  sky130_fd_sc_hd__nor4_1 U21633 ( .A(n17600), .B(n18418), .C(n17611), .D(
        n18395), .Y(n16712) );
  sky130_fd_sc_hd__a31oi_1 U21634 ( .A1(n18400), .A2(n16712), .A3(n17923), 
        .B1(n18439), .Y(n16719) );
  sky130_fd_sc_hd__nand2_1 U21635 ( .A(n16737), .B(n17756), .Y(n18444) );
  sky130_fd_sc_hd__nor2_1 U21636 ( .A(n17784), .B(n18444), .Y(n17846) );
  sky130_fd_sc_hd__nand2_1 U21637 ( .A(n17868), .B(n17548), .Y(n17597) );
  sky130_fd_sc_hd__nor4_1 U21638 ( .A(n18392), .B(n17752), .C(n17619), .D(
        n17597), .Y(n16713) );
  sky130_fd_sc_hd__a31oi_1 U21639 ( .A1(n17846), .A2(n16714), .A3(n16713), 
        .B1(n18445), .Y(n16718) );
  sky130_fd_sc_hd__nand2_1 U21640 ( .A(n16737), .B(n17534), .Y(n18391) );
  sky130_fd_sc_hd__nor2_1 U21641 ( .A(n17865), .B(n17847), .Y(n17907) );
  sky130_fd_sc_hd__nor2_1 U21642 ( .A(n17842), .B(n16769), .Y(n17523) );
  sky130_fd_sc_hd__nand2_1 U21643 ( .A(n17907), .B(n17523), .Y(n18442) );
  sky130_fd_sc_hd__nor4b_1 U21644 ( .D_N(n16739), .A(n17867), .B(n18391), .C(
        n18442), .Y(n17595) );
  sky130_fd_sc_hd__nor2_1 U21645 ( .A(n17944), .B(n18444), .Y(n17770) );
  sky130_fd_sc_hd__nand2_1 U21646 ( .A(n17863), .B(n18347), .Y(n17549) );
  sky130_fd_sc_hd__nor2_1 U21647 ( .A(n18397), .B(n17549), .Y(n18388) );
  sky130_fd_sc_hd__nand2_1 U21648 ( .A(n17779), .B(n17676), .Y(n17472) );
  sky130_fd_sc_hd__nor2_1 U21649 ( .A(n17472), .B(n17670), .Y(n17657) );
  sky130_fd_sc_hd__nand4_1 U21650 ( .A(n17770), .B(n18388), .C(n17657), .D(
        n17875), .Y(n16715) );
  sky130_fd_sc_hd__nor3_1 U21651 ( .A(n17945), .B(n17915), .C(n16715), .Y(
        n16716) );
  sky130_fd_sc_hd__o22ai_1 U21652 ( .A1(n17595), .A2(n18423), .B1(n16716), 
        .B2(n18437), .Y(n16717) );
  sky130_fd_sc_hd__nor3_1 U21653 ( .A(n16719), .B(n16718), .C(n16717), .Y(
        n16735) );
  sky130_fd_sc_hd__a22o_1 U21654 ( .A1(n18367), .A2(
        j202_soc_core_memory0_ram_dout0[10]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[74]), .X(n16720) );
  sky130_fd_sc_hd__a21oi_1 U21655 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[106]), .B1(n16720), .Y(n16722) );
  sky130_fd_sc_hd__a22oi_1 U21656 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[170]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[138]), .Y(n16721) );
  sky130_fd_sc_hd__a21oi_1 U21657 ( .A1(n16722), .A2(n16721), .B1(n18736), .Y(
        n16733) );
  sky130_fd_sc_hd__a22oi_1 U21658 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[266]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[42]), .Y(n16731) );
  sky130_fd_sc_hd__a22o_1 U21659 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[298]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[330]), .X(n16723) );
  sky130_fd_sc_hd__a21oi_1 U21660 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[362]), .B1(n16723), .Y(n16730) );
  sky130_fd_sc_hd__nand2_1 U21661 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[234]), .Y(n16727) );
  sky130_fd_sc_hd__a21oi_1 U21662 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[458]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n16726) );
  sky130_fd_sc_hd__nand2_1 U21663 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[394]), .Y(n16725) );
  sky130_fd_sc_hd__nand2_1 U21664 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[426]), .Y(n16724) );
  sky130_fd_sc_hd__nand4_1 U21665 ( .A(n16727), .B(n16726), .C(n16725), .D(
        n16724), .Y(n16728) );
  sky130_fd_sc_hd__a21oi_1 U21666 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[202]), .B1(n16728), .Y(n16729) );
  sky130_fd_sc_hd__nand3_1 U21667 ( .A(n16731), .B(n16730), .C(n16729), .Y(
        n16732) );
  sky130_fd_sc_hd__o22ai_1 U21668 ( .A1(j202_soc_core_memory0_ram_dout0[490]), 
        .A2(n18758), .B1(n16733), .B2(n16732), .Y(n16734) );
  sky130_fd_sc_hd__o22ai_1 U21669 ( .A1(n16735), .A2(n18666), .B1(n18761), 
        .B2(n16734), .Y(n16781) );
  sky130_fd_sc_hd__nand2_1 U21670 ( .A(n16764), .B(n16736), .Y(n18386) );
  sky130_fd_sc_hd__nor2_1 U21671 ( .A(n17795), .B(n17611), .Y(n17480) );
  sky130_fd_sc_hd__nand2_1 U21672 ( .A(n17480), .B(n18399), .Y(n18443) );
  sky130_fd_sc_hd__nand2_1 U21673 ( .A(n17923), .B(n16737), .Y(n16738) );
  sky130_fd_sc_hd__nor4_1 U21674 ( .A(n17865), .B(n18386), .C(n18443), .D(
        n16738), .Y(n16752) );
  sky130_fd_sc_hd__nand3_1 U21676 ( .A(n17478), .B(n17911), .C(n17771), .Y(
        n18441) );
  sky130_fd_sc_hd__nor2_1 U21677 ( .A(n17915), .B(n18441), .Y(n17851) );
  sky130_fd_sc_hd__nand2_1 U21678 ( .A(n17770), .B(n17875), .Y(n16742) );
  sky130_fd_sc_hd__nor4_1 U21679 ( .A(n18397), .B(n17472), .C(n17669), .D(
        n16742), .Y(n16743) );
  sky130_fd_sc_hd__a21oi_1 U21680 ( .A1(n17851), .A2(n16743), .B1(n18439), .Y(
        n16749) );
  sky130_fd_sc_hd__nand2_1 U21681 ( .A(n17596), .B(n18345), .Y(n17940) );
  sky130_fd_sc_hd__nand2_1 U21682 ( .A(n17869), .B(n17771), .Y(n17677) );
  sky130_fd_sc_hd__nor3_1 U21683 ( .A(n17910), .B(n17746), .C(n16767), .Y(
        n16759) );
  sky130_fd_sc_hd__a211oi_1 U21684 ( .A1(n17469), .A2(n16744), .B1(n17677), 
        .C1(n17843), .Y(n16745) );
  sky130_fd_sc_hd__a31oi_1 U21685 ( .A1(n16747), .A2(n16746), .A3(n16745), 
        .B1(n18445), .Y(n16748) );
  sky130_fd_sc_hd__a211oi_1 U21686 ( .A1(n17543), .A2(n16750), .B1(n16749), 
        .C1(n16748), .Y(n16751) );
  sky130_fd_sc_hd__nand2_1 U21688 ( .A(n18629), .B(
        j202_soc_core_bldc_core_00_pwm_period[10]), .Y(n16756) );
  sky130_fd_sc_hd__a22oi_1 U21689 ( .A1(n18724), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[106]), .B1(n18725), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[10]), .Y(n16755) );
  sky130_fd_sc_hd__nand2_1 U21690 ( .A(n18726), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[42]), .Y(n16754) );
  sky130_fd_sc_hd__nand2_1 U21691 ( .A(n18727), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[74]), .Y(n16753) );
  sky130_fd_sc_hd__nand4_1 U21692 ( .A(n16756), .B(n16755), .C(n16754), .D(
        n16753), .Y(n16757) );
  sky130_fd_sc_hd__a21oi_1 U21693 ( .A1(n16758), .A2(n18605), .B1(n16757), .Y(
        n16780) );
  sky130_fd_sc_hd__nand3_1 U21694 ( .A(n18400), .B(n18519), .C(n18446), .Y(
        n17660) );
  sky130_fd_sc_hd__nor2_1 U21695 ( .A(n17945), .B(n18354), .Y(n17793) );
  sky130_fd_sc_hd__a21oi_1 U21696 ( .A1(n18428), .A2(n17793), .B1(n18423), .Y(
        n16763) );
  sky130_fd_sc_hd__nand2_1 U21697 ( .A(n16759), .B(n17618), .Y(n17905) );
  sky130_fd_sc_hd__nor4_1 U21698 ( .A(n17619), .B(n17420), .C(n16769), .D(
        n17905), .Y(n16761) );
  sky130_fd_sc_hd__nand2_1 U21699 ( .A(n17793), .B(n16759), .Y(n17926) );
  sky130_fd_sc_hd__nand2_1 U21700 ( .A(n17678), .B(n17548), .Y(n17852) );
  sky130_fd_sc_hd__nand2b_1 U21701 ( .A_N(n17852), .B(n18388), .Y(n17917) );
  sky130_fd_sc_hd__nor3_1 U21702 ( .A(n17784), .B(n17926), .C(n17917), .Y(
        n16760) );
  sky130_fd_sc_hd__o22ai_1 U21703 ( .A1(n16761), .A2(n18445), .B1(n16760), 
        .B2(n18439), .Y(n16762) );
  sky130_fd_sc_hd__a211oi_1 U21704 ( .A1(n17543), .A2(n17660), .B1(n16763), 
        .C1(n16762), .Y(n16778) );
  sky130_fd_sc_hd__nand4_1 U21705 ( .A(n16765), .B(n16764), .C(n18345), .D(
        n18446), .Y(n17902) );
  sky130_fd_sc_hd__nor2_1 U21706 ( .A(n17910), .B(n17752), .Y(n17481) );
  sky130_fd_sc_hd__a31oi_1 U21707 ( .A1(n18388), .A2(n16766), .A3(n17674), 
        .B1(n18445), .Y(n16776) );
  sky130_fd_sc_hd__nor2_1 U21708 ( .A(n17915), .B(n16767), .Y(n18424) );
  sky130_fd_sc_hd__nand2_1 U21709 ( .A(n17771), .B(n18341), .Y(n17605) );
  sky130_fd_sc_hd__nor4_1 U21710 ( .A(n17624), .B(n18354), .C(n18444), .D(
        n17605), .Y(n16768) );
  sky130_fd_sc_hd__a21oi_1 U21711 ( .A1(n18424), .A2(n16768), .B1(n18437), .Y(
        n16775) );
  sky130_fd_sc_hd__nor2_1 U21712 ( .A(n17746), .B(n16769), .Y(n18389) );
  sky130_fd_sc_hd__nor3_1 U21713 ( .A(n17945), .B(n17910), .C(n17727), .Y(
        n17769) );
  sky130_fd_sc_hd__nor3_1 U21714 ( .A(n17593), .B(n17592), .C(n17942), .Y(
        n16770) );
  sky130_fd_sc_hd__a31oi_1 U21715 ( .A1(n18389), .A2(n17769), .A3(n16770), 
        .B1(n18423), .Y(n16774) );
  sky130_fd_sc_hd__nand3_1 U21716 ( .A(n17869), .B(n17618), .C(n17676), .Y(
        n18353) );
  sky130_fd_sc_hd__nor2_1 U21717 ( .A(n18354), .B(n18353), .Y(n16772) );
  sky130_fd_sc_hd__nor2_1 U21718 ( .A(n17746), .B(n17727), .Y(n17761) );
  sky130_fd_sc_hd__nor2_1 U21719 ( .A(n18392), .B(n17619), .Y(n16771) );
  sky130_fd_sc_hd__a31oi_1 U21720 ( .A1(n16772), .A2(n17761), .A3(n16771), 
        .B1(n18439), .Y(n16773) );
  sky130_fd_sc_hd__nor4_1 U21721 ( .A(n16776), .B(n16775), .C(n16774), .D(
        n16773), .Y(n16777) );
  sky130_fd_sc_hd__o22a_1 U21722 ( .A1(n16778), .A2(n18552), .B1(n16777), .B2(
        n18720), .X(n16779) );
  sky130_fd_sc_hd__nand3b_1 U21723 ( .A_N(n16781), .B(n16780), .C(n16779), .Y(
        n25314) );
  sky130_fd_sc_hd__nand2_1 U21724 ( .A(n18853), .B(n16782), .Y(n16786) );
  sky130_fd_sc_hd__a21oi_1 U21725 ( .A1(n16785), .A2(n16784), .B1(n16783), .Y(
        n19945) );
  sky130_fd_sc_hd__xnor2_1 U21727 ( .A(n16786), .B(n18854), .Y(n21692) );
  sky130_fd_sc_hd__nand2_1 U21728 ( .A(n21692), .B(n20030), .Y(n16801) );
  sky130_fd_sc_hd__a21oi_1 U21730 ( .A1(n19951), .A2(n19950), .B1(n16792), .Y(
        n16797) );
  sky130_fd_sc_hd__nand2_1 U21731 ( .A(n16795), .B(n16794), .Y(n16796) );
  sky130_fd_sc_hd__xor2_1 U21732 ( .A(n16797), .B(n16796), .X(n19566) );
  sky130_fd_sc_hd__o22ai_1 U21733 ( .A1(n20007), .A2(n21799), .B1(n16798), 
        .B2(n20005), .Y(n16799) );
  sky130_fd_sc_hd__a21oi_1 U21734 ( .A1(n19566), .A2(n20025), .B1(n16799), .Y(
        n16800) );
  sky130_fd_sc_hd__nand2_1 U21735 ( .A(n16801), .B(n16800), .Y(n21793) );
  sky130_fd_sc_hd__nand2_1 U21736 ( .A(n21793), .B(n22125), .Y(n16811) );
  sky130_fd_sc_hd__nand2_1 U21737 ( .A(n16804), .B(n16803), .Y(n16807) );
  sky130_fd_sc_hd__xnor2_1 U21739 ( .A(n16807), .B(n16806), .Y(n21797) );
  sky130_fd_sc_hd__o22ai_1 U21740 ( .A1(n20014), .A2(n21799), .B1(n16808), 
        .B2(n20012), .Y(n16809) );
  sky130_fd_sc_hd__a21oi_1 U21741 ( .A1(n21797), .A2(n20016), .B1(n16809), .Y(
        n16810) );
  sky130_fd_sc_hd__nand2_1 U21742 ( .A(n16811), .B(n16810), .Y(n20735) );
  sky130_fd_sc_hd__nand2_1 U21743 ( .A(n20735), .B(n20019), .Y(n16888) );
  sky130_fd_sc_hd__a22oi_1 U21744 ( .A1(n16812), .A2(
        j202_soc_core_j22_cpu_pc[2]), .B1(n19985), .B2(
        j202_soc_core_j22_cpu_rf_vbr[2]), .Y(n16819) );
  sky130_fd_sc_hd__o22a_1 U21745 ( .A1(n16814), .A2(n19971), .B1(n16813), .B2(
        n19975), .X(n16818) );
  sky130_fd_sc_hd__a2bb2oi_1 U21746 ( .B1(j202_soc_core_j22_cpu_rf_tmp[2]), 
        .B2(n19843), .A1_N(n16815), .A2_N(n19986), .Y(n16817) );
  sky130_fd_sc_hd__nand2_1 U21747 ( .A(n19842), .B(
        j202_soc_core_j22_cpu_rf_gpr[2]), .Y(n16816) );
  sky130_fd_sc_hd__nand4_1 U21748 ( .A(n16819), .B(n16818), .C(n16817), .D(
        n16816), .Y(n16820) );
  sky130_fd_sc_hd__a21oi_1 U21749 ( .A1(n16821), .A2(n19969), .B1(n16820), .Y(
        n19506) );
  sky130_fd_sc_hd__nand2_1 U21750 ( .A(n16824), .B(n16823), .Y(n16828) );
  sky130_fd_sc_hd__a21oi_1 U21751 ( .A1(n19216), .A2(n16826), .B1(n16825), .Y(
        n19854) );
  sky130_fd_sc_hd__xnor2_1 U21753 ( .A(n16828), .B(n16827), .Y(n21703) );
  sky130_fd_sc_hd__nand2_1 U21754 ( .A(n21703), .B(n20030), .Y(n16838) );
  sky130_fd_sc_hd__nand2_1 U21755 ( .A(n16831), .B(n16830), .Y(n16834) );
  sky130_fd_sc_hd__xnor2_1 U21757 ( .A(n16834), .B(n16833), .Y(n19451) );
  sky130_fd_sc_hd__o22ai_1 U21758 ( .A1(n20007), .A2(n22238), .B1(n16835), 
        .B2(n20005), .Y(n16836) );
  sky130_fd_sc_hd__a21oi_1 U21759 ( .A1(n19451), .A2(n20025), .B1(n16836), .Y(
        n16837) );
  sky130_fd_sc_hd__nand2_1 U21760 ( .A(n16838), .B(n16837), .Y(n22210) );
  sky130_fd_sc_hd__nand2_1 U21761 ( .A(n22210), .B(n22125), .Y(n16846) );
  sky130_fd_sc_hd__nand2_1 U21762 ( .A(n16840), .B(n16839), .Y(n16842) );
  sky130_fd_sc_hd__xnor2_1 U21763 ( .A(n16842), .B(n16841), .Y(n22236) );
  sky130_fd_sc_hd__o22ai_1 U21764 ( .A1(n20014), .A2(n22238), .B1(n16843), 
        .B2(n20012), .Y(n16844) );
  sky130_fd_sc_hd__a21oi_1 U21765 ( .A1(n22236), .A2(n20016), .B1(n16844), .Y(
        n16845) );
  sky130_fd_sc_hd__nand2_1 U21766 ( .A(n16846), .B(n16845), .Y(n19503) );
  sky130_fd_sc_hd__nand2_1 U21767 ( .A(n19503), .B(n21137), .Y(n16874) );
  sky130_fd_sc_hd__nand2_1 U21768 ( .A(n22262), .B(n21178), .Y(n16869) );
  sky130_fd_sc_hd__nand2_1 U21769 ( .A(n20711), .B(n21775), .Y(n16848) );
  sky130_fd_sc_hd__a2bb2oi_1 U21770 ( .B1(n23304), .B2(n20716), .A1_N(n21807), 
        .A2_N(n20712), .Y(n16847) );
  sky130_fd_sc_hd__o211ai_1 U21771 ( .A1(n22647), .A2(n21163), .B1(n16848), 
        .C1(n16847), .Y(n16856) );
  sky130_fd_sc_hd__o22ai_1 U21772 ( .A1(n20805), .A2(n21155), .B1(n22488), 
        .B2(n21154), .Y(n16849) );
  sky130_fd_sc_hd__a21oi_1 U21773 ( .A1(n21164), .A2(n22584), .B1(n16849), .Y(
        n16854) );
  sky130_fd_sc_hd__nand2_1 U21774 ( .A(n22264), .B(n22487), .Y(n22430) );
  sky130_fd_sc_hd__nand2_1 U21775 ( .A(n22181), .B(n21019), .Y(n22620) );
  sky130_fd_sc_hd__o22ai_1 U21776 ( .A1(n22181), .A2(n21145), .B1(n21150), 
        .B2(n22620), .Y(n16850) );
  sky130_fd_sc_hd__a31oi_1 U21777 ( .A1(n21147), .A2(n22430), .A3(n22620), 
        .B1(n16850), .Y(n16853) );
  sky130_fd_sc_hd__nand2_1 U21778 ( .A(n19884), .B(n22181), .Y(n16852) );
  sky130_fd_sc_hd__nand2_1 U21779 ( .A(n21156), .B(n20935), .Y(n16851) );
  sky130_fd_sc_hd__nand4_1 U21780 ( .A(n16854), .B(n16853), .C(n16852), .D(
        n16851), .Y(n16855) );
  sky130_fd_sc_hd__nor2_1 U21781 ( .A(n16856), .B(n16855), .Y(n16868) );
  sky130_fd_sc_hd__nand2_1 U21782 ( .A(j202_soc_core_j22_cpu_ma_M_address[0]), 
        .B(j202_soc_core_j22_cpu_ma_M_address[1]), .Y(n16857) );
  sky130_fd_sc_hd__nand2_1 U21783 ( .A(n25246), .B(n19895), .Y(n16864) );
  sky130_fd_sc_hd__nor2_1 U21784 ( .A(n16859), .B(
        j202_soc_core_j22_cpu_ma_M_address[1]), .Y(n19239) );
  sky130_fd_sc_hd__a22oi_1 U21785 ( .A1(n19239), .A2(n20825), .B1(n25314), 
        .B2(n19889), .Y(n16863) );
  sky130_fd_sc_hd__nand2_1 U21786 ( .A(n20616), .B(n16861), .Y(n19893) );
  sky130_fd_sc_hd__nand2_1 U21787 ( .A(n22523), .B(n19893), .Y(n16862) );
  sky130_fd_sc_hd__nand2_1 U21788 ( .A(n21019), .B(n21170), .Y(n16865) );
  sky130_fd_sc_hd__o211ai_1 U21789 ( .A1(n21027), .A2(n21019), .B1(n16865), 
        .C1(n21174), .Y(n16866) );
  sky130_fd_sc_hd__nand2_1 U21790 ( .A(n22547), .B(n16866), .Y(n16867) );
  sky130_fd_sc_hd__and3_1 U21791 ( .A(n16869), .B(n16868), .C(n16867), .X(
        n16873) );
  sky130_fd_sc_hd__nand2_1 U21792 ( .A(n20839), .B(n22691), .Y(n16870) );
  sky130_fd_sc_hd__nand2_1 U21794 ( .A(n16871), .B(n21019), .Y(n16872) );
  sky130_fd_sc_hd__nand2_1 U21795 ( .A(n22258), .B(n19905), .Y(n19504) );
  sky130_fd_sc_hd__o21a_1 U21796 ( .A1(n19506), .A2(n19967), .B1(n19504), .X(
        n19584) );
  sky130_fd_sc_hd__nand2_1 U21797 ( .A(n16875), .B(n19969), .Y(n16886) );
  sky130_fd_sc_hd__o22ai_1 U21798 ( .A1(n16877), .A2(n19977), .B1(n19971), 
        .B2(n16876), .Y(n16878) );
  sky130_fd_sc_hd__a21oi_1 U21799 ( .A1(n19842), .A2(
        j202_soc_core_j22_cpu_rf_gpr[10]), .B1(n16878), .Y(n16885) );
  sky130_fd_sc_hd__o22ai_1 U21800 ( .A1(n16880), .A2(n19975), .B1(n16879), 
        .B2(n19986), .Y(n16883) );
  sky130_fd_sc_hd__o2bb2ai_1 U21801 ( .B1(n16881), .B2(n19981), .A1_N(
        j202_soc_core_j22_cpu_rf_vbr[10]), .A2_N(n19985), .Y(n16882) );
  sky130_fd_sc_hd__nor2_1 U21802 ( .A(n16883), .B(n16882), .Y(n16884) );
  sky130_fd_sc_hd__nand3_1 U21803 ( .A(n16886), .B(n16885), .C(n16884), .Y(
        n19582) );
  sky130_fd_sc_hd__nand2_1 U21804 ( .A(n19582), .B(n20020), .Y(n16887) );
  sky130_fd_sc_hd__nand3_1 U21805 ( .A(n16888), .B(n19584), .C(n16887), .Y(
        n25342) );
  sky130_fd_sc_hd__nand2_1 U21806 ( .A(n25731), .B(
        j202_soc_core_qspi_wb_wdat[10]), .Y(n24422) );
  sky130_fd_sc_hd__nor2_1 U21807 ( .A(n16996), .B(n18543), .Y(n18320) );
  sky130_fd_sc_hd__a31oi_1 U21808 ( .A1(n18264), .A2(n16907), .A3(n18320), 
        .B1(n18779), .Y(n16894) );
  sky130_fd_sc_hd__a31oi_1 U21809 ( .A1(n16889), .A2(n18270), .A3(n18680), 
        .B1(n18771), .Y(n16893) );
  sky130_fd_sc_hd__nor2_1 U21810 ( .A(n18645), .B(n17508), .Y(n18318) );
  sky130_fd_sc_hd__a31oi_1 U21811 ( .A1(n16890), .A2(n18318), .A3(n18593), 
        .B1(n18783), .Y(n16892) );
  sky130_fd_sc_hd__nor4_1 U21812 ( .A(n16894), .B(n16893), .C(n16892), .D(
        n16891), .Y(n16900) );
  sky130_fd_sc_hd__or4_1 U21813 ( .A(n16926), .B(n18248), .C(n18703), .D(
        n18644), .X(n16895) );
  sky130_fd_sc_hd__o31ai_1 U21815 ( .A1(n18527), .A2(n16898), .A3(n16897), 
        .B1(n18651), .Y(n16899) );
  sky130_fd_sc_hd__a31oi_1 U21816 ( .A1(n16900), .A2(n18302), .A3(n16899), 
        .B1(n18722), .Y(n16941) );
  sky130_fd_sc_hd__nand2_1 U21817 ( .A(n18593), .B(n16901), .Y(n18708) );
  sky130_fd_sc_hd__nand3_1 U21818 ( .A(n18662), .B(n18522), .C(n18569), .Y(
        n18316) );
  sky130_fd_sc_hd__nor2_1 U21819 ( .A(n18708), .B(n18316), .Y(n18258) );
  sky130_fd_sc_hd__nor4b_1 U21820 ( .D_N(n18270), .A(n18702), .B(n18641), .C(
        n16908), .Y(n16902) );
  sky130_fd_sc_hd__a21oi_1 U21821 ( .A1(n18258), .A2(n16902), .B1(n18771), .Y(
        n16913) );
  sky130_fd_sc_hd__nor3_1 U21822 ( .A(n18687), .B(n18638), .C(n18511), .Y(
        n18297) );
  sky130_fd_sc_hd__nor2_1 U21823 ( .A(n18709), .B(n18512), .Y(n18542) );
  sky130_fd_sc_hd__nand2_1 U21824 ( .A(n18593), .B(n18592), .Y(n16903) );
  sky130_fd_sc_hd__nor3b_1 U21825 ( .C_N(n16915), .A(n16908), .B(n16903), .Y(
        n16904) );
  sky130_fd_sc_hd__a31oi_1 U21826 ( .A1(n18297), .A2(n18542), .A3(n16904), 
        .B1(n18783), .Y(n16912) );
  sky130_fd_sc_hd__nor4_1 U21827 ( .A(n18673), .B(n18702), .C(n16906), .D(
        n16905), .Y(n16910) );
  sky130_fd_sc_hd__nand2_1 U21828 ( .A(n18661), .B(n18518), .Y(n18591) );
  sky130_fd_sc_hd__nor4_1 U21829 ( .A(n16908), .B(n18688), .C(n18591), .D(
        n18315), .Y(n16909) );
  sky130_fd_sc_hd__o22ai_1 U21830 ( .A1(n16910), .A2(n18792), .B1(n16909), 
        .B2(n18779), .Y(n16911) );
  sky130_fd_sc_hd__nor3_1 U21831 ( .A(n16913), .B(n16912), .C(n16911), .Y(
        n16914) );
  sky130_fd_sc_hd__o22ai_1 U21832 ( .A1(n16914), .A2(n18552), .B1(n18759), 
        .B2(n25174), .Y(n16940) );
  sky130_fd_sc_hd__a31oi_1 U21833 ( .A1(n16915), .A2(n18252), .A3(n18569), 
        .B1(n18779), .Y(n16923) );
  sky130_fd_sc_hd__nor2_1 U21834 ( .A(n18709), .B(n18638), .Y(n16917) );
  sky130_fd_sc_hd__a31oi_1 U21835 ( .A1(n16917), .A2(n16916), .A3(n18522), 
        .B1(n18792), .Y(n16922) );
  sky130_fd_sc_hd__o21ai_1 U21836 ( .A1(n16919), .A2(n18771), .B1(n16918), .Y(
        n16920) );
  sky130_fd_sc_hd__nor4_1 U21837 ( .A(n16923), .B(n16922), .C(n16921), .D(
        n16920), .Y(n16938) );
  sky130_fd_sc_hd__nor2_1 U21838 ( .A(n18703), .B(n16924), .Y(n18714) );
  sky130_fd_sc_hd__nand2_1 U21839 ( .A(n18642), .B(n18521), .Y(n18563) );
  sky130_fd_sc_hd__nand2_1 U21840 ( .A(n16925), .B(n18698), .Y(n16927) );
  sky130_fd_sc_hd__nor4_1 U21841 ( .A(n18563), .B(n16927), .C(n16926), .D(
        n18299), .Y(n16928) );
  sky130_fd_sc_hd__a31oi_1 U21842 ( .A1(n18714), .A2(n16928), .A3(n16977), 
        .B1(n18792), .Y(n16936) );
  sky130_fd_sc_hd__a31oi_1 U21843 ( .A1(n18297), .A2(n16929), .A3(n18593), 
        .B1(n18779), .Y(n16935) );
  sky130_fd_sc_hd__nor4_1 U21844 ( .A(n18687), .B(n18511), .C(n16931), .D(
        n16930), .Y(n16932) );
  sky130_fd_sc_hd__o22ai_1 U21845 ( .A1(n16933), .A2(n18771), .B1(n16932), 
        .B2(n18783), .Y(n16934) );
  sky130_fd_sc_hd__nor3_1 U21846 ( .A(n16936), .B(n16935), .C(n16934), .Y(
        n16937) );
  sky130_fd_sc_hd__o22ai_1 U21847 ( .A1(n16938), .A2(n18666), .B1(n16937), 
        .B2(n18720), .Y(n16939) );
  sky130_fd_sc_hd__nor3_1 U21848 ( .A(n16941), .B(n16940), .C(n16939), .Y(
        n16967) );
  sky130_fd_sc_hd__a22oi_1 U21849 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[260]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[36]), .Y(n16955) );
  sky130_fd_sc_hd__a22o_1 U21850 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[292]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[324]), .X(n16942) );
  sky130_fd_sc_hd__a21oi_1 U21851 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[356]), .B1(n16942), .Y(n16954) );
  sky130_fd_sc_hd__nand2_1 U21852 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[228]), .Y(n16946) );
  sky130_fd_sc_hd__a21oi_1 U21853 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[452]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n16945) );
  sky130_fd_sc_hd__nand2_1 U21854 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[388]), .Y(n16944) );
  sky130_fd_sc_hd__nand2_1 U21855 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[420]), .Y(n16943) );
  sky130_fd_sc_hd__nand4_1 U21856 ( .A(n16946), .B(n16945), .C(n16944), .D(
        n16943), .Y(n16947) );
  sky130_fd_sc_hd__a21oi_1 U21857 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[196]), .B1(n16947), .Y(n16953) );
  sky130_fd_sc_hd__a22o_1 U21858 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[4]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[68]), .X(n16948) );
  sky130_fd_sc_hd__a21oi_1 U21859 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[100]), .B1(n16948), .Y(n16950) );
  sky130_fd_sc_hd__a22oi_1 U21860 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[164]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[132]), .Y(n16949) );
  sky130_fd_sc_hd__nand2_1 U21861 ( .A(n16950), .B(n16949), .Y(n16951) );
  sky130_fd_sc_hd__nand2_1 U21862 ( .A(n16951), .B(n17639), .Y(n16952) );
  sky130_fd_sc_hd__nand4_1 U21863 ( .A(n16955), .B(n16954), .C(n16953), .D(
        n16952), .Y(n16965) );
  sky130_fd_sc_hd__nor2_1 U21864 ( .A(j202_soc_core_memory0_ram_dout0[484]), 
        .B(n18758), .Y(n16956) );
  sky130_fd_sc_hd__nor2_1 U21865 ( .A(n16956), .B(n18761), .Y(n16964) );
  sky130_fd_sc_hd__a22oi_1 U21866 ( .A1(n18241), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[28]), .B1(n18243), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[4]), .Y(n16958) );
  sky130_fd_sc_hd__a22oi_1 U21867 ( .A1(n18242), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[12]), .B1(n18244), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[20]), .Y(n16957) );
  sky130_fd_sc_hd__a21oi_1 U21868 ( .A1(n16958), .A2(n16957), .B1(n18245), .Y(
        n16959) );
  sky130_fd_sc_hd__a21oi_1 U21869 ( .A1(
        j202_soc_core_ahblite_interconnect_s_hrdata[100]), .A2(n18724), .B1(
        n16959), .Y(n16962) );
  sky130_fd_sc_hd__a22oi_1 U21870 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[4]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[36]), .Y(n16961) );
  sky130_fd_sc_hd__nand2_1 U21871 ( .A(n18727), .B(
        j202_soc_core_ahblite_interconnect_s_hrdata[68]), .Y(n16960) );
  sky130_fd_sc_hd__nand3_1 U21872 ( .A(n16962), .B(n16961), .C(n16960), .Y(
        n16963) );
  sky130_fd_sc_hd__a21oi_1 U21873 ( .A1(n16965), .A2(n16964), .B1(n16963), .Y(
        n16966) );
  sky130_fd_sc_hd__nand2_1 U21874 ( .A(n16967), .B(n16966), .Y(n25256) );
  sky130_fd_sc_hd__a22oi_1 U21875 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[76]), .B1(n18725), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[12]), .Y(n17027) );
  sky130_fd_sc_hd__a22oi_1 U21876 ( .A1(n18724), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[108]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[44]), .Y(n17026) );
  sky130_fd_sc_hd__nor2_1 U21877 ( .A(n16968), .B(n18645), .Y(n18536) );
  sky130_fd_sc_hd__a31oi_1 U21878 ( .A1(n18536), .A2(n18559), .A3(n18519), 
        .B1(n18771), .Y(n16969) );
  sky130_fd_sc_hd__a21oi_1 U21879 ( .A1(n18513), .A2(n18563), .B1(n16969), .Y(
        n16972) );
  sky130_fd_sc_hd__nor2b_1 U21880 ( .B_N(n18556), .A(n18703), .Y(n18545) );
  sky130_fd_sc_hd__o21bai_1 U21881 ( .A1(n18651), .A2(n18655), .B1_N(n18545), 
        .Y(n16971) );
  sky130_fd_sc_hd__a31oi_1 U21883 ( .A1(n16972), .A2(n16971), .A3(n16970), 
        .B1(n18666), .Y(n16973) );
  sky130_fd_sc_hd__a21oi_1 U21884 ( .A1(j202_soc_core_bldc_core_00_pwm_duty[0]), .A2(n18629), .B1(n16973), .Y(n17025) );
  sky130_fd_sc_hd__nand2_1 U21885 ( .A(n16974), .B(n18514), .Y(n18701) );
  sky130_fd_sc_hd__nor4_1 U21886 ( .A(n18564), .B(n18527), .C(n18701), .D(
        n16978), .Y(n18654) );
  sky130_fd_sc_hd__nor2_1 U21887 ( .A(n18654), .B(n18783), .Y(n18532) );
  sky130_fd_sc_hd__nand2_1 U21888 ( .A(n18593), .B(n16975), .Y(n18789) );
  sky130_fd_sc_hd__nor2_1 U21889 ( .A(n16976), .B(n18789), .Y(n18706) );
  sky130_fd_sc_hd__a31oi_1 U21890 ( .A1(n18706), .A2(n18560), .A3(n18559), 
        .B1(n18779), .Y(n16982) );
  sky130_fd_sc_hd__nor4_1 U21891 ( .A(n18703), .B(n18312), .C(n18790), .D(
        n18323), .Y(n16980) );
  sky130_fd_sc_hd__nor4_1 U21892 ( .A(n16978), .B(n18708), .C(n18568), .D(
        n16986), .Y(n16979) );
  sky130_fd_sc_hd__o22ai_1 U21893 ( .A1(n16980), .A2(n18771), .B1(n16979), 
        .B2(n18792), .Y(n16981) );
  sky130_fd_sc_hd__nor3_1 U21894 ( .A(n18532), .B(n16982), .C(n16981), .Y(
        n16995) );
  sky130_fd_sc_hd__nand4b_1 U21895 ( .A_N(n16986), .B(n18533), .C(n16985), .D(
        n16984), .Y(n16993) );
  sky130_fd_sc_hd__nor3_1 U21896 ( .A(n18645), .B(n18702), .C(n16987), .Y(
        n18712) );
  sky130_fd_sc_hd__a21oi_1 U21897 ( .A1(n16988), .A2(n18712), .B1(n18792), .Y(
        n16992) );
  sky130_fd_sc_hd__nor2_1 U21898 ( .A(n18673), .B(n16989), .Y(n18587) );
  sky130_fd_sc_hd__nand2_1 U21899 ( .A(n16990), .B(n18661), .Y(n16997) );
  sky130_fd_sc_hd__nor3_1 U21900 ( .A(n18527), .B(n16997), .C(n18322), .Y(
        n18572) );
  sky130_fd_sc_hd__o22ai_1 U21901 ( .A1(n18587), .A2(n18771), .B1(n18572), 
        .B2(n18783), .Y(n16991) );
  sky130_fd_sc_hd__a211oi_1 U21902 ( .A1(n18655), .A2(n16993), .B1(n16992), 
        .C1(n16991), .Y(n16994) );
  sky130_fd_sc_hd__o22ai_1 U21903 ( .A1(n16995), .A2(n18552), .B1(n16994), 
        .B2(n18722), .Y(n17023) );
  sky130_fd_sc_hd__nor2_1 U21904 ( .A(n16996), .B(n18701), .Y(n16999) );
  sky130_fd_sc_hd__a31oi_1 U21905 ( .A1(n16999), .A2(n18648), .A3(n18555), 
        .B1(n18792), .Y(n17005) );
  sky130_fd_sc_hd__a21oi_1 U21906 ( .A1(n16999), .A2(n16998), .B1(n18783), .Y(
        n17004) );
  sky130_fd_sc_hd__nor3_1 U21907 ( .A(n18564), .B(n17001), .C(n17000), .Y(
        n17002) );
  sky130_fd_sc_hd__nor3_1 U21908 ( .A(n18253), .B(n18585), .C(n18511), .Y(
        n18647) );
  sky130_fd_sc_hd__o22ai_1 U21909 ( .A1(n17002), .A2(n18771), .B1(n18647), 
        .B2(n18779), .Y(n17003) );
  sky130_fd_sc_hd__nor3_1 U21910 ( .A(n17005), .B(n17004), .C(n17003), .Y(
        n17021) );
  sky130_fd_sc_hd__a22oi_1 U21911 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[236]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[204]), .Y(n17009) );
  sky130_fd_sc_hd__a22oi_1 U21912 ( .A1(n18734), .A2(
        j202_soc_core_memory0_ram_dout0[140]), .B1(n18733), .B2(
        j202_soc_core_memory0_ram_dout0[108]), .Y(n17008) );
  sky130_fd_sc_hd__a22oi_1 U21913 ( .A1(n18361), .A2(
        j202_soc_core_memory0_ram_dout0[44]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[76]), .Y(n17007) );
  sky130_fd_sc_hd__nand2_1 U21914 ( .A(n18735), .B(
        j202_soc_core_memory0_ram_dout0[172]), .Y(n17006) );
  sky130_fd_sc_hd__nand4_1 U21915 ( .A(n17009), .B(n17008), .C(n17007), .D(
        n17006), .Y(n17010) );
  sky130_fd_sc_hd__a21oi_1 U21916 ( .A1(n18367), .A2(
        j202_soc_core_memory0_ram_dout0[12]), .B1(n17010), .Y(n17018) );
  sky130_fd_sc_hd__a22oi_1 U21917 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[300]), .B1(n18062), .B2(
        j202_soc_core_memory0_ram_dout0[268]), .Y(n17017) );
  sky130_fd_sc_hd__nand2_1 U21918 ( .A(n18743), .B(
        j202_soc_core_memory0_ram_dout0[364]), .Y(n17014) );
  sky130_fd_sc_hd__a21oi_1 U21919 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[460]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n17013) );
  sky130_fd_sc_hd__nand2_1 U21920 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[396]), .Y(n17012) );
  sky130_fd_sc_hd__nand2_1 U21921 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[428]), .Y(n17011) );
  sky130_fd_sc_hd__nand4_1 U21922 ( .A(n17014), .B(n17013), .C(n17012), .D(
        n17011), .Y(n17015) );
  sky130_fd_sc_hd__a21oi_1 U21923 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[332]), .B1(n17015), .Y(n17016) );
  sky130_fd_sc_hd__o211ai_1 U21924 ( .A1(n18736), .A2(n17018), .B1(n17017), 
        .C1(n17016), .Y(n17019) );
  sky130_fd_sc_hd__o21ai_1 U21925 ( .A1(j202_soc_core_memory0_ram_dout0[492]), 
        .A2(n18758), .B1(n17019), .Y(n17020) );
  sky130_fd_sc_hd__o22ai_1 U21926 ( .A1(n17021), .A2(n18720), .B1(n18761), 
        .B2(n17020), .Y(n17022) );
  sky130_fd_sc_hd__nor2_1 U21927 ( .A(n17023), .B(n17022), .Y(n17024) );
  sky130_fd_sc_hd__nand4_1 U21928 ( .A(n17027), .B(n17026), .C(n17025), .D(
        n17024), .Y(n25312) );
  sky130_fd_sc_hd__nand2_1 U21929 ( .A(n17028), .B(n19095), .Y(n17029) );
  sky130_fd_sc_hd__xnor2_1 U21930 ( .A(n17029), .B(n19920), .Y(n21700) );
  sky130_fd_sc_hd__a21oi_1 U21932 ( .A1(n18859), .A2(n18861), .B1(n17033), .Y(
        n17038) );
  sky130_fd_sc_hd__nand2_1 U21933 ( .A(n17036), .B(n17035), .Y(n17037) );
  sky130_fd_sc_hd__xor2_1 U21934 ( .A(n17038), .B(n17037), .X(n19777) );
  sky130_fd_sc_hd__o22ai_1 U21935 ( .A1(n20007), .A2(n22098), .B1(n17039), 
        .B2(n20005), .Y(n17040) );
  sky130_fd_sc_hd__a21oi_1 U21936 ( .A1(n19777), .A2(n20025), .B1(n17040), .Y(
        n17041) );
  sky130_fd_sc_hd__a21oi_1 U21937 ( .A1(n18867), .A2(n18866), .B1(n17043), .Y(
        n17047) );
  sky130_fd_sc_hd__nand2_1 U21938 ( .A(n17045), .B(n17044), .Y(n17046) );
  sky130_fd_sc_hd__xor2_1 U21939 ( .A(n17047), .B(n17046), .X(n22096) );
  sky130_fd_sc_hd__o22ai_1 U21940 ( .A1(n20014), .A2(n22098), .B1(n17048), 
        .B2(n20012), .Y(n17049) );
  sky130_fd_sc_hd__a21oi_1 U21941 ( .A1(n22096), .A2(n20016), .B1(n17049), .Y(
        n17050) );
  sky130_fd_sc_hd__o21a_1 U21942 ( .A1(j202_soc_core_j22_cpu_macop_MAC_[0]), 
        .A2(n22095), .B1(n17050), .X(n20637) );
  sky130_fd_sc_hd__nand2_1 U21943 ( .A(n17051), .B(n19969), .Y(n17062) );
  sky130_fd_sc_hd__o22ai_1 U21944 ( .A1(n17053), .A2(n19977), .B1(n19971), 
        .B2(n17052), .Y(n17054) );
  sky130_fd_sc_hd__a21oi_1 U21945 ( .A1(n19842), .A2(
        j202_soc_core_j22_cpu_rf_gpr[12]), .B1(n17054), .Y(n17061) );
  sky130_fd_sc_hd__o22ai_1 U21946 ( .A1(n17056), .A2(n19975), .B1(n17055), 
        .B2(n19986), .Y(n17059) );
  sky130_fd_sc_hd__o2bb2ai_1 U21947 ( .B1(n17057), .B2(n19981), .A1_N(
        j202_soc_core_j22_cpu_rf_vbr[12]), .A2_N(n19985), .Y(n17058) );
  sky130_fd_sc_hd__nor2_1 U21948 ( .A(n17059), .B(n17058), .Y(n17060) );
  sky130_fd_sc_hd__nand3_1 U21949 ( .A(n17062), .B(n17061), .C(n17060), .Y(
        n19792) );
  sky130_fd_sc_hd__nand2_1 U21950 ( .A(n19792), .B(n20020), .Y(n17134) );
  sky130_fd_sc_hd__o22ai_1 U21951 ( .A1(n17064), .A2(n19973), .B1(n17063), 
        .B2(n19971), .Y(n17068) );
  sky130_fd_sc_hd__o22ai_1 U21952 ( .A1(n17066), .A2(n19977), .B1(n17065), 
        .B2(n19975), .Y(n17067) );
  sky130_fd_sc_hd__nor2_1 U21953 ( .A(n17068), .B(n17067), .Y(n17073) );
  sky130_fd_sc_hd__a2bb2oi_1 U21954 ( .B1(j202_soc_core_j22_cpu_rf_vbr[4]), 
        .B2(n19985), .A1_N(n17069), .A2_N(n19986), .Y(n17072) );
  sky130_fd_sc_hd__nand2_1 U21955 ( .A(n19842), .B(
        j202_soc_core_j22_cpu_rf_gpr[4]), .Y(n17071) );
  sky130_fd_sc_hd__nand2_1 U21956 ( .A(n19843), .B(
        j202_soc_core_j22_cpu_rf_tmp[4]), .Y(n17070) );
  sky130_fd_sc_hd__nand4_1 U21957 ( .A(n17073), .B(n17072), .C(n17071), .D(
        n17070), .Y(n17074) );
  sky130_fd_sc_hd__a21oi_1 U21958 ( .A1(n17075), .A2(n19969), .B1(n17074), .Y(
        n19476) );
  sky130_fd_sc_hd__nand2_1 U21959 ( .A(n17078), .B(n17077), .Y(n17081) );
  sky130_fd_sc_hd__o21ai_1 U21960 ( .A1(n18873), .A2(n17079), .B1(n18874), .Y(
        n17080) );
  sky130_fd_sc_hd__xnor2_1 U21961 ( .A(n17081), .B(n17080), .Y(n21704) );
  sky130_fd_sc_hd__nand2_1 U21962 ( .A(n22204), .B(
        j202_soc_core_j22_cpu_ml_bufa[4]), .Y(n17091) );
  sky130_fd_sc_hd__a21oi_1 U21963 ( .A1(n19007), .A2(n18879), .B1(n17084), .Y(
        n17089) );
  sky130_fd_sc_hd__nand2_1 U21964 ( .A(n17087), .B(n17086), .Y(n17088) );
  sky130_fd_sc_hd__xor2_1 U21965 ( .A(n17089), .B(n17088), .X(n19429) );
  sky130_fd_sc_hd__nand2_1 U21966 ( .A(n19429), .B(n20025), .Y(n17090) );
  sky130_fd_sc_hd__o211ai_1 U21967 ( .A1(n20005), .A2(n17092), .B1(n17091), 
        .C1(n17090), .Y(n17093) );
  sky130_fd_sc_hd__a21oi_1 U21968 ( .A1(n21704), .A2(n20030), .B1(n17093), .Y(
        n21992) );
  sky130_fd_sc_hd__nand2_1 U21969 ( .A(n17096), .B(n17095), .Y(n17098) );
  sky130_fd_sc_hd__xor2_1 U21970 ( .A(n17098), .B(n17097), .X(n19431) );
  sky130_fd_sc_hd__nand2_1 U21971 ( .A(n19431), .B(n20040), .Y(n17102) );
  sky130_fd_sc_hd__nand2_1 U21972 ( .A(n17099), .B(
        j202_soc_core_j22_cpu_ml_macl[4]), .Y(n17101) );
  sky130_fd_sc_hd__nand2_1 U21973 ( .A(n22225), .B(
        j202_soc_core_j22_cpu_ml_bufa[4]), .Y(n17100) );
  sky130_fd_sc_hd__nand3_1 U21974 ( .A(n17102), .B(n17101), .C(n17100), .Y(
        n21994) );
  sky130_fd_sc_hd__nor2_1 U21975 ( .A(n22125), .B(n21994), .Y(n17103) );
  sky130_fd_sc_hd__a21oi_1 U21976 ( .A1(n21992), .A2(n22125), .B1(n17103), .Y(
        n19473) );
  sky130_fd_sc_hd__nand2_1 U21977 ( .A(n19473), .B(n21137), .Y(n17133) );
  sky130_fd_sc_hd__nand2_1 U21978 ( .A(n25256), .B(n19895), .Y(n17106) );
  sky130_fd_sc_hd__a2bb2oi_1 U21979 ( .B1(n19889), .B2(n25312), .A1_N(n22525), 
        .A2_N(n19891), .Y(n17105) );
  sky130_fd_sc_hd__nand2_1 U21980 ( .A(n22540), .B(n19893), .Y(n17104) );
  sky130_fd_sc_hd__nand2_1 U21981 ( .A(n20839), .B(n17108), .Y(n17109) );
  sky130_fd_sc_hd__nand2_1 U21982 ( .A(n21139), .B(n17109), .Y(n21010) );
  sky130_fd_sc_hd__o21ai_1 U21983 ( .A1(n20908), .A2(n22483), .B1(n21010), .Y(
        n17120) );
  sky130_fd_sc_hd__nand3_1 U21984 ( .A(n22484), .B(n21170), .C(n22483), .Y(
        n17118) );
  sky130_fd_sc_hd__a2bb2oi_1 U21985 ( .B1(n21019), .B2(n21164), .A1_N(n22612), 
        .A2_N(n21163), .Y(n17117) );
  sky130_fd_sc_hd__a2bb2oi_1 U21986 ( .B1(n23310), .B2(n20716), .A1_N(n22064), 
        .A2_N(n20712), .Y(n17116) );
  sky130_fd_sc_hd__o22ai_1 U21987 ( .A1(n21145), .A2(n22705), .B1(n19028), 
        .B2(n22641), .Y(n17113) );
  sky130_fd_sc_hd__xnor2_1 U21988 ( .A(n22483), .B(n22705), .Y(n22444) );
  sky130_fd_sc_hd__o22a_1 U21989 ( .A1(n21108), .A2(n22444), .B1(n22641), .B2(
        n19875), .X(n17112) );
  sky130_fd_sc_hd__nand2_1 U21990 ( .A(n21029), .B(n19173), .Y(n17111) );
  sky130_fd_sc_hd__a2bb2oi_1 U21991 ( .B1(n21156), .B2(n20720), .A1_N(n22488), 
        .A2_N(n21155), .Y(n17110) );
  sky130_fd_sc_hd__nand4b_1 U21992 ( .A_N(n17113), .B(n17112), .C(n17111), .D(
        n17110), .Y(n17114) );
  sky130_fd_sc_hd__a21oi_1 U21993 ( .A1(n19884), .A2(n22705), .B1(n17114), .Y(
        n17115) );
  sky130_fd_sc_hd__nand4_1 U21994 ( .A(n17118), .B(n17117), .C(n17116), .D(
        n17115), .Y(n17119) );
  sky130_fd_sc_hd__a21oi_1 U21995 ( .A1(n22484), .A2(n17120), .B1(n17119), .Y(
        n17132) );
  sky130_fd_sc_hd__a21oi_1 U21996 ( .A1(n22705), .A2(n21089), .B1(n20641), .Y(
        n17121) );
  sky130_fd_sc_hd__a21oi_1 U21998 ( .A1(n19045), .A2(n17834), .B1(n17124), .Y(
        n17129) );
  sky130_fd_sc_hd__nand2_1 U21999 ( .A(n17127), .B(n17126), .Y(n17128) );
  sky130_fd_sc_hd__xor2_1 U22000 ( .A(n17129), .B(n17128), .X(n22053) );
  sky130_fd_sc_hd__a22oi_1 U22001 ( .A1(n22483), .A2(n17130), .B1(n22053), 
        .B2(n21178), .Y(n17131) );
  sky130_fd_sc_hd__nand2_1 U22002 ( .A(n22057), .B(n19905), .Y(n19474) );
  sky130_fd_sc_hd__o21a_1 U22003 ( .A1(n19476), .A2(n19967), .B1(n19474), .X(
        n19794) );
  sky130_fd_sc_hd__o211ai_1 U22004 ( .A1(n20637), .A2(n20067), .B1(n17134), 
        .C1(n19794), .Y(n25302) );
  sky130_fd_sc_hd__nand2_1 U22005 ( .A(j202_soc_core_intc_core_00_rg_itgt[11]), 
        .B(j202_soc_core_intc_core_00_in_intreq[11]), .Y(n17135) );
  sky130_fd_sc_hd__nand2_1 U22006 ( .A(
        j202_soc_core_intc_core_00_in_intreq[10]), .B(
        j202_soc_core_intc_core_00_rg_itgt[10]), .Y(n17182) );
  sky130_fd_sc_hd__nand2_1 U22007 ( .A(n17135), .B(n17182), .Y(n17177) );
  sky130_fd_sc_hd__nand2_1 U22008 ( .A(j202_soc_core_intc_core_00_in_intreq[9]), .B(j202_soc_core_intc_core_00_rg_itgt[9]), .Y(n17169) );
  sky130_fd_sc_hd__nand2_1 U22009 ( .A(j202_soc_core_intc_core_00_in_intreq[8]), .B(j202_soc_core_intc_core_00_rg_itgt[8]), .Y(n17173) );
  sky130_fd_sc_hd__nand2_1 U22010 ( .A(n17169), .B(n17173), .Y(n17194) );
  sky130_fd_sc_hd__nor2_1 U22011 ( .A(n17177), .B(n17194), .Y(n17225) );
  sky130_fd_sc_hd__nand2_1 U22012 ( .A(j202_soc_core_intc_core_00_rg_itgt[13]), 
        .B(j202_soc_core_intc_core_00_in_intreq[13]), .Y(n17136) );
  sky130_fd_sc_hd__nand2_1 U22013 ( .A(j202_soc_core_intc_core_00_rg_itgt[12]), 
        .B(j202_soc_core_intc_core_00_in_intreq[12]), .Y(n17152) );
  sky130_fd_sc_hd__nand2_1 U22014 ( .A(n17136), .B(n17152), .Y(n17222) );
  sky130_fd_sc_hd__nand2_1 U22015 ( .A(j202_soc_core_intc_core_00_rg_itgt[15]), 
        .B(j202_soc_core_intc_core_00_in_intreq[15]), .Y(n17146) );
  sky130_fd_sc_hd__nand2_1 U22016 ( .A(j202_soc_core_intc_core_00_rg_itgt[14]), 
        .B(j202_soc_core_intc_core_00_in_intreq[14]), .Y(n17137) );
  sky130_fd_sc_hd__nand2_1 U22017 ( .A(n17146), .B(n17137), .Y(n17223) );
  sky130_fd_sc_hd__nor2_1 U22018 ( .A(n17222), .B(n17223), .Y(n17138) );
  sky130_fd_sc_hd__nand2_1 U22019 ( .A(n17225), .B(n17138), .Y(n17342) );
  sky130_fd_sc_hd__nand2_1 U22020 ( .A(j202_soc_core_intc_core_00_rg_itgt[3]), 
        .B(j202_soc_core_intc_core_00_in_intreq[3]), .Y(n17232) );
  sky130_fd_sc_hd__nand2_1 U22021 ( .A(j202_soc_core_intc_core_00_rg_itgt[2]), 
        .B(j202_soc_core_intc_core_00_in_intreq[2]), .Y(n17139) );
  sky130_fd_sc_hd__nand2_1 U22022 ( .A(n17232), .B(n17139), .Y(n17311) );
  sky130_fd_sc_hd__nand2_1 U22023 ( .A(j202_soc_core_intc_core_00_rg_itgt[1]), 
        .B(j202_soc_core_intc_core_00_in_intreq[1]), .Y(n17235) );
  sky130_fd_sc_hd__nand2_1 U22024 ( .A(j202_soc_core_intc_core_00_in_intreq[0]), .B(j202_soc_core_intc_core_00_rg_itgt[0]), .Y(n17239) );
  sky130_fd_sc_hd__nand2_1 U22025 ( .A(n17235), .B(n17239), .Y(n17310) );
  sky130_fd_sc_hd__nor2_1 U22026 ( .A(n17311), .B(n17310), .Y(n17142) );
  sky130_fd_sc_hd__nand2_1 U22027 ( .A(j202_soc_core_intc_core_00_rg_itgt[5]), 
        .B(j202_soc_core_intc_core_00_in_intreq[5]), .Y(n17265) );
  sky130_fd_sc_hd__nand2_1 U22028 ( .A(j202_soc_core_intc_core_00_rg_itgt[4]), 
        .B(j202_soc_core_intc_core_00_in_intreq[4]), .Y(n17140) );
  sky130_fd_sc_hd__nand2_1 U22029 ( .A(n17265), .B(n17140), .Y(n17286) );
  sky130_fd_sc_hd__nand2_1 U22030 ( .A(j202_soc_core_intc_core_00_rg_itgt[7]), 
        .B(j202_soc_core_intc_core_00_in_intreq[7]), .Y(n17272) );
  sky130_fd_sc_hd__nand2_1 U22031 ( .A(j202_soc_core_intc_core_00_rg_itgt[6]), 
        .B(j202_soc_core_intc_core_00_in_intreq[6]), .Y(n17141) );
  sky130_fd_sc_hd__nand2_1 U22032 ( .A(n17272), .B(n17141), .Y(n17284) );
  sky130_fd_sc_hd__nor2_1 U22033 ( .A(n17286), .B(n17284), .Y(n17313) );
  sky130_fd_sc_hd__nand2_1 U22034 ( .A(n17142), .B(n17313), .Y(n17341) );
  sky130_fd_sc_hd__nor2_1 U22035 ( .A(n17342), .B(n17341), .Y(n17414) );
  sky130_fd_sc_hd__a22oi_1 U22036 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[18]), .A2(
        j202_soc_core_intc_core_00_rg_itgt[18]), .B1(
        j202_soc_core_intc_core_00_in_intreq[19]), .B2(
        j202_soc_core_intc_core_00_rg_itgt[19]), .Y(n17371) );
  sky130_fd_sc_hd__a22oi_1 U22037 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[17]), .A2(
        j202_soc_core_intc_core_00_rg_itgt[17]), .B1(
        j202_soc_core_intc_core_00_in_intreq[16]), .B2(
        j202_soc_core_intc_core_00_rg_itgt[16]), .Y(n17368) );
  sky130_fd_sc_hd__nand2_1 U22038 ( .A(n17371), .B(n17368), .Y(n17389) );
  sky130_fd_sc_hd__a21oi_1 U22039 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[20]), .A2(
        j202_soc_core_intc_core_00_rg_itgt[20]), .B1(n17389), .Y(n17413) );
  sky130_fd_sc_hd__nand2_1 U22040 ( .A(n17414), .B(n17413), .Y(n21397) );
  sky130_fd_sc_hd__nor2_1 U22041 ( .A(j202_soc_core_rst), .B(n21397), .Y(
        n25370) );
  sky130_fd_sc_hd__nand2_1 U22042 ( .A(n21397), .B(n25731), .Y(n21343) );
  sky130_fd_sc_hd__a22oi_1 U22043 ( .A1(j202_soc_core_intc_core_00_rg_ipr[57]), 
        .A2(n24373), .B1(j202_soc_core_intc_core_00_rg_ipr[56]), .B2(n24743), 
        .Y(n17144) );
  sky130_fd_sc_hd__o22ai_1 U22044 ( .A1(j202_soc_core_intc_core_00_rg_ipr[57]), 
        .A2(n24373), .B1(j202_soc_core_intc_core_00_rg_ipr[58]), .B2(n24374), 
        .Y(n17143) );
  sky130_fd_sc_hd__o22ai_1 U22045 ( .A1(j202_soc_core_intc_core_00_rg_ipr[62]), 
        .A2(n24371), .B1(n17144), .B2(n17143), .Y(n17145) );
  sky130_fd_sc_hd__maj3_1 U22046 ( .A(j202_soc_core_intc_core_00_rg_ipr[59]), 
        .B(n24377), .C(n17145), .X(n17147) );
  sky130_fd_sc_hd__a31oi_1 U22047 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[14]), .A2(
        j202_soc_core_intc_core_00_rg_itgt[14]), .A3(n17147), .B1(n17146), .Y(
        n21348) );
  sky130_fd_sc_hd__nand2_1 U22048 ( .A(n21348), .B(
        j202_soc_core_intc_core_00_rg_ipr[63]), .Y(n17148) );
  sky130_fd_sc_hd__o21ai_1 U22050 ( .A1(j202_soc_core_intc_core_00_rg_ipr[49]), 
        .A2(n24368), .B1(j202_soc_core_intc_core_00_rg_ipr[48]), .Y(n17149) );
  sky130_fd_sc_hd__o22ai_1 U22051 ( .A1(j202_soc_core_intc_core_00_rg_ipr[52]), 
        .A2(n17149), .B1(j202_soc_core_intc_core_00_rg_ipr[53]), .B2(n24665), 
        .Y(n17150) );
  sky130_fd_sc_hd__a222oi_1 U22052 ( .A1(j202_soc_core_intc_core_00_rg_ipr[50]), .A2(n24702), .B1(j202_soc_core_intc_core_00_rg_ipr[50]), .B2(n17150), .C1(
        n24702), .C2(n17150), .Y(n17151) );
  sky130_fd_sc_hd__maj3_1 U22053 ( .A(j202_soc_core_intc_core_00_rg_ipr[55]), 
        .B(n17151), .C(n24366), .X(n17153) );
  sky130_fd_sc_hd__a31oi_1 U22054 ( .A1(j202_soc_core_intc_core_00_rg_itgt[13]), .A2(j202_soc_core_intc_core_00_in_intreq[13]), .A3(n17153), .B1(n17152), .Y(
        n21349) );
  sky130_fd_sc_hd__nand2_1 U22055 ( .A(n21349), .B(n24366), .Y(n17154) );
  sky130_fd_sc_hd__nand2_1 U22057 ( .A(n21349), .B(n24365), .Y(n17155) );
  sky130_fd_sc_hd__nand2_1 U22059 ( .A(n21348), .B(
        j202_soc_core_intc_core_00_rg_ipr[60]), .Y(n17156) );
  sky130_fd_sc_hd__o21ai_1 U22060 ( .A1(n24719), .A2(n21348), .B1(n17156), .Y(
        n17214) );
  sky130_fd_sc_hd__nand2_1 U22061 ( .A(n21349), .B(n24364), .Y(n17157) );
  sky130_fd_sc_hd__o21ai_1 U22062 ( .A1(j202_soc_core_intc_core_00_rg_ipr[52]), 
        .A2(n21349), .B1(n17157), .Y(n17212) );
  sky130_fd_sc_hd__nand2_1 U22063 ( .A(n21349), .B(n24665), .Y(n17158) );
  sky130_fd_sc_hd__nand2_1 U22065 ( .A(n21348), .B(
        j202_soc_core_intc_core_00_rg_ipr[61]), .Y(n17159) );
  sky130_fd_sc_hd__o22ai_1 U22067 ( .A1(n17214), .A2(n17212), .B1(n17208), 
        .B2(n17206), .Y(n17161) );
  sky130_fd_sc_hd__nand2_1 U22068 ( .A(n17208), .B(n17206), .Y(n17160) );
  sky130_fd_sc_hd__nand2_1 U22069 ( .A(n17161), .B(n17160), .Y(n17163) );
  sky130_fd_sc_hd__nand2_1 U22070 ( .A(n21348), .B(
        j202_soc_core_intc_core_00_rg_ipr[62]), .Y(n17162) );
  sky130_fd_sc_hd__o21ai_1 U22071 ( .A1(n24371), .A2(n21348), .B1(n17162), .Y(
        n17200) );
  sky130_fd_sc_hd__maj3_1 U22072 ( .A(n17202), .B(n17163), .C(n17200), .X(
        n17164) );
  sky130_fd_sc_hd__maj3_1 U22073 ( .A(n17166), .B(n17168), .C(n17164), .X(
        n17165) );
  sky130_fd_sc_hd__nand2_1 U22074 ( .A(n21382), .B(n17166), .Y(n17167) );
  sky130_fd_sc_hd__a21oi_1 U22076 ( .A1(j202_soc_core_intc_core_00_rg_ipr[35]), 
        .A2(n24357), .B1(n17169), .Y(n17175) );
  sky130_fd_sc_hd__a22oi_1 U22077 ( .A1(j202_soc_core_intc_core_00_rg_ipr[32]), 
        .A2(n24355), .B1(j202_soc_core_intc_core_00_rg_ipr[33]), .B2(n24559), 
        .Y(n17171) );
  sky130_fd_sc_hd__o22ai_1 U22078 ( .A1(j202_soc_core_intc_core_00_rg_ipr[34]), 
        .A2(n24356), .B1(j202_soc_core_intc_core_00_rg_ipr[33]), .B2(n24559), 
        .Y(n17170) );
  sky130_fd_sc_hd__o22ai_1 U22079 ( .A1(n17171), .A2(n17170), .B1(
        j202_soc_core_intc_core_00_rg_ipr[38]), .B2(n24353), .Y(n17172) );
  sky130_fd_sc_hd__o21ai_1 U22080 ( .A1(j202_soc_core_intc_core_00_rg_ipr[35]), 
        .A2(n24357), .B1(n17172), .Y(n17174) );
  sky130_fd_sc_hd__a21oi_1 U22081 ( .A1(n17175), .A2(n17174), .B1(n17173), .Y(
        n21345) );
  sky130_fd_sc_hd__nand2_1 U22082 ( .A(n21345), .B(
        j202_soc_core_intc_core_00_rg_ipr[35]), .Y(n17176) );
  sky130_fd_sc_hd__o22ai_1 U22084 ( .A1(j202_soc_core_intc_core_00_rg_ipr[44]), 
        .A2(n24358), .B1(j202_soc_core_intc_core_00_rg_ipr[45]), .B2(n24359), 
        .Y(n17178) );
  sky130_fd_sc_hd__o21ai_1 U22085 ( .A1(j202_soc_core_intc_core_00_rg_ipr[42]), 
        .A2(n24363), .B1(n17178), .Y(n17179) );
  sky130_fd_sc_hd__a21oi_1 U22086 ( .A1(j202_soc_core_intc_core_00_rg_ipr[45]), 
        .A2(n24359), .B1(n17179), .Y(n17181) );
  sky130_fd_sc_hd__o22ai_1 U22087 ( .A1(j202_soc_core_intc_core_00_rg_ipr[46]), 
        .A2(n24360), .B1(j202_soc_core_intc_core_00_rg_ipr[47]), .B2(n24615), 
        .Y(n17180) );
  sky130_fd_sc_hd__o22ai_1 U22088 ( .A1(j202_soc_core_intc_core_00_rg_ipr[43]), 
        .A2(n24651), .B1(n17181), .B2(n17180), .Y(n17183) );
  sky130_fd_sc_hd__a31oi_1 U22089 ( .A1(j202_soc_core_intc_core_00_rg_itgt[11]), .A2(j202_soc_core_intc_core_00_in_intreq[11]), .A3(n17183), .B1(n17182), .Y(
        n21346) );
  sky130_fd_sc_hd__nand2_1 U22090 ( .A(n21346), .B(n24615), .Y(n17184) );
  sky130_fd_sc_hd__nand2_1 U22092 ( .A(n21346), .B(n24360), .Y(n17185) );
  sky130_fd_sc_hd__o21ai_1 U22093 ( .A1(j202_soc_core_intc_core_00_rg_ipr[46]), 
        .A2(n21346), .B1(n17185), .Y(n17203) );
  sky130_fd_sc_hd__nand2_1 U22094 ( .A(n21345), .B(n24351), .Y(n17186) );
  sky130_fd_sc_hd__o21ai_1 U22095 ( .A1(j202_soc_core_intc_core_00_rg_ipr[36]), 
        .A2(n21345), .B1(n17186), .Y(n17215) );
  sky130_fd_sc_hd__nand2_1 U22096 ( .A(n21346), .B(n24359), .Y(n17187) );
  sky130_fd_sc_hd__o21ai_1 U22097 ( .A1(j202_soc_core_intc_core_00_rg_ipr[45]), 
        .A2(n21346), .B1(n17187), .Y(n17209) );
  sky130_fd_sc_hd__nand2_1 U22098 ( .A(n21345), .B(
        j202_soc_core_intc_core_00_rg_ipr[33]), .Y(n17188) );
  sky130_fd_sc_hd__o21ai_1 U22099 ( .A1(n24559), .A2(n21345), .B1(n17188), .Y(
        n17211) );
  sky130_fd_sc_hd__nand2_1 U22100 ( .A(n21346), .B(n24358), .Y(n17189) );
  sky130_fd_sc_hd__o21ai_1 U22101 ( .A1(j202_soc_core_intc_core_00_rg_ipr[44]), 
        .A2(n21346), .B1(n17189), .Y(n17217) );
  sky130_fd_sc_hd__o21ai_1 U22102 ( .A1(n17209), .A2(n17211), .B1(n17217), .Y(
        n17190) );
  sky130_fd_sc_hd__o2bb2ai_1 U22103 ( .B1(n17215), .B2(n17190), .A1_N(n17209), 
        .A2_N(n17211), .Y(n17192) );
  sky130_fd_sc_hd__nand2_1 U22104 ( .A(n21345), .B(
        j202_soc_core_intc_core_00_rg_ipr[34]), .Y(n17191) );
  sky130_fd_sc_hd__o21ai_1 U22105 ( .A1(n24356), .A2(n21345), .B1(n17191), .Y(
        n17205) );
  sky130_fd_sc_hd__maj3_1 U22106 ( .A(n17203), .B(n17192), .C(n17205), .X(
        n17193) );
  sky130_fd_sc_hd__maj3_1 U22107 ( .A(n17197), .B(n17199), .C(n17193), .X(
        n17195) );
  sky130_fd_sc_hd__nand2_1 U22109 ( .A(n17197), .B(n21379), .Y(n17198) );
  sky130_fd_sc_hd__nand2_1 U22111 ( .A(n17200), .B(n21350), .Y(n17201) );
  sky130_fd_sc_hd__o21ai_1 U22112 ( .A1(n17202), .A2(n21350), .B1(n17201), .Y(
        n17320) );
  sky130_fd_sc_hd__nand2_1 U22113 ( .A(n17203), .B(n21379), .Y(n17204) );
  sky130_fd_sc_hd__nand2_1 U22115 ( .A(n17206), .B(n21350), .Y(n17207) );
  sky130_fd_sc_hd__o21ai_1 U22116 ( .A1(n17208), .A2(n21350), .B1(n17207), .Y(
        n17330) );
  sky130_fd_sc_hd__nand2_1 U22117 ( .A(n17209), .B(n21379), .Y(n17210) );
  sky130_fd_sc_hd__o21ai_1 U22118 ( .A1(n17211), .A2(n21379), .B1(n17210), .Y(
        n17331) );
  sky130_fd_sc_hd__nand2_1 U22119 ( .A(n21382), .B(n17212), .Y(n17213) );
  sky130_fd_sc_hd__nand2b_1 U22121 ( .A_N(n17215), .B(n21347), .Y(n17216) );
  sky130_fd_sc_hd__o21ai_1 U22122 ( .A1(n17217), .A2(n21347), .B1(n17216), .Y(
        n17324) );
  sky130_fd_sc_hd__nand2_1 U22123 ( .A(n17326), .B(n17324), .Y(n17218) );
  sky130_fd_sc_hd__fa_1 U22124 ( .A(n17330), .B(n17331), .CIN(n17218), .COUT(
        n17219), .SUM() );
  sky130_fd_sc_hd__maj3_1 U22125 ( .A(n17221), .B(n17226), .C(n17220), .X(
        n17224) );
  sky130_fd_sc_hd__o22ai_1 U22126 ( .A1(n17225), .A2(n17224), .B1(n17223), 
        .B2(n17222), .Y(n21381) );
  sky130_fd_sc_hd__nand2b_1 U22127 ( .A_N(n17226), .B(n21381), .Y(n17227) );
  sky130_fd_sc_hd__o21ai_1 U22128 ( .A1(n17228), .A2(n21381), .B1(n17227), .Y(
        n17346) );
  sky130_fd_sc_hd__a22oi_1 U22129 ( .A1(j202_soc_core_intc_core_00_rg_ipr[9]), 
        .A2(n24632), .B1(j202_soc_core_intc_core_00_rg_ipr[8]), .B2(n24623), 
        .Y(n17230) );
  sky130_fd_sc_hd__o22ai_1 U22130 ( .A1(j202_soc_core_intc_core_00_rg_ipr[9]), 
        .A2(n24632), .B1(j202_soc_core_intc_core_00_rg_ipr[10]), .B2(n24641), 
        .Y(n17229) );
  sky130_fd_sc_hd__o22ai_1 U22131 ( .A1(j202_soc_core_intc_core_00_rg_ipr[14]), 
        .A2(n24609), .B1(n17230), .B2(n17229), .Y(n17231) );
  sky130_fd_sc_hd__maj3_1 U22132 ( .A(j202_soc_core_intc_core_00_rg_ipr[11]), 
        .B(n24653), .C(n17231), .X(n17233) );
  sky130_fd_sc_hd__a31oi_1 U22133 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[2]), .A2(
        j202_soc_core_intc_core_00_rg_itgt[2]), .A3(n17233), .B1(n17232), .Y(
        n21357) );
  sky130_fd_sc_hd__nand2_1 U22134 ( .A(n21357), .B(n24653), .Y(n17234) );
  sky130_fd_sc_hd__a21oi_1 U22136 ( .A1(j202_soc_core_intc_core_00_rg_ipr[3]), 
        .A2(n24382), .B1(n17235), .Y(n17241) );
  sky130_fd_sc_hd__o21ai_1 U22137 ( .A1(j202_soc_core_intc_core_00_rg_ipr[1]), 
        .A2(n24381), .B1(j202_soc_core_intc_core_00_rg_ipr[0]), .Y(n17236) );
  sky130_fd_sc_hd__o22ai_1 U22138 ( .A1(j202_soc_core_intc_core_00_rg_ipr[4]), 
        .A2(n17236), .B1(j202_soc_core_intc_core_00_rg_ipr[5]), .B2(n24510), 
        .Y(n17237) );
  sky130_fd_sc_hd__maj3_1 U22139 ( .A(j202_soc_core_intc_core_00_rg_ipr[2]), 
        .B(n24561), .C(n17237), .X(n17238) );
  sky130_fd_sc_hd__o21ai_1 U22140 ( .A1(j202_soc_core_intc_core_00_rg_ipr[3]), 
        .A2(n24382), .B1(n17238), .Y(n17240) );
  sky130_fd_sc_hd__a21oi_1 U22141 ( .A1(n17241), .A2(n17240), .B1(n17239), .Y(
        n21358) );
  sky130_fd_sc_hd__nand2_1 U22142 ( .A(n21358), .B(n24530), .Y(n17242) );
  sky130_fd_sc_hd__nand2_1 U22144 ( .A(n21358), .B(n24520), .Y(n17243) );
  sky130_fd_sc_hd__o21ai_1 U22145 ( .A1(j202_soc_core_intc_core_00_rg_ipr[6]), 
        .A2(n21358), .B1(n17243), .Y(n17259) );
  sky130_fd_sc_hd__nand2_1 U22146 ( .A(n21357), .B(
        j202_soc_core_intc_core_00_rg_ipr[12]), .Y(n17244) );
  sky130_fd_sc_hd__o21ai_1 U22147 ( .A1(n24588), .A2(n21357), .B1(n17244), .Y(
        n17300) );
  sky130_fd_sc_hd__nand2_1 U22148 ( .A(n21358), .B(n24500), .Y(n17245) );
  sky130_fd_sc_hd__o21ai_1 U22149 ( .A1(j202_soc_core_intc_core_00_rg_ipr[4]), 
        .A2(n21358), .B1(n17245), .Y(n17301) );
  sky130_fd_sc_hd__nand2_1 U22150 ( .A(n21358), .B(n24510), .Y(n17246) );
  sky130_fd_sc_hd__o21ai_1 U22151 ( .A1(j202_soc_core_intc_core_00_rg_ipr[5]), 
        .A2(n21358), .B1(n17246), .Y(n17294) );
  sky130_fd_sc_hd__nand2_1 U22152 ( .A(n21357), .B(
        j202_soc_core_intc_core_00_rg_ipr[13]), .Y(n17247) );
  sky130_fd_sc_hd__o21ai_1 U22153 ( .A1(n24600), .A2(n21357), .B1(n17247), .Y(
        n17293) );
  sky130_fd_sc_hd__o22ai_1 U22154 ( .A1(n17300), .A2(n17301), .B1(n17294), 
        .B2(n17293), .Y(n17249) );
  sky130_fd_sc_hd__nand2_1 U22155 ( .A(n17294), .B(n17293), .Y(n17248) );
  sky130_fd_sc_hd__nand2_1 U22156 ( .A(n17249), .B(n17248), .Y(n17251) );
  sky130_fd_sc_hd__nand2_1 U22157 ( .A(n21357), .B(
        j202_soc_core_intc_core_00_rg_ipr[14]), .Y(n17250) );
  sky130_fd_sc_hd__o21ai_1 U22158 ( .A1(n24609), .A2(n21357), .B1(n17250), .Y(
        n17258) );
  sky130_fd_sc_hd__maj3_1 U22159 ( .A(n17259), .B(n17251), .C(n17258), .X(
        n17252) );
  sky130_fd_sc_hd__maj3_1 U22160 ( .A(n17255), .B(n17253), .C(n17252), .X(
        n17254) );
  sky130_fd_sc_hd__nand2b_1 U22161 ( .A_N(n17255), .B(n21375), .Y(n17256) );
  sky130_fd_sc_hd__nand2b_1 U22163 ( .A_N(n17259), .B(n21375), .Y(n17260) );
  sky130_fd_sc_hd__o21ai_1 U22164 ( .A1(n17261), .A2(n21375), .B1(n17260), .Y(
        n17319) );
  sky130_fd_sc_hd__a22oi_1 U22165 ( .A1(j202_soc_core_intc_core_00_rg_ipr[17]), 
        .A2(n24388), .B1(j202_soc_core_intc_core_00_rg_ipr[16]), .B2(n24386), 
        .Y(n17263) );
  sky130_fd_sc_hd__o22ai_1 U22166 ( .A1(j202_soc_core_intc_core_00_rg_ipr[17]), 
        .A2(n24388), .B1(j202_soc_core_intc_core_00_rg_ipr[18]), .B2(n24706), 
        .Y(n17262) );
  sky130_fd_sc_hd__o22ai_1 U22167 ( .A1(j202_soc_core_intc_core_00_rg_ipr[22]), 
        .A2(n24385), .B1(n17263), .B2(n17262), .Y(n17264) );
  sky130_fd_sc_hd__maj3_1 U22168 ( .A(j202_soc_core_intc_core_00_rg_ipr[19]), 
        .B(n24391), .C(n17264), .X(n17266) );
  sky130_fd_sc_hd__a31oi_1 U22169 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[4]), .A2(
        j202_soc_core_intc_core_00_rg_itgt[4]), .A3(n17266), .B1(n17265), .Y(
        n21355) );
  sky130_fd_sc_hd__nand2_1 U22170 ( .A(n21355), .B(
        j202_soc_core_intc_core_00_rg_ipr[22]), .Y(n17267) );
  sky130_fd_sc_hd__nand2_1 U22172 ( .A(n21355), .B(
        j202_soc_core_intc_core_00_rg_ipr[23]), .Y(n17268) );
  sky130_fd_sc_hd__o21ai_1 U22173 ( .A1(n24680), .A2(n21355), .B1(n17268), .Y(
        n17308) );
  sky130_fd_sc_hd__a22oi_1 U22174 ( .A1(j202_soc_core_intc_core_00_rg_ipr[25]), 
        .A2(n24401), .B1(j202_soc_core_intc_core_00_rg_ipr[24]), .B2(n24747), 
        .Y(n17270) );
  sky130_fd_sc_hd__o22ai_1 U22175 ( .A1(j202_soc_core_intc_core_00_rg_ipr[25]), 
        .A2(n24401), .B1(j202_soc_core_intc_core_00_rg_ipr[26]), .B2(n24403), 
        .Y(n17269) );
  sky130_fd_sc_hd__o22ai_1 U22176 ( .A1(n17270), .A2(n17269), .B1(
        j202_soc_core_intc_core_00_rg_ipr[30]), .B2(n24396), .Y(n17271) );
  sky130_fd_sc_hd__maj3_1 U22177 ( .A(j202_soc_core_intc_core_00_rg_ipr[27]), 
        .B(n24407), .C(n17271), .X(n17273) );
  sky130_fd_sc_hd__a31oi_1 U22178 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[6]), .A2(
        j202_soc_core_intc_core_00_rg_itgt[6]), .A3(n17273), .B1(n17272), .Y(
        n21356) );
  sky130_fd_sc_hd__nand2_1 U22179 ( .A(n21356), .B(n24403), .Y(n17274) );
  sky130_fd_sc_hd__nand2_1 U22181 ( .A(n21355), .B(n24386), .Y(n17275) );
  sky130_fd_sc_hd__o21ai_1 U22182 ( .A1(j202_soc_core_intc_core_00_rg_ipr[16]), 
        .A2(n21355), .B1(n17275), .Y(n17292) );
  sky130_fd_sc_hd__nand2_1 U22183 ( .A(n21356), .B(n24401), .Y(n17276) );
  sky130_fd_sc_hd__o21ai_1 U22184 ( .A1(j202_soc_core_intc_core_00_rg_ipr[25]), 
        .A2(n21356), .B1(n17276), .Y(n17297) );
  sky130_fd_sc_hd__nand2_1 U22185 ( .A(n21355), .B(
        j202_soc_core_intc_core_00_rg_ipr[21]), .Y(n17277) );
  sky130_fd_sc_hd__o21ai_1 U22186 ( .A1(n24666), .A2(n21355), .B1(n17277), .Y(
        n17299) );
  sky130_fd_sc_hd__nand2_1 U22187 ( .A(n21356), .B(n24747), .Y(n17278) );
  sky130_fd_sc_hd__o21ai_1 U22189 ( .A1(n17297), .A2(n17299), .B1(n17290), .Y(
        n17279) );
  sky130_fd_sc_hd__o2bb2ai_1 U22190 ( .B1(n17292), .B2(n17279), .A1_N(n17297), 
        .A2_N(n17299), .Y(n17280) );
  sky130_fd_sc_hd__maj3_1 U22191 ( .A(n17287), .B(n17289), .C(n17280), .X(
        n17282) );
  sky130_fd_sc_hd__nand2_1 U22192 ( .A(n21356), .B(n24407), .Y(n17281) );
  sky130_fd_sc_hd__nand2_1 U22195 ( .A(n17308), .B(n17282), .Y(n17283) );
  sky130_fd_sc_hd__nand3_1 U22196 ( .A(n17285), .B(n17284), .C(n17283), .Y(
        n21354) );
  sky130_fd_sc_hd__nand2_1 U22197 ( .A(n17286), .B(n21354), .Y(n21378) );
  sky130_fd_sc_hd__nand2_1 U22198 ( .A(n21378), .B(n17287), .Y(n17288) );
  sky130_fd_sc_hd__o21ai_1 U22199 ( .A1(n17289), .A2(n21378), .B1(n17288), .Y(
        n17317) );
  sky130_fd_sc_hd__nand2b_1 U22200 ( .A_N(n17290), .B(n21378), .Y(n17291) );
  sky130_fd_sc_hd__o21ai_1 U22201 ( .A1(n17292), .A2(n21378), .B1(n17291), .Y(
        n17327) );
  sky130_fd_sc_hd__nand2b_1 U22202 ( .A_N(n17294), .B(n21375), .Y(n17295) );
  sky130_fd_sc_hd__o21ai_1 U22203 ( .A1(n17296), .A2(n21375), .B1(n17295), .Y(
        n17336) );
  sky130_fd_sc_hd__nand2_1 U22204 ( .A(n21378), .B(n17297), .Y(n17298) );
  sky130_fd_sc_hd__o21ai_1 U22205 ( .A1(n17299), .A2(n21378), .B1(n17298), .Y(
        n17334) );
  sky130_fd_sc_hd__nand2b_1 U22206 ( .A_N(n17301), .B(n21375), .Y(n17302) );
  sky130_fd_sc_hd__o21ai_1 U22208 ( .A1(n17336), .A2(n17334), .B1(n17329), .Y(
        n17304) );
  sky130_fd_sc_hd__o2bb2ai_1 U22209 ( .B1(n17327), .B2(n17304), .A1_N(n17334), 
        .A2_N(n17336), .Y(n17305) );
  sky130_fd_sc_hd__maj3_1 U22210 ( .A(n17319), .B(n17317), .C(n17305), .X(
        n17309) );
  sky130_fd_sc_hd__nand2_1 U22211 ( .A(n21378), .B(n17306), .Y(n17307) );
  sky130_fd_sc_hd__o21ai_1 U22212 ( .A1(n17308), .A2(n21378), .B1(n17307), .Y(
        n17314) );
  sky130_fd_sc_hd__maj3_1 U22213 ( .A(n17309), .B(n17316), .C(n17314), .X(
        n17312) );
  sky130_fd_sc_hd__o22ai_1 U22214 ( .A1(n17313), .A2(n17312), .B1(n17311), 
        .B2(n17310), .Y(n21361) );
  sky130_fd_sc_hd__nand2_1 U22215 ( .A(n21361), .B(n17314), .Y(n17315) );
  sky130_fd_sc_hd__nand2_1 U22217 ( .A(n21361), .B(n17317), .Y(n17318) );
  sky130_fd_sc_hd__o21ai_1 U22218 ( .A1(n17319), .A2(n21361), .B1(n17318), .Y(
        n17394) );
  sky130_fd_sc_hd__nand2b_1 U22219 ( .A_N(n17321), .B(n21381), .Y(n17322) );
  sky130_fd_sc_hd__o21ai_1 U22220 ( .A1(n17323), .A2(n21381), .B1(n17322), .Y(
        n17396) );
  sky130_fd_sc_hd__nand2_1 U22221 ( .A(n21381), .B(n17324), .Y(n17325) );
  sky130_fd_sc_hd__nand2b_1 U22223 ( .A_N(n17327), .B(n21361), .Y(n17328) );
  sky130_fd_sc_hd__o21ai_1 U22224 ( .A1(n17329), .A2(n21361), .B1(n17328), .Y(
        n17399) );
  sky130_fd_sc_hd__nand2b_1 U22225 ( .A_N(n17331), .B(n21381), .Y(n17332) );
  sky130_fd_sc_hd__o21ai_1 U22226 ( .A1(n17333), .A2(n21381), .B1(n17332), .Y(
        n17404) );
  sky130_fd_sc_hd__nand2_1 U22227 ( .A(n21361), .B(n17334), .Y(n17335) );
  sky130_fd_sc_hd__o21ai_1 U22228 ( .A1(n17336), .A2(n21361), .B1(n17335), .Y(
        n17402) );
  sky130_fd_sc_hd__o22ai_1 U22229 ( .A1(n17401), .A2(n17399), .B1(n17404), 
        .B2(n17402), .Y(n17338) );
  sky130_fd_sc_hd__nand2_1 U22230 ( .A(n17404), .B(n17402), .Y(n17337) );
  sky130_fd_sc_hd__nand2_1 U22231 ( .A(n17338), .B(n17337), .Y(n17339) );
  sky130_fd_sc_hd__maj3_1 U22232 ( .A(n17394), .B(n17396), .C(n17339), .X(
        n17340) );
  sky130_fd_sc_hd__maj3_1 U22233 ( .A(n17346), .B(n17344), .C(n17340), .X(
        n17343) );
  sky130_fd_sc_hd__nand2_1 U22234 ( .A(n21365), .B(n17344), .Y(n17345) );
  sky130_fd_sc_hd__o21ai_1 U22235 ( .A1(n17346), .A2(n21365), .B1(n17345), .Y(
        n22786) );
  sky130_fd_sc_hd__o21ai_1 U22236 ( .A1(j202_soc_core_intc_core_00_rg_ipr[65]), 
        .A2(n24329), .B1(j202_soc_core_intc_core_00_rg_ipr[64]), .Y(n17347) );
  sky130_fd_sc_hd__o22ai_1 U22237 ( .A1(j202_soc_core_intc_core_00_rg_ipr[68]), 
        .A2(n17347), .B1(j202_soc_core_intc_core_00_rg_ipr[69]), .B2(n24511), 
        .Y(n17348) );
  sky130_fd_sc_hd__a222oi_1 U22238 ( .A1(j202_soc_core_intc_core_00_rg_ipr[66]), .A2(n24562), .B1(j202_soc_core_intc_core_00_rg_ipr[66]), .B2(n17348), .C1(
        n24562), .C2(n17348), .Y(n17349) );
  sky130_fd_sc_hd__maj3_1 U22239 ( .A(j202_soc_core_intc_core_00_rg_ipr[71]), 
        .B(n24531), .C(n17349), .X(n17351) );
  sky130_fd_sc_hd__nand2_1 U22240 ( .A(
        j202_soc_core_intc_core_00_in_intreq[16]), .B(
        j202_soc_core_intc_core_00_rg_itgt[16]), .Y(n17350) );
  sky130_fd_sc_hd__a31oi_1 U22241 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[17]), .A2(
        j202_soc_core_intc_core_00_rg_itgt[17]), .A3(n17351), .B1(n17350), .Y(
        n21368) );
  sky130_fd_sc_hd__nand2_1 U22242 ( .A(n21368), .B(
        j202_soc_core_intc_core_00_rg_ipr[67]), .Y(n17352) );
  sky130_fd_sc_hd__o21ai_1 U22243 ( .A1(n24330), .A2(n21368), .B1(n17352), .Y(
        n17374) );
  sky130_fd_sc_hd__o22ai_1 U22245 ( .A1(j202_soc_core_intc_core_00_rg_ipr[77]), 
        .A2(n24597), .B1(j202_soc_core_intc_core_00_rg_ipr[76]), .B2(n17353), 
        .Y(n17354) );
  sky130_fd_sc_hd__a222oi_1 U22246 ( .A1(j202_soc_core_intc_core_00_rg_ipr[74]), .A2(n24642), .B1(j202_soc_core_intc_core_00_rg_ipr[74]), .B2(n17354), .C1(
        n24642), .C2(n17354), .Y(n17355) );
  sky130_fd_sc_hd__maj3_1 U22247 ( .A(j202_soc_core_intc_core_00_rg_ipr[79]), 
        .B(n24616), .C(n17355), .X(n17357) );
  sky130_fd_sc_hd__nand2_1 U22248 ( .A(
        j202_soc_core_intc_core_00_in_intreq[18]), .B(
        j202_soc_core_intc_core_00_rg_itgt[18]), .Y(n17356) );
  sky130_fd_sc_hd__a31oi_1 U22249 ( .A1(j202_soc_core_intc_core_00_rg_itgt[19]), .A2(j202_soc_core_intc_core_00_in_intreq[19]), .A3(n17357), .B1(n17356), .Y(
        n21369) );
  sky130_fd_sc_hd__nand2_1 U22250 ( .A(n21369), .B(n24616), .Y(n17358) );
  sky130_fd_sc_hd__o21ai_1 U22251 ( .A1(j202_soc_core_intc_core_00_rg_ipr[79]), 
        .A2(n21369), .B1(n17358), .Y(n17372) );
  sky130_fd_sc_hd__nand2_1 U22252 ( .A(n21369), .B(n24606), .Y(n17359) );
  sky130_fd_sc_hd__o21ai_1 U22253 ( .A1(j202_soc_core_intc_core_00_rg_ipr[78]), 
        .A2(n21369), .B1(n17359), .Y(n17375) );
  sky130_fd_sc_hd__nand2_1 U22254 ( .A(n21368), .B(
        j202_soc_core_intc_core_00_rg_ipr[66]), .Y(n17360) );
  sky130_fd_sc_hd__nand2_1 U22256 ( .A(n21368), .B(n24501), .Y(n17361) );
  sky130_fd_sc_hd__o21ai_1 U22257 ( .A1(j202_soc_core_intc_core_00_rg_ipr[68]), 
        .A2(n21368), .B1(n17361), .Y(n17378) );
  sky130_fd_sc_hd__nand2_1 U22258 ( .A(n21369), .B(n24597), .Y(n17362) );
  sky130_fd_sc_hd__o21ai_1 U22259 ( .A1(j202_soc_core_intc_core_00_rg_ipr[77]), 
        .A2(n21369), .B1(n17362), .Y(n17382) );
  sky130_fd_sc_hd__nand2_1 U22260 ( .A(n21368), .B(
        j202_soc_core_intc_core_00_rg_ipr[65]), .Y(n17363) );
  sky130_fd_sc_hd__o21ai_1 U22261 ( .A1(n24329), .A2(n21368), .B1(n17363), .Y(
        n17384) );
  sky130_fd_sc_hd__nand2_1 U22262 ( .A(n21369), .B(n24589), .Y(n17364) );
  sky130_fd_sc_hd__o2bb2ai_1 U22265 ( .B1(n17378), .B2(n17365), .A1_N(n17382), 
        .A2_N(n17384), .Y(n17366) );
  sky130_fd_sc_hd__maj3_1 U22266 ( .A(n17375), .B(n17377), .C(n17366), .X(
        n17367) );
  sky130_fd_sc_hd__maj3_1 U22267 ( .A(n17372), .B(n17367), .C(n17374), .X(
        n17370) );
  sky130_fd_sc_hd__o21ai_1 U22268 ( .A1(n17371), .A2(n17370), .B1(n17369), .Y(
        n21387) );
  sky130_fd_sc_hd__nand2_1 U22269 ( .A(n17372), .B(n21387), .Y(n17373) );
  sky130_fd_sc_hd__o21ai_1 U22270 ( .A1(n17374), .A2(n21387), .B1(n17373), .Y(
        n17393) );
  sky130_fd_sc_hd__nand2_1 U22271 ( .A(
        j202_soc_core_intc_core_00_in_intreq[20]), .B(
        j202_soc_core_intc_core_00_rg_itgt[20]), .Y(n17391) );
  sky130_fd_sc_hd__nand2_1 U22272 ( .A(n17375), .B(n21387), .Y(n17376) );
  sky130_fd_sc_hd__o21ai_1 U22273 ( .A1(n17377), .A2(n21387), .B1(n17376), .Y(
        n17410) );
  sky130_fd_sc_hd__nand2_1 U22274 ( .A(n17379), .B(n21387), .Y(n17380) );
  sky130_fd_sc_hd__nand2_1 U22276 ( .A(n17382), .B(n21387), .Y(n17383) );
  sky130_fd_sc_hd__o22ai_1 U22278 ( .A1(j202_soc_core_intc_core_00_rg_ipr[80]), 
        .A2(n17398), .B1(j202_soc_core_intc_core_00_rg_ipr[81]), .B2(n17406), 
        .Y(n17386) );
  sky130_fd_sc_hd__nand2_1 U22279 ( .A(j202_soc_core_intc_core_00_rg_ipr[81]), 
        .B(n17406), .Y(n17385) );
  sky130_fd_sc_hd__nand2_1 U22280 ( .A(n17386), .B(n17385), .Y(n17387) );
  sky130_fd_sc_hd__maj3_1 U22281 ( .A(n17410), .B(
        j202_soc_core_intc_core_00_rg_ipr[82]), .C(n17387), .X(n17388) );
  sky130_fd_sc_hd__a222oi_1 U22282 ( .A1(j202_soc_core_intc_core_00_rg_ipr[83]), .A2(n17393), .B1(j202_soc_core_intc_core_00_rg_ipr[83]), .B2(n17388), .C1(
        n17393), .C2(n17388), .Y(n17390) );
  sky130_fd_sc_hd__o21ai_1 U22283 ( .A1(n17391), .A2(n17390), .B1(n17389), .Y(
        n21366) );
  sky130_fd_sc_hd__nand2_1 U22284 ( .A(j202_soc_core_intc_core_00_rg_ipr[83]), 
        .B(n21366), .Y(n17392) );
  sky130_fd_sc_hd__nand2_1 U22286 ( .A(n21365), .B(n17394), .Y(n17395) );
  sky130_fd_sc_hd__nand2_1 U22288 ( .A(j202_soc_core_intc_core_00_rg_ipr[80]), 
        .B(n21366), .Y(n17397) );
  sky130_fd_sc_hd__nand2_1 U22290 ( .A(n21365), .B(n17399), .Y(n17400) );
  sky130_fd_sc_hd__nand2_1 U22292 ( .A(n21365), .B(n17402), .Y(n17403) );
  sky130_fd_sc_hd__nand2_1 U22294 ( .A(j202_soc_core_intc_core_00_rg_ipr[81]), 
        .B(n21366), .Y(n17405) );
  sky130_fd_sc_hd__o22ai_1 U22296 ( .A1(n22061), .A2(n22063), .B1(n22044), 
        .B2(n22042), .Y(n17408) );
  sky130_fd_sc_hd__nand2_1 U22297 ( .A(n22044), .B(n22042), .Y(n17407) );
  sky130_fd_sc_hd__nand2_1 U22298 ( .A(n17408), .B(n17407), .Y(n17411) );
  sky130_fd_sc_hd__nand2_1 U22299 ( .A(j202_soc_core_intc_core_00_rg_ipr[82]), 
        .B(n21366), .Y(n17409) );
  sky130_fd_sc_hd__o21ai_1 U22300 ( .A1(n17410), .A2(n21366), .B1(n17409), .Y(
        n21854) );
  sky130_fd_sc_hd__maj3_1 U22301 ( .A(n21856), .B(n17411), .C(n21854), .X(
        n17412) );
  sky130_fd_sc_hd__maj3_1 U22302 ( .A(n22786), .B(n22783), .C(n17412), .X(
        n17416) );
  sky130_fd_sc_hd__a21oi_1 U22303 ( .A1(n17416), .A2(n17415), .B1(n17414), .Y(
        n21388) );
  sky130_fd_sc_hd__nor2_1 U22304 ( .A(n21343), .B(n21388), .Y(n25390) );
  sky130_fd_sc_hd__nor3_1 U22305 ( .A(n17916), .B(n17509), .C(n17530), .Y(
        n17754) );
  sky130_fd_sc_hd__a31oi_1 U22306 ( .A1(n17418), .A2(n17754), .A3(n17417), 
        .B1(n18437), .Y(n17426) );
  sky130_fd_sc_hd__nor2_1 U22307 ( .A(n17744), .B(n17420), .Y(n17527) );
  sky130_fd_sc_hd__nand2_1 U22308 ( .A(n17868), .B(n17675), .Y(n18434) );
  sky130_fd_sc_hd__nor3_1 U22309 ( .A(n17530), .B(n17605), .C(n18434), .Y(
        n17419) );
  sky130_fd_sc_hd__a31oi_1 U22310 ( .A1(n17527), .A2(n17613), .A3(n17419), 
        .B1(n18423), .Y(n17425) );
  sky130_fd_sc_hd__nand2_1 U22311 ( .A(n17480), .B(n17761), .Y(n18351) );
  sky130_fd_sc_hd__nand2b_1 U22312 ( .A_N(n17420), .B(n17676), .Y(n18396) );
  sky130_fd_sc_hd__nor4_1 U22313 ( .A(n17783), .B(n17677), .C(n18351), .D(
        n18396), .Y(n17423) );
  sky130_fd_sc_hd__nand3b_1 U22314 ( .A_N(n17552), .B(n18402), .C(n17528), .Y(
        n17421) );
  sky130_fd_sc_hd__nor3_1 U22315 ( .A(n18354), .B(n17508), .C(n17421), .Y(
        n17422) );
  sky130_fd_sc_hd__o22ai_1 U22316 ( .A1(n17423), .A2(n18439), .B1(n17422), 
        .B2(n18445), .Y(n17424) );
  sky130_fd_sc_hd__nor3_1 U22317 ( .A(n17426), .B(n17425), .C(n17424), .Y(
        n17431) );
  sky130_fd_sc_hd__a22oi_1 U22318 ( .A1(n17715), .A2(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[1]), .B1(j202_soc_core_bldc_core_00_comm[1]), .B2(n17427), .Y(n17428) );
  sky130_fd_sc_hd__o21ai_1 U22319 ( .A1(n18282), .A2(n25156), .B1(n17428), .Y(
        n17429) );
  sky130_fd_sc_hd__a31oi_1 U22320 ( .A1(n20430), .A2(
        j202_soc_core_bldc_core_00_adc_en), .A3(n17711), .B1(n17429), .Y(
        n17430) );
  sky130_fd_sc_hd__o22ai_1 U22321 ( .A1(n17431), .A2(n18666), .B1(n17430), 
        .B2(n17717), .Y(n17494) );
  sky130_fd_sc_hd__nand2_1 U22322 ( .A(
        j202_soc_core_ahblite_interconnect_s_hrdata[1]), .B(n18725), .Y(n17437) );
  sky130_fd_sc_hd__a22oi_1 U22323 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[65]), .B1(n18724), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[97]), .Y(n17436) );
  sky130_fd_sc_hd__a22oi_1 U22324 ( .A1(n18241), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[25]), .B1(n18243), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[1]), .Y(n17433) );
  sky130_fd_sc_hd__a22oi_1 U22325 ( .A1(n18242), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[9]), .B1(n18244), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[17]), .Y(n17432) );
  sky130_fd_sc_hd__a21oi_1 U22326 ( .A1(n17433), .A2(n17432), .B1(n18245), .Y(
        n17434) );
  sky130_fd_sc_hd__a21oi_1 U22327 ( .A1(n18726), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[33]), .B1(n17434), .Y(
        n17435) );
  sky130_fd_sc_hd__nand3_1 U22328 ( .A(n17437), .B(n17436), .C(n17435), .Y(
        n17493) );
  sky130_fd_sc_hd__nand3_1 U22329 ( .A(n17672), .B(n17863), .C(n17791), .Y(
        n17531) );
  sky130_fd_sc_hd__nand2_1 U22330 ( .A(n17470), .B(n18430), .Y(n17559) );
  sky130_fd_sc_hd__nand2_1 U22331 ( .A(n17618), .B(n18346), .Y(n17939) );
  sky130_fd_sc_hd__nor4_1 U22332 ( .A(n17531), .B(n18434), .C(n17559), .D(
        n17939), .Y(n17438) );
  sky130_fd_sc_hd__nand2_1 U22333 ( .A(n17923), .B(n17596), .Y(n17748) );
  sky130_fd_sc_hd__a31oi_1 U22334 ( .A1(n17438), .A2(n17937), .A3(n18399), 
        .B1(n18437), .Y(n17450) );
  sky130_fd_sc_hd__nand2_1 U22335 ( .A(n17554), .B(n17756), .Y(n18412) );
  sky130_fd_sc_hd__nand2_1 U22336 ( .A(n17654), .B(n17771), .Y(n17720) );
  sky130_fd_sc_hd__nor4_1 U22337 ( .A(n18354), .B(n17944), .C(n18412), .D(
        n17720), .Y(n17439) );
  sky130_fd_sc_hd__a31oi_1 U22338 ( .A1(n17440), .A2(n17750), .A3(n17439), 
        .B1(n18439), .Y(n17449) );
  sky130_fd_sc_hd__nor2_1 U22339 ( .A(n17442), .B(n17441), .Y(n17929) );
  sky130_fd_sc_hd__nand4_1 U22340 ( .A(n17618), .B(n17676), .C(n17548), .D(
        n18346), .Y(n17745) );
  sky130_fd_sc_hd__nor2_1 U22341 ( .A(n17745), .B(n17526), .Y(n17736) );
  sky130_fd_sc_hd__nand2_1 U22342 ( .A(n17736), .B(n17675), .Y(n17726) );
  sky130_fd_sc_hd__nor4_1 U22343 ( .A(n17929), .B(n17726), .C(n17444), .D(
        n17443), .Y(n17447) );
  sky130_fd_sc_hd__nor4bb_1 U22344 ( .C_N(n17445), .D_N(n17756), .A(n17509), 
        .B(n17915), .Y(n17484) );
  sky130_fd_sc_hd__nand2_1 U22345 ( .A(n17724), .B(n17875), .Y(n17511) );
  sky130_fd_sc_hd__nor4b_1 U22346 ( .D_N(n17484), .A(n18397), .B(n17530), .C(
        n17511), .Y(n17446) );
  sky130_fd_sc_hd__o22ai_1 U22347 ( .A1(n17447), .A2(n18445), .B1(n17446), 
        .B2(n18423), .Y(n17448) );
  sky130_fd_sc_hd__nor3_1 U22348 ( .A(n17450), .B(n17449), .C(n17448), .Y(
        n17466) );
  sky130_fd_sc_hd__a22o_1 U22349 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[1]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[65]), .X(n17451) );
  sky130_fd_sc_hd__a21oi_1 U22350 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[97]), .B1(n17451), .Y(n17453) );
  sky130_fd_sc_hd__a22oi_1 U22351 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[161]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[129]), .Y(n17452) );
  sky130_fd_sc_hd__a21oi_1 U22352 ( .A1(n17453), .A2(n17452), .B1(n18736), .Y(
        n17464) );
  sky130_fd_sc_hd__a22oi_1 U22353 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[257]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[33]), .Y(n17462) );
  sky130_fd_sc_hd__a22o_1 U22354 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[289]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[321]), .X(n17454) );
  sky130_fd_sc_hd__a21oi_1 U22355 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[353]), .B1(n17454), .Y(n17461) );
  sky130_fd_sc_hd__nand2_1 U22356 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[225]), .Y(n17458) );
  sky130_fd_sc_hd__a21oi_1 U22357 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[449]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n17457) );
  sky130_fd_sc_hd__nand2_1 U22358 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[385]), .Y(n17456) );
  sky130_fd_sc_hd__nand2_1 U22359 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[417]), .Y(n17455) );
  sky130_fd_sc_hd__nand4_1 U22360 ( .A(n17458), .B(n17457), .C(n17456), .D(
        n17455), .Y(n17459) );
  sky130_fd_sc_hd__a21oi_1 U22361 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[193]), .B1(n17459), .Y(n17460) );
  sky130_fd_sc_hd__nand3_1 U22362 ( .A(n17462), .B(n17461), .C(n17460), .Y(
        n17463) );
  sky130_fd_sc_hd__o22ai_1 U22363 ( .A1(j202_soc_core_memory0_ram_dout0[481]), 
        .A2(n18758), .B1(n17464), .B2(n17463), .Y(n17465) );
  sky130_fd_sc_hd__o22ai_1 U22364 ( .A1(n17466), .A2(n18722), .B1(n18761), 
        .B2(n17465), .Y(n17492) );
  sky130_fd_sc_hd__nand2_1 U22365 ( .A(n17876), .B(n17678), .Y(n17721) );
  sky130_fd_sc_hd__nor2_1 U22366 ( .A(n17721), .B(n17745), .Y(n17513) );
  sky130_fd_sc_hd__nor3_1 U22367 ( .A(n17945), .B(n17916), .C(n17531), .Y(
        n17729) );
  sky130_fd_sc_hd__nor4_1 U22368 ( .A(n17600), .B(n17737), .C(n18397), .D(
        n17516), .Y(n17467) );
  sky130_fd_sc_hd__a31oi_1 U22369 ( .A1(n17513), .A2(n17729), .A3(n17467), 
        .B1(n18439), .Y(n17477) );
  sky130_fd_sc_hd__nor2_1 U22370 ( .A(n17721), .B(n17943), .Y(n17780) );
  sky130_fd_sc_hd__nand3_1 U22371 ( .A(n17469), .B(
        j202_soc_core_bootrom_00_address_w[10]), .C(n17468), .Y(n17850) );
  sky130_fd_sc_hd__nand4_1 U22372 ( .A(n17672), .B(n17653), .C(n17850), .D(
        n18345), .Y(n17782) );
  sky130_fd_sc_hd__nor2_1 U22373 ( .A(n17746), .B(n17782), .Y(n17776) );
  sky130_fd_sc_hd__nand2_1 U22374 ( .A(n17470), .B(n17868), .Y(n17794) );
  sky130_fd_sc_hd__nor3_1 U22375 ( .A(n17794), .B(n17549), .C(n17529), .Y(
        n17471) );
  sky130_fd_sc_hd__a31oi_1 U22376 ( .A1(n17780), .A2(n17776), .A3(n17471), 
        .B1(n18445), .Y(n17476) );
  sky130_fd_sc_hd__nor4_1 U22377 ( .A(n18392), .B(n17600), .C(n17783), .D(
        n17794), .Y(n17474) );
  sky130_fd_sc_hd__nor4_1 U22378 ( .A(n18444), .B(n17748), .C(n17472), .D(
        n17517), .Y(n17473) );
  sky130_fd_sc_hd__o22ai_1 U22379 ( .A1(n17474), .A2(n18423), .B1(n17473), 
        .B2(n18437), .Y(n17475) );
  sky130_fd_sc_hd__nor3_1 U22380 ( .A(n17477), .B(n17476), .C(n17475), .Y(
        n17490) );
  sky130_fd_sc_hd__a31oi_1 U22381 ( .A1(n17480), .A2(n17479), .A3(n17478), 
        .B1(n18423), .Y(n17488) );
  sky130_fd_sc_hd__a31oi_1 U22382 ( .A1(n17802), .A2(n17481), .A3(n17527), 
        .B1(n18445), .Y(n17487) );
  sky130_fd_sc_hd__nor2_1 U22383 ( .A(n17509), .B(n17941), .Y(n17722) );
  sky130_fd_sc_hd__nor4_1 U22384 ( .A(n18354), .B(n17944), .C(n17751), .D(
        n17482), .Y(n17483) );
  sky130_fd_sc_hd__a31oi_1 U22385 ( .A1(n17722), .A2(n17483), .A3(n17676), 
        .B1(n18439), .Y(n17486) );
  sky130_fd_sc_hd__nor2_1 U22386 ( .A(n17737), .B(n17847), .Y(n18429) );
  sky130_fd_sc_hd__a31oi_1 U22387 ( .A1(n17735), .A2(n18429), .A3(n17484), 
        .B1(n18437), .Y(n17485) );
  sky130_fd_sc_hd__nor4_1 U22388 ( .A(n17488), .B(n17487), .C(n17486), .D(
        n17485), .Y(n17489) );
  sky130_fd_sc_hd__o22ai_1 U22389 ( .A1(n17490), .A2(n18720), .B1(n17489), 
        .B2(n18552), .Y(n17491) );
  sky130_fd_sc_hd__nor2_1 U22390 ( .A(n17915), .B(n17619), .Y(n17497) );
  sky130_fd_sc_hd__nor2_1 U22391 ( .A(n18398), .B(n18354), .Y(n17938) );
  sky130_fd_sc_hd__nor4_1 U22392 ( .A(n17941), .B(n17746), .C(n17508), .D(
        n17495), .Y(n17496) );
  sky130_fd_sc_hd__a31oi_1 U22393 ( .A1(n17497), .A2(n17938), .A3(n17496), 
        .B1(n18423), .Y(n17506) );
  sky130_fd_sc_hd__nor4_1 U22394 ( .A(n17498), .B(n17509), .C(n17621), .D(
        n17531), .Y(n17499) );
  sky130_fd_sc_hd__a21oi_1 U22395 ( .A1(n17770), .A2(n17499), .B1(n18437), .Y(
        n17505) );
  sky130_fd_sc_hd__nor2_1 U22396 ( .A(n18397), .B(n17611), .Y(n17551) );
  sky130_fd_sc_hd__nor2_1 U22397 ( .A(n17910), .B(n17662), .Y(n17925) );
  sky130_fd_sc_hd__nor3b_1 U22398 ( .C_N(n17925), .A(n18412), .B(n18390), .Y(
        n17798) );
  sky130_fd_sc_hd__a31oi_1 U22399 ( .A1(n17551), .A2(n17500), .A3(n17798), 
        .B1(n18439), .Y(n17504) );
  sky130_fd_sc_hd__nor4_1 U22400 ( .A(n18354), .B(n17624), .C(n17556), .D(
        n17661), .Y(n17501) );
  sky130_fd_sc_hd__a31oi_1 U22401 ( .A1(n17502), .A2(n17501), .A3(n17771), 
        .B1(n18445), .Y(n17503) );
  sky130_fd_sc_hd__nor4_1 U22402 ( .A(n17506), .B(n17505), .C(n17504), .D(
        n17503), .Y(n17507) );
  sky130_fd_sc_hd__nor2_1 U22403 ( .A(n17507), .B(n18552), .Y(n17547) );
  sky130_fd_sc_hd__nor2_1 U22404 ( .A(n17945), .B(n17916), .Y(n17510) );
  sky130_fd_sc_hd__nor2_1 U22405 ( .A(n17509), .B(n17508), .Y(n17914) );
  sky130_fd_sc_hd__nand2_1 U22406 ( .A(n18399), .B(n17914), .Y(n17805) );
  sky130_fd_sc_hd__a31oi_1 U22407 ( .A1(n17527), .A2(n17510), .A3(n17801), 
        .B1(n18437), .Y(n17522) );
  sky130_fd_sc_hd__nor3_1 U22408 ( .A(n17945), .B(n18435), .C(n17511), .Y(
        n17512) );
  sky130_fd_sc_hd__a31oi_1 U22409 ( .A1(n17514), .A2(n17513), .A3(n17512), 
        .B1(n18439), .Y(n17521) );
  sky130_fd_sc_hd__nand2_1 U22410 ( .A(n18430), .B(n17875), .Y(n17515) );
  sky130_fd_sc_hd__nor4_1 U22411 ( .A(n17944), .B(n17795), .C(n17516), .D(
        n17515), .Y(n17519) );
  sky130_fd_sc_hd__nand2_1 U22412 ( .A(n17849), .B(n17911), .Y(n17804) );
  sky130_fd_sc_hd__nor3_1 U22413 ( .A(n17517), .B(n17804), .C(n17555), .Y(
        n17518) );
  sky130_fd_sc_hd__o22ai_1 U22414 ( .A1(n17519), .A2(n18423), .B1(n17518), 
        .B2(n18445), .Y(n17520) );
  sky130_fd_sc_hd__nor3_1 U22415 ( .A(n17522), .B(n17521), .C(n17520), .Y(
        n17545) );
  sky130_fd_sc_hd__nand4_1 U22416 ( .A(n17801), .B(n17525), .C(n17524), .D(
        n17523), .Y(n17542) );
  sky130_fd_sc_hd__nor2_1 U22417 ( .A(n17860), .B(n17526), .Y(n17800) );
  sky130_fd_sc_hd__a31oi_1 U22418 ( .A1(n17528), .A2(n17527), .A3(n17800), 
        .B1(n18439), .Y(n17541) );
  sky130_fd_sc_hd__nor4b_1 U22419 ( .D_N(n17729), .A(n17624), .B(n17529), .C(
        n17852), .Y(n17539) );
  sky130_fd_sc_hd__nor3_1 U22420 ( .A(n17944), .B(n17531), .C(n17530), .Y(
        n17535) );
  sky130_fd_sc_hd__nand2_1 U22421 ( .A(n17533), .B(n17532), .Y(n18413) );
  sky130_fd_sc_hd__nand3_1 U22422 ( .A(n17535), .B(n17534), .C(n18413), .Y(
        n17732) );
  sky130_fd_sc_hd__nor4_1 U22423 ( .A(n18397), .B(n17537), .C(n17536), .D(
        n17732), .Y(n17538) );
  sky130_fd_sc_hd__o22ai_1 U22424 ( .A1(n17539), .A2(n18423), .B1(n17538), 
        .B2(n18445), .Y(n17540) );
  sky130_fd_sc_hd__a211oi_1 U22425 ( .A1(n17543), .A2(n17542), .B1(n17541), 
        .C1(n17540), .Y(n17544) );
  sky130_fd_sc_hd__o22ai_1 U22426 ( .A1(n17545), .A2(n18666), .B1(n17544), 
        .B2(n18722), .Y(n17546) );
  sky130_fd_sc_hd__a211oi_1 U22427 ( .A1(
        j202_soc_core_bldc_core_00_pwm_period[3]), .A2(n18629), .B1(n17547), 
        .C1(n17546), .Y(n17589) );
  sky130_fd_sc_hd__nand2_1 U22428 ( .A(n17925), .B(n17548), .Y(n18405) );
  sky130_fd_sc_hd__nor4_1 U22429 ( .A(n17784), .B(n17782), .C(n17549), .D(
        n18405), .Y(n17550) );
  sky130_fd_sc_hd__a31oi_1 U22430 ( .A1(n17914), .A2(n17550), .A3(n17757), 
        .B1(n18439), .Y(n17564) );
  sky130_fd_sc_hd__nor4_1 U22431 ( .A(n18354), .B(n17552), .C(n17939), .D(
        n17747), .Y(n17553) );
  sky130_fd_sc_hd__a31oi_1 U22432 ( .A1(n17761), .A2(n17557), .A3(n17553), 
        .B1(n18445), .Y(n17563) );
  sky130_fd_sc_hd__nand3_1 U22433 ( .A(n17554), .B(n18347), .C(n18341), .Y(
        n17719) );
  sky130_fd_sc_hd__nand2_1 U22434 ( .A(n17868), .B(n17875), .Y(n17755) );
  sky130_fd_sc_hd__nor4_1 U22435 ( .A(n17719), .B(n17755), .C(n17556), .D(
        n17555), .Y(n17561) );
  sky130_fd_sc_hd__nand2_1 U22436 ( .A(n17557), .B(n17761), .Y(n17558) );
  sky130_fd_sc_hd__nor4_1 U22437 ( .A(n17604), .B(n17751), .C(n17559), .D(
        n17558), .Y(n17560) );
  sky130_fd_sc_hd__o22ai_1 U22438 ( .A1(n17561), .A2(n18437), .B1(n17560), 
        .B2(n18423), .Y(n17562) );
  sky130_fd_sc_hd__o31a_1 U22439 ( .A1(n17564), .A2(n17563), .A3(n17562), .B1(
        n17609), .X(n17587) );
  sky130_fd_sc_hd__a22oi_1 U22440 ( .A1(n18244), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[19]), .B1(n18241), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[27]), .Y(n17566) );
  sky130_fd_sc_hd__a22oi_1 U22441 ( .A1(n18242), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[11]), .B1(n18243), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[3]), .Y(n17565) );
  sky130_fd_sc_hd__a21oi_1 U22442 ( .A1(n17566), .A2(n17565), .B1(n18245), .Y(
        n17568) );
  sky130_fd_sc_hd__a22oi_1 U22443 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[3]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[35]), .Y(n17567) );
  sky130_fd_sc_hd__nand2b_1 U22444 ( .A_N(n17568), .B(n17567), .Y(n17586) );
  sky130_fd_sc_hd__a22o_1 U22445 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[3]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[67]), .X(n17569) );
  sky130_fd_sc_hd__a21oi_1 U22446 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[99]), .B1(n17569), .Y(n17571) );
  sky130_fd_sc_hd__a22oi_1 U22447 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[163]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[131]), .Y(n17570) );
  sky130_fd_sc_hd__a21oi_1 U22448 ( .A1(n17571), .A2(n17570), .B1(n18736), .Y(
        n17582) );
  sky130_fd_sc_hd__a22oi_1 U22449 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[259]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[35]), .Y(n17580) );
  sky130_fd_sc_hd__a22o_1 U22450 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[291]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[323]), .X(n17572) );
  sky130_fd_sc_hd__a21oi_1 U22451 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[355]), .B1(n17572), .Y(n17579) );
  sky130_fd_sc_hd__nand2_1 U22452 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[227]), .Y(n17576) );
  sky130_fd_sc_hd__a21oi_1 U22453 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[451]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n17575) );
  sky130_fd_sc_hd__nand2_1 U22454 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[387]), .Y(n17574) );
  sky130_fd_sc_hd__nand2_1 U22455 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[419]), .Y(n17573) );
  sky130_fd_sc_hd__nand4_1 U22456 ( .A(n17576), .B(n17575), .C(n17574), .D(
        n17573), .Y(n17577) );
  sky130_fd_sc_hd__a21oi_1 U22457 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[195]), .B1(n17577), .Y(n17578) );
  sky130_fd_sc_hd__nand3_1 U22458 ( .A(n17580), .B(n17579), .C(n17578), .Y(
        n17581) );
  sky130_fd_sc_hd__o22ai_1 U22459 ( .A1(j202_soc_core_memory0_ram_dout0[483]), 
        .A2(n18758), .B1(n17582), .B2(n17581), .Y(n17584) );
  sky130_fd_sc_hd__a22oi_1 U22460 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[67]), .B1(n18724), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[99]), .Y(n17583) );
  sky130_fd_sc_hd__nor3_1 U22462 ( .A(n17587), .B(n17586), .C(n17585), .Y(
        n17588) );
  sky130_fd_sc_hd__nand2_1 U22463 ( .A(n17589), .B(n17588), .Y(n25253) );
  sky130_fd_sc_hd__nand2_1 U22464 ( .A(n17722), .B(n17791), .Y(n18433) );
  sky130_fd_sc_hd__a31oi_1 U22465 ( .A1(n17591), .A2(n17590), .A3(n17674), 
        .B1(n18445), .Y(n18359) );
  sky130_fd_sc_hd__nor2_1 U22466 ( .A(n17593), .B(n17592), .Y(n17594) );
  sky130_fd_sc_hd__a31oi_1 U22467 ( .A1(n17595), .A2(n17938), .A3(n17594), 
        .B1(n18439), .Y(n17603) );
  sky130_fd_sc_hd__nand2_1 U22468 ( .A(n17596), .B(n17617), .Y(n17927) );
  sky130_fd_sc_hd__nand2_1 U22469 ( .A(n17912), .B(n17850), .Y(n17862) );
  sky130_fd_sc_hd__nor3_1 U22470 ( .A(n17927), .B(n17862), .C(n17597), .Y(
        n17598) );
  sky130_fd_sc_hd__a21oi_1 U22471 ( .A1(n17599), .A2(n17598), .B1(n18437), .Y(
        n17602) );
  sky130_fd_sc_hd__nor3_1 U22472 ( .A(n17600), .B(n18397), .C(n18441), .Y(
        n17664) );
  sky130_fd_sc_hd__a31oi_1 U22473 ( .A1(n17876), .A2(n17664), .A3(n17672), 
        .B1(n18445), .Y(n17601) );
  sky130_fd_sc_hd__nor4_1 U22474 ( .A(n18359), .B(n17603), .C(n17602), .D(
        n17601), .Y(n17608) );
  sky130_fd_sc_hd__nor2_1 U22475 ( .A(n17604), .B(n17619), .Y(n17792) );
  sky130_fd_sc_hd__nand4b_1 U22476 ( .A_N(n17605), .B(n17792), .C(n18347), .D(
        n18345), .Y(n17673) );
  sky130_fd_sc_hd__nor2_1 U22477 ( .A(n18395), .B(n17673), .Y(n17679) );
  sky130_fd_sc_hd__nand2b_1 U22478 ( .A_N(n17842), .B(n17679), .Y(n17873) );
  sky130_fd_sc_hd__o31ai_1 U22479 ( .A1(n18349), .A2(n17852), .A3(n17873), 
        .B1(n17606), .Y(n17607) );
  sky130_fd_sc_hd__nand2_1 U22480 ( .A(n17608), .B(n17607), .Y(n17610) );
  sky130_fd_sc_hd__nand2_1 U22481 ( .A(n17610), .B(n17609), .Y(n17690) );
  sky130_fd_sc_hd__nor4_1 U22482 ( .A(n17860), .B(n17737), .C(n17746), .D(
        n17611), .Y(n17612) );
  sky130_fd_sc_hd__a21oi_1 U22483 ( .A1(n17613), .A2(n17612), .B1(n18423), .Y(
        n18422) );
  sky130_fd_sc_hd__a21oi_1 U22484 ( .A1(n17615), .A2(n17614), .B1(n18437), .Y(
        n17629) );
  sky130_fd_sc_hd__o31a_1 U22485 ( .A1(n17910), .A2(n17616), .A3(n17927), .B1(
        n17812), .X(n17628) );
  sky130_fd_sc_hd__nand2_1 U22486 ( .A(n17849), .B(n17676), .Y(n17903) );
  sky130_fd_sc_hd__nand2_1 U22487 ( .A(n17618), .B(n17617), .Y(n17909) );
  sky130_fd_sc_hd__nor4_1 U22488 ( .A(n17915), .B(n17619), .C(n17903), .D(
        n17909), .Y(n17626) );
  sky130_fd_sc_hd__nand2_1 U22489 ( .A(n17756), .B(n17620), .Y(n17934) );
  sky130_fd_sc_hd__nor2_1 U22490 ( .A(n17621), .B(n18397), .Y(n17874) );
  sky130_fd_sc_hd__nand4b_1 U22491 ( .A_N(n17934), .B(n17623), .C(n17622), .D(
        n17874), .Y(n18417) );
  sky130_fd_sc_hd__nor4_1 U22492 ( .A(n18392), .B(n17916), .C(n17624), .D(
        n18417), .Y(n17625) );
  sky130_fd_sc_hd__o22ai_1 U22493 ( .A1(n17626), .A2(n18423), .B1(n17625), 
        .B2(n18439), .Y(n17627) );
  sky130_fd_sc_hd__nor4_1 U22494 ( .A(n18422), .B(n17629), .C(n17628), .D(
        n17627), .Y(n17652) );
  sky130_fd_sc_hd__a22oi_1 U22495 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[267]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[43]), .Y(n17644) );
  sky130_fd_sc_hd__a22o_1 U22496 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[299]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[331]), .X(n17630) );
  sky130_fd_sc_hd__a21oi_1 U22497 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[363]), .B1(n17630), .Y(n17643) );
  sky130_fd_sc_hd__nand2_1 U22498 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[235]), .Y(n17634) );
  sky130_fd_sc_hd__a21oi_1 U22499 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[459]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n17633) );
  sky130_fd_sc_hd__nand2_1 U22500 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[395]), .Y(n17632) );
  sky130_fd_sc_hd__nand2_1 U22501 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[427]), .Y(n17631) );
  sky130_fd_sc_hd__nand4_1 U22502 ( .A(n17634), .B(n17633), .C(n17632), .D(
        n17631), .Y(n17635) );
  sky130_fd_sc_hd__a21oi_1 U22503 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[203]), .B1(n17635), .Y(n17642) );
  sky130_fd_sc_hd__a22o_1 U22504 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[11]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[75]), .X(n17636) );
  sky130_fd_sc_hd__a21oi_1 U22505 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[107]), .B1(n17636), .Y(n17638) );
  sky130_fd_sc_hd__a22oi_1 U22506 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[171]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[139]), .Y(n17637) );
  sky130_fd_sc_hd__nand2_1 U22507 ( .A(n17638), .B(n17637), .Y(n17640) );
  sky130_fd_sc_hd__nand2_1 U22508 ( .A(n17640), .B(n17639), .Y(n17641) );
  sky130_fd_sc_hd__nand4_1 U22509 ( .A(n17644), .B(n17643), .C(n17642), .D(
        n17641), .Y(n17650) );
  sky130_fd_sc_hd__nor2_1 U22510 ( .A(j202_soc_core_memory0_ram_dout0[491]), 
        .B(n18758), .Y(n17645) );
  sky130_fd_sc_hd__nor2_1 U22511 ( .A(n17645), .B(n18761), .Y(n17649) );
  sky130_fd_sc_hd__a22oi_1 U22512 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[11]), .B1(n18724), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[107]), .Y(n17647) );
  sky130_fd_sc_hd__a22oi_1 U22513 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[75]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[43]), .Y(n17646) );
  sky130_fd_sc_hd__o211ai_1 U22514 ( .A1(n18759), .A2(n25184), .B1(n17647), 
        .C1(n17646), .Y(n17648) );
  sky130_fd_sc_hd__a21oi_1 U22515 ( .A1(n17650), .A2(n17649), .B1(n17648), .Y(
        n17651) );
  sky130_fd_sc_hd__o21a_1 U22516 ( .A1(n18722), .A2(n17652), .B1(n17651), .X(
        n17689) );
  sky130_fd_sc_hd__and3_1 U22517 ( .A(n17653), .B(n18446), .C(n17938), .X(
        n17655) );
  sky130_fd_sc_hd__a31oi_1 U22518 ( .A1(n17654), .A2(n17937), .A3(n17655), 
        .B1(n18423), .Y(n17668) );
  sky130_fd_sc_hd__a31oi_1 U22519 ( .A1(n17656), .A2(n17722), .A3(n17655), 
        .B1(n18437), .Y(n17667) );
  sky130_fd_sc_hd__nor2_1 U22520 ( .A(n18398), .B(n18386), .Y(n17659) );
  sky130_fd_sc_hd__a31oi_1 U22521 ( .A1(n17659), .A2(n17658), .A3(n17657), 
        .B1(n18439), .Y(n17666) );
  sky130_fd_sc_hd__nor4_1 U22522 ( .A(n17662), .B(n18444), .C(n17661), .D(
        n17660), .Y(n17663) );
  sky130_fd_sc_hd__a21oi_1 U22523 ( .A1(n17664), .A2(n17663), .B1(n18445), .Y(
        n17665) );
  sky130_fd_sc_hd__nor4_1 U22524 ( .A(n17668), .B(n17667), .C(n17666), .D(
        n17665), .Y(n17687) );
  sky130_fd_sc_hd__nor4_1 U22525 ( .A(n17746), .B(n17670), .C(n17669), .D(
        n18441), .Y(n17671) );
  sky130_fd_sc_hd__a31oi_1 U22526 ( .A1(n18430), .A2(n17671), .A3(n17768), 
        .B1(n18445), .Y(n17685) );
  sky130_fd_sc_hd__nor3_1 U22527 ( .A(n17935), .B(n18390), .C(n17673), .Y(
        n17853) );
  sky130_fd_sc_hd__a31oi_1 U22528 ( .A1(n17853), .A2(n17674), .A3(n17911), 
        .B1(n18423), .Y(n17684) );
  sky130_fd_sc_hd__nand3_1 U22529 ( .A(n17912), .B(n17676), .C(n17675), .Y(
        n18432) );
  sky130_fd_sc_hd__nor3_1 U22530 ( .A(n17677), .B(n18442), .C(n18432), .Y(
        n17682) );
  sky130_fd_sc_hd__nand3_1 U22531 ( .A(n17679), .B(n17678), .C(n17875), .Y(
        n17680) );
  sky130_fd_sc_hd__nor4_1 U22532 ( .A(n17943), .B(n17939), .C(n17927), .D(
        n17680), .Y(n17681) );
  sky130_fd_sc_hd__o22ai_1 U22533 ( .A1(n17682), .A2(n18439), .B1(n17681), 
        .B2(n18437), .Y(n17683) );
  sky130_fd_sc_hd__nor3_1 U22534 ( .A(n17685), .B(n17684), .C(n17683), .Y(
        n17686) );
  sky130_fd_sc_hd__o22a_1 U22535 ( .A1(n18552), .A2(n17687), .B1(n18666), .B2(
        n17686), .X(n17688) );
  sky130_fd_sc_hd__nand3_1 U22536 ( .A(n17690), .B(n17689), .C(n17688), .Y(
        n25311) );
  sky130_fd_sc_hd__a22oi_1 U22537 ( .A1(n18244), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[16]), .B1(n18243), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[0]), .Y(n17692) );
  sky130_fd_sc_hd__a22oi_1 U22538 ( .A1(n18242), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[8]), .B1(n18241), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[24]), .Y(n17691) );
  sky130_fd_sc_hd__a21oi_1 U22539 ( .A1(n17692), .A2(n17691), .B1(n18245), .Y(
        n17693) );
  sky130_fd_sc_hd__a21oi_1 U22540 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[0]), .B1(n17693), .Y(
        n17821) );
  sky130_fd_sc_hd__a22oi_1 U22541 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[64]), .B1(n18724), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[96]), .Y(n17820) );
  sky130_fd_sc_hd__a22oi_1 U22542 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[224]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[192]), .Y(n17697) );
  sky130_fd_sc_hd__a22oi_1 U22543 ( .A1(n18734), .A2(
        j202_soc_core_memory0_ram_dout0[128]), .B1(n18733), .B2(
        j202_soc_core_memory0_ram_dout0[96]), .Y(n17696) );
  sky130_fd_sc_hd__a22oi_1 U22544 ( .A1(n18361), .A2(
        j202_soc_core_memory0_ram_dout0[32]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[64]), .Y(n17695) );
  sky130_fd_sc_hd__nand2_1 U22545 ( .A(n18735), .B(
        j202_soc_core_memory0_ram_dout0[160]), .Y(n17694) );
  sky130_fd_sc_hd__nand4_1 U22546 ( .A(n17697), .B(n17696), .C(n17695), .D(
        n17694), .Y(n17698) );
  sky130_fd_sc_hd__a21oi_1 U22547 ( .A1(n18367), .A2(
        j202_soc_core_memory0_ram_dout0[0]), .B1(n17698), .Y(n17706) );
  sky130_fd_sc_hd__a22oi_1 U22548 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[288]), .B1(n18062), .B2(
        j202_soc_core_memory0_ram_dout0[256]), .Y(n17705) );
  sky130_fd_sc_hd__nand2_1 U22549 ( .A(n18743), .B(
        j202_soc_core_memory0_ram_dout0[352]), .Y(n17702) );
  sky130_fd_sc_hd__a21oi_1 U22550 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[448]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n17701) );
  sky130_fd_sc_hd__nand2_1 U22551 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[384]), .Y(n17700) );
  sky130_fd_sc_hd__nand2_1 U22552 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[416]), .Y(n17699) );
  sky130_fd_sc_hd__nand4_1 U22553 ( .A(n17702), .B(n17701), .C(n17700), .D(
        n17699), .Y(n17703) );
  sky130_fd_sc_hd__a21oi_1 U22554 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[320]), .B1(n17703), .Y(n17704) );
  sky130_fd_sc_hd__o211ai_1 U22555 ( .A1(n18736), .A2(n17706), .B1(n17705), 
        .C1(n17704), .Y(n17707) );
  sky130_fd_sc_hd__a2bb2oi_1 U22557 ( .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[32]), .A1_N(n18761), 
        .A2_N(n17708), .Y(n17819) );
  sky130_fd_sc_hd__nand2b_1 U22558 ( .A_N(n17710), .B(n17709), .Y(n19741) );
  sky130_fd_sc_hd__nor2b_1 U22559 ( .B_N(n19742), .A(n19741), .Y(n25165) );
  sky130_fd_sc_hd__a222oi_1 U22560 ( .A1(n20430), .A2(
        j202_soc_core_bldc_core_00_pwm_en), .B1(n25159), .B2(
        j202_soc_core_bldc_core_00_comm[0]), .C1(n25165), .C2(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_), .Y(n17713) );
  sky130_fd_sc_hd__o22ai_1 U22561 ( .A1(n17713), .A2(n17712), .B1(n18282), 
        .B2(n25172), .Y(n17714) );
  sky130_fd_sc_hd__a21oi_1 U22562 ( .A1(n17715), .A2(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_hsvr_00_latch_status[0]), .B1(n17714), .Y(n17718) );
  sky130_fd_sc_hd__nand3_1 U22563 ( .A(n17716), .B(n25165), .C(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_0_), .Y(n23809) );
  sky130_fd_sc_hd__a21oi_1 U22564 ( .A1(n17718), .A2(n23809), .B1(n17717), .Y(
        n17817) );
  sky130_fd_sc_hd__nor4b_1 U22565 ( .D_N(n17722), .A(n17721), .B(n17720), .C(
        n17719), .Y(n17723) );
  sky130_fd_sc_hd__a21oi_1 U22566 ( .A1(n17724), .A2(n17723), .B1(n18439), .Y(
        n17743) );
  sky130_fd_sc_hd__nor4_1 U22567 ( .A(n17727), .B(n18435), .C(n17726), .D(
        n17725), .Y(n17728) );
  sky130_fd_sc_hd__a31oi_1 U22568 ( .A1(n17914), .A2(n17729), .A3(n17728), 
        .B1(n18423), .Y(n17742) );
  sky130_fd_sc_hd__nor2_1 U22569 ( .A(n17731), .B(n17730), .Y(n17733) );
  sky130_fd_sc_hd__nor3_1 U22570 ( .A(n17860), .B(n17733), .C(n17732), .Y(
        n17734) );
  sky130_fd_sc_hd__a31oi_1 U22571 ( .A1(n17736), .A2(n17735), .A3(n17734), 
        .B1(n18445), .Y(n17741) );
  sky130_fd_sc_hd__nor4_1 U22572 ( .A(n17737), .B(n18434), .C(n17927), .D(
        n18386), .Y(n17738) );
  sky130_fd_sc_hd__a31oi_1 U22573 ( .A1(n17739), .A2(n17776), .A3(n17738), 
        .B1(n18437), .Y(n17740) );
  sky130_fd_sc_hd__nor4_1 U22574 ( .A(n17743), .B(n17742), .C(n17741), .D(
        n17740), .Y(n17767) );
  sky130_fd_sc_hd__nor3_1 U22575 ( .A(n17746), .B(n17745), .C(n17744), .Y(
        n17797) );
  sky130_fd_sc_hd__nor2_1 U22576 ( .A(n17748), .B(n17747), .Y(n17749) );
  sky130_fd_sc_hd__a31oi_1 U22577 ( .A1(n17797), .A2(n17750), .A3(n17749), 
        .B1(n18439), .Y(n17765) );
  sky130_fd_sc_hd__nor3_1 U22578 ( .A(n17752), .B(n17944), .C(n17751), .Y(
        n17753) );
  sky130_fd_sc_hd__a31oi_1 U22579 ( .A1(n17754), .A2(n18402), .A3(n17753), 
        .B1(n18445), .Y(n17764) );
  sky130_fd_sc_hd__nor4_1 U22580 ( .A(n17910), .B(n17795), .C(n17944), .D(
        n17755), .Y(n17758) );
  sky130_fd_sc_hd__a31oi_1 U22581 ( .A1(n17758), .A2(n17757), .A3(n17756), 
        .B1(n18423), .Y(n17763) );
  sky130_fd_sc_hd__nor3b_1 U22582 ( .C_N(n17907), .A(n17794), .B(n17759), .Y(
        n17760) );
  sky130_fd_sc_hd__a31oi_1 U22583 ( .A1(n17793), .A2(n17761), .A3(n17760), 
        .B1(n18437), .Y(n17762) );
  sky130_fd_sc_hd__nor4_1 U22584 ( .A(n17765), .B(n17764), .C(n17763), .D(
        n17762), .Y(n17766) );
  sky130_fd_sc_hd__o22ai_1 U22585 ( .A1(n17767), .A2(n18722), .B1(n17766), 
        .B2(n18666), .Y(n17816) );
  sky130_fd_sc_hd__a31oi_1 U22586 ( .A1(n17770), .A2(n17769), .A3(n17768), 
        .B1(n18437), .Y(n17790) );
  sky130_fd_sc_hd__nand2_1 U22587 ( .A(n17923), .B(n17771), .Y(n17772) );
  sky130_fd_sc_hd__nor4_1 U22588 ( .A(n17774), .B(n17773), .C(n17772), .D(
        n18391), .Y(n17775) );
  sky130_fd_sc_hd__a21oi_1 U22589 ( .A1(n17776), .A2(n17775), .B1(n18445), .Y(
        n17789) );
  sky130_fd_sc_hd__nand2b_1 U22590 ( .A_N(n17778), .B(n17777), .Y(n18344) );
  sky130_fd_sc_hd__nand3_1 U22591 ( .A(n17780), .B(n17914), .C(n17779), .Y(
        n17781) );
  sky130_fd_sc_hd__nor4b_1 U22592 ( .D_N(n18344), .A(n17784), .B(n17782), .C(
        n17781), .Y(n17787) );
  sky130_fd_sc_hd__nor4_1 U22593 ( .A(n17785), .B(n17784), .C(n17783), .D(
        n17864), .Y(n17786) );
  sky130_fd_sc_hd__o22ai_1 U22594 ( .A1(n17787), .A2(n18439), .B1(n17786), 
        .B2(n18423), .Y(n17788) );
  sky130_fd_sc_hd__nor3_1 U22595 ( .A(n17790), .B(n17789), .C(n17788), .Y(
        n17814) );
  sky130_fd_sc_hd__nand4_1 U22596 ( .A(n17797), .B(n17793), .C(n17792), .D(
        n17791), .Y(n17811) );
  sky130_fd_sc_hd__nor3_1 U22597 ( .A(n17795), .B(n17794), .C(n18391), .Y(
        n17796) );
  sky130_fd_sc_hd__a31oi_1 U22598 ( .A1(n17798), .A2(n17797), .A3(n17796), 
        .B1(n18437), .Y(n17810) );
  sky130_fd_sc_hd__nand4_1 U22599 ( .A(n17802), .B(n17801), .C(n17800), .D(
        n17799), .Y(n17803) );
  sky130_fd_sc_hd__nor3_1 U22600 ( .A(n18435), .B(n18412), .C(n17803), .Y(
        n17808) );
  sky130_fd_sc_hd__nor4_1 U22601 ( .A(n17806), .B(n17940), .C(n17805), .D(
        n17804), .Y(n17807) );
  sky130_fd_sc_hd__o22ai_1 U22602 ( .A1(n17808), .A2(n18423), .B1(n17807), 
        .B2(n18439), .Y(n17809) );
  sky130_fd_sc_hd__a211oi_1 U22603 ( .A1(n17812), .A2(n17811), .B1(n17810), 
        .C1(n17809), .Y(n17813) );
  sky130_fd_sc_hd__o22ai_1 U22604 ( .A1(n17814), .A2(n18720), .B1(n17813), 
        .B2(n18552), .Y(n17815) );
  sky130_fd_sc_hd__nor3_1 U22605 ( .A(n17817), .B(n17816), .C(n17815), .Y(
        n17818) );
  sky130_fd_sc_hd__nand4_1 U22606 ( .A(n17821), .B(n17820), .C(n17819), .D(
        n17818), .Y(n25259) );
  sky130_fd_sc_hd__nand2_1 U22607 ( .A(n17826), .B(n17825), .Y(n17827) );
  sky130_fd_sc_hd__xor2_1 U22608 ( .A(n17828), .B(n17827), .X(n22750) );
  sky130_fd_sc_hd__nand2_1 U22609 ( .A(n22750), .B(n19729), .Y(n17831) );
  sky130_fd_sc_hd__o22ai_1 U22610 ( .A1(n20805), .A2(n19731), .B1(
        j202_soc_core_j22_cpu_pc[1]), .B2(n19734), .Y(n17829) );
  sky130_fd_sc_hd__a21oi_1 U22611 ( .A1(n19736), .A2(n22183), .B1(n17829), .Y(
        n17830) );
  sky130_fd_sc_hd__nand2_1 U22612 ( .A(n17831), .B(n17830), .Y(n17832) );
  sky130_fd_sc_hd__nand2_1 U22613 ( .A(n17834), .B(n17833), .Y(n17835) );
  sky130_fd_sc_hd__xnor2_1 U22614 ( .A(n17835), .B(n19045), .Y(n22010) );
  sky130_fd_sc_hd__nand2_1 U22615 ( .A(n22010), .B(n19729), .Y(n17841) );
  sky130_fd_sc_hd__o22a_1 U22616 ( .A1(n22711), .A2(n18948), .B1(n22488), .B2(
        n19731), .X(n17838) );
  sky130_fd_sc_hd__ha_1 U22617 ( .A(j202_soc_core_j22_cpu_pc[3]), .B(n17836), 
        .COUT(n19194), .SUM(n22009) );
  sky130_fd_sc_hd__nand2_1 U22618 ( .A(n19661), .B(n22009), .Y(n17837) );
  sky130_fd_sc_hd__o211ai_1 U22619 ( .A1(n22711), .A2(n19083), .B1(n17838), 
        .C1(n17837), .Y(n17839) );
  sky130_fd_sc_hd__a21oi_1 U22620 ( .A1(n25253), .A2(n19737), .B1(n17839), .Y(
        n17840) );
  sky130_fd_sc_hd__nand2_1 U22621 ( .A(n17841), .B(n17840), .Y(n25334) );
  sky130_fd_sc_hd__nor3_1 U22622 ( .A(n17945), .B(n17842), .C(n18435), .Y(
        n18425) );
  sky130_fd_sc_hd__nor4b_1 U22623 ( .D_N(n18425), .A(n18392), .B(n18354), .C(
        n17843), .Y(n17844) );
  sky130_fd_sc_hd__a31oi_1 U22624 ( .A1(n17846), .A2(n17845), .A3(n17844), 
        .B1(n18437), .Y(n17857) );
  sky130_fd_sc_hd__nor2_1 U22625 ( .A(n17847), .B(n18349), .Y(n17872) );
  sky130_fd_sc_hd__a31oi_1 U22626 ( .A1(n17849), .A2(n17848), .A3(n17872), 
        .B1(n18439), .Y(n17856) );
  sky130_fd_sc_hd__a31oi_1 U22627 ( .A1(n17851), .A2(n17850), .A3(n18344), 
        .B1(n18445), .Y(n17855) );
  sky130_fd_sc_hd__nor2_1 U22628 ( .A(n18354), .B(n17852), .Y(n18394) );
  sky130_fd_sc_hd__a31oi_1 U22629 ( .A1(n17853), .A2(n18401), .A3(n18394), 
        .B1(n18423), .Y(n17854) );
  sky130_fd_sc_hd__nor4_1 U22630 ( .A(n17857), .B(n17856), .C(n17855), .D(
        n17854), .Y(n17858) );
  sky130_fd_sc_hd__o22ai_1 U22631 ( .A1(n17858), .A2(n18666), .B1(n18759), 
        .B2(n25182), .Y(n17901) );
  sky130_fd_sc_hd__a22o_1 U22632 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[72]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[40]), .X(n17900) );
  sky130_fd_sc_hd__clkinv_1 U22633 ( .A(j202_soc_core_uart_TOP_rx_fifo_wp[0]), 
        .Y(n25234) );
  sky130_fd_sc_hd__clkinv_1 U22634 ( .A(j202_soc_core_uart_TOP_rx_fifo_wp[1]), 
        .Y(n25232) );
  sky130_fd_sc_hd__o22ai_1 U22635 ( .A1(j202_soc_core_uart_TOP_rx_fifo_rp[1]), 
        .A2(j202_soc_core_uart_TOP_rx_fifo_wp[1]), .B1(n25203), .B2(n25232), 
        .Y(n23261) );
  sky130_fd_sc_hd__o221ai_1 U22636 ( .A1(j202_soc_core_uart_TOP_rx_fifo_wp[0]), 
        .A2(n25206), .B1(n25234), .B2(j202_soc_core_uart_TOP_rx_fifo_rp[0]), 
        .C1(n23261), .Y(n20073) );
  sky130_fd_sc_hd__a22oi_1 U22637 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[8]), .B1(n18724), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[104]), .Y(n17859) );
  sky130_fd_sc_hd__o31ai_1 U22638 ( .A1(j202_soc_core_uart_TOP_rx_fifo_gb), 
        .A2(n18245), .A3(n20073), .B1(n17859), .Y(n17899) );
  sky130_fd_sc_hd__nor4_1 U22639 ( .A(n17860), .B(n17866), .C(n17915), .D(
        n18353), .Y(n17861) );
  sky130_fd_sc_hd__a31oi_1 U22640 ( .A1(n18389), .A2(n18394), .A3(n17861), 
        .B1(n18439), .Y(n17881) );
  sky130_fd_sc_hd__nor2_1 U22641 ( .A(n17940), .B(n17862), .Y(n18342) );
  sky130_fd_sc_hd__a31oi_1 U22642 ( .A1(n17874), .A2(n18342), .A3(n17863), 
        .B1(n18437), .Y(n17880) );
  sky130_fd_sc_hd__nor3_1 U22643 ( .A(n17866), .B(n17865), .C(n17864), .Y(
        n18427) );
  sky130_fd_sc_hd__nor2_1 U22644 ( .A(n17915), .B(n17867), .Y(n17947) );
  sky130_fd_sc_hd__nand2_1 U22645 ( .A(n17869), .B(n17868), .Y(n18411) );
  sky130_fd_sc_hd__nor4_1 U22646 ( .A(n17870), .B(n18395), .C(n18411), .D(
        n18433), .Y(n17871) );
  sky130_fd_sc_hd__a31oi_1 U22647 ( .A1(n18427), .A2(n17947), .A3(n17871), 
        .B1(n18445), .Y(n17879) );
  sky130_fd_sc_hd__nor3b_1 U22648 ( .C_N(n17874), .A(n18352), .B(n17873), .Y(
        n17877) );
  sky130_fd_sc_hd__a31oi_1 U22649 ( .A1(n17877), .A2(n17876), .A3(n17875), 
        .B1(n18423), .Y(n17878) );
  sky130_fd_sc_hd__nor4_1 U22650 ( .A(n17881), .B(n17880), .C(n17879), .D(
        n17878), .Y(n17897) );
  sky130_fd_sc_hd__a22o_1 U22651 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[8]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[72]), .X(n17882) );
  sky130_fd_sc_hd__a21oi_1 U22652 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[104]), .B1(n17882), .Y(n17884) );
  sky130_fd_sc_hd__a22oi_1 U22653 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[168]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[136]), .Y(n17883) );
  sky130_fd_sc_hd__a21oi_1 U22654 ( .A1(n17884), .A2(n17883), .B1(n18736), .Y(
        n17895) );
  sky130_fd_sc_hd__a22oi_1 U22655 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[264]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[40]), .Y(n17893) );
  sky130_fd_sc_hd__a22o_1 U22656 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[296]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[328]), .X(n17885) );
  sky130_fd_sc_hd__a21oi_1 U22657 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[360]), .B1(n17885), .Y(n17892) );
  sky130_fd_sc_hd__nand2_1 U22658 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[232]), .Y(n17889) );
  sky130_fd_sc_hd__a21oi_1 U22659 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[456]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n17888) );
  sky130_fd_sc_hd__nand2_1 U22660 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[392]), .Y(n17887) );
  sky130_fd_sc_hd__nand2_1 U22661 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[424]), .Y(n17886) );
  sky130_fd_sc_hd__nand4_1 U22662 ( .A(n17889), .B(n17888), .C(n17887), .D(
        n17886), .Y(n17890) );
  sky130_fd_sc_hd__a21oi_1 U22663 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[200]), .B1(n17890), .Y(n17891) );
  sky130_fd_sc_hd__nand3_1 U22664 ( .A(n17893), .B(n17892), .C(n17891), .Y(
        n17894) );
  sky130_fd_sc_hd__o22ai_1 U22665 ( .A1(j202_soc_core_memory0_ram_dout0[488]), 
        .A2(n18758), .B1(n17895), .B2(n17894), .Y(n17896) );
  sky130_fd_sc_hd__o22ai_1 U22666 ( .A1(n17897), .A2(n18720), .B1(n18761), 
        .B2(n17896), .Y(n17898) );
  sky130_fd_sc_hd__nor4_1 U22667 ( .A(n17901), .B(n17900), .C(n17899), .D(
        n17898), .Y(n17955) );
  sky130_fd_sc_hd__nor3_1 U22668 ( .A(n17926), .B(n17903), .C(n17902), .Y(
        n17904) );
  sky130_fd_sc_hd__a31oi_1 U22669 ( .A1(n18429), .A2(n17904), .A3(n18347), 
        .B1(n18423), .Y(n17922) );
  sky130_fd_sc_hd__nor4_1 U22670 ( .A(n18412), .B(n18404), .C(n17905), .D(
        n18349), .Y(n17906) );
  sky130_fd_sc_hd__a31oi_1 U22671 ( .A1(n17908), .A2(n17907), .A3(n17906), 
        .B1(n18445), .Y(n17921) );
  sky130_fd_sc_hd__nor2_1 U22672 ( .A(n17910), .B(n17909), .Y(n18415) );
  sky130_fd_sc_hd__nand4_1 U22673 ( .A(n18415), .B(n17912), .C(n17911), .D(
        n18399), .Y(n17913) );
  sky130_fd_sc_hd__nor4b_1 U22674 ( .D_N(n17914), .A(n18392), .B(n18442), .C(
        n17913), .Y(n17919) );
  sky130_fd_sc_hd__nor2_1 U22675 ( .A(n17916), .B(n17915), .Y(n18343) );
  sky130_fd_sc_hd__nor4_1 U22676 ( .A(n18441), .B(n18395), .C(n17917), .D(
        n18416), .Y(n17918) );
  sky130_fd_sc_hd__o22ai_1 U22677 ( .A1(n17919), .A2(n18437), .B1(n17918), 
        .B2(n18439), .Y(n17920) );
  sky130_fd_sc_hd__nor3_1 U22678 ( .A(n17922), .B(n17921), .C(n17920), .Y(
        n17953) );
  sky130_fd_sc_hd__nand2_1 U22679 ( .A(n18425), .B(n18399), .Y(n18350) );
  sky130_fd_sc_hd__nor3_1 U22680 ( .A(n18417), .B(n18353), .C(n18350), .Y(
        n17924) );
  sky130_fd_sc_hd__a31oi_1 U22681 ( .A1(n17925), .A2(n17924), .A3(n17923), 
        .B1(n18439), .Y(n17951) );
  sky130_fd_sc_hd__nor4_1 U22682 ( .A(n17929), .B(n17928), .C(n17927), .D(
        n17926), .Y(n17933) );
  sky130_fd_sc_hd__nand2_1 U22683 ( .A(n17931), .B(n17930), .Y(n17932) );
  sky130_fd_sc_hd__a31oi_1 U22684 ( .A1(n17933), .A2(n17932), .A3(n18413), 
        .B1(n18445), .Y(n17950) );
  sky130_fd_sc_hd__nor4_1 U22685 ( .A(n17935), .B(n18392), .C(n17934), .D(
        n18443), .Y(n17936) );
  sky130_fd_sc_hd__a31oi_1 U22686 ( .A1(n17938), .A2(n17937), .A3(n17936), 
        .B1(n18423), .Y(n17949) );
  sky130_fd_sc_hd__nor3_1 U22687 ( .A(n17941), .B(n17940), .C(n17939), .Y(
        n18426) );
  sky130_fd_sc_hd__nor4_1 U22688 ( .A(n17945), .B(n17944), .C(n17943), .D(
        n17942), .Y(n17946) );
  sky130_fd_sc_hd__a31oi_1 U22689 ( .A1(n17947), .A2(n18426), .A3(n17946), 
        .B1(n18437), .Y(n17948) );
  sky130_fd_sc_hd__nor4_1 U22690 ( .A(n17951), .B(n17950), .C(n17949), .D(
        n17948), .Y(n17952) );
  sky130_fd_sc_hd__o22a_1 U22691 ( .A1(n17953), .A2(n18552), .B1(n18722), .B2(
        n17952), .X(n17954) );
  sky130_fd_sc_hd__nand2_1 U22692 ( .A(n17955), .B(n17954), .Y(n25308) );
  sky130_fd_sc_hd__nor2_1 U22693 ( .A(n17957), .B(n17956), .Y(n18175) );
  sky130_fd_sc_hd__nand4_1 U22694 ( .A(n18175), .B(n17959), .C(n18120), .D(
        n17958), .Y(n17967) );
  sky130_fd_sc_hd__nor2_1 U22695 ( .A(n17960), .B(n18114), .Y(n18171) );
  sky130_fd_sc_hd__nand2_1 U22696 ( .A(n17961), .B(n18149), .Y(n18138) );
  sky130_fd_sc_hd__nor4_1 U22697 ( .A(n17968), .B(n17963), .C(n18138), .D(
        n17962), .Y(n17964) );
  sky130_fd_sc_hd__a31oi_1 U22698 ( .A1(n17965), .A2(n18171), .A3(n17964), 
        .B1(n18147), .Y(n17966) );
  sky130_fd_sc_hd__a21oi_1 U22699 ( .A1(n18161), .A2(n17967), .B1(n17966), .Y(
        n17980) );
  sky130_fd_sc_hd__nor2_1 U22700 ( .A(n17969), .B(n17968), .Y(n18160) );
  sky130_fd_sc_hd__nand4_1 U22701 ( .A(n17972), .B(n18160), .C(n17971), .D(
        n17970), .Y(n17973) );
  sky130_fd_sc_hd__o21ai_1 U22702 ( .A1(n17974), .A2(n17973), .B1(n18155), .Y(
        n17979) );
  sky130_fd_sc_hd__nor2_1 U22703 ( .A(n17975), .B(n18101), .Y(n17976) );
  sky130_fd_sc_hd__nand4_1 U22704 ( .A(n17976), .B(n18095), .C(n18144), .D(
        n18158), .Y(n17977) );
  sky130_fd_sc_hd__o21ai_1 U22705 ( .A1(n18131), .A2(n17977), .B1(n18189), .Y(
        n17978) );
  sky130_fd_sc_hd__a31oi_1 U22706 ( .A1(n17980), .A2(n17979), .A3(n17978), 
        .B1(n18164), .Y(n18056) );
  sky130_fd_sc_hd__nand4_1 U22707 ( .A(n17992), .B(n17983), .C(n17982), .D(
        n17981), .Y(n17987) );
  sky130_fd_sc_hd__nor3_1 U22708 ( .A(n17984), .B(n18101), .C(n18009), .Y(
        n18082) );
  sky130_fd_sc_hd__a31oi_1 U22709 ( .A1(n18082), .A2(n18181), .A3(n17985), 
        .B1(n18147), .Y(n17986) );
  sky130_fd_sc_hd__a21oi_1 U22710 ( .A1(n18161), .A2(n17987), .B1(n17986), .Y(
        n18002) );
  sky130_fd_sc_hd__nand2_1 U22711 ( .A(n18115), .B(n17988), .Y(n18163) );
  sky130_fd_sc_hd__nand2_1 U22712 ( .A(n18119), .B(n18032), .Y(n18025) );
  sky130_fd_sc_hd__nor3_1 U22713 ( .A(n17991), .B(n17990), .C(n17989), .Y(
        n18088) );
  sky130_fd_sc_hd__nand4b_1 U22714 ( .A_N(n18025), .B(n18088), .C(n17993), .D(
        n17992), .Y(n17994) );
  sky130_fd_sc_hd__o21ai_1 U22715 ( .A1(n18163), .A2(n17994), .B1(n18155), .Y(
        n18001) );
  sky130_fd_sc_hd__nor3_1 U22716 ( .A(n17997), .B(n17996), .C(n17995), .Y(
        n18186) );
  sky130_fd_sc_hd__nand4_1 U22717 ( .A(n17998), .B(n18186), .C(n18180), .D(
        n18081), .Y(n17999) );
  sky130_fd_sc_hd__o21ai_1 U22718 ( .A1(n18010), .A2(n17999), .B1(n18189), .Y(
        n18000) );
  sky130_fd_sc_hd__a31oi_1 U22719 ( .A1(n18002), .A2(n18001), .A3(n18000), 
        .B1(n18190), .Y(n18055) );
  sky130_fd_sc_hd__nand2_1 U22720 ( .A(n18135), .B(n18003), .Y(n18157) );
  sky130_fd_sc_hd__nor4_1 U22721 ( .A(n18006), .B(n18005), .C(n18004), .D(
        n18157), .Y(n18008) );
  sky130_fd_sc_hd__a21oi_1 U22722 ( .A1(n18008), .A2(n18007), .B1(n18172), .Y(
        n18023) );
  sky130_fd_sc_hd__nor4_1 U22723 ( .A(n18112), .B(n18099), .C(n18010), .D(
        n18009), .Y(n18011) );
  sky130_fd_sc_hd__a31oi_1 U22724 ( .A1(n18011), .A2(n18125), .A3(n18086), 
        .B1(n18147), .Y(n18022) );
  sky130_fd_sc_hd__nor4_1 U22725 ( .A(n18015), .B(n18014), .C(n18013), .D(
        n18012), .Y(n18020) );
  sky130_fd_sc_hd__nor4b_1 U22726 ( .D_N(n18018), .A(n18025), .B(n18017), .C(
        n18016), .Y(n18019) );
  sky130_fd_sc_hd__o22ai_1 U22727 ( .A1(n18020), .A2(n18183), .B1(n18019), 
        .B2(n18047), .Y(n18021) );
  sky130_fd_sc_hd__nor3_1 U22728 ( .A(n18023), .B(n18022), .C(n18021), .Y(
        n18053) );
  sky130_fd_sc_hd__nor4_1 U22729 ( .A(n18026), .B(n18025), .C(n18024), .D(
        n18117), .Y(n18027) );
  sky130_fd_sc_hd__a31oi_1 U22730 ( .A1(n18029), .A2(n18028), .A3(n18027), 
        .B1(n18183), .Y(n18051) );
  sky130_fd_sc_hd__nor2_1 U22731 ( .A(n18031), .B(n18030), .Y(n18184) );
  sky130_fd_sc_hd__a31oi_1 U22732 ( .A1(n18184), .A2(n18033), .A3(n18032), 
        .B1(n18172), .Y(n18050) );
  sky130_fd_sc_hd__nor2_1 U22733 ( .A(n18034), .B(n18123), .Y(n18036) );
  sky130_fd_sc_hd__nand4_1 U22734 ( .A(n18037), .B(n18036), .C(n18035), .D(
        n18154), .Y(n18038) );
  sky130_fd_sc_hd__nor4_1 U22735 ( .A(n18041), .B(n18040), .C(n18039), .D(
        n18038), .Y(n18048) );
  sky130_fd_sc_hd__nor4_1 U22736 ( .A(n18045), .B(n18044), .C(n18043), .D(
        n18042), .Y(n18046) );
  sky130_fd_sc_hd__o22ai_1 U22737 ( .A1(n18048), .A2(n18047), .B1(n18046), 
        .B2(n18147), .Y(n18049) );
  sky130_fd_sc_hd__nor3_1 U22738 ( .A(n18051), .B(n18050), .C(n18049), .Y(
        n18052) );
  sky130_fd_sc_hd__o22ai_1 U22739 ( .A1(n18053), .A2(n18139), .B1(n18052), 
        .B2(n18107), .Y(n18054) );
  sky130_fd_sc_hd__nor3_1 U22740 ( .A(n18056), .B(n18055), .C(n18054), .Y(
        n18073) );
  sky130_fd_sc_hd__a22oi_1 U22741 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[240]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[208]), .Y(n18060) );
  sky130_fd_sc_hd__a22oi_1 U22742 ( .A1(n18734), .A2(
        j202_soc_core_memory0_ram_dout0[144]), .B1(n18733), .B2(
        j202_soc_core_memory0_ram_dout0[112]), .Y(n18059) );
  sky130_fd_sc_hd__a22oi_1 U22743 ( .A1(n18361), .A2(
        j202_soc_core_memory0_ram_dout0[48]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[80]), .Y(n18058) );
  sky130_fd_sc_hd__nand2_1 U22744 ( .A(n18735), .B(
        j202_soc_core_memory0_ram_dout0[176]), .Y(n18057) );
  sky130_fd_sc_hd__nand4_1 U22745 ( .A(n18060), .B(n18059), .C(n18058), .D(
        n18057), .Y(n18061) );
  sky130_fd_sc_hd__a21oi_1 U22746 ( .A1(n18367), .A2(
        j202_soc_core_memory0_ram_dout0[16]), .B1(n18061), .Y(n18070) );
  sky130_fd_sc_hd__a22oi_1 U22747 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[304]), .B1(n18062), .B2(
        j202_soc_core_memory0_ram_dout0[272]), .Y(n18069) );
  sky130_fd_sc_hd__nand2_1 U22748 ( .A(n18743), .B(
        j202_soc_core_memory0_ram_dout0[368]), .Y(n18066) );
  sky130_fd_sc_hd__a21oi_1 U22749 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[464]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n18065) );
  sky130_fd_sc_hd__nand2_1 U22750 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[400]), .Y(n18064) );
  sky130_fd_sc_hd__nand2_1 U22751 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[432]), .Y(n18063) );
  sky130_fd_sc_hd__nand4_1 U22752 ( .A(n18066), .B(n18065), .C(n18064), .D(
        n18063), .Y(n18067) );
  sky130_fd_sc_hd__a21oi_1 U22753 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[336]), .B1(n18067), .Y(n18068) );
  sky130_fd_sc_hd__o211ai_1 U22754 ( .A1(n18736), .A2(n18070), .B1(n18069), 
        .C1(n18068), .Y(n18071) );
  sky130_fd_sc_hd__o22ai_1 U22756 ( .A1(n18073), .A2(n18212), .B1(n18761), 
        .B2(n18072), .Y(n18074) );
  sky130_fd_sc_hd__a21oi_1 U22757 ( .A1(n18629), .A2(
        j202_soc_core_bldc_core_00_pwm_duty[4]), .B1(n18074), .Y(n18077) );
  sky130_fd_sc_hd__a22oi_1 U22758 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[16]), .B1(n18727), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[80]), .Y(n18076) );
  sky130_fd_sc_hd__a22oi_1 U22759 ( .A1(n18726), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[48]), .B1(n18379), .B2(
        j202_soc_core_uart_div1[0]), .Y(n18075) );
  sky130_fd_sc_hd__nand3_1 U22760 ( .A(n18077), .B(n18076), .C(n18075), .Y(
        n22516) );
  sky130_fd_sc_hd__nand2_1 U22761 ( .A(n22516), .B(n19089), .Y(n18080) );
  sky130_fd_sc_hd__a22oi_1 U22762 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__0_), .B1(n19088), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__0_), .Y(n18079) );
  sky130_fd_sc_hd__nand2_1 U22763 ( .A(n25259), .B(n19087), .Y(n18078) );
  sky130_fd_sc_hd__nand3_1 U22764 ( .A(n18080), .B(n18079), .C(n18078), .Y(
        n25372) );
  sky130_fd_sc_hd__nand4_1 U22765 ( .A(n18144), .B(n18083), .C(n18082), .D(
        n18081), .Y(n18090) );
  sky130_fd_sc_hd__nor2_1 U22766 ( .A(n18085), .B(n18084), .Y(n18087) );
  sky130_fd_sc_hd__a31oi_1 U22767 ( .A1(n18088), .A2(n18087), .A3(n18086), 
        .B1(n18147), .Y(n18089) );
  sky130_fd_sc_hd__a21oi_1 U22768 ( .A1(n18155), .A2(n18090), .B1(n18089), .Y(
        n18110) );
  sky130_fd_sc_hd__nor2_1 U22769 ( .A(n18092), .B(n18091), .Y(n18094) );
  sky130_fd_sc_hd__nand4_1 U22770 ( .A(n18095), .B(n18094), .C(n18093), .D(
        n18134), .Y(n18096) );
  sky130_fd_sc_hd__o21ai_1 U22771 ( .A1(n18097), .A2(n18096), .B1(n18189), .Y(
        n18109) );
  sky130_fd_sc_hd__nor4_1 U22772 ( .A(n18101), .B(n18100), .C(n18099), .D(
        n18098), .Y(n18103) );
  sky130_fd_sc_hd__nand4_1 U22773 ( .A(n18104), .B(n18103), .C(n18179), .D(
        n18102), .Y(n18105) );
  sky130_fd_sc_hd__a31oi_1 U22775 ( .A1(n18110), .A2(n18109), .A3(n18108), 
        .B1(n18107), .Y(n18196) );
  sky130_fd_sc_hd__nor4_1 U22776 ( .A(n18114), .B(n18113), .C(n18112), .D(
        n18111), .Y(n18116) );
  sky130_fd_sc_hd__nand4b_1 U22777 ( .A_N(n18117), .B(n18160), .C(n18116), .D(
        n18115), .Y(n18129) );
  sky130_fd_sc_hd__nand2_1 U22778 ( .A(n18118), .B(n18133), .Y(n18122) );
  sky130_fd_sc_hd__nand4_1 U22779 ( .A(n18121), .B(n18120), .C(n18154), .D(
        n18119), .Y(n18146) );
  sky130_fd_sc_hd__nor4_1 U22780 ( .A(n18124), .B(n18123), .C(n18122), .D(
        n18146), .Y(n18126) );
  sky130_fd_sc_hd__a31oi_1 U22781 ( .A1(n18127), .A2(n18126), .A3(n18125), 
        .B1(n18147), .Y(n18128) );
  sky130_fd_sc_hd__a21oi_1 U22782 ( .A1(n18189), .A2(n18129), .B1(n18128), .Y(
        n18142) );
  sky130_fd_sc_hd__o31ai_1 U22783 ( .A1(n18132), .A2(n18131), .A3(n18130), 
        .B1(n18161), .Y(n18141) );
  sky130_fd_sc_hd__nand4_1 U22784 ( .A(n18136), .B(n18135), .C(n18134), .D(
        n18133), .Y(n18137) );
  sky130_fd_sc_hd__o21ai_1 U22785 ( .A1(n18138), .A2(n18137), .B1(n18155), .Y(
        n18140) );
  sky130_fd_sc_hd__a31oi_1 U22786 ( .A1(n18142), .A2(n18141), .A3(n18140), 
        .B1(n18139), .Y(n18195) );
  sky130_fd_sc_hd__nand4_1 U22787 ( .A(n18145), .B(n18144), .C(n18143), .D(
        n18174), .Y(n18151) );
  sky130_fd_sc_hd__a21oi_1 U22788 ( .A1(n18149), .A2(n18148), .B1(n18147), .Y(
        n18150) );
  sky130_fd_sc_hd__a21oi_1 U22789 ( .A1(n18189), .A2(n18151), .B1(n18150), .Y(
        n18167) );
  sky130_fd_sc_hd__nand3_1 U22790 ( .A(n18154), .B(n18153), .C(n18152), .Y(
        n18156) );
  sky130_fd_sc_hd__o21ai_1 U22791 ( .A1(n18157), .A2(n18156), .B1(n18155), .Y(
        n18166) );
  sky130_fd_sc_hd__nand4_1 U22792 ( .A(n18160), .B(n18159), .C(n18179), .D(
        n18158), .Y(n18162) );
  sky130_fd_sc_hd__a31oi_1 U22794 ( .A1(n18167), .A2(n18166), .A3(n18165), 
        .B1(n18164), .Y(n18194) );
  sky130_fd_sc_hd__nand4_1 U22795 ( .A(n18171), .B(n18170), .C(n18169), .D(
        n18168), .Y(n18177) );
  sky130_fd_sc_hd__a31oi_1 U22796 ( .A1(n18175), .A2(n18174), .A3(n18173), 
        .B1(n18172), .Y(n18176) );
  sky130_fd_sc_hd__a21oi_1 U22797 ( .A1(n18178), .A2(n18177), .B1(n18176), .Y(
        n18192) );
  sky130_fd_sc_hd__nand4_1 U22798 ( .A(n18182), .B(n18181), .C(n18180), .D(
        n18179), .Y(n18188) );
  sky130_fd_sc_hd__a31oi_1 U22799 ( .A1(n18186), .A2(n18185), .A3(n18184), 
        .B1(n18183), .Y(n18187) );
  sky130_fd_sc_hd__a21oi_1 U22800 ( .A1(n18189), .A2(n18188), .B1(n18187), .Y(
        n18191) );
  sky130_fd_sc_hd__a21oi_1 U22801 ( .A1(n18192), .A2(n18191), .B1(n18190), .Y(
        n18193) );
  sky130_fd_sc_hd__nor4_1 U22802 ( .A(n18196), .B(n18195), .C(n18194), .D(
        n18193), .Y(n18213) );
  sky130_fd_sc_hd__a22o_1 U22803 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[17]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[81]), .X(n18197) );
  sky130_fd_sc_hd__a21oi_1 U22804 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[113]), .B1(n18197), .Y(n18199) );
  sky130_fd_sc_hd__a22oi_1 U22805 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[177]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[145]), .Y(n18198) );
  sky130_fd_sc_hd__a21oi_1 U22806 ( .A1(n18199), .A2(n18198), .B1(n18736), .Y(
        n18210) );
  sky130_fd_sc_hd__a22oi_1 U22807 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[273]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[49]), .Y(n18208) );
  sky130_fd_sc_hd__a22o_1 U22808 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[305]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[337]), .X(n18200) );
  sky130_fd_sc_hd__a21oi_1 U22809 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[369]), .B1(n18200), .Y(n18207) );
  sky130_fd_sc_hd__nand2_1 U22810 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[241]), .Y(n18204) );
  sky130_fd_sc_hd__a21oi_1 U22811 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[465]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n18203) );
  sky130_fd_sc_hd__nand2_1 U22812 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[401]), .Y(n18202) );
  sky130_fd_sc_hd__nand2_1 U22813 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[433]), .Y(n18201) );
  sky130_fd_sc_hd__nand4_1 U22814 ( .A(n18204), .B(n18203), .C(n18202), .D(
        n18201), .Y(n18205) );
  sky130_fd_sc_hd__a21oi_1 U22815 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[209]), .B1(n18205), .Y(n18206) );
  sky130_fd_sc_hd__nand3_1 U22816 ( .A(n18208), .B(n18207), .C(n18206), .Y(
        n18209) );
  sky130_fd_sc_hd__o22ai_1 U22817 ( .A1(j202_soc_core_memory0_ram_dout0[497]), 
        .A2(n18758), .B1(n18210), .B2(n18209), .Y(n18211) );
  sky130_fd_sc_hd__o22ai_1 U22818 ( .A1(n18213), .A2(n18212), .B1(n18761), 
        .B2(n18211), .Y(n18214) );
  sky130_fd_sc_hd__a21oi_1 U22819 ( .A1(n18629), .A2(
        j202_soc_core_bldc_core_00_pwm_duty[5]), .B1(n18214), .Y(n18217) );
  sky130_fd_sc_hd__a22oi_1 U22820 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[17]), .B1(n18727), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[81]), .Y(n18216) );
  sky130_fd_sc_hd__a22oi_1 U22821 ( .A1(n18726), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[49]), .B1(n18379), .B2(
        j202_soc_core_uart_div1[1]), .Y(n18215) );
  sky130_fd_sc_hd__nand3_1 U22822 ( .A(n18217), .B(n18216), .C(n18215), .Y(
        n22521) );
  sky130_fd_sc_hd__a22oi_1 U22823 ( .A1(n19089), .A2(n22521), .B1(n25274), 
        .B2(n19087), .Y(n18219) );
  sky130_fd_sc_hd__a22oi_1 U22824 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__1_), .B1(n19088), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__1_), .Y(n18218) );
  sky130_fd_sc_hd__nand2_1 U22825 ( .A(n25246), .B(n19087), .Y(n18222) );
  sky130_fd_sc_hd__a22oi_1 U22826 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__2_), .B1(n19088), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__2_), .Y(n18221) );
  sky130_fd_sc_hd__nand2_1 U22827 ( .A(n22523), .B(n19089), .Y(n18220) );
  sky130_fd_sc_hd__nand2_1 U22828 ( .A(n22522), .B(n19089), .Y(n18225) );
  sky130_fd_sc_hd__a22oi_1 U22829 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__3_), .B1(n19088), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__3_), .Y(n18224) );
  sky130_fd_sc_hd__nand2_1 U22830 ( .A(n25253), .B(n19087), .Y(n18223) );
  sky130_fd_sc_hd__a22o_1 U22831 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[6]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[70]), .X(n18226) );
  sky130_fd_sc_hd__a21oi_1 U22832 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[102]), .B1(n18226), .Y(n18228) );
  sky130_fd_sc_hd__a22oi_1 U22833 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[166]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[134]), .Y(n18227) );
  sky130_fd_sc_hd__a21oi_1 U22834 ( .A1(n18228), .A2(n18227), .B1(n18736), .Y(
        n18239) );
  sky130_fd_sc_hd__a22oi_1 U22835 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[262]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[38]), .Y(n18237) );
  sky130_fd_sc_hd__a22o_1 U22836 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[294]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[326]), .X(n18229) );
  sky130_fd_sc_hd__a21oi_1 U22837 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[358]), .B1(n18229), .Y(n18236) );
  sky130_fd_sc_hd__nand2_1 U22838 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[230]), .Y(n18233) );
  sky130_fd_sc_hd__a21oi_1 U22839 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[454]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n18232) );
  sky130_fd_sc_hd__nand2_1 U22840 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[390]), .Y(n18231) );
  sky130_fd_sc_hd__nand2_1 U22841 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[422]), .Y(n18230) );
  sky130_fd_sc_hd__nand4_1 U22842 ( .A(n18233), .B(n18232), .C(n18231), .D(
        n18230), .Y(n18234) );
  sky130_fd_sc_hd__a21oi_1 U22843 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[198]), .B1(n18234), .Y(n18235) );
  sky130_fd_sc_hd__nand3_1 U22844 ( .A(n18237), .B(n18236), .C(n18235), .Y(
        n18238) );
  sky130_fd_sc_hd__o22ai_1 U22845 ( .A1(j202_soc_core_memory0_ram_dout0[486]), 
        .A2(n18758), .B1(n18239), .B2(n18238), .Y(n18240) );
  sky130_fd_sc_hd__nor2_1 U22846 ( .A(n18761), .B(n18240), .Y(n18311) );
  sky130_fd_sc_hd__a22oi_1 U22847 ( .A1(n18242), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[14]), .B1(n18241), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[30]), .Y(n18247) );
  sky130_fd_sc_hd__a22oi_1 U22848 ( .A1(n18244), .A2(
        j202_soc_core_uart_TOP_rx_fifo_mem[22]), .B1(n18243), .B2(
        j202_soc_core_uart_TOP_rx_fifo_mem[6]), .Y(n18246) );
  sky130_fd_sc_hd__a21oi_1 U22849 ( .A1(n18247), .A2(n18246), .B1(n18245), .Y(
        n18310) );
  sky130_fd_sc_hd__nor2_1 U22850 ( .A(n18248), .B(n18703), .Y(n18249) );
  sky130_fd_sc_hd__a31oi_1 U22851 ( .A1(n18249), .A2(n18544), .A3(n18252), 
        .B1(n18779), .Y(n18262) );
  sky130_fd_sc_hd__nor3_1 U22852 ( .A(n18250), .B(n18776), .C(n18679), .Y(
        n18251) );
  sky130_fd_sc_hd__a31oi_1 U22853 ( .A1(n18252), .A2(n18542), .A3(n18251), 
        .B1(n18792), .Y(n18261) );
  sky130_fd_sc_hd__o31a_1 U22854 ( .A1(n18254), .A2(n18253), .A3(n18312), .B1(
        n18664), .X(n18260) );
  sky130_fd_sc_hd__nor3_1 U22855 ( .A(n18256), .B(n18524), .C(n18255), .Y(
        n18257) );
  sky130_fd_sc_hd__a31oi_1 U22856 ( .A1(n18258), .A2(n18683), .A3(n18257), 
        .B1(n18783), .Y(n18259) );
  sky130_fd_sc_hd__nor4_1 U22857 ( .A(n18262), .B(n18261), .C(n18260), .D(
        n18259), .Y(n18275) );
  sky130_fd_sc_hd__a21oi_1 U22858 ( .A1(n18265), .A2(n18264), .B1(n18779), .Y(
        n18272) );
  sky130_fd_sc_hd__nand2_1 U22859 ( .A(n18267), .B(n18266), .Y(n18690) );
  sky130_fd_sc_hd__nand2_1 U22860 ( .A(n18698), .B(n18681), .Y(n18319) );
  sky130_fd_sc_hd__nor4_1 U22861 ( .A(n18673), .B(n18268), .C(n18690), .D(
        n18319), .Y(n18269) );
  sky130_fd_sc_hd__o22ai_1 U22862 ( .A1(n18270), .A2(n18783), .B1(n18269), 
        .B2(n18792), .Y(n18271) );
  sky130_fd_sc_hd__a211oi_1 U22863 ( .A1(n18664), .A2(n18273), .B1(n18272), 
        .C1(n18271), .Y(n18274) );
  sky130_fd_sc_hd__o22ai_1 U22864 ( .A1(n18275), .A2(n18666), .B1(n18274), 
        .B2(n18720), .Y(n18309) );
  sky130_fd_sc_hd__a21oi_1 U22865 ( .A1(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[2]), .A2(j202_soc_core_ahblite_interconnect_s_hrdata[38]), .B1(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[3]), .Y(n18279) );
  sky130_fd_sc_hd__nand3_1 U22866 ( .A(n18277), .B(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[1]), .C(j202_soc_core_ahblite_interconnect_s_hrdata[70]), .Y(n18278) );
  sky130_fd_sc_hd__nand2_1 U22867 ( .A(n18279), .B(n18278), .Y(n18280) );
  sky130_fd_sc_hd__a21oi_1 U22868 ( .A1(n18281), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[102]), .B1(n18280), .Y(
        n18286) );
  sky130_fd_sc_hd__a21oi_1 U22869 ( .A1(n18284), .A2(
        j202_soc_core_bldc_core_00_pwm_period[6]), .B1(n18283), .Y(n18285) );
  sky130_fd_sc_hd__o31ai_1 U22870 ( .A1(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[4]), .A2(n18286), .A3(n18285), .B1(n18288), .Y(n18287) );
  sky130_fd_sc_hd__nand4_1 U22872 ( .A(n18712), .B(n18321), .C(n18290), .D(
        n18289), .Y(n18304) );
  sky130_fd_sc_hd__nand4_1 U22873 ( .A(n18292), .B(n18555), .C(n18291), .D(
        n18662), .Y(n18293) );
  sky130_fd_sc_hd__o21ai_1 U22874 ( .A1(n18294), .A2(n18293), .B1(n18513), .Y(
        n18301) );
  sky130_fd_sc_hd__nor2_1 U22875 ( .A(n18296), .B(n18295), .Y(n18598) );
  sky130_fd_sc_hd__nand4b_1 U22876 ( .A_N(n18598), .B(n18594), .C(n18320), .D(
        n18297), .Y(n18298) );
  sky130_fd_sc_hd__nand3_1 U22878 ( .A(n18302), .B(n18301), .C(n18300), .Y(
        n18303) );
  sky130_fd_sc_hd__a21oi_1 U22879 ( .A1(n18651), .A2(n18304), .B1(n18303), .Y(
        n18305) );
  sky130_fd_sc_hd__o22ai_1 U22880 ( .A1(n18307), .A2(n18306), .B1(n18305), 
        .B2(n18722), .Y(n18308) );
  sky130_fd_sc_hd__nor4_1 U22881 ( .A(n18311), .B(n18310), .C(n18309), .D(
        n18308), .Y(n18331) );
  sky130_fd_sc_hd__nor2_1 U22882 ( .A(n18645), .B(n18585), .Y(n18577) );
  sky130_fd_sc_hd__nor2_1 U22883 ( .A(n18527), .B(n18312), .Y(n18313) );
  sky130_fd_sc_hd__a31oi_1 U22884 ( .A1(n18314), .A2(n18577), .A3(n18313), 
        .B1(n18792), .Y(n18328) );
  sky130_fd_sc_hd__nor4_1 U22885 ( .A(n18710), .B(n18638), .C(n18316), .D(
        n18315), .Y(n18317) );
  sky130_fd_sc_hd__a31oi_1 U22886 ( .A1(n18318), .A2(n18542), .A3(n18317), 
        .B1(n18779), .Y(n18327) );
  sky130_fd_sc_hd__nor4bb_1 U22887 ( .C_N(n18321), .D_N(n18320), .A(n18770), 
        .B(n18319), .Y(n18325) );
  sky130_fd_sc_hd__nor3_1 U22888 ( .A(n18766), .B(n18323), .C(n18322), .Y(
        n18324) );
  sky130_fd_sc_hd__o22ai_1 U22889 ( .A1(n18325), .A2(n18771), .B1(n18324), 
        .B2(n18783), .Y(n18326) );
  sky130_fd_sc_hd__nor3_1 U22890 ( .A(n18328), .B(n18327), .C(n18326), .Y(
        n18329) );
  sky130_fd_sc_hd__nand2b_1 U22891 ( .A_N(n18329), .B(n18798), .Y(n18330) );
  sky130_fd_sc_hd__nand2_1 U22892 ( .A(n18331), .B(n18330), .Y(n25276) );
  sky130_fd_sc_hd__nand2_1 U22893 ( .A(n25276), .B(n19087), .Y(n18334) );
  sky130_fd_sc_hd__a22oi_1 U22894 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__6_), .B1(n19088), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__6_), .Y(n18333) );
  sky130_fd_sc_hd__nand2_1 U22895 ( .A(n21135), .B(n19089), .Y(n18332) );
  sky130_fd_sc_hd__nand3_1 U22896 ( .A(n18334), .B(n18333), .C(n18332), .Y(
        n25384) );
  sky130_fd_sc_hd__nand2_1 U22897 ( .A(n22531), .B(n19089), .Y(n18337) );
  sky130_fd_sc_hd__a22oi_1 U22898 ( .A1(j202_soc_core_j22_cpu_id_opn_inst__7_), 
        .A2(n19088), .B1(j202_soc_core_j22_cpu_id_op2_v_), .B2(
        j202_soc_core_j22_cpu_id_op2_inst__7_), .Y(n18336) );
  sky130_fd_sc_hd__nand2_1 U22899 ( .A(n25247), .B(n19087), .Y(n18335) );
  sky130_fd_sc_hd__nand3_1 U22900 ( .A(n18337), .B(n18336), .C(n18335), .Y(
        n25383) );
  sky130_fd_sc_hd__nand2_1 U22901 ( .A(n25308), .B(n19087), .Y(n18340) );
  sky130_fd_sc_hd__a22oi_1 U22902 ( .A1(j202_soc_core_j22_cpu_id_opn_inst__8_), 
        .A2(n19088), .B1(j202_soc_core_j22_cpu_id_op2_v_), .B2(
        j202_soc_core_j22_cpu_id_op2_inst__8_), .Y(n18339) );
  sky130_fd_sc_hd__nand2_1 U22903 ( .A(n22524), .B(n19089), .Y(n18338) );
  sky130_fd_sc_hd__a31oi_1 U22904 ( .A1(n18343), .A2(n18342), .A3(n18341), 
        .B1(n18437), .Y(n18358) );
  sky130_fd_sc_hd__nand4_1 U22905 ( .A(n18347), .B(n18346), .C(n18345), .D(
        n18344), .Y(n18348) );
  sky130_fd_sc_hd__nor4_1 U22906 ( .A(n18351), .B(n18350), .C(n18349), .D(
        n18348), .Y(n18356) );
  sky130_fd_sc_hd__nor3_1 U22907 ( .A(n18354), .B(n18353), .C(n18352), .Y(
        n18355) );
  sky130_fd_sc_hd__o22ai_1 U22908 ( .A1(n18356), .A2(n18423), .B1(n18355), 
        .B2(n18439), .Y(n18357) );
  sky130_fd_sc_hd__nor3_1 U22909 ( .A(n18359), .B(n18358), .C(n18357), .Y(
        n18378) );
  sky130_fd_sc_hd__a22oi_1 U22910 ( .A1(j202_soc_core_memory0_ram_dout0_sel[7]), .A2(j202_soc_core_memory0_ram_dout0[233]), .B1(n18360), .B2(
        j202_soc_core_memory0_ram_dout0[201]), .Y(n18365) );
  sky130_fd_sc_hd__a22oi_1 U22911 ( .A1(n18734), .A2(
        j202_soc_core_memory0_ram_dout0[137]), .B1(n18733), .B2(
        j202_soc_core_memory0_ram_dout0[105]), .Y(n18364) );
  sky130_fd_sc_hd__a22oi_1 U22912 ( .A1(n18361), .A2(
        j202_soc_core_memory0_ram_dout0[41]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[73]), .Y(n18363) );
  sky130_fd_sc_hd__nand2_1 U22913 ( .A(n18735), .B(
        j202_soc_core_memory0_ram_dout0[169]), .Y(n18362) );
  sky130_fd_sc_hd__nand4_1 U22914 ( .A(n18365), .B(n18364), .C(n18363), .D(
        n18362), .Y(n18366) );
  sky130_fd_sc_hd__a21oi_1 U22915 ( .A1(n18367), .A2(
        j202_soc_core_memory0_ram_dout0[9]), .B1(n18366), .Y(n18375) );
  sky130_fd_sc_hd__a22oi_1 U22916 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[297]), .B1(n18062), .B2(
        j202_soc_core_memory0_ram_dout0[265]), .Y(n18374) );
  sky130_fd_sc_hd__nand2_1 U22917 ( .A(n18743), .B(
        j202_soc_core_memory0_ram_dout0[361]), .Y(n18371) );
  sky130_fd_sc_hd__a21oi_1 U22918 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[457]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n18370) );
  sky130_fd_sc_hd__nand2_1 U22919 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[393]), .Y(n18369) );
  sky130_fd_sc_hd__nand2_1 U22920 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[425]), .Y(n18368) );
  sky130_fd_sc_hd__nand4_1 U22921 ( .A(n18371), .B(n18370), .C(n18369), .D(
        n18368), .Y(n18372) );
  sky130_fd_sc_hd__a21oi_1 U22922 ( .A1(n18740), .A2(
        j202_soc_core_memory0_ram_dout0[329]), .B1(n18372), .Y(n18373) );
  sky130_fd_sc_hd__o211ai_1 U22923 ( .A1(n18736), .A2(n18375), .B1(n18374), 
        .C1(n18373), .Y(n18376) );
  sky130_fd_sc_hd__o22ai_1 U22925 ( .A1(n18378), .A2(n18720), .B1(n18761), 
        .B2(n18377), .Y(n18384) );
  sky130_fd_sc_hd__a22oi_1 U22926 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[9]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[41]), .Y(n18382) );
  sky130_fd_sc_hd__a22oi_1 U22927 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[73]), .B1(n18724), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[105]), .Y(n18381) );
  sky130_fd_sc_hd__clkinv_1 U22928 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[1]), 
        .Y(n23812) );
  sky130_fd_sc_hd__clkinv_1 U22929 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[1]), 
        .Y(n23831) );
  sky130_fd_sc_hd__o22ai_1 U22930 ( .A1(j202_soc_core_uart_TOP_tx_fifo_wp[1]), 
        .A2(j202_soc_core_uart_TOP_tx_fifo_rp[1]), .B1(n23812), .B2(n23831), 
        .Y(n23256) );
  sky130_fd_sc_hd__a21oi_1 U22932 ( .A1(j202_soc_core_uart_TOP_tx_fifo_wp[0]), 
        .A2(n25123), .B1(n23255), .Y(n23862) );
  sky130_fd_sc_hd__nand3_1 U22933 ( .A(n18379), .B(n23862), .C(
        j202_soc_core_uart_TOP_tx_fifo_gb), .Y(n18380) );
  sky130_fd_sc_hd__nand3_1 U22934 ( .A(n18382), .B(n18381), .C(n18380), .Y(
        n18383) );
  sky130_fd_sc_hd__a211oi_1 U22935 ( .A1(n18629), .A2(
        j202_soc_core_bldc_core_00_pwm_period[9]), .B1(n18384), .C1(n18383), 
        .Y(n18455) );
  sky130_fd_sc_hd__nand2_1 U22936 ( .A(n18401), .B(n18399), .Y(n18385) );
  sky130_fd_sc_hd__nor4_1 U22937 ( .A(n18398), .B(n18386), .C(n18411), .D(
        n18385), .Y(n18387) );
  sky130_fd_sc_hd__a31oi_1 U22938 ( .A1(n18389), .A2(n18388), .A3(n18387), 
        .B1(n18437), .Y(n18410) );
  sky130_fd_sc_hd__nor4_1 U22939 ( .A(n18392), .B(n18391), .C(n18390), .D(
        n18441), .Y(n18393) );
  sky130_fd_sc_hd__a21oi_1 U22940 ( .A1(n18394), .A2(n18393), .B1(n18445), .Y(
        n18409) );
  sky130_fd_sc_hd__nor4_1 U22941 ( .A(n18398), .B(n18397), .C(n18396), .D(
        n18395), .Y(n18407) );
  sky130_fd_sc_hd__nand4_1 U22942 ( .A(n18402), .B(n18401), .C(n18400), .D(
        n18399), .Y(n18403) );
  sky130_fd_sc_hd__nor3_1 U22943 ( .A(n18405), .B(n18404), .C(n18403), .Y(
        n18406) );
  sky130_fd_sc_hd__o22ai_1 U22944 ( .A1(n18407), .A2(n18439), .B1(n18406), 
        .B2(n18423), .Y(n18408) );
  sky130_fd_sc_hd__o31a_1 U22945 ( .A1(n18410), .A2(n18409), .A3(n18408), .B1(
        n18610), .X(n18453) );
  sky130_fd_sc_hd__nor2_1 U22946 ( .A(n18412), .B(n18411), .Y(n18414) );
  sky130_fd_sc_hd__a31oi_1 U22947 ( .A1(n18415), .A2(n18414), .A3(n18413), 
        .B1(n18445), .Y(n18421) );
  sky130_fd_sc_hd__nor3_1 U22948 ( .A(n18418), .B(n18417), .C(n18416), .Y(
        n18419) );
  sky130_fd_sc_hd__o22ai_1 U22949 ( .A1(n18427), .A2(n18437), .B1(n18419), 
        .B2(n18439), .Y(n18420) );
  sky130_fd_sc_hd__o31a_1 U22950 ( .A1(n18422), .A2(n18421), .A3(n18420), .B1(
        n18605), .X(n18452) );
  sky130_fd_sc_hd__a31oi_1 U22951 ( .A1(n18426), .A2(n18425), .A3(n18424), 
        .B1(n18423), .Y(n18450) );
  sky130_fd_sc_hd__nand4_1 U22952 ( .A(n18430), .B(n18429), .C(n18428), .D(
        n18427), .Y(n18431) );
  sky130_fd_sc_hd__nor2_1 U22953 ( .A(n18432), .B(n18431), .Y(n18440) );
  sky130_fd_sc_hd__nor4_1 U22954 ( .A(n18436), .B(n18435), .C(n18434), .D(
        n18433), .Y(n18438) );
  sky130_fd_sc_hd__o22ai_1 U22955 ( .A1(n18440), .A2(n18439), .B1(n18438), 
        .B2(n18437), .Y(n18449) );
  sky130_fd_sc_hd__nor4_1 U22956 ( .A(n18444), .B(n18443), .C(n18442), .D(
        n18441), .Y(n18447) );
  sky130_fd_sc_hd__a31oi_1 U22957 ( .A1(n18447), .A2(n18519), .A3(n18446), 
        .B1(n18445), .Y(n18448) );
  sky130_fd_sc_hd__o31a_1 U22958 ( .A1(n18450), .A2(n18449), .A3(n18448), .B1(
        n18798), .X(n18451) );
  sky130_fd_sc_hd__nor3_1 U22959 ( .A(n18453), .B(n18452), .C(n18451), .Y(
        n18454) );
  sky130_fd_sc_hd__nand2_1 U22960 ( .A(n18455), .B(n18454), .Y(n25313) );
  sky130_fd_sc_hd__nand2_1 U22961 ( .A(n25313), .B(n19087), .Y(n18458) );
  sky130_fd_sc_hd__a22oi_1 U22962 ( .A1(j202_soc_core_j22_cpu_id_opn_inst__9_), 
        .A2(n19088), .B1(j202_soc_core_j22_cpu_id_op2_v_), .B2(
        j202_soc_core_j22_cpu_id_op2_inst__9_), .Y(n18457) );
  sky130_fd_sc_hd__nand2_1 U22963 ( .A(n22541), .B(n19089), .Y(n18456) );
  sky130_fd_sc_hd__nand3_1 U22964 ( .A(n18458), .B(n18457), .C(n18456), .Y(
        n25385) );
  sky130_fd_sc_hd__nand2_1 U22965 ( .A(n25314), .B(n19087), .Y(n18461) );
  sky130_fd_sc_hd__a22oi_1 U22966 ( .A1(j202_soc_core_j22_cpu_id_opn_inst__10_), .A2(n19088), .B1(j202_soc_core_j22_cpu_id_op2_v_), .B2(
        j202_soc_core_j22_cpu_id_op2_inst__10_), .Y(n18460) );
  sky130_fd_sc_hd__nand2_1 U22967 ( .A(n20825), .B(n19089), .Y(n18459) );
  sky130_fd_sc_hd__nand3_1 U22968 ( .A(n18461), .B(n18460), .C(n18459), .Y(
        n25369) );
  sky130_fd_sc_hd__nand2b_1 U22969 ( .A_N(n22538), .B(n19089), .Y(n18464) );
  sky130_fd_sc_hd__a22oi_1 U22970 ( .A1(j202_soc_core_j22_cpu_id_opn_inst__11_), .A2(n19088), .B1(j202_soc_core_j22_cpu_id_op2_v_), .B2(
        j202_soc_core_j22_cpu_id_op2_inst__11_), .Y(n18463) );
  sky130_fd_sc_hd__nand2_1 U22971 ( .A(n25311), .B(n19087), .Y(n18462) );
  sky130_fd_sc_hd__nand3_1 U22972 ( .A(n18464), .B(n18463), .C(n18462), .Y(
        n25258) );
  sky130_fd_sc_hd__nand2_1 U22973 ( .A(n25312), .B(n19087), .Y(n18468) );
  sky130_fd_sc_hd__a22oi_1 U22974 ( .A1(j202_soc_core_j22_cpu_id_opn_inst__12_), .A2(n19088), .B1(j202_soc_core_j22_cpu_id_op2_v_), .B2(
        j202_soc_core_j22_cpu_id_op2_inst__12_), .Y(n18467) );
  sky130_fd_sc_hd__nand2_1 U22975 ( .A(n18465), .B(n19089), .Y(n18466) );
  sky130_fd_sc_hd__nand3_1 U22976 ( .A(n18468), .B(n18467), .C(n18466), .Y(
        n25315) );
  sky130_fd_sc_hd__nand2b_1 U22977 ( .A_N(n22542), .B(n19089), .Y(n18471) );
  sky130_fd_sc_hd__a22oi_1 U22978 ( .A1(j202_soc_core_j22_cpu_id_opn_inst__15_), .A2(n19088), .B1(j202_soc_core_j22_cpu_id_op2_v_), .B2(
        j202_soc_core_j22_cpu_id_op2_inst__15_), .Y(n18470) );
  sky130_fd_sc_hd__nand2_1 U22979 ( .A(n25388), .B(n19087), .Y(n18469) );
  sky130_fd_sc_hd__nand3_1 U22980 ( .A(n18471), .B(n18470), .C(n18469), .Y(
        n25316) );
  sky130_fd_sc_hd__xnor2_1 U22981 ( .A(n18473), .B(n18472), .Y(n18474) );
  sky130_fd_sc_hd__nand3_1 U22982 ( .A(n18476), .B(n18475), .C(n18474), .Y(
        n18477) );
  sky130_fd_sc_hd__nand2_1 U22983 ( .A(n22099), .B(n25731), .Y(n21904) );
  sky130_fd_sc_hd__nor2b_1 U22984 ( .B_N(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[2]), .Y(n23592) );
  sky130_fd_sc_hd__nand3_1 U22985 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[2]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_sck), .C(n25731), .Y(n23610) );
  sky130_fd_sc_hd__nand2_1 U22986 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[0]), .B(n20116), .Y(n23752) );
  sky130_fd_sc_hd__nand3_1 U22987 ( .A(n18479), .B(n23697), .C(n20116), .Y(
        n22862) );
  sky130_fd_sc_hd__nor2_1 U22988 ( .A(n22880), .B(n25392), .Y(n23734) );
  sky130_fd_sc_hd__nor2_1 U22989 ( .A(n23396), .B(
        j202_soc_core_wbqspiflash_00_spi_busy), .Y(n23590) );
  sky130_fd_sc_hd__nand2_1 U22990 ( .A(n23740), .B(n23590), .Y(n23591) );
  sky130_fd_sc_hd__nor2_1 U22991 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .B(
        j202_soc_core_wbqspiflash_00_lldriver_state[2]), .Y(n18480) );
  sky130_fd_sc_hd__nand3_1 U22992 ( .A(n18480), .B(
        j202_soc_core_wbqspiflash_00_lldriver_state[0]), .C(n25731), .Y(n21234) );
  sky130_fd_sc_hd__nor2_1 U22993 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[0]), .B(n23731), .Y(n22860) );
  sky130_fd_sc_hd__nor2_1 U22994 ( .A(n21324), .B(n22860), .Y(n23612) );
  sky130_fd_sc_hd__o21ai_1 U22995 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .A2(n23752), .B1(
        n23598), .Y(n25396) );
  sky130_fd_sc_hd__clkinv_1 U22996 ( .A(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[0]), .Y(n20431) );
  sky130_fd_sc_hd__nor2_1 U22997 ( .A(j202_soc_core_ahb2apb_00_state[0]), .B(
        n22767), .Y(n22766) );
  sky130_fd_sc_hd__nand2_1 U22998 ( .A(n22766), .B(n22768), .Y(n24781) );
  sky130_fd_sc_hd__nand2_1 U22999 ( .A(n18483), .B(n18482), .Y(n18484) );
  sky130_fd_sc_hd__xor2_1 U23000 ( .A(n18485), .B(n18484), .X(n22373) );
  sky130_fd_sc_hd__nand2_1 U23001 ( .A(n22373), .B(n19729), .Y(n18492) );
  sky130_fd_sc_hd__ha_1 U23002 ( .A(j202_soc_core_j22_cpu_pc[16]), .B(n18486), 
        .COUT(n18496), .SUM(n22377) );
  sky130_fd_sc_hd__nand2_1 U23003 ( .A(n22516), .B(n19737), .Y(n18488) );
  sky130_fd_sc_hd__a22oi_1 U23004 ( .A1(n19657), .A2(n22133), .B1(n19736), 
        .B2(n23298), .Y(n18487) );
  sky130_fd_sc_hd__nand2_1 U23005 ( .A(n18488), .B(n18487), .Y(n18489) );
  sky130_fd_sc_hd__a21oi_1 U23006 ( .A1(n22377), .A2(n19517), .B1(n18489), .Y(
        n18491) );
  sky130_fd_sc_hd__nand2_1 U23007 ( .A(n22377), .B(n19732), .Y(n18490) );
  sky130_fd_sc_hd__nand3_1 U23008 ( .A(n18492), .B(n18491), .C(n18490), .Y(
        n25260) );
  sky130_fd_sc_hd__nand2_1 U23009 ( .A(n11181), .B(n18493), .Y(n18495) );
  sky130_fd_sc_hd__xnor2_1 U23010 ( .A(n18495), .B(n18494), .Y(n22115) );
  sky130_fd_sc_hd__nand2_1 U23011 ( .A(n22115), .B(n19729), .Y(n18501) );
  sky130_fd_sc_hd__ha_1 U23012 ( .A(j202_soc_core_j22_cpu_pc[17]), .B(n18496), 
        .COUT(n13546), .SUM(n22118) );
  sky130_fd_sc_hd__nand2_1 U23013 ( .A(n22521), .B(n19737), .Y(n18498) );
  sky130_fd_sc_hd__a22oi_1 U23014 ( .A1(n19657), .A2(n21683), .B1(n19736), 
        .B2(n23301), .Y(n18497) );
  sky130_fd_sc_hd__nand2_1 U23015 ( .A(n18498), .B(n18497), .Y(n18499) );
  sky130_fd_sc_hd__a21oi_1 U23016 ( .A1(n22118), .A2(n19661), .B1(n18499), .Y(
        n18500) );
  sky130_fd_sc_hd__nand2_1 U23017 ( .A(n18501), .B(n18500), .Y(n25254) );
  sky130_fd_sc_hd__nand4_1 U23018 ( .A(n18504), .B(n18503), .C(n18502), .D(
        n25251), .Y(n18505) );
  sky130_fd_sc_hd__nor3_1 U23019 ( .A(n18506), .B(n18505), .C(n21074), .Y(
        n18507) );
  sky130_fd_sc_hd__nand3b_1 U23020 ( .A_N(n18509), .B(n18508), .C(n18507), .Y(
        n18510) );
  sky130_fd_sc_hd__nor3_1 U23021 ( .A(n18703), .B(n18511), .C(n18602), .Y(
        n18774) );
  sky130_fd_sc_hd__o31ai_1 U23022 ( .A1(n18585), .A2(n18516), .A3(n18526), 
        .B1(n18513), .Y(n18791) );
  sky130_fd_sc_hd__nand2_1 U23023 ( .A(n18514), .B(n18661), .Y(n18515) );
  sky130_fd_sc_hd__nor4_1 U23024 ( .A(n18562), .B(n18516), .C(n18672), .D(
        n18515), .Y(n18517) );
  sky130_fd_sc_hd__a31oi_1 U23025 ( .A1(n18573), .A2(n18517), .A3(n18569), 
        .B1(n18779), .Y(n18531) );
  sky130_fd_sc_hd__nand4_1 U23026 ( .A(n18545), .B(n18520), .C(n18519), .D(
        n18518), .Y(n18788) );
  sky130_fd_sc_hd__nand3_1 U23027 ( .A(n18566), .B(n18522), .C(n18521), .Y(
        n18523) );
  sky130_fd_sc_hd__nor4_1 U23028 ( .A(n18767), .B(n18777), .C(n18788), .D(
        n18523), .Y(n18529) );
  sky130_fd_sc_hd__nor2_1 U23029 ( .A(n18524), .B(n18584), .Y(n18700) );
  sky130_fd_sc_hd__nor4_1 U23030 ( .A(n18527), .B(n18768), .C(n18526), .D(
        n18525), .Y(n18528) );
  sky130_fd_sc_hd__o22ai_1 U23031 ( .A1(n18529), .A2(n18792), .B1(n18528), 
        .B2(n18771), .Y(n18530) );
  sky130_fd_sc_hd__nor4b_1 U23032 ( .D_N(n18791), .A(n18532), .B(n18531), .C(
        n18530), .Y(n18553) );
  sky130_fd_sc_hd__nand2_1 U23033 ( .A(n18533), .B(n18680), .Y(n18657) );
  sky130_fd_sc_hd__nor3_1 U23034 ( .A(n18534), .B(n18562), .C(n18657), .Y(
        n18535) );
  sky130_fd_sc_hd__a21oi_1 U23035 ( .A1(n18536), .A2(n18535), .B1(n18783), .Y(
        n18550) );
  sky130_fd_sc_hd__a31oi_1 U23036 ( .A1(n18538), .A2(n18537), .A3(n18566), 
        .B1(n18792), .Y(n18549) );
  sky130_fd_sc_hd__nand2_1 U23037 ( .A(n18574), .B(n18662), .Y(n18539) );
  sky130_fd_sc_hd__nor2_1 U23038 ( .A(n18768), .B(n18539), .Y(n18567) );
  sky130_fd_sc_hd__nor3b_1 U23039 ( .C_N(n18567), .A(n18540), .B(n18777), .Y(
        n18541) );
  sky130_fd_sc_hd__a31oi_1 U23040 ( .A1(n18542), .A2(n18604), .A3(n18541), 
        .B1(n18779), .Y(n18548) );
  sky130_fd_sc_hd__nor3_1 U23041 ( .A(n18564), .B(n18543), .C(n18673), .Y(
        n18786) );
  sky130_fd_sc_hd__and4_1 U23042 ( .A(n18569), .B(n18545), .C(n18589), .D(
        n18544), .X(n18546) );
  sky130_fd_sc_hd__a31oi_1 U23043 ( .A1(n18786), .A2(n18647), .A3(n18546), 
        .B1(n18771), .Y(n18547) );
  sky130_fd_sc_hd__nor4_1 U23044 ( .A(n18550), .B(n18549), .C(n18548), .D(
        n18547), .Y(n18551) );
  sky130_fd_sc_hd__o22a_1 U23045 ( .A1(n18553), .A2(n18552), .B1(n18551), .B2(
        n18720), .X(n18634) );
  sky130_fd_sc_hd__nor3_1 U23046 ( .A(n18673), .B(n18777), .C(n18657), .Y(
        n18684) );
  sky130_fd_sc_hd__nand2_1 U23047 ( .A(n18684), .B(n18569), .Y(n18576) );
  sky130_fd_sc_hd__nand4_1 U23048 ( .A(n18556), .B(n18555), .C(n18554), .D(
        n18660), .Y(n18590) );
  sky130_fd_sc_hd__nor2_1 U23049 ( .A(n18557), .B(n18702), .Y(n18785) );
  sky130_fd_sc_hd__nand4_1 U23050 ( .A(n18560), .B(n18785), .C(n18559), .D(
        n18558), .Y(n18561) );
  sky130_fd_sc_hd__nor3_1 U23051 ( .A(n18576), .B(n18590), .C(n18561), .Y(
        n18582) );
  sky130_fd_sc_hd__nor4_1 U23052 ( .A(n18564), .B(n18563), .C(n18562), .D(
        n18602), .Y(n18565) );
  sky130_fd_sc_hd__a31oi_1 U23053 ( .A1(n18567), .A2(n18566), .A3(n18565), 
        .B1(n18783), .Y(n18580) );
  sky130_fd_sc_hd__nor3_1 U23054 ( .A(n18687), .B(n18638), .C(n18568), .Y(
        n18658) );
  sky130_fd_sc_hd__nand2_1 U23055 ( .A(n18573), .B(n18569), .Y(n18570) );
  sky130_fd_sc_hd__nor3_1 U23056 ( .A(n18643), .B(n18697), .C(n18570), .Y(
        n18571) );
  sky130_fd_sc_hd__a31oi_1 U23057 ( .A1(n18658), .A2(n18572), .A3(n18571), 
        .B1(n18771), .Y(n18579) );
  sky130_fd_sc_hd__nand3_1 U23058 ( .A(n18574), .B(n18573), .C(n18593), .Y(
        n18575) );
  sky130_fd_sc_hd__nor3_1 U23059 ( .A(n18679), .B(n18576), .C(n18575), .Y(
        n18640) );
  sky130_fd_sc_hd__a31oi_1 U23060 ( .A1(n18640), .A2(n18577), .A3(n18675), 
        .B1(n18792), .Y(n18578) );
  sky130_fd_sc_hd__nor3_1 U23061 ( .A(n18580), .B(n18579), .C(n18578), .Y(
        n18581) );
  sky130_fd_sc_hd__nor2_1 U23063 ( .A(n18767), .B(n18583), .Y(n18715) );
  sky130_fd_sc_hd__nor4_1 U23064 ( .A(n18770), .B(n18710), .C(n18585), .D(
        n18584), .Y(n18586) );
  sky130_fd_sc_hd__a31oi_1 U23065 ( .A1(n18715), .A2(n18587), .A3(n18586), 
        .B1(n18792), .Y(n18608) );
  sky130_fd_sc_hd__nand3_1 U23066 ( .A(n18589), .B(n18648), .C(n18588), .Y(
        n18671) );
  sky130_fd_sc_hd__nor4_1 U23067 ( .A(n18701), .B(n18671), .C(n18591), .D(
        n18590), .Y(n18600) );
  sky130_fd_sc_hd__nand3_1 U23068 ( .A(n18594), .B(n18593), .C(n18592), .Y(
        n18689) );
  sky130_fd_sc_hd__nand3b_1 U23069 ( .A_N(n18657), .B(n18786), .C(n18595), .Y(
        n18596) );
  sky130_fd_sc_hd__nor4_1 U23070 ( .A(n18598), .B(n18597), .C(n18689), .D(
        n18596), .Y(n18599) );
  sky130_fd_sc_hd__o22ai_1 U23071 ( .A1(n18600), .A2(n18783), .B1(n18599), 
        .B2(n18779), .Y(n18607) );
  sky130_fd_sc_hd__nor3_1 U23072 ( .A(n18766), .B(n18602), .C(n18601), .Y(
        n18603) );
  sky130_fd_sc_hd__a31oi_1 U23073 ( .A1(n18604), .A2(n18658), .A3(n18603), 
        .B1(n18771), .Y(n18606) );
  sky130_fd_sc_hd__o31a_1 U23074 ( .A1(n18608), .A2(n18607), .A3(n18606), .B1(
        n18605), .X(n18609) );
  sky130_fd_sc_hd__a21oi_1 U23075 ( .A1(n18611), .A2(n18610), .B1(n18609), .Y(
        n18633) );
  sky130_fd_sc_hd__a22o_1 U23076 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[14]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[78]), .X(n18612) );
  sky130_fd_sc_hd__a21oi_1 U23077 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[110]), .B1(n18612), .Y(n18614) );
  sky130_fd_sc_hd__a22oi_1 U23078 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[174]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[142]), .Y(n18613) );
  sky130_fd_sc_hd__a21oi_1 U23079 ( .A1(n18614), .A2(n18613), .B1(n18736), .Y(
        n18625) );
  sky130_fd_sc_hd__a22oi_1 U23080 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[270]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[46]), .Y(n18623) );
  sky130_fd_sc_hd__a22o_1 U23081 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[302]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[334]), .X(n18615) );
  sky130_fd_sc_hd__a21oi_1 U23082 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[366]), .B1(n18615), .Y(n18622) );
  sky130_fd_sc_hd__nand2_1 U23083 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[238]), .Y(n18619) );
  sky130_fd_sc_hd__a21oi_1 U23084 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[462]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n18618) );
  sky130_fd_sc_hd__nand2_1 U23085 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[398]), .Y(n18617) );
  sky130_fd_sc_hd__nand2_1 U23086 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[430]), .Y(n18616) );
  sky130_fd_sc_hd__nand4_1 U23087 ( .A(n18619), .B(n18618), .C(n18617), .D(
        n18616), .Y(n18620) );
  sky130_fd_sc_hd__a21oi_1 U23088 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[206]), .B1(n18620), .Y(n18621) );
  sky130_fd_sc_hd__nand3_1 U23089 ( .A(n18623), .B(n18622), .C(n18621), .Y(
        n18624) );
  sky130_fd_sc_hd__o22ai_1 U23090 ( .A1(j202_soc_core_memory0_ram_dout0[494]), 
        .A2(n18758), .B1(n18625), .B2(n18624), .Y(n18627) );
  sky130_fd_sc_hd__a22oi_1 U23091 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[78]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[46]), .Y(n18626) );
  sky130_fd_sc_hd__a21oi_1 U23093 ( .A1(n18629), .A2(
        j202_soc_core_bldc_core_00_pwm_duty[2]), .B1(n18628), .Y(n18631) );
  sky130_fd_sc_hd__a22oi_1 U23094 ( .A1(n18724), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[110]), .B1(n18725), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[14]), .Y(n18630) );
  sky130_fd_sc_hd__nand3_1 U23095 ( .A(n18634), .B(n18633), .C(n18632), .Y(
        n25310) );
  sky130_fd_sc_hd__nand2_1 U23096 ( .A(n25310), .B(n19087), .Y(n18637) );
  sky130_fd_sc_hd__a22oi_1 U23097 ( .A1(j202_soc_core_j22_cpu_id_opn_inst__14_), .A2(n19088), .B1(j202_soc_core_j22_cpu_id_op2_v_), .B2(
        j202_soc_core_j22_cpu_id_op2_inst__14_), .Y(n18636) );
  sky130_fd_sc_hd__nand2_1 U23098 ( .A(n22517), .B(n19089), .Y(n18635) );
  sky130_fd_sc_hd__nand3_1 U23099 ( .A(n18637), .B(n18636), .C(n18635), .Y(
        n25304) );
  sky130_fd_sc_hd__nor2_1 U23100 ( .A(n18766), .B(n18638), .Y(n18653) );
  sky130_fd_sc_hd__nand4_1 U23101 ( .A(n18640), .B(n18653), .C(n18642), .D(
        n18639), .Y(n18650) );
  sky130_fd_sc_hd__nand3_1 U23102 ( .A(n18700), .B(n18782), .C(n18642), .Y(
        n18787) );
  sky130_fd_sc_hd__nor4_1 U23103 ( .A(n18645), .B(n18644), .C(n18643), .D(
        n18787), .Y(n18646) );
  sky130_fd_sc_hd__a31oi_1 U23104 ( .A1(n18648), .A2(n18647), .A3(n18646), 
        .B1(n18783), .Y(n18649) );
  sky130_fd_sc_hd__a21oi_1 U23105 ( .A1(n18651), .A2(n18650), .B1(n18649), .Y(
        n18669) );
  sky130_fd_sc_hd__nand4_1 U23106 ( .A(n18654), .B(n18653), .C(n18652), .D(
        n18660), .Y(n18656) );
  sky130_fd_sc_hd__o21ai_1 U23107 ( .A1(n18657), .A2(n18656), .B1(n18655), .Y(
        n18668) );
  sky130_fd_sc_hd__nand2_1 U23108 ( .A(n18659), .B(n18658), .Y(n18707) );
  sky130_fd_sc_hd__nand4_1 U23109 ( .A(n18663), .B(n18662), .C(n18661), .D(
        n18660), .Y(n18665) );
  sky130_fd_sc_hd__a31oi_1 U23111 ( .A1(n18669), .A2(n18668), .A3(n18667), 
        .B1(n18666), .Y(n18765) );
  sky130_fd_sc_hd__nor4_1 U23112 ( .A(n18674), .B(n18673), .C(n18672), .D(
        n18671), .Y(n18676) );
  sky130_fd_sc_hd__a31oi_1 U23113 ( .A1(n18677), .A2(n18676), .A3(n18675), 
        .B1(n18783), .Y(n18696) );
  sky130_fd_sc_hd__nor3_1 U23114 ( .A(n18703), .B(n18679), .C(n18678), .Y(
        n18682) );
  sky130_fd_sc_hd__a31oi_1 U23115 ( .A1(n18682), .A2(n18681), .A3(n18680), 
        .B1(n18771), .Y(n18695) );
  sky130_fd_sc_hd__nand2_1 U23116 ( .A(n18684), .B(n18683), .Y(n18691) );
  sky130_fd_sc_hd__nor4_1 U23117 ( .A(n18687), .B(n18691), .C(n18686), .D(
        n18685), .Y(n18693) );
  sky130_fd_sc_hd__nor4_1 U23118 ( .A(n18691), .B(n18690), .C(n18689), .D(
        n18688), .Y(n18692) );
  sky130_fd_sc_hd__o22ai_1 U23119 ( .A1(n18693), .A2(n18792), .B1(n18692), 
        .B2(n18779), .Y(n18694) );
  sky130_fd_sc_hd__nor3_1 U23120 ( .A(n18696), .B(n18695), .C(n18694), .Y(
        n18723) );
  sky130_fd_sc_hd__nor3_1 U23121 ( .A(n18701), .B(n18708), .C(n18697), .Y(
        n18699) );
  sky130_fd_sc_hd__a31oi_1 U23122 ( .A1(n18700), .A2(n18699), .A3(n18698), 
        .B1(n18771), .Y(n18719) );
  sky130_fd_sc_hd__nor4_1 U23123 ( .A(n18704), .B(n18703), .C(n18702), .D(
        n18701), .Y(n18705) );
  sky130_fd_sc_hd__a21oi_1 U23124 ( .A1(n18706), .A2(n18705), .B1(n18792), .Y(
        n18718) );
  sky130_fd_sc_hd__nor4_1 U23125 ( .A(n18710), .B(n18709), .C(n18708), .D(
        n18707), .Y(n18711) );
  sky130_fd_sc_hd__a21oi_1 U23126 ( .A1(n18712), .A2(n18711), .B1(n18779), .Y(
        n18717) );
  sky130_fd_sc_hd__a31oi_1 U23127 ( .A1(n18715), .A2(n18714), .A3(n18713), 
        .B1(n18783), .Y(n18716) );
  sky130_fd_sc_hd__nor4_1 U23128 ( .A(n18719), .B(n18718), .C(n18717), .D(
        n18716), .Y(n18721) );
  sky130_fd_sc_hd__o22ai_1 U23129 ( .A1(n18723), .A2(n18722), .B1(n18721), 
        .B2(n18720), .Y(n18764) );
  sky130_fd_sc_hd__a22oi_1 U23130 ( .A1(n18725), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[13]), .B1(n18724), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[109]), .Y(n18729) );
  sky130_fd_sc_hd__a22oi_1 U23131 ( .A1(n18727), .A2(
        j202_soc_core_ahblite_interconnect_s_hrdata[77]), .B1(n18726), .B2(
        j202_soc_core_ahblite_interconnect_s_hrdata[45]), .Y(n18728) );
  sky130_fd_sc_hd__nand2_1 U23132 ( .A(n18729), .B(n18728), .Y(n18763) );
  sky130_fd_sc_hd__a22o_1 U23133 ( .A1(n18731), .A2(
        j202_soc_core_memory0_ram_dout0[13]), .B1(n18730), .B2(
        j202_soc_core_memory0_ram_dout0[77]), .X(n18732) );
  sky130_fd_sc_hd__a21oi_1 U23134 ( .A1(n18733), .A2(
        j202_soc_core_memory0_ram_dout0[109]), .B1(n18732), .Y(n18738) );
  sky130_fd_sc_hd__a22oi_1 U23135 ( .A1(n18735), .A2(
        j202_soc_core_memory0_ram_dout0[173]), .B1(n18734), .B2(
        j202_soc_core_memory0_ram_dout0[141]), .Y(n18737) );
  sky130_fd_sc_hd__a21oi_1 U23136 ( .A1(n18738), .A2(n18737), .B1(n18736), .Y(
        n18757) );
  sky130_fd_sc_hd__a22oi_1 U23137 ( .A1(n18062), .A2(
        j202_soc_core_memory0_ram_dout0[269]), .B1(n18739), .B2(
        j202_soc_core_memory0_ram_dout0[45]), .Y(n18755) );
  sky130_fd_sc_hd__a22o_1 U23138 ( .A1(n18741), .A2(
        j202_soc_core_memory0_ram_dout0[301]), .B1(n18740), .B2(
        j202_soc_core_memory0_ram_dout0[333]), .X(n18742) );
  sky130_fd_sc_hd__a21oi_1 U23139 ( .A1(n18743), .A2(
        j202_soc_core_memory0_ram_dout0[365]), .B1(n18742), .Y(n18754) );
  sky130_fd_sc_hd__nand2_1 U23140 ( .A(n18744), .B(
        j202_soc_core_memory0_ram_dout0[237]), .Y(n18750) );
  sky130_fd_sc_hd__a21oi_1 U23141 ( .A1(
        j202_soc_core_memory0_ram_dout0_sel[14]), .A2(
        j202_soc_core_memory0_ram_dout0[461]), .B1(
        j202_soc_core_memory0_ram_dout0_sel[15]), .Y(n18749) );
  sky130_fd_sc_hd__nand2_1 U23142 ( .A(n18745), .B(
        j202_soc_core_memory0_ram_dout0[397]), .Y(n18748) );
  sky130_fd_sc_hd__nand2_1 U23143 ( .A(n18746), .B(
        j202_soc_core_memory0_ram_dout0[429]), .Y(n18747) );
  sky130_fd_sc_hd__nand4_1 U23144 ( .A(n18750), .B(n18749), .C(n18748), .D(
        n18747), .Y(n18751) );
  sky130_fd_sc_hd__a21oi_1 U23145 ( .A1(n18752), .A2(
        j202_soc_core_memory0_ram_dout0[205]), .B1(n18751), .Y(n18753) );
  sky130_fd_sc_hd__nand3_1 U23146 ( .A(n18755), .B(n18754), .C(n18753), .Y(
        n18756) );
  sky130_fd_sc_hd__o22ai_1 U23147 ( .A1(j202_soc_core_memory0_ram_dout0[493]), 
        .A2(n18758), .B1(n18757), .B2(n18756), .Y(n18760) );
  sky130_fd_sc_hd__o22ai_1 U23148 ( .A1(n18761), .A2(n18760), .B1(n18759), 
        .B2(n25186), .Y(n18762) );
  sky130_fd_sc_hd__nor4_1 U23149 ( .A(n18765), .B(n18764), .C(n18763), .D(
        n18762), .Y(n18801) );
  sky130_fd_sc_hd__nor2_1 U23150 ( .A(n18766), .B(n18790), .Y(n18773) );
  sky130_fd_sc_hd__nor4_1 U23151 ( .A(n18770), .B(n18769), .C(n18768), .D(
        n18767), .Y(n18772) );
  sky130_fd_sc_hd__a31oi_1 U23152 ( .A1(n18774), .A2(n18773), .A3(n18772), 
        .B1(n18771), .Y(n18797) );
  sky130_fd_sc_hd__nor4_1 U23153 ( .A(n18778), .B(n18777), .C(n18776), .D(
        n18775), .Y(n18780) );
  sky130_fd_sc_hd__a31oi_1 U23154 ( .A1(n18782), .A2(n18781), .A3(n18780), 
        .B1(n18779), .Y(n18796) );
  sky130_fd_sc_hd__a31oi_1 U23155 ( .A1(n18786), .A2(n18785), .A3(n18784), 
        .B1(n18783), .Y(n18795) );
  sky130_fd_sc_hd__nor4_1 U23156 ( .A(n18790), .B(n18789), .C(n18788), .D(
        n18787), .Y(n18793) );
  sky130_fd_sc_hd__nor4_1 U23158 ( .A(n18797), .B(n18796), .C(n18795), .D(
        n18794), .Y(n18799) );
  sky130_fd_sc_hd__nand2b_1 U23159 ( .A_N(n18799), .B(n18798), .Y(n18800) );
  sky130_fd_sc_hd__nand2_1 U23160 ( .A(n18801), .B(n18800), .Y(n25309) );
  sky130_fd_sc_hd__nand2_1 U23161 ( .A(n25309), .B(n19087), .Y(n18804) );
  sky130_fd_sc_hd__a22oi_1 U23162 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        j202_soc_core_j22_cpu_id_op2_inst__13_), .B1(n19088), .B2(
        j202_soc_core_j22_cpu_id_opn_inst__13_), .Y(n18803) );
  sky130_fd_sc_hd__nand2_1 U23163 ( .A(n20546), .B(n19089), .Y(n18802) );
  sky130_fd_sc_hd__nand3_1 U23164 ( .A(n18804), .B(n18803), .C(n18802), .Y(
        n25303) );
  sky130_fd_sc_hd__nand2_1 U23165 ( .A(n18807), .B(n18806), .Y(n18808) );
  sky130_fd_sc_hd__xor2_1 U23166 ( .A(n18809), .B(n18808), .X(n21861) );
  sky130_fd_sc_hd__nand2_1 U23167 ( .A(n21861), .B(n19729), .Y(n18816) );
  sky130_fd_sc_hd__ha_1 U23168 ( .A(j202_soc_core_j22_cpu_pc[14]), .B(n18810), 
        .COUT(n19656), .SUM(n21864) );
  sky130_fd_sc_hd__nand2_1 U23169 ( .A(n25310), .B(n19737), .Y(n18812) );
  sky130_fd_sc_hd__a22oi_1 U23170 ( .A1(n19657), .A2(n21152), .B1(n19736), 
        .B2(n22156), .Y(n18811) );
  sky130_fd_sc_hd__nand2_1 U23171 ( .A(n18812), .B(n18811), .Y(n18813) );
  sky130_fd_sc_hd__a21oi_1 U23172 ( .A1(n21864), .A2(n19517), .B1(n18813), .Y(
        n18815) );
  sky130_fd_sc_hd__nand2_1 U23173 ( .A(n21864), .B(n19732), .Y(n18814) );
  sky130_fd_sc_hd__nand3_1 U23174 ( .A(n18816), .B(n18815), .C(n18814), .Y(
        n25273) );
  sky130_fd_sc_hd__nand2_1 U23175 ( .A(n18819), .B(n18818), .Y(n18820) );
  sky130_fd_sc_hd__xor2_1 U23176 ( .A(n18821), .B(n18820), .X(n22066) );
  sky130_fd_sc_hd__nand2_1 U23177 ( .A(n22066), .B(n19729), .Y(n18827) );
  sky130_fd_sc_hd__ha_1 U23178 ( .A(j202_soc_core_j22_cpu_pc[12]), .B(n18822), 
        .COUT(n18831), .SUM(n22070) );
  sky130_fd_sc_hd__o22a_1 U23179 ( .A1(n22064), .A2(n18948), .B1(n22560), .B2(
        n19731), .X(n18824) );
  sky130_fd_sc_hd__nand2_1 U23180 ( .A(n25312), .B(n19737), .Y(n18823) );
  sky130_fd_sc_hd__o211ai_1 U23181 ( .A1(n22064), .A2(n19083), .B1(n18824), 
        .C1(n18823), .Y(n18825) );
  sky130_fd_sc_hd__a21oi_1 U23182 ( .A1(n22070), .A2(n19661), .B1(n18825), .Y(
        n18826) );
  sky130_fd_sc_hd__nand2_1 U23183 ( .A(n18827), .B(n18826), .Y(n25272) );
  sky130_fd_sc_hd__nand2_1 U23184 ( .A(n11195), .B(n18828), .Y(n18830) );
  sky130_fd_sc_hd__xnor2_1 U23185 ( .A(n18830), .B(n18829), .Y(n22302) );
  sky130_fd_sc_hd__nand2_1 U23186 ( .A(n22302), .B(n19729), .Y(n18836) );
  sky130_fd_sc_hd__ha_1 U23187 ( .A(j202_soc_core_j22_cpu_pc[13]), .B(n18831), 
        .COUT(n18810), .SUM(n22298) );
  sky130_fd_sc_hd__o22a_1 U23188 ( .A1(n22300), .A2(n18948), .B1(n22561), .B2(
        n19731), .X(n18833) );
  sky130_fd_sc_hd__nand2_1 U23189 ( .A(n25309), .B(n19737), .Y(n18832) );
  sky130_fd_sc_hd__o211ai_1 U23190 ( .A1(n22300), .A2(n19083), .B1(n18833), 
        .C1(n18832), .Y(n18834) );
  sky130_fd_sc_hd__a21oi_1 U23191 ( .A1(n22298), .A2(n19661), .B1(n18834), .Y(
        n18835) );
  sky130_fd_sc_hd__nand2_1 U23192 ( .A(n18839), .B(n18838), .Y(n18843) );
  sky130_fd_sc_hd__xnor2_1 U23194 ( .A(n18843), .B(n18842), .Y(n22353) );
  sky130_fd_sc_hd__nand2_1 U23195 ( .A(n22353), .B(n19729), .Y(n18851) );
  sky130_fd_sc_hd__ha_1 U23196 ( .A(j202_soc_core_j22_cpu_pc[11]), .B(n18844), 
        .COUT(n18822), .SUM(n22349) );
  sky130_fd_sc_hd__nand2_1 U23197 ( .A(n22349), .B(n19732), .Y(n18849) );
  sky130_fd_sc_hd__nand2_1 U23198 ( .A(n22349), .B(n19517), .Y(n18848) );
  sky130_fd_sc_hd__o22a_1 U23199 ( .A1(n22351), .A2(n18948), .B1(n22564), .B2(
        n19731), .X(n18845) );
  sky130_fd_sc_hd__a21oi_1 U23201 ( .A1(n25311), .A2(n19737), .B1(n18846), .Y(
        n18847) );
  sky130_fd_sc_hd__and3_1 U23202 ( .A(n18849), .B(n18848), .C(n18847), .X(
        n18850) );
  sky130_fd_sc_hd__nor2_1 U23203 ( .A(n25272), .B(n25271), .Y(n21244) );
  sky130_fd_sc_hd__nand2_1 U23204 ( .A(n23241), .B(n24894), .Y(n22827) );
  sky130_fd_sc_hd__nand2b_1 U23205 ( .A_N(n11036), .B(n22827), .Y(n21208) );
  sky130_fd_sc_hd__nand3_1 U23206 ( .A(n19833), .B(n21245), .C(n19832), .Y(
        n19802) );
  sky130_fd_sc_hd__nor2_1 U23207 ( .A(n19836), .B(n19802), .Y(n25321) );
  sky130_fd_sc_hd__a21oi_1 U23208 ( .A1(n18854), .A2(n18853), .B1(n18852), .Y(
        n18858) );
  sky130_fd_sc_hd__nand2_1 U23209 ( .A(n18856), .B(n18855), .Y(n18857) );
  sky130_fd_sc_hd__xor2_1 U23210 ( .A(n18858), .B(n18857), .X(n21721) );
  sky130_fd_sc_hd__nand2_1 U23211 ( .A(n21721), .B(n20030), .Y(n18864) );
  sky130_fd_sc_hd__nand2_1 U23212 ( .A(n18861), .B(n18860), .Y(n18862) );
  sky130_fd_sc_hd__xor2_1 U23213 ( .A(n18975), .B(n18862), .X(n19810) );
  sky130_fd_sc_hd__a22oi_1 U23214 ( .A1(j202_soc_core_j22_cpu_ml_mach[11]), 
        .A2(n20032), .B1(n19810), .B2(n20025), .Y(n18863) );
  sky130_fd_sc_hd__nand2_1 U23215 ( .A(n18864), .B(n18863), .Y(n21961) );
  sky130_fd_sc_hd__nand2_1 U23216 ( .A(n21961), .B(n22125), .Y(n18872) );
  sky130_fd_sc_hd__nand2_1 U23217 ( .A(n18866), .B(n18865), .Y(n18868) );
  sky130_fd_sc_hd__xnor2_1 U23218 ( .A(n18868), .B(n18867), .Y(n21958) );
  sky130_fd_sc_hd__o22ai_1 U23219 ( .A1(n20043), .A2(n21960), .B1(n18869), 
        .B2(n20012), .Y(n18870) );
  sky130_fd_sc_hd__a21oi_1 U23220 ( .A1(n21958), .A2(n20016), .B1(n18870), .Y(
        n18871) );
  sky130_fd_sc_hd__nand2_1 U23221 ( .A(n18872), .B(n18871), .Y(n20594) );
  sky130_fd_sc_hd__nand2_1 U23222 ( .A(n20594), .B(n20019), .Y(n18938) );
  sky130_fd_sc_hd__nand2_1 U23223 ( .A(n18875), .B(n18874), .Y(n18877) );
  sky130_fd_sc_hd__xnor2_1 U23224 ( .A(n18877), .B(n18876), .Y(n21698) );
  sky130_fd_sc_hd__nand2_1 U23225 ( .A(n21698), .B(n20030), .Y(n18882) );
  sky130_fd_sc_hd__nand2_1 U23226 ( .A(n18879), .B(n18878), .Y(n18880) );
  sky130_fd_sc_hd__xnor2_1 U23227 ( .A(n18880), .B(n19007), .Y(n20041) );
  sky130_fd_sc_hd__a22oi_1 U23228 ( .A1(j202_soc_core_j22_cpu_ml_mach[3]), 
        .A2(n20032), .B1(n20041), .B2(n20025), .Y(n18881) );
  sky130_fd_sc_hd__nand2_1 U23229 ( .A(n18882), .B(n18881), .Y(n22003) );
  sky130_fd_sc_hd__nand2_1 U23230 ( .A(n22003), .B(n22125), .Y(n18891) );
  sky130_fd_sc_hd__nand2_1 U23231 ( .A(n18885), .B(n18884), .Y(n18887) );
  sky130_fd_sc_hd__xor2_1 U23232 ( .A(n18887), .B(n18886), .X(n22000) );
  sky130_fd_sc_hd__o22ai_1 U23233 ( .A1(n20043), .A2(n22002), .B1(n18888), 
        .B2(n20012), .Y(n18889) );
  sky130_fd_sc_hd__a21oi_1 U23234 ( .A1(n22000), .A2(n20016), .B1(n18889), .Y(
        n18890) );
  sky130_fd_sc_hd__nand2_1 U23235 ( .A(n18891), .B(n18890), .Y(n19318) );
  sky130_fd_sc_hd__nand2_1 U23236 ( .A(n19318), .B(n21137), .Y(n18911) );
  sky130_fd_sc_hd__nand2_1 U23237 ( .A(n22522), .B(n19893), .Y(n18894) );
  sky130_fd_sc_hd__a2bb2oi_1 U23238 ( .B1(n19889), .B2(n25311), .A1_N(n19891), 
        .A2_N(n22538), .Y(n18893) );
  sky130_fd_sc_hd__nand2_1 U23239 ( .A(n25253), .B(n19895), .Y(n18892) );
  sky130_fd_sc_hd__nand2_1 U23240 ( .A(n22583), .B(n21170), .Y(n18895) );
  sky130_fd_sc_hd__o211ai_1 U23241 ( .A1(n21027), .A2(n22583), .B1(n21174), 
        .C1(n18895), .Y(n18907) );
  sky130_fd_sc_hd__nand2_1 U23242 ( .A(n22010), .B(n21178), .Y(n18905) );
  sky130_fd_sc_hd__a22oi_1 U23243 ( .A1(n20711), .A2(n21963), .B1(n21164), 
        .B2(n22141), .Y(n18904) );
  sky130_fd_sc_hd__a2bb2oi_1 U23244 ( .B1(n23307), .B2(n20716), .A1_N(n22351), 
        .A2_N(n20712), .Y(n18903) );
  sky130_fd_sc_hd__nor2_1 U23245 ( .A(n22711), .B(n22488), .Y(n22441) );
  sky130_fd_sc_hd__nand2_1 U23246 ( .A(n22488), .B(n22711), .Y(n22436) );
  sky130_fd_sc_hd__nand3_1 U23247 ( .A(n22651), .B(n22436), .C(n21147), .Y(
        n18897) );
  sky130_fd_sc_hd__nand2_1 U23248 ( .A(n22441), .B(n21089), .Y(n18896) );
  sky130_fd_sc_hd__o211ai_1 U23249 ( .A1(n21145), .A2(n22179), .B1(n18897), 
        .C1(n18896), .Y(n18898) );
  sky130_fd_sc_hd__a21oi_1 U23250 ( .A1(n21029), .A2(n22483), .B1(n18898), .Y(
        n18900) );
  sky130_fd_sc_hd__a2bb2oi_1 U23251 ( .B1(n21156), .B2(n20689), .A1_N(n22487), 
        .A2_N(n21155), .Y(n18899) );
  sky130_fd_sc_hd__o211ai_1 U23252 ( .A1(n22580), .A2(n21163), .B1(n18900), 
        .C1(n18899), .Y(n18901) );
  sky130_fd_sc_hd__a21oi_1 U23253 ( .A1(n19884), .A2(n22179), .B1(n18901), .Y(
        n18902) );
  sky130_fd_sc_hd__nand4_1 U23254 ( .A(n18905), .B(n18904), .C(n18903), .D(
        n18902), .Y(n18906) );
  sky130_fd_sc_hd__a21oi_1 U23255 ( .A1(n22013), .A2(n18907), .B1(n18906), .Y(
        n18910) );
  sky130_fd_sc_hd__nand2_1 U23257 ( .A(n18908), .B(n22583), .Y(n18909) );
  sky130_fd_sc_hd__nand2_1 U23258 ( .A(n22006), .B(n19905), .Y(n20065) );
  sky130_fd_sc_hd__nand2_1 U23259 ( .A(n18912), .B(n19969), .Y(n18923) );
  sky130_fd_sc_hd__o22ai_1 U23260 ( .A1(n18914), .A2(n19971), .B1(n18913), 
        .B2(n19975), .Y(n18915) );
  sky130_fd_sc_hd__a21oi_1 U23261 ( .A1(n19842), .A2(
        j202_soc_core_j22_cpu_rf_gpr[3]), .B1(n18915), .Y(n18922) );
  sky130_fd_sc_hd__o22ai_1 U23262 ( .A1(n18917), .A2(n19981), .B1(n18916), 
        .B2(n19986), .Y(n18920) );
  sky130_fd_sc_hd__o2bb2ai_1 U23263 ( .B1(n18918), .B2(n19977), .A1_N(
        j202_soc_core_j22_cpu_rf_vbr[3]), .A2_N(n19985), .Y(n18919) );
  sky130_fd_sc_hd__nor2_1 U23264 ( .A(n18920), .B(n18919), .Y(n18921) );
  sky130_fd_sc_hd__nand3_1 U23265 ( .A(n18923), .B(n18922), .C(n18921), .Y(
        n20063) );
  sky130_fd_sc_hd__nand2_1 U23266 ( .A(n20063), .B(n19285), .Y(n18924) );
  sky130_fd_sc_hd__nand2_1 U23267 ( .A(n18925), .B(n19969), .Y(n18936) );
  sky130_fd_sc_hd__o22ai_1 U23268 ( .A1(n18927), .A2(n19977), .B1(n19971), 
        .B2(n18926), .Y(n18928) );
  sky130_fd_sc_hd__a21oi_1 U23269 ( .A1(n19842), .A2(
        j202_soc_core_j22_cpu_rf_gpr[11]), .B1(n18928), .Y(n18935) );
  sky130_fd_sc_hd__o22ai_1 U23270 ( .A1(n18930), .A2(n19975), .B1(n18929), 
        .B2(n19986), .Y(n18933) );
  sky130_fd_sc_hd__o2bb2ai_1 U23271 ( .B1(n18931), .B2(n19981), .A1_N(
        j202_soc_core_j22_cpu_rf_vbr[11]), .A2_N(n19985), .Y(n18932) );
  sky130_fd_sc_hd__nor2_1 U23272 ( .A(n18933), .B(n18932), .Y(n18934) );
  sky130_fd_sc_hd__nand3_1 U23273 ( .A(n18936), .B(n18935), .C(n18934), .Y(
        n19828) );
  sky130_fd_sc_hd__nand2_1 U23274 ( .A(n19828), .B(n20020), .Y(n18937) );
  sky130_fd_sc_hd__nand3_1 U23275 ( .A(n18938), .B(n19830), .C(n18937), .Y(
        n25343) );
  sky130_fd_sc_hd__nand2_1 U23276 ( .A(n19509), .B(n19507), .Y(n18944) );
  sky130_fd_sc_hd__o21ai_1 U23277 ( .A1(n18943), .A2(n19725), .B1(n18942), .Y(
        n19510) );
  sky130_fd_sc_hd__xnor2_1 U23278 ( .A(n18944), .B(n19510), .Y(n22316) );
  sky130_fd_sc_hd__nand2_1 U23279 ( .A(n22316), .B(n19729), .Y(n18951) );
  sky130_fd_sc_hd__ha_1 U23280 ( .A(j202_soc_core_j22_cpu_pc[9]), .B(n18945), 
        .COUT(n19516), .SUM(n22313) );
  sky130_fd_sc_hd__a2bb2oi_1 U23281 ( .B1(n19517), .B2(n22313), .A1_N(n22314), 
        .A2_N(n19083), .Y(n18947) );
  sky130_fd_sc_hd__a22oi_1 U23282 ( .A1(n19657), .A2(n20699), .B1(n22313), 
        .B2(n19732), .Y(n18946) );
  sky130_fd_sc_hd__o211ai_1 U23283 ( .A1(n22314), .A2(n18948), .B1(n18947), 
        .C1(n18946), .Y(n18949) );
  sky130_fd_sc_hd__a21oi_1 U23284 ( .A1(n25313), .A2(n19737), .B1(n18949), .Y(
        n18950) );
  sky130_fd_sc_hd__nand2_1 U23285 ( .A(n18951), .B(n18950), .Y(n25375) );
  sky130_fd_sc_hd__o22ai_1 U23286 ( .A1(n18953), .A2(n19977), .B1(n19971), 
        .B2(n18952), .Y(n18954) );
  sky130_fd_sc_hd__a21oi_1 U23287 ( .A1(n19842), .A2(
        j202_soc_core_j22_cpu_rf_gpr[14]), .B1(n18954), .Y(n18960) );
  sky130_fd_sc_hd__a22oi_1 U23288 ( .A1(n19843), .A2(
        j202_soc_core_j22_cpu_rf_tmp[14]), .B1(n19985), .B2(
        j202_soc_core_j22_cpu_rf_vbr[14]), .Y(n18959) );
  sky130_fd_sc_hd__clkinv_1 U23289 ( .A(n19986), .Y(n18955) );
  sky130_fd_sc_hd__nand2_1 U23290 ( .A(n18955), .B(
        j202_soc_core_j22_cpu_rf_gpr[494]), .Y(n18958) );
  sky130_fd_sc_hd__clkinv_1 U23291 ( .A(n19975), .Y(n18956) );
  sky130_fd_sc_hd__nand2_1 U23292 ( .A(n18956), .B(
        j202_soc_core_j22_cpu_rf_gbr[14]), .Y(n18957) );
  sky130_fd_sc_hd__nand4_1 U23293 ( .A(n18960), .B(n18959), .C(n18958), .D(
        n18957), .Y(n18961) );
  sky130_fd_sc_hd__a21oi_1 U23294 ( .A1(n18962), .A2(n19969), .B1(n18961), .Y(
        n19765) );
  sky130_fd_sc_hd__a21oi_1 U23295 ( .A1(n19920), .A2(n18966), .B1(n18965), .Y(
        n18971) );
  sky130_fd_sc_hd__nand2_1 U23296 ( .A(n18969), .B(n18968), .Y(n18970) );
  sky130_fd_sc_hd__xor2_1 U23297 ( .A(n18971), .B(n18970), .X(n21699) );
  sky130_fd_sc_hd__nand2_1 U23298 ( .A(n21699), .B(n20030), .Y(n18985) );
  sky130_fd_sc_hd__o21ai_1 U23299 ( .A1(n18976), .A2(n18975), .B1(n18974), .Y(
        n19102) );
  sky130_fd_sc_hd__a21oi_1 U23300 ( .A1(n19102), .A2(n19101), .B1(n18978), .Y(
        n18983) );
  sky130_fd_sc_hd__nand2_1 U23301 ( .A(n18981), .B(n18980), .Y(n18982) );
  sky130_fd_sc_hd__xor2_1 U23302 ( .A(n18983), .B(n18982), .X(n19751) );
  sky130_fd_sc_hd__a22oi_1 U23303 ( .A1(j202_soc_core_j22_cpu_ml_mach[14]), 
        .A2(n20032), .B1(n19751), .B2(n20025), .Y(n18984) );
  sky130_fd_sc_hd__nand2_1 U23304 ( .A(n18985), .B(n18984), .Y(n21901) );
  sky130_fd_sc_hd__nand2_1 U23305 ( .A(n21901), .B(n22125), .Y(n18995) );
  sky130_fd_sc_hd__nand2_1 U23306 ( .A(n18988), .B(n18987), .Y(n18991) );
  sky130_fd_sc_hd__xnor2_1 U23308 ( .A(n18991), .B(n18990), .Y(n21898) );
  sky130_fd_sc_hd__o22ai_1 U23309 ( .A1(n20043), .A2(n21900), .B1(n18992), 
        .B2(n20012), .Y(n18993) );
  sky130_fd_sc_hd__a21oi_1 U23310 ( .A1(n21898), .A2(n20016), .B1(n18993), .Y(
        n18994) );
  sky130_fd_sc_hd__nand2_1 U23311 ( .A(n18995), .B(n18994), .Y(n20571) );
  sky130_fd_sc_hd__nand2_1 U23312 ( .A(n20571), .B(n20019), .Y(n19065) );
  sky130_fd_sc_hd__nand2_1 U23313 ( .A(n18997), .B(n18996), .Y(n19001) );
  sky130_fd_sc_hd__xnor2_1 U23315 ( .A(n19001), .B(n19000), .Y(n21708) );
  sky130_fd_sc_hd__nand2_1 U23316 ( .A(n21708), .B(n20030), .Y(n19011) );
  sky130_fd_sc_hd__nand2_1 U23317 ( .A(n19004), .B(n19003), .Y(n19009) );
  sky130_fd_sc_hd__a21oi_1 U23318 ( .A1(n19007), .A2(n19006), .B1(n19005), .Y(
        n19135) );
  sky130_fd_sc_hd__xnor2_1 U23320 ( .A(n19009), .B(n19008), .Y(n19535) );
  sky130_fd_sc_hd__a22oi_1 U23321 ( .A1(j202_soc_core_j22_cpu_ml_mach[6]), 
        .A2(n20032), .B1(n19535), .B2(n20025), .Y(n19010) );
  sky130_fd_sc_hd__nand2_1 U23322 ( .A(n19011), .B(n19010), .Y(n22050) );
  sky130_fd_sc_hd__nand2_1 U23323 ( .A(n22050), .B(n22125), .Y(n19020) );
  sky130_fd_sc_hd__nand2_1 U23324 ( .A(n19014), .B(n19013), .Y(n19016) );
  sky130_fd_sc_hd__xor2_1 U23325 ( .A(n19016), .B(n19015), .X(n22047) );
  sky130_fd_sc_hd__o22ai_1 U23326 ( .A1(n20043), .A2(n22049), .B1(n19017), 
        .B2(n20012), .Y(n19018) );
  sky130_fd_sc_hd__a21oi_1 U23327 ( .A1(n22047), .A2(n20016), .B1(n19018), .Y(
        n19019) );
  sky130_fd_sc_hd__nand2_1 U23328 ( .A(n19020), .B(n19019), .Y(n19467) );
  sky130_fd_sc_hd__nand2_1 U23329 ( .A(n19467), .B(n21137), .Y(n19050) );
  sky130_fd_sc_hd__nand2_1 U23330 ( .A(n25276), .B(n19895), .Y(n19023) );
  sky130_fd_sc_hd__a2bb2oi_1 U23331 ( .B1(n21135), .B2(n19893), .A1_N(n19891), 
        .A2_N(n21045), .Y(n19022) );
  sky130_fd_sc_hd__nand2_1 U23332 ( .A(n25310), .B(n19889), .Y(n19021) );
  sky130_fd_sc_hd__a21oi_1 U23333 ( .A1(n22708), .A2(n21089), .B1(n20641), .Y(
        n19025) );
  sky130_fd_sc_hd__nand2_1 U23334 ( .A(n22045), .B(n21170), .Y(n19024) );
  sky130_fd_sc_hd__o211ai_1 U23335 ( .A1(n20908), .A2(n22045), .B1(n19025), 
        .C1(n19024), .Y(n19039) );
  sky130_fd_sc_hd__o2bb2ai_1 U23337 ( .B1(n21862), .B2(n20712), .A1_N(n23316), 
        .A2_N(n20716), .Y(n19027) );
  sky130_fd_sc_hd__o2bb2ai_1 U23338 ( .B1(n22558), .B2(n21163), .A1_N(n21164), 
        .A2_N(n22483), .Y(n19026) );
  sky130_fd_sc_hd__nor2_1 U23339 ( .A(n19027), .B(n19026), .Y(n19035) );
  sky130_fd_sc_hd__xor2_1 U23340 ( .A(n20530), .B(n22708), .X(n22433) );
  sky130_fd_sc_hd__a22oi_1 U23341 ( .A1(n21156), .A2(n21152), .B1(n22433), 
        .B2(n21147), .Y(n19034) );
  sky130_fd_sc_hd__o22ai_1 U23342 ( .A1(n21145), .A2(n22708), .B1(n19028), 
        .B2(n22567), .Y(n19031) );
  sky130_fd_sc_hd__nor2_1 U23343 ( .A(n22567), .B(n19875), .Y(n19030) );
  sky130_fd_sc_hd__o22ai_1 U23344 ( .A1(n22580), .A2(n21155), .B1(n22645), 
        .B2(n21154), .Y(n19029) );
  sky130_fd_sc_hd__nor3_1 U23345 ( .A(n19031), .B(n19030), .C(n19029), .Y(
        n19033) );
  sky130_fd_sc_hd__nand2_1 U23346 ( .A(n19884), .B(n22708), .Y(n19032) );
  sky130_fd_sc_hd__nand4_1 U23347 ( .A(n19035), .B(n19034), .C(n19033), .D(
        n19032), .Y(n19036) );
  sky130_fd_sc_hd__a21oi_1 U23348 ( .A1(n22045), .A2(n19037), .B1(n19036), .Y(
        n19038) );
  sky130_fd_sc_hd__nand2_1 U23349 ( .A(n19042), .B(n19041), .Y(n19047) );
  sky130_fd_sc_hd__a21oi_1 U23350 ( .A1(n19045), .A2(n19044), .B1(n19043), .Y(
        n19076) );
  sky130_fd_sc_hd__o21ai_1 U23351 ( .A1(n19072), .A2(n19076), .B1(n19073), .Y(
        n19046) );
  sky130_fd_sc_hd__xnor2_1 U23352 ( .A(n19047), .B(n19046), .Y(n21846) );
  sky130_fd_sc_hd__nand2_1 U23353 ( .A(n21846), .B(n21178), .Y(n19048) );
  sky130_fd_sc_hd__nand2_1 U23354 ( .A(n21850), .B(n19905), .Y(n19547) );
  sky130_fd_sc_hd__o22ai_1 U23355 ( .A1(n19052), .A2(n19973), .B1(n19051), 
        .B2(n19971), .Y(n19056) );
  sky130_fd_sc_hd__o22ai_1 U23356 ( .A1(n19054), .A2(n19977), .B1(n19053), 
        .B2(n19975), .Y(n19055) );
  sky130_fd_sc_hd__nor2_1 U23357 ( .A(n19056), .B(n19055), .Y(n19061) );
  sky130_fd_sc_hd__a2bb2oi_1 U23358 ( .B1(j202_soc_core_j22_cpu_rf_vbr[6]), 
        .B2(n19985), .A1_N(n19057), .A2_N(n19986), .Y(n19060) );
  sky130_fd_sc_hd__nand2_1 U23359 ( .A(n19842), .B(
        j202_soc_core_j22_cpu_rf_gpr[6]), .Y(n19059) );
  sky130_fd_sc_hd__nand2_1 U23360 ( .A(n19843), .B(
        j202_soc_core_j22_cpu_rf_tmp[6]), .Y(n19058) );
  sky130_fd_sc_hd__nand4_1 U23361 ( .A(n19061), .B(n19060), .C(n19059), .D(
        n19058), .Y(n19062) );
  sky130_fd_sc_hd__a21oi_1 U23362 ( .A1(n19063), .A2(n19969), .B1(n19062), .Y(
        n19546) );
  sky130_fd_sc_hd__nand2b_1 U23363 ( .A_N(n19546), .B(n19285), .Y(n19064) );
  sky130_fd_sc_hd__o211ai_1 U23364 ( .A1(n19317), .A2(n19765), .B1(n19065), 
        .C1(n19767), .Y(n25301) );
  sky130_fd_sc_hd__nand2_1 U23365 ( .A(n21846), .B(n19729), .Y(n19071) );
  sky130_fd_sc_hd__ha_1 U23366 ( .A(j202_soc_core_j22_cpu_pc[6]), .B(n19066), 
        .COUT(n16706), .SUM(n21851) );
  sky130_fd_sc_hd__nand2_1 U23367 ( .A(n19661), .B(n21851), .Y(n19068) );
  sky130_fd_sc_hd__nand2_1 U23368 ( .A(n19736), .B(n22708), .Y(n19067) );
  sky130_fd_sc_hd__o211ai_1 U23369 ( .A1(n22612), .A2(n19731), .B1(n19068), 
        .C1(n19067), .Y(n19069) );
  sky130_fd_sc_hd__a21oi_1 U23370 ( .A1(n25276), .A2(n19737), .B1(n19069), .Y(
        n19070) );
  sky130_fd_sc_hd__nand2_1 U23371 ( .A(n19071), .B(n19070), .Y(n25337) );
  sky130_fd_sc_hd__nand2_1 U23372 ( .A(n19074), .B(n19073), .Y(n19075) );
  sky130_fd_sc_hd__xor2_1 U23373 ( .A(n19076), .B(n19075), .X(n22039) );
  sky130_fd_sc_hd__nand2_1 U23374 ( .A(n22039), .B(n19729), .Y(n19086) );
  sky130_fd_sc_hd__ha_1 U23375 ( .A(j202_soc_core_j22_cpu_pc[5]), .B(n19077), 
        .COUT(n19066), .SUM(n22034) );
  sky130_fd_sc_hd__o22ai_1 U23376 ( .A1(n22041), .A2(n19078), .B1(n22580), 
        .B2(n19731), .Y(n19079) );
  sky130_fd_sc_hd__a21oi_1 U23377 ( .A1(n19080), .A2(n22176), .B1(n19079), .Y(
        n19082) );
  sky130_fd_sc_hd__nand2_1 U23378 ( .A(n19517), .B(n22034), .Y(n19081) );
  sky130_fd_sc_hd__o211ai_1 U23379 ( .A1(n22037), .A2(n19083), .B1(n19082), 
        .C1(n19081), .Y(n19084) );
  sky130_fd_sc_hd__a21oi_1 U23380 ( .A1(n25255), .A2(n19737), .B1(n19084), .Y(
        n19085) );
  sky130_fd_sc_hd__nand2_1 U23381 ( .A(n19086), .B(n19085), .Y(n25336) );
  sky130_fd_sc_hd__nand2_1 U23382 ( .A(n25256), .B(n19087), .Y(n19092) );
  sky130_fd_sc_hd__a22oi_1 U23383 ( .A1(j202_soc_core_j22_cpu_id_opn_inst__4_), 
        .A2(n19088), .B1(j202_soc_core_j22_cpu_id_op2_v_), .B2(
        j202_soc_core_j22_cpu_id_op2_inst__4_), .Y(n19091) );
  sky130_fd_sc_hd__nand2_1 U23384 ( .A(n22540), .B(n19089), .Y(n19090) );
  sky130_fd_sc_hd__nand3_1 U23385 ( .A(n19092), .B(n19091), .C(n19090), .Y(
        n25386) );
  sky130_fd_sc_hd__clkinv_1 U23386 ( .A(j202_soc_core_uart_BRG_br_clr), .Y(
        n24823) );
  sky130_fd_sc_hd__nor2_1 U23387 ( .A(j202_soc_core_uart_BRG_sio_ce_x4_r), .B(
        n24823), .Y(n25400) );
  sky130_fd_sc_hd__nor2b_1 U23388 ( .B_N(j202_soc_core_uart_TOP_dpll_state[0]), 
        .A(j202_soc_core_uart_TOP_dpll_state[1]), .Y(n25405) );
  sky130_fd_sc_hd__nand2_1 U23389 ( .A(n19094), .B(n19093), .Y(n19099) );
  sky130_fd_sc_hd__xnor2_1 U23391 ( .A(n19099), .B(n19098), .Y(n21696) );
  sky130_fd_sc_hd__nand2_1 U23392 ( .A(n19101), .B(n19100), .Y(n19103) );
  sky130_fd_sc_hd__xnor2_1 U23393 ( .A(n19103), .B(n19102), .Y(n19601) );
  sky130_fd_sc_hd__o22ai_1 U23394 ( .A1(n20007), .A2(n22232), .B1(n19104), 
        .B2(n20005), .Y(n19105) );
  sky130_fd_sc_hd__a21oi_1 U23395 ( .A1(n19601), .A2(n20025), .B1(n19105), .Y(
        n19106) );
  sky130_fd_sc_hd__nand2_1 U23396 ( .A(n19109), .B(n19108), .Y(n19110) );
  sky130_fd_sc_hd__xor2_1 U23397 ( .A(n19111), .B(n19110), .X(n22230) );
  sky130_fd_sc_hd__o22ai_1 U23398 ( .A1(n20014), .A2(n22232), .B1(n19112), 
        .B2(n20012), .Y(n19113) );
  sky130_fd_sc_hd__a21oi_1 U23399 ( .A1(n22230), .A2(n20016), .B1(n19113), .Y(
        n19114) );
  sky130_fd_sc_hd__o21a_1 U23400 ( .A1(j202_soc_core_j22_cpu_macop_MAC_[0]), 
        .A2(n22207), .B1(n19114), .X(n20568) );
  sky130_fd_sc_hd__nand2_1 U23401 ( .A(n19115), .B(n19969), .Y(n19126) );
  sky130_fd_sc_hd__o22ai_1 U23402 ( .A1(n19117), .A2(n19971), .B1(n19116), 
        .B2(n19975), .Y(n19118) );
  sky130_fd_sc_hd__a21oi_1 U23403 ( .A1(n19842), .A2(
        j202_soc_core_j22_cpu_rf_gpr[13]), .B1(n19118), .Y(n19125) );
  sky130_fd_sc_hd__o22ai_1 U23404 ( .A1(n19120), .A2(n19981), .B1(n19119), 
        .B2(n19986), .Y(n19123) );
  sky130_fd_sc_hd__o2bb2ai_1 U23405 ( .B1(n19121), .B2(n19977), .A1_N(
        j202_soc_core_j22_cpu_rf_vbr[13]), .A2_N(n19985), .Y(n19122) );
  sky130_fd_sc_hd__nor2_1 U23406 ( .A(n19123), .B(n19122), .Y(n19124) );
  sky130_fd_sc_hd__nand3_1 U23407 ( .A(n19126), .B(n19125), .C(n19124), .Y(
        n19617) );
  sky130_fd_sc_hd__nand2_1 U23408 ( .A(n19617), .B(n20020), .Y(n19193) );
  sky130_fd_sc_hd__nand2_1 U23409 ( .A(n19128), .B(n19127), .Y(n19130) );
  sky130_fd_sc_hd__xnor2_1 U23410 ( .A(n19130), .B(n19129), .Y(n21709) );
  sky130_fd_sc_hd__nand2_1 U23411 ( .A(n21709), .B(n20030), .Y(n19139) );
  sky130_fd_sc_hd__nand2_1 U23412 ( .A(n19133), .B(n19132), .Y(n19134) );
  sky130_fd_sc_hd__xor2_1 U23413 ( .A(n19135), .B(n19134), .X(n19399) );
  sky130_fd_sc_hd__o22ai_1 U23414 ( .A1(n20007), .A2(n22031), .B1(n19136), 
        .B2(n20005), .Y(n19137) );
  sky130_fd_sc_hd__a21oi_1 U23415 ( .A1(n19399), .A2(n20025), .B1(n19137), .Y(
        n19138) );
  sky130_fd_sc_hd__nand2_1 U23416 ( .A(n19139), .B(n19138), .Y(n22027) );
  sky130_fd_sc_hd__nand2_1 U23417 ( .A(n22027), .B(n22125), .Y(n19147) );
  sky130_fd_sc_hd__nand2_1 U23418 ( .A(n19141), .B(n19140), .Y(n19142) );
  sky130_fd_sc_hd__xnor2_1 U23419 ( .A(n19143), .B(n19142), .Y(n22029) );
  sky130_fd_sc_hd__o22ai_1 U23420 ( .A1(n20014), .A2(n22031), .B1(n19144), 
        .B2(n20012), .Y(n19145) );
  sky130_fd_sc_hd__a21oi_1 U23421 ( .A1(n22029), .A2(n20016), .B1(n19145), .Y(
        n19146) );
  sky130_fd_sc_hd__nand2_1 U23422 ( .A(n19147), .B(n19146), .Y(n19469) );
  sky130_fd_sc_hd__nand2_1 U23423 ( .A(n19469), .B(n21137), .Y(n19178) );
  sky130_fd_sc_hd__nand2_1 U23424 ( .A(n25309), .B(n19889), .Y(n19151) );
  sky130_fd_sc_hd__o22a_1 U23425 ( .A1(n22527), .A2(n19891), .B1(n19148), .B2(
        n22526), .X(n19150) );
  sky130_fd_sc_hd__nand2_1 U23426 ( .A(n25255), .B(n19895), .Y(n19149) );
  sky130_fd_sc_hd__nand3_1 U23427 ( .A(n22555), .B(n21170), .C(n19173), .Y(
        n19166) );
  sky130_fd_sc_hd__nand2_1 U23428 ( .A(n22441), .B(n19152), .Y(n19879) );
  sky130_fd_sc_hd__nor2_1 U23429 ( .A(n19153), .B(n19879), .Y(n19156) );
  sky130_fd_sc_hd__nand2_1 U23430 ( .A(n22176), .B(n19173), .Y(n22649) );
  sky130_fd_sc_hd__a2bb2oi_1 U23431 ( .B1(n20641), .B2(n19173), .A1_N(n21145), 
        .A2_N(n22176), .Y(n19154) );
  sky130_fd_sc_hd__a211o_1 U23433 ( .A1(n19157), .A2(n22578), .B1(n19156), 
        .C1(n19155), .X(n19158) );
  sky130_fd_sc_hd__a21oi_1 U23434 ( .A1(n20716), .A2(n23313), .B1(n19158), .Y(
        n19165) );
  sky130_fd_sc_hd__o2bb2ai_1 U23435 ( .B1(n22647), .B2(n21155), .A1_N(n21156), 
        .A2_N(n20648), .Y(n19162) );
  sky130_fd_sc_hd__nand2_1 U23436 ( .A(n22037), .B(n22580), .Y(n19159) );
  sky130_fd_sc_hd__nand2_1 U23437 ( .A(n19159), .B(n22649), .Y(n22432) );
  sky130_fd_sc_hd__o22ai_1 U23438 ( .A1(n21108), .A2(n22432), .B1(n22612), 
        .B2(n21154), .Y(n19161) );
  sky130_fd_sc_hd__o22ai_1 U23439 ( .A1(n22300), .A2(n20712), .B1(n22645), 
        .B2(n21163), .Y(n19160) );
  sky130_fd_sc_hd__nor3_1 U23440 ( .A(n19162), .B(n19161), .C(n19160), .Y(
        n19164) );
  sky130_fd_sc_hd__nand2_1 U23441 ( .A(n19884), .B(n22176), .Y(n19163) );
  sky130_fd_sc_hd__nand4_1 U23442 ( .A(n19166), .B(n19165), .C(n19164), .D(
        n19163), .Y(n19171) );
  sky130_fd_sc_hd__nand2_1 U23443 ( .A(n22039), .B(n21178), .Y(n19169) );
  sky130_fd_sc_hd__nand2_1 U23444 ( .A(n22555), .B(n19167), .Y(n19168) );
  sky130_fd_sc_hd__nand2_1 U23445 ( .A(n19169), .B(n19168), .Y(n19170) );
  sky130_fd_sc_hd__nor2_1 U23446 ( .A(n19171), .B(n19170), .Y(n19177) );
  sky130_fd_sc_hd__xnor2_1 U23447 ( .A(n19173), .B(n22555), .Y(n19174) );
  sky130_fd_sc_hd__o22ai_1 U23448 ( .A1(n22600), .A2(n21017), .B1(n22509), 
        .B2(n19174), .Y(n19175) );
  sky130_fd_sc_hd__nand2_1 U23449 ( .A(n19175), .B(n21139), .Y(n19176) );
  sky130_fd_sc_hd__nand2_1 U23450 ( .A(n22033), .B(n19905), .Y(n19470) );
  sky130_fd_sc_hd__o22ai_1 U23451 ( .A1(n19180), .A2(n19973), .B1(n19179), 
        .B2(n19971), .Y(n19184) );
  sky130_fd_sc_hd__o22ai_1 U23452 ( .A1(n19182), .A2(n19977), .B1(n19181), 
        .B2(n19975), .Y(n19183) );
  sky130_fd_sc_hd__nor2_1 U23453 ( .A(n19184), .B(n19183), .Y(n19189) );
  sky130_fd_sc_hd__a2bb2oi_1 U23454 ( .B1(j202_soc_core_j22_cpu_rf_vbr[5]), 
        .B2(n19985), .A1_N(n19185), .A2_N(n19986), .Y(n19188) );
  sky130_fd_sc_hd__nand2_1 U23455 ( .A(n19842), .B(
        j202_soc_core_j22_cpu_rf_gpr[5]), .Y(n19187) );
  sky130_fd_sc_hd__nand2_1 U23456 ( .A(n19843), .B(
        j202_soc_core_j22_cpu_rf_tmp[5]), .Y(n19186) );
  sky130_fd_sc_hd__nand4_1 U23457 ( .A(n19189), .B(n19188), .C(n19187), .D(
        n19186), .Y(n19190) );
  sky130_fd_sc_hd__a21oi_1 U23458 ( .A1(n19191), .A2(n19969), .B1(n19190), .Y(
        n19472) );
  sky130_fd_sc_hd__nand2b_1 U23459 ( .A_N(n19472), .B(n19285), .Y(n19192) );
  sky130_fd_sc_hd__o211ai_1 U23460 ( .A1(n20568), .A2(n20067), .B1(n19193), 
        .C1(n19619), .Y(n25344) );
  sky130_fd_sc_hd__nand2_1 U23461 ( .A(n22053), .B(n19729), .Y(n19199) );
  sky130_fd_sc_hd__ha_1 U23462 ( .A(j202_soc_core_j22_cpu_pc[4]), .B(n19194), 
        .COUT(n19077), .SUM(n22058) );
  sky130_fd_sc_hd__nand2_1 U23463 ( .A(n19661), .B(n22058), .Y(n19196) );
  sky130_fd_sc_hd__nand2_1 U23464 ( .A(n19736), .B(n22705), .Y(n19195) );
  sky130_fd_sc_hd__o211ai_1 U23465 ( .A1(n22647), .A2(n19731), .B1(n19196), 
        .C1(n19195), .Y(n19197) );
  sky130_fd_sc_hd__a21oi_1 U23466 ( .A1(n25256), .A2(n19737), .B1(n19197), .Y(
        n19198) );
  sky130_fd_sc_hd__nand2_1 U23467 ( .A(n19199), .B(n19198), .Y(n25335) );
  sky130_fd_sc_hd__o22ai_1 U23468 ( .A1(n19201), .A2(n19973), .B1(n19200), 
        .B2(n19971), .Y(n19205) );
  sky130_fd_sc_hd__o22ai_1 U23469 ( .A1(n19203), .A2(n19977), .B1(n19202), 
        .B2(n19975), .Y(n19204) );
  sky130_fd_sc_hd__nor2_1 U23470 ( .A(n19205), .B(n19204), .Y(n19210) );
  sky130_fd_sc_hd__a2bb2oi_1 U23471 ( .B1(j202_soc_core_j22_cpu_rf_vbr[8]), 
        .B2(n19985), .A1_N(n19206), .A2_N(n19986), .Y(n19209) );
  sky130_fd_sc_hd__nand2_1 U23472 ( .A(n19842), .B(
        j202_soc_core_j22_cpu_rf_gpr[8]), .Y(n19208) );
  sky130_fd_sc_hd__nand2_1 U23473 ( .A(n19843), .B(
        j202_soc_core_j22_cpu_rf_tmp[8]), .Y(n19207) );
  sky130_fd_sc_hd__nand4_1 U23474 ( .A(n19210), .B(n19209), .C(n19208), .D(
        n19207), .Y(n19211) );
  sky130_fd_sc_hd__a21oi_1 U23475 ( .A1(n19212), .A2(n19969), .B1(n19211), .Y(
        n19717) );
  sky130_fd_sc_hd__a21oi_1 U23476 ( .A1(n19216), .A2(n19215), .B1(n19214), .Y(
        n19221) );
  sky130_fd_sc_hd__nand2_1 U23477 ( .A(n19219), .B(n19218), .Y(n19220) );
  sky130_fd_sc_hd__xor2_1 U23478 ( .A(n19221), .B(n19220), .X(n21702) );
  sky130_fd_sc_hd__nand2_1 U23479 ( .A(n21702), .B(n20030), .Y(n19231) );
  sky130_fd_sc_hd__a21oi_1 U23480 ( .A1(n19224), .A2(n19223), .B1(n19222), .Y(
        n19228) );
  sky130_fd_sc_hd__nand2_1 U23481 ( .A(n19226), .B(n19225), .Y(n19227) );
  sky130_fd_sc_hd__xor2_1 U23482 ( .A(n19228), .B(n19227), .X(n19675) );
  sky130_fd_sc_hd__o2bb2ai_1 U23483 ( .B1(n20007), .B2(n22247), .A1_N(
        j202_soc_core_j22_cpu_ml_mach[0]), .A2_N(n20032), .Y(n19229) );
  sky130_fd_sc_hd__a21oi_1 U23484 ( .A1(n19675), .A2(n20025), .B1(n19229), .Y(
        n19230) );
  sky130_fd_sc_hd__nand2_1 U23485 ( .A(n19231), .B(n19230), .Y(n22215) );
  sky130_fd_sc_hd__nand2_1 U23486 ( .A(n22215), .B(n22125), .Y(n19238) );
  sky130_fd_sc_hd__xnor2_1 U23487 ( .A(n19234), .B(n19233), .Y(n22242) );
  sky130_fd_sc_hd__o22ai_1 U23488 ( .A1(n22247), .A2(n20014), .B1(n19235), 
        .B2(n20012), .Y(n19236) );
  sky130_fd_sc_hd__a21oi_1 U23489 ( .A1(n22242), .A2(n20016), .B1(n19236), .Y(
        n19237) );
  sky130_fd_sc_hd__nand2_1 U23490 ( .A(n19238), .B(n19237), .Y(n19499) );
  sky130_fd_sc_hd__nand2_1 U23491 ( .A(n19499), .B(n21137), .Y(n19271) );
  sky130_fd_sc_hd__nand2_1 U23492 ( .A(n22516), .B(n19893), .Y(n19242) );
  sky130_fd_sc_hd__a22oi_1 U23493 ( .A1(n19239), .A2(n22524), .B1(n25259), 
        .B2(n19895), .Y(n19241) );
  sky130_fd_sc_hd__nand2_1 U23494 ( .A(n25308), .B(n19889), .Y(n19240) );
  sky130_fd_sc_hd__o21ai_1 U23495 ( .A1(n20908), .A2(n22584), .B1(n21010), .Y(
        n19266) );
  sky130_fd_sc_hd__nand2_1 U23496 ( .A(n19245), .B(n19244), .Y(n19246) );
  sky130_fd_sc_hd__xnor2_1 U23497 ( .A(n19247), .B(n19246), .Y(n21625) );
  sky130_fd_sc_hd__nand2_1 U23498 ( .A(n22037), .B(n22608), .Y(n19249) );
  sky130_fd_sc_hd__nand2_1 U23499 ( .A(n22176), .B(n11202), .Y(n19248) );
  sky130_fd_sc_hd__nand4_1 U23500 ( .A(n22592), .B(n19249), .C(n22181), .D(
        n19248), .Y(n19251) );
  sky130_fd_sc_hd__nand2_1 U23501 ( .A(n21627), .B(n22146), .Y(n22437) );
  sky130_fd_sc_hd__nand2_1 U23502 ( .A(n22185), .B(n22584), .Y(n22619) );
  sky130_fd_sc_hd__nand3_1 U23503 ( .A(n22437), .B(n21147), .C(n22619), .Y(
        n19250) );
  sky130_fd_sc_hd__o211ai_1 U23504 ( .A1(n20805), .A2(n21154), .B1(n19251), 
        .C1(n19250), .Y(n19252) );
  sky130_fd_sc_hd__a21oi_1 U23505 ( .A1(n20716), .A2(n23298), .B1(n19252), .Y(
        n19263) );
  sky130_fd_sc_hd__nand3_1 U23506 ( .A(n21139), .B(n19255), .C(n19254), .Y(
        n19256) );
  sky130_fd_sc_hd__o21a_1 U23507 ( .A1(n21145), .A2(n22185), .B1(n19256), .X(
        n19257) );
  sky130_fd_sc_hd__a21oi_1 U23509 ( .A1(n21156), .A2(n20721), .B1(n19258), .Y(
        n19259) );
  sky130_fd_sc_hd__o21a_1 U23510 ( .A1(n22487), .A2(n21163), .B1(n19259), .X(
        n19262) );
  sky130_fd_sc_hd__a2bb2oi_1 U23511 ( .B1(n22133), .B2(n20711), .A1_N(n21929), 
        .A2_N(n20712), .Y(n19261) );
  sky130_fd_sc_hd__nand2_1 U23512 ( .A(n19884), .B(n22185), .Y(n19260) );
  sky130_fd_sc_hd__nand4_1 U23513 ( .A(n19263), .B(n19262), .C(n19261), .D(
        n19260), .Y(n19264) );
  sky130_fd_sc_hd__a21oi_1 U23514 ( .A1(n21625), .A2(n21178), .B1(n19264), .Y(
        n19265) );
  sky130_fd_sc_hd__nand2_1 U23515 ( .A(n22725), .B(n21170), .Y(n19267) );
  sky130_fd_sc_hd__o211ai_1 U23516 ( .A1(n20908), .A2(n22725), .B1(n20905), 
        .C1(n19267), .Y(n19268) );
  sky130_fd_sc_hd__nand2_1 U23517 ( .A(n19268), .B(n22584), .Y(n19269) );
  sky130_fd_sc_hd__nand2_1 U23518 ( .A(n21613), .B(n19905), .Y(n19691) );
  sky130_fd_sc_hd__nand2_1 U23519 ( .A(n19272), .B(n19969), .Y(n19284) );
  sky130_fd_sc_hd__o22ai_1 U23520 ( .A1(n11202), .A2(n19973), .B1(n19273), 
        .B2(n19971), .Y(n19276) );
  sky130_fd_sc_hd__o22ai_1 U23521 ( .A1(n21630), .A2(n19977), .B1(n19274), 
        .B2(n19975), .Y(n19275) );
  sky130_fd_sc_hd__nor2_1 U23522 ( .A(n19276), .B(n19275), .Y(n19283) );
  sky130_fd_sc_hd__o22ai_1 U23523 ( .A1(n19278), .A2(n19983), .B1(n19277), 
        .B2(n19981), .Y(n19281) );
  sky130_fd_sc_hd__o2bb2ai_1 U23524 ( .B1(n19279), .B2(n19986), .A1_N(
        j202_soc_core_j22_cpu_rf_vbr[0]), .A2_N(n19985), .Y(n19280) );
  sky130_fd_sc_hd__nor2_1 U23525 ( .A(n19281), .B(n19280), .Y(n19282) );
  sky130_fd_sc_hd__nand3_1 U23526 ( .A(n19284), .B(n19283), .C(n19282), .Y(
        n19690) );
  sky130_fd_sc_hd__nand2_1 U23527 ( .A(n19690), .B(n19285), .Y(n19286) );
  sky130_fd_sc_hd__nand2_1 U23528 ( .A(n19289), .B(n19288), .Y(n19294) );
  sky130_fd_sc_hd__xnor2_1 U23530 ( .A(n19294), .B(n19293), .Y(n21717) );
  sky130_fd_sc_hd__nand2_1 U23531 ( .A(n21717), .B(n20030), .Y(n19306) );
  sky130_fd_sc_hd__nand2_1 U23532 ( .A(n19297), .B(n19296), .Y(n19302) );
  sky130_fd_sc_hd__o21ai_1 U23533 ( .A1(n19300), .A2(n19299), .B1(n19298), .Y(
        n19301) );
  sky130_fd_sc_hd__xnor2_1 U23534 ( .A(n19302), .B(n19301), .Y(n19703) );
  sky130_fd_sc_hd__o22ai_1 U23535 ( .A1(n20007), .A2(n21922), .B1(n19303), 
        .B2(n20005), .Y(n19304) );
  sky130_fd_sc_hd__a21oi_1 U23536 ( .A1(n19703), .A2(n20025), .B1(n19304), .Y(
        n19305) );
  sky130_fd_sc_hd__nand2_1 U23537 ( .A(n19306), .B(n19305), .Y(n21918) );
  sky130_fd_sc_hd__nand2_1 U23538 ( .A(n21918), .B(n22125), .Y(n19315) );
  sky130_fd_sc_hd__nand2_1 U23539 ( .A(n19309), .B(n19308), .Y(n19311) );
  sky130_fd_sc_hd__xor2_1 U23540 ( .A(n19311), .B(n19310), .X(n21920) );
  sky130_fd_sc_hd__o22ai_1 U23541 ( .A1(n20014), .A2(n21922), .B1(n19312), 
        .B2(n20012), .Y(n19313) );
  sky130_fd_sc_hd__a21oi_1 U23542 ( .A1(n21920), .A2(n20016), .B1(n19313), .Y(
        n19314) );
  sky130_fd_sc_hd__nand2_1 U23543 ( .A(n19315), .B(n19314), .Y(n20521) );
  sky130_fd_sc_hd__nand2_1 U23544 ( .A(n20521), .B(n20019), .Y(n19316) );
  sky130_fd_sc_hd__o211ai_1 U23545 ( .A1(n19317), .A2(n19717), .B1(n19719), 
        .C1(n19316), .Y(n25367) );
  sky130_fd_sc_hd__nand3_1 U23546 ( .A(n19833), .B(n21245), .C(n25374), .Y(
        n20069) );
  sky130_fd_sc_hd__nor2_1 U23547 ( .A(n19836), .B(n20069), .Y(n25324) );
  sky130_fd_sc_hd__nand2_1 U23548 ( .A(n20063), .B(n19500), .Y(n19320) );
  sky130_fd_sc_hd__nand2_1 U23549 ( .A(n19318), .B(n20019), .Y(n19319) );
  sky130_fd_sc_hd__nand3_1 U23550 ( .A(n20065), .B(n19320), .C(n19319), .Y(
        n25363) );
  sky130_fd_sc_hd__nand2_1 U23551 ( .A(n19479), .B(n24872), .Y(n21586) );
  sky130_fd_sc_hd__nand2_1 U23552 ( .A(n25381), .B(n21420), .Y(n20983) );
  sky130_fd_sc_hd__nor2_1 U23553 ( .A(n25377), .B(n22330), .Y(n21435) );
  sky130_fd_sc_hd__nand2_1 U23554 ( .A(n22734), .B(n21435), .Y(n21568) );
  sky130_fd_sc_hd__nor3_1 U23555 ( .A(n25315), .B(n21586), .C(n21568), .Y(
        n21427) );
  sky130_fd_sc_hd__nand2_1 U23556 ( .A(n19480), .B(n25303), .Y(n20327) );
  sky130_fd_sc_hd__nor2_1 U23557 ( .A(n21586), .B(n20327), .Y(n21635) );
  sky130_fd_sc_hd__nand2_1 U23558 ( .A(n22330), .B(n21635), .Y(n21457) );
  sky130_fd_sc_hd__nor2_1 U23559 ( .A(n25303), .B(n19480), .Y(n21735) );
  sky130_fd_sc_hd__nor2_1 U23560 ( .A(n21586), .B(n20341), .Y(n21464) );
  sky130_fd_sc_hd__nand2_1 U23561 ( .A(n22330), .B(n22734), .Y(n22385) );
  sky130_fd_sc_hd__nor2_1 U23562 ( .A(n25303), .B(n25315), .Y(n24873) );
  sky130_fd_sc_hd__nor2_1 U23563 ( .A(n21418), .B(n21586), .Y(n20737) );
  sky130_fd_sc_hd__nand3_1 U23564 ( .A(n25304), .B(n24873), .C(n24872), .Y(
        n20335) );
  sky130_fd_sc_hd__nor2_1 U23565 ( .A(n25383), .B(n25384), .Y(n19321) );
  sky130_fd_sc_hd__nand2_1 U23566 ( .A(n19483), .B(n19321), .Y(n20752) );
  sky130_fd_sc_hd__nor2_1 U23567 ( .A(n20752), .B(n25386), .Y(n20736) );
  sky130_fd_sc_hd__nand2_1 U23568 ( .A(n19322), .B(n20736), .Y(n19493) );
  sky130_fd_sc_hd__nand2_1 U23569 ( .A(n21420), .B(n25377), .Y(n22743) );
  sky130_fd_sc_hd__nor2_1 U23570 ( .A(n25381), .B(n22743), .Y(n20336) );
  sky130_fd_sc_hd__nand2_1 U23571 ( .A(n25372), .B(n20336), .Y(n20759) );
  sky130_fd_sc_hd__nor2_1 U23572 ( .A(n19493), .B(n20759), .Y(n21518) );
  sky130_fd_sc_hd__nor4_1 U23573 ( .A(n19483), .B(n25383), .C(n25384), .D(
        n25386), .Y(n21640) );
  sky130_fd_sc_hd__nand2_1 U23574 ( .A(n19322), .B(n21640), .Y(n21480) );
  sky130_fd_sc_hd__nand2_1 U23575 ( .A(n21403), .B(n20336), .Y(n21555) );
  sky130_fd_sc_hd__nand2_1 U23576 ( .A(n21487), .B(n19322), .Y(n21505) );
  sky130_fd_sc_hd__nor2_1 U23577 ( .A(n21505), .B(n24827), .Y(n20331) );
  sky130_fd_sc_hd__nand2_1 U23578 ( .A(n20331), .B(n21331), .Y(n21333) );
  sky130_fd_sc_hd__nand2_1 U23579 ( .A(n21555), .B(n21333), .Y(n21540) );
  sky130_fd_sc_hd__nor2_1 U23580 ( .A(n21518), .B(n21540), .Y(n20750) );
  sky130_fd_sc_hd__a211oi_1 U23582 ( .A1(n21420), .A2(n20995), .B1(n21464), 
        .C1(n19323), .Y(n21436) );
  sky130_fd_sc_hd__nor3_1 U23583 ( .A(n25380), .B(n25377), .C(n25381), .Y(
        n20766) );
  sky130_fd_sc_hd__nand2_1 U23584 ( .A(n20766), .B(n21635), .Y(n21402) );
  sky130_fd_sc_hd__nand3b_1 U23585 ( .A_N(n21427), .B(n21436), .C(n21402), .Y(
        n21509) );
  sky130_fd_sc_hd__nand4_1 U23586 ( .A(j202_soc_core_j22_cpu_opst[4]), .B(
        n20773), .C(n21441), .D(n22417), .Y(n22803) );
  sky130_fd_sc_hd__nand2_1 U23587 ( .A(n24879), .B(n19325), .Y(n21644) );
  sky130_fd_sc_hd__a21o_1 U23588 ( .A1(n21509), .A2(n24858), .B1(n24863), .X(
        n25371) );
  sky130_fd_sc_hd__nor2_1 U23589 ( .A(n19326), .B(n21592), .Y(n25393) );
  sky130_fd_sc_hd__nor2_1 U23590 ( .A(n19623), .B(n19327), .Y(n19329) );
  sky130_fd_sc_hd__nor2_1 U23591 ( .A(n19623), .B(n19328), .Y(n19629) );
  sky130_fd_sc_hd__nand2_1 U23592 ( .A(n19596), .B(n19329), .Y(n19550) );
  sky130_fd_sc_hd__nand2_1 U23593 ( .A(n19552), .B(n19550), .Y(n19371) );
  sky130_fd_sc_hd__nor2_1 U23594 ( .A(n19623), .B(n19330), .Y(n19370) );
  sky130_fd_sc_hd__nor2_1 U23595 ( .A(n19370), .B(n19596), .Y(n19523) );
  sky130_fd_sc_hd__nor2_1 U23596 ( .A(n19623), .B(n19427), .Y(n19366) );
  sky130_fd_sc_hd__nor2_1 U23597 ( .A(n19366), .B(n19596), .Y(n19419) );
  sky130_fd_sc_hd__nor2_1 U23598 ( .A(n19623), .B(n19331), .Y(n19356) );
  sky130_fd_sc_hd__nor2_1 U23599 ( .A(n19356), .B(n19596), .Y(n19441) );
  sky130_fd_sc_hd__a222oi_1 U23600 ( .A1(n19334), .A2(n11170), .B1(n19333), 
        .B2(n11170), .C1(n19332), .C2(n11170), .Y(n19335) );
  sky130_fd_sc_hd__xnor2_1 U23602 ( .A(j202_soc_core_j22_cpu_ml_bufa[32]), .B(
        n19337), .Y(n19346) );
  sky130_fd_sc_hd__fa_1 U23604 ( .A(n19342), .B(n19341), .CIN(n19340), .COUT(
        n19353), .SUM(n16587) );
  sky130_fd_sc_hd__nor2_1 U23605 ( .A(n19352), .B(n19353), .Y(n19668) );
  sky130_fd_sc_hd__nand2_1 U23606 ( .A(n19343), .B(n19350), .Y(n19664) );
  sky130_fd_sc_hd__nor2_1 U23607 ( .A(n19668), .B(n19664), .Y(n19919) );
  sky130_fd_sc_hd__fa_1 U23608 ( .A(n19346), .B(n19345), .CIN(n19344), .COUT(
        n19354), .SUM(n19352) );
  sky130_fd_sc_hd__nand2_1 U23609 ( .A(n19919), .B(n19922), .Y(n19437) );
  sky130_fd_sc_hd__nor2_1 U23610 ( .A(n19441), .B(n19437), .Y(n19358) );
  sky130_fd_sc_hd__nand2_1 U23611 ( .A(n19347), .B(n19358), .Y(n19362) );
  sky130_fd_sc_hd__a21oi_1 U23612 ( .A1(n19351), .A2(n19350), .B1(n19349), .Y(
        n19665) );
  sky130_fd_sc_hd__nand2_1 U23613 ( .A(n19353), .B(n19352), .Y(n19669) );
  sky130_fd_sc_hd__nand2_1 U23615 ( .A(n19354), .B(n19596), .Y(n19921) );
  sky130_fd_sc_hd__a21oi_1 U23616 ( .A1(n19918), .A2(n19922), .B1(n19355), .Y(
        n19438) );
  sky130_fd_sc_hd__nand2_1 U23617 ( .A(n19596), .B(n19356), .Y(n19442) );
  sky130_fd_sc_hd__o21ai_1 U23618 ( .A1(n19441), .A2(n19438), .B1(n19442), .Y(
        n19357) );
  sky130_fd_sc_hd__a21oi_1 U23619 ( .A1(n19359), .A2(n19358), .B1(n19357), .Y(
        n19360) );
  sky130_fd_sc_hd__nor2_1 U23621 ( .A(n19623), .B(n19363), .Y(n19364) );
  sky130_fd_sc_hd__nand2_1 U23622 ( .A(n19596), .B(n19364), .Y(n20026) );
  sky130_fd_sc_hd__a21oi_1 U23623 ( .A1(n20028), .A2(n20027), .B1(n19365), .Y(
        n19423) );
  sky130_fd_sc_hd__nand2_1 U23624 ( .A(n19596), .B(n19366), .Y(n19420) );
  sky130_fd_sc_hd__nor2_1 U23626 ( .A(n19623), .B(n19367), .Y(n19368) );
  sky130_fd_sc_hd__nand2_1 U23627 ( .A(n19596), .B(n19368), .Y(n19389) );
  sky130_fd_sc_hd__a21oi_1 U23628 ( .A1(n19391), .A2(n19390), .B1(n19369), .Y(
        n19527) );
  sky130_fd_sc_hd__nand2_1 U23629 ( .A(n19596), .B(n19370), .Y(n19524) );
  sky130_fd_sc_hd__xnor2_1 U23631 ( .A(n19371), .B(n19553), .Y(n19372) );
  sky130_fd_sc_hd__a22oi_1 U23632 ( .A1(j202_soc_core_j22_cpu_ml_mach[23]), 
        .A2(n20032), .B1(n19372), .B2(n20030), .Y(n19374) );
  sky130_fd_sc_hd__nand2_1 U23633 ( .A(n21694), .B(n20025), .Y(n19373) );
  sky130_fd_sc_hd__nand2_1 U23634 ( .A(n19374), .B(n19373), .Y(n21830) );
  sky130_fd_sc_hd__a22oi_1 U23635 ( .A1(j202_soc_core_j22_cpu_ml_macl[23]), 
        .A2(n19953), .B1(n22233), .B2(n19959), .Y(n19375) );
  sky130_fd_sc_hd__o22ai_1 U23636 ( .A1(n20043), .A2(n19377), .B1(n22125), 
        .B2(n21833), .Y(n19378) );
  sky130_fd_sc_hd__a21oi_1 U23637 ( .A1(n21830), .A2(n22125), .B1(n19378), .Y(
        n20881) );
  sky130_fd_sc_hd__nor2_1 U23638 ( .A(j202_soc_core_j22_cpu_regop_Rs__1_), .B(
        n21212), .Y(n20053) );
  sky130_fd_sc_hd__nor2_1 U23639 ( .A(n21212), .B(n19981), .Y(n20047) );
  sky130_fd_sc_hd__nor2_1 U23640 ( .A(n21212), .B(n19986), .Y(n20048) );
  sky130_fd_sc_hd__a22oi_1 U23641 ( .A1(n20047), .A2(
        j202_soc_core_j22_cpu_rf_tmp[23]), .B1(n20048), .B2(
        j202_soc_core_j22_cpu_rf_gpr[503]), .Y(n19384) );
  sky130_fd_sc_hd__nor2_1 U23642 ( .A(n19971), .B(n21212), .Y(n20056) );
  sky130_fd_sc_hd__nor2_1 U23643 ( .A(n19975), .B(n21212), .Y(n20055) );
  sky130_fd_sc_hd__a22oi_1 U23644 ( .A1(n20056), .A2(
        j202_soc_core_j22_cpu_rf_pr[23]), .B1(j202_soc_core_j22_cpu_rf_gbr[23]), .B2(n20055), .Y(n19383) );
  sky130_fd_sc_hd__nor2_1 U23645 ( .A(n19977), .B(n21212), .Y(n20046) );
  sky130_fd_sc_hd__nand2_1 U23646 ( .A(n19985), .B(n19379), .Y(n19908) );
  sky130_fd_sc_hd__a2bb2oi_1 U23647 ( .B1(j202_soc_core_j22_cpu_pc[23]), .B2(
        n20046), .A1_N(n19380), .A2_N(n19908), .Y(n19382) );
  sky130_fd_sc_hd__nor2_1 U23648 ( .A(n19983), .B(n21212), .Y(n20057) );
  sky130_fd_sc_hd__nand2_1 U23649 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[23]), .Y(n19381) );
  sky130_fd_sc_hd__nand4_1 U23650 ( .A(n19384), .B(n19383), .C(n19382), .D(
        n19381), .Y(n19385) );
  sky130_fd_sc_hd__a21oi_1 U23651 ( .A1(n20053), .A2(n19386), .B1(n19385), .Y(
        n19387) );
  sky130_fd_sc_hd__o21a_1 U23652 ( .A1(n19466), .A2(n19917), .B1(n19387), .X(
        n19388) );
  sky130_fd_sc_hd__o211ai_1 U23653 ( .A1(n20067), .A2(n20881), .B1(n19388), 
        .C1(n19464), .Y(n25353) );
  sky130_fd_sc_hd__nand2_1 U23654 ( .A(n21709), .B(n20025), .Y(n19395) );
  sky130_fd_sc_hd__nand2_1 U23655 ( .A(n19390), .B(n19389), .Y(n19392) );
  sky130_fd_sc_hd__xnor2_1 U23656 ( .A(n19392), .B(n19391), .Y(n19393) );
  sky130_fd_sc_hd__a22oi_1 U23657 ( .A1(j202_soc_core_j22_cpu_ml_mach[21]), 
        .A2(n20032), .B1(n19393), .B2(n20030), .Y(n19394) );
  sky130_fd_sc_hd__nand2_1 U23658 ( .A(n19395), .B(n19394), .Y(n21748) );
  sky130_fd_sc_hd__nand2_1 U23659 ( .A(n22029), .B(n19959), .Y(n19397) );
  sky130_fd_sc_hd__a22oi_1 U23660 ( .A1(j202_soc_core_j22_cpu_ml_bufa[21]), 
        .A2(n22225), .B1(n19953), .B2(j202_soc_core_j22_cpu_ml_macl[21]), .Y(
        n19396) );
  sky130_fd_sc_hd__nand2_1 U23661 ( .A(n19397), .B(n19396), .Y(n19398) );
  sky130_fd_sc_hd__a21oi_1 U23662 ( .A1(n19399), .A2(n20040), .B1(n19398), .Y(
        n21750) );
  sky130_fd_sc_hd__o22ai_1 U23663 ( .A1(n19565), .A2(n19400), .B1(n22125), 
        .B2(n21750), .Y(n19401) );
  sky130_fd_sc_hd__a21oi_1 U23664 ( .A1(n21748), .A2(n22125), .B1(n19401), .Y(
        n20857) );
  sky130_fd_sc_hd__a22oi_1 U23665 ( .A1(n20047), .A2(
        j202_soc_core_j22_cpu_rf_tmp[21]), .B1(n20048), .B2(
        j202_soc_core_j22_cpu_rf_gpr[501]), .Y(n19406) );
  sky130_fd_sc_hd__a22oi_1 U23666 ( .A1(n20056), .A2(
        j202_soc_core_j22_cpu_rf_pr[21]), .B1(j202_soc_core_j22_cpu_rf_gbr[21]), .B2(n20055), .Y(n19405) );
  sky130_fd_sc_hd__a2bb2oi_1 U23667 ( .B1(j202_soc_core_j22_cpu_pc[21]), .B2(
        n20046), .A1_N(n19402), .A2_N(n19908), .Y(n19404) );
  sky130_fd_sc_hd__nand2_1 U23668 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[21]), .Y(n19403) );
  sky130_fd_sc_hd__nand4_1 U23669 ( .A(n19406), .B(n19405), .C(n19404), .D(
        n19403), .Y(n19407) );
  sky130_fd_sc_hd__a21oi_1 U23670 ( .A1(n20053), .A2(n19408), .B1(n19407), .Y(
        n19409) );
  sky130_fd_sc_hd__o21a_1 U23671 ( .A1(n19472), .A2(n19917), .B1(n19409), .X(
        n19410) );
  sky130_fd_sc_hd__o211ai_1 U23672 ( .A1(n20857), .A2(n20067), .B1(n19410), 
        .C1(n19470), .Y(n25351) );
  sky130_fd_sc_hd__a22oi_1 U23673 ( .A1(n20047), .A2(
        j202_soc_core_j22_cpu_rf_tmp[20]), .B1(n20048), .B2(
        j202_soc_core_j22_cpu_rf_gpr[500]), .Y(n19415) );
  sky130_fd_sc_hd__a22oi_1 U23674 ( .A1(n20056), .A2(
        j202_soc_core_j22_cpu_rf_pr[20]), .B1(j202_soc_core_j22_cpu_rf_gbr[20]), .B2(n20055), .Y(n19414) );
  sky130_fd_sc_hd__a2bb2oi_1 U23675 ( .B1(j202_soc_core_j22_cpu_pc[20]), .B2(
        n20046), .A1_N(n19411), .A2_N(n19908), .Y(n19413) );
  sky130_fd_sc_hd__nand2_1 U23676 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[20]), .Y(n19412) );
  sky130_fd_sc_hd__nand4_1 U23677 ( .A(n19415), .B(n19414), .C(n19413), .D(
        n19412), .Y(n19416) );
  sky130_fd_sc_hd__a21oi_1 U23678 ( .A1(n20053), .A2(n19417), .B1(n19416), .Y(
        n19418) );
  sky130_fd_sc_hd__o21a_1 U23679 ( .A1(n19476), .A2(n19917), .B1(n19418), .X(
        n19436) );
  sky130_fd_sc_hd__nand2_1 U23680 ( .A(n22204), .B(
        j202_soc_core_j22_cpu_ml_bufa[20]), .Y(n19426) );
  sky130_fd_sc_hd__nand2_1 U23681 ( .A(n19421), .B(n19420), .Y(n19422) );
  sky130_fd_sc_hd__xor2_1 U23682 ( .A(n19423), .B(n19422), .X(n19424) );
  sky130_fd_sc_hd__nand2_1 U23683 ( .A(n19424), .B(n20030), .Y(n19425) );
  sky130_fd_sc_hd__o211ai_1 U23684 ( .A1(n20005), .A2(n19427), .B1(n19426), 
        .C1(n19425), .Y(n19428) );
  sky130_fd_sc_hd__a21oi_1 U23685 ( .A1(n21704), .A2(n20025), .B1(n19428), .Y(
        n21737) );
  sky130_fd_sc_hd__nand2_1 U23686 ( .A(n19429), .B(n20040), .Y(n19433) );
  sky130_fd_sc_hd__a22o_1 U23687 ( .A1(j202_soc_core_j22_cpu_ml_bufa[20]), 
        .A2(n22225), .B1(n19953), .B2(j202_soc_core_j22_cpu_ml_macl[20]), .X(
        n19430) );
  sky130_fd_sc_hd__a21oi_1 U23688 ( .A1(n19431), .A2(n19959), .B1(n19430), .Y(
        n19432) );
  sky130_fd_sc_hd__nand2_1 U23689 ( .A(n19433), .B(n19432), .Y(n21739) );
  sky130_fd_sc_hd__nor2_1 U23690 ( .A(n22125), .B(n21739), .Y(n19434) );
  sky130_fd_sc_hd__a21oi_1 U23691 ( .A1(n21737), .A2(n22125), .B1(n19434), .Y(
        n20407) );
  sky130_fd_sc_hd__nand2_1 U23692 ( .A(n20407), .B(n20019), .Y(n19435) );
  sky130_fd_sc_hd__nand3_1 U23693 ( .A(n19474), .B(n19436), .C(n19435), .Y(
        n25350) );
  sky130_fd_sc_hd__a21oi_1 U23694 ( .A1(n19920), .A2(n19440), .B1(n19439), .Y(
        n19445) );
  sky130_fd_sc_hd__nand2_1 U23695 ( .A(n19443), .B(n19442), .Y(n19444) );
  sky130_fd_sc_hd__xor2_1 U23696 ( .A(n19445), .B(n19444), .X(n19446) );
  sky130_fd_sc_hd__nand2_1 U23697 ( .A(n19446), .B(n20030), .Y(n19449) );
  sky130_fd_sc_hd__nand2_1 U23698 ( .A(n21703), .B(n20025), .Y(n19448) );
  sky130_fd_sc_hd__nand2b_1 U23699 ( .A_N(n20005), .B(
        j202_soc_core_j22_cpu_ml_mach[18]), .Y(n19447) );
  sky130_fd_sc_hd__nand3_1 U23700 ( .A(n19449), .B(n19448), .C(n19447), .Y(
        n21777) );
  sky130_fd_sc_hd__a22oi_1 U23701 ( .A1(j202_soc_core_j22_cpu_ml_macl[18]), 
        .A2(n19953), .B1(n22236), .B2(n19959), .Y(n19450) );
  sky130_fd_sc_hd__o22ai_1 U23702 ( .A1(n20043), .A2(n19452), .B1(n22125), 
        .B2(n21780), .Y(n19453) );
  sky130_fd_sc_hd__a21oi_1 U23703 ( .A1(n21777), .A2(n22125), .B1(n19453), .Y(
        n20930) );
  sky130_fd_sc_hd__a22oi_1 U23704 ( .A1(n20047), .A2(
        j202_soc_core_j22_cpu_rf_tmp[18]), .B1(n20048), .B2(
        j202_soc_core_j22_cpu_rf_gpr[498]), .Y(n19458) );
  sky130_fd_sc_hd__a22oi_1 U23705 ( .A1(n20056), .A2(
        j202_soc_core_j22_cpu_rf_pr[18]), .B1(j202_soc_core_j22_cpu_rf_gbr[18]), .B2(n20055), .Y(n19457) );
  sky130_fd_sc_hd__a2bb2oi_1 U23706 ( .B1(j202_soc_core_j22_cpu_pc[18]), .B2(
        n20046), .A1_N(n19454), .A2_N(n19908), .Y(n19456) );
  sky130_fd_sc_hd__nand2_1 U23707 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[18]), .Y(n19455) );
  sky130_fd_sc_hd__nand4_1 U23708 ( .A(n19458), .B(n19457), .C(n19456), .D(
        n19455), .Y(n19459) );
  sky130_fd_sc_hd__a21oi_1 U23709 ( .A1(n20053), .A2(n19460), .B1(n19459), .Y(
        n19461) );
  sky130_fd_sc_hd__o21a_1 U23710 ( .A1(n19506), .A2(n19917), .B1(n19461), .X(
        n19462) );
  sky130_fd_sc_hd__o211ai_1 U23711 ( .A1(n20930), .A2(n20067), .B1(n19462), 
        .C1(n19504), .Y(n25348) );
  sky130_fd_sc_hd__nand2_1 U23712 ( .A(n19463), .B(n20019), .Y(n19465) );
  sky130_fd_sc_hd__o211ai_1 U23713 ( .A1(n19907), .A2(n19466), .B1(n19465), 
        .C1(n19464), .Y(n25366) );
  sky130_fd_sc_hd__nand2_1 U23714 ( .A(n19467), .B(n20019), .Y(n19468) );
  sky130_fd_sc_hd__o211ai_1 U23715 ( .A1(n19907), .A2(n19546), .B1(n19468), 
        .C1(n19547), .Y(n25300) );
  sky130_fd_sc_hd__nand2_1 U23716 ( .A(n19469), .B(n20019), .Y(n19471) );
  sky130_fd_sc_hd__o211ai_1 U23717 ( .A1(n19907), .A2(n19472), .B1(n19471), 
        .C1(n19470), .Y(n25365) );
  sky130_fd_sc_hd__nand2_1 U23718 ( .A(n19473), .B(n20019), .Y(n19475) );
  sky130_fd_sc_hd__o211ai_1 U23719 ( .A1(n19907), .A2(n19476), .B1(n19475), 
        .C1(n19474), .Y(n25364) );
  sky130_fd_sc_hd__nor2_1 U23720 ( .A(n21443), .B(
        j202_soc_core_j22_cpu_opst[3]), .Y(n20500) );
  sky130_fd_sc_hd__nand2_1 U23721 ( .A(n24879), .B(n20500), .Y(n22416) );
  sky130_fd_sc_hd__nor2_1 U23722 ( .A(n23229), .B(n24858), .Y(n21607) );
  sky130_fd_sc_hd__nand2_1 U23723 ( .A(n25304), .B(n25316), .Y(n20326) );
  sky130_fd_sc_hd__nor2_1 U23724 ( .A(n21418), .B(n20326), .Y(n21533) );
  sky130_fd_sc_hd__nor2_1 U23725 ( .A(n25258), .B(n20343), .Y(n20981) );
  sky130_fd_sc_hd__nand2_1 U23726 ( .A(n22342), .B(n24826), .Y(n21536) );
  sky130_fd_sc_hd__nand2_1 U23727 ( .A(n25387), .B(n21461), .Y(n24860) );
  sky130_fd_sc_hd__nor2_1 U23728 ( .A(n20343), .B(n22762), .Y(n21336) );
  sky130_fd_sc_hd__nor2_1 U23729 ( .A(n22342), .B(n21534), .Y(n24867) );
  sky130_fd_sc_hd__nor2b_1 U23730 ( .B_N(n24860), .A(n24867), .Y(n20753) );
  sky130_fd_sc_hd__nor2_1 U23731 ( .A(n25372), .B(n25377), .Y(n22733) );
  sky130_fd_sc_hd__nand2_1 U23732 ( .A(n25380), .B(n25381), .Y(n20985) );
  sky130_fd_sc_hd__nor2_1 U23733 ( .A(n25377), .B(n20985), .Y(n21454) );
  sky130_fd_sc_hd__a31oi_1 U23734 ( .A1(n22733), .A2(n25381), .A3(n25386), 
        .B1(n21454), .Y(n19478) );
  sky130_fd_sc_hd__nor2_1 U23735 ( .A(n22330), .B(n22333), .Y(n20986) );
  sky130_fd_sc_hd__nor2_1 U23736 ( .A(n21487), .B(n21640), .Y(n20328) );
  sky130_fd_sc_hd__a21oi_1 U23738 ( .A1(n19478), .A2(n19477), .B1(n20335), .Y(
        n19492) );
  sky130_fd_sc_hd__nand2_1 U23739 ( .A(n25316), .B(n19479), .Y(n21734) );
  sky130_fd_sc_hd__nor2_1 U23740 ( .A(n21418), .B(n21734), .Y(n20339) );
  sky130_fd_sc_hd__nor2_1 U23741 ( .A(n22762), .B(n22309), .Y(n20979) );
  sky130_fd_sc_hd__nor3b_1 U23742 ( .C_N(n20339), .A(n20761), .B(n20979), .Y(
        n19491) );
  sky130_fd_sc_hd__nor3b_1 U23743 ( .C_N(n25303), .A(n21586), .B(n19480), .Y(
        n22735) );
  sky130_fd_sc_hd__nor2_1 U23744 ( .A(n20742), .B(n22742), .Y(n20989) );
  sky130_fd_sc_hd__a31oi_1 U23745 ( .A1(n24872), .A2(n24873), .A3(n20328), 
        .B1(n20989), .Y(n19482) );
  sky130_fd_sc_hd__nand2_1 U23746 ( .A(n25303), .B(n25315), .Y(n19481) );
  sky130_fd_sc_hd__o22ai_1 U23747 ( .A1(n19482), .A2(n25381), .B1(n20326), 
        .B2(n19481), .Y(n19490) );
  sky130_fd_sc_hd__nor2_1 U23748 ( .A(n25380), .B(n25381), .Y(n20996) );
  sky130_fd_sc_hd__o21ai_0 U23749 ( .A1(n22330), .A2(n24827), .B1(n25377), .Y(
        n19486) );
  sky130_fd_sc_hd__nor2_1 U23750 ( .A(n25385), .B(n25387), .Y(n24869) );
  sky130_fd_sc_hd__nand3_1 U23751 ( .A(n22762), .B(n22342), .C(n24869), .Y(
        n20330) );
  sky130_fd_sc_hd__o21ai_0 U23752 ( .A1(n22330), .A2(n19483), .B1(n22328), .Y(
        n19484) );
  sky130_fd_sc_hd__nand2_1 U23753 ( .A(n25380), .B(n22328), .Y(n21573) );
  sky130_fd_sc_hd__nor2_1 U23754 ( .A(n21574), .B(n21573), .Y(n21564) );
  sky130_fd_sc_hd__a22oi_1 U23756 ( .A1(n20996), .A2(n19486), .B1(n20330), 
        .B2(n19485), .Y(n19488) );
  sky130_fd_sc_hd__nand2_1 U23757 ( .A(n25258), .B(n20339), .Y(n22389) );
  sky130_fd_sc_hd__nor2_1 U23758 ( .A(n22342), .B(n25387), .Y(n24825) );
  sky130_fd_sc_hd__a22oi_1 U23759 ( .A1(n21635), .A2(n21331), .B1(n21424), 
        .B2(n24825), .Y(n19487) );
  sky130_fd_sc_hd__o21ai_1 U23760 ( .A1(n19488), .A2(n21455), .B1(n19487), .Y(
        n19489) );
  sky130_fd_sc_hd__nor4_1 U23761 ( .A(n19492), .B(n19491), .C(n19490), .D(
        n19489), .Y(n24861) );
  sky130_fd_sc_hd__nor2_1 U23762 ( .A(n25372), .B(n22333), .Y(n21416) );
  sky130_fd_sc_hd__nand2_1 U23763 ( .A(n21416), .B(n21575), .Y(n21474) );
  sky130_fd_sc_hd__nand2_1 U23764 ( .A(n21480), .B(n19493), .Y(n21330) );
  sky130_fd_sc_hd__nand2_1 U23765 ( .A(n20331), .B(n21564), .Y(n24884) );
  sky130_fd_sc_hd__nor2_1 U23766 ( .A(n20327), .B(n25316), .Y(n21609) );
  sky130_fd_sc_hd__nand2_1 U23767 ( .A(n21609), .B(n25304), .Y(n22390) );
  sky130_fd_sc_hd__nand2_1 U23768 ( .A(n21420), .B(n21563), .Y(n20998) );
  sky130_fd_sc_hd__nor2_1 U23769 ( .A(n20986), .B(n20998), .Y(n24833) );
  sky130_fd_sc_hd__a21oi_1 U23770 ( .A1(n24833), .A2(n25381), .B1(n23229), .Y(
        n21493) );
  sky130_fd_sc_hd__and4_1 U23771 ( .A(n20753), .B(n24861), .C(n21537), .D(
        n21493), .X(n19494) );
  sky130_fd_sc_hd__o22ai_1 U23772 ( .A1(j202_soc_core_j22_cpu_opst[2]), .A2(
        n22416), .B1(n21607), .B2(n19494), .Y(n25305) );
  sky130_fd_sc_hd__nand2_1 U23773 ( .A(j202_soc_core_aquc_SEL__0_), .B(
        j202_soc_core_aquc_CE__1_), .Y(n19495) );
  sky130_fd_sc_hd__nor2_1 U23774 ( .A(j202_soc_core_aquc_WE_), .B(n19495), .Y(
        n25394) );
  sky130_fd_sc_hd__nand2_1 U23775 ( .A(n25259), .B(n19737), .Y(n19498) );
  sky130_fd_sc_hd__a22oi_1 U23776 ( .A1(n19657), .A2(n22584), .B1(n19736), 
        .B2(n22185), .Y(n19497) );
  sky130_fd_sc_hd__a22oi_1 U23777 ( .A1(j202_soc_core_j22_cpu_pc[0]), .A2(
        n19661), .B1(n21625), .B2(n19729), .Y(n19496) );
  sky130_fd_sc_hd__nand2_1 U23778 ( .A(n19690), .B(n19500), .Y(n19501) );
  sky130_fd_sc_hd__o211ai_1 U23779 ( .A1(n19502), .A2(n20067), .B1(n19501), 
        .C1(n19691), .Y(n25341) );
  sky130_fd_sc_hd__nand2_1 U23780 ( .A(n19503), .B(n20019), .Y(n19505) );
  sky130_fd_sc_hd__o211ai_1 U23781 ( .A1(n19907), .A2(n19506), .B1(n19505), 
        .C1(n19504), .Y(n25360) );
  sky130_fd_sc_hd__a21oi_1 U23782 ( .A1(n19510), .A2(n19509), .B1(n19508), .Y(
        n19515) );
  sky130_fd_sc_hd__nand2_1 U23783 ( .A(n19513), .B(n19512), .Y(n19514) );
  sky130_fd_sc_hd__xor2_1 U23784 ( .A(n19515), .B(n19514), .X(n21809) );
  sky130_fd_sc_hd__nand2_1 U23785 ( .A(n21809), .B(n19729), .Y(n19522) );
  sky130_fd_sc_hd__ha_1 U23786 ( .A(j202_soc_core_j22_cpu_pc[10]), .B(n19516), 
        .COUT(n18844), .SUM(n21806) );
  sky130_fd_sc_hd__a22oi_1 U23787 ( .A1(n19657), .A2(n20935), .B1(n21806), 
        .B2(n19517), .Y(n19519) );
  sky130_fd_sc_hd__a22oi_1 U23788 ( .A1(n25314), .A2(n19737), .B1(n21806), 
        .B2(n19732), .Y(n19518) );
  sky130_fd_sc_hd__o211a_2 U23789 ( .A1(n19520), .A2(n21807), .B1(n19519), 
        .C1(n19518), .X(n19521) );
  sky130_fd_sc_hd__nand2_1 U23790 ( .A(n19522), .B(n19521), .Y(n25373) );
  sky130_fd_sc_hd__nand2_1 U23791 ( .A(n21708), .B(n20025), .Y(n19531) );
  sky130_fd_sc_hd__nand2_1 U23792 ( .A(n19525), .B(n19524), .Y(n19526) );
  sky130_fd_sc_hd__xor2_1 U23793 ( .A(n19527), .B(n19526), .X(n19528) );
  sky130_fd_sc_hd__nand2_1 U23794 ( .A(n19528), .B(n20030), .Y(n19530) );
  sky130_fd_sc_hd__nand2b_1 U23795 ( .A_N(n20005), .B(
        j202_soc_core_j22_cpu_ml_mach[22]), .Y(n19529) );
  sky130_fd_sc_hd__nand3_1 U23796 ( .A(n19531), .B(n19530), .C(n19529), .Y(
        n21869) );
  sky130_fd_sc_hd__o22ai_1 U23797 ( .A1(n20038), .A2(n19533), .B1(n20036), 
        .B2(n19532), .Y(n19534) );
  sky130_fd_sc_hd__a21oi_1 U23798 ( .A1(n19535), .A2(n20040), .B1(n19534), .Y(
        n21872) );
  sky130_fd_sc_hd__o22ai_1 U23799 ( .A1(n20043), .A2(n19536), .B1(n22125), 
        .B2(n21872), .Y(n19537) );
  sky130_fd_sc_hd__a21oi_1 U23800 ( .A1(n21869), .A2(n22125), .B1(n19537), .Y(
        n21138) );
  sky130_fd_sc_hd__a22oi_1 U23801 ( .A1(n20047), .A2(
        j202_soc_core_j22_cpu_rf_tmp[22]), .B1(n20048), .B2(
        j202_soc_core_j22_cpu_rf_gpr[502]), .Y(n19542) );
  sky130_fd_sc_hd__a22oi_1 U23802 ( .A1(n20056), .A2(
        j202_soc_core_j22_cpu_rf_pr[22]), .B1(j202_soc_core_j22_cpu_rf_gbr[22]), .B2(n20055), .Y(n19541) );
  sky130_fd_sc_hd__a2bb2oi_1 U23803 ( .B1(j202_soc_core_j22_cpu_pc[22]), .B2(
        n20046), .A1_N(n19538), .A2_N(n19908), .Y(n19540) );
  sky130_fd_sc_hd__nand2_1 U23804 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[22]), .Y(n19539) );
  sky130_fd_sc_hd__nand4_1 U23805 ( .A(n19542), .B(n19541), .C(n19540), .D(
        n19539), .Y(n19543) );
  sky130_fd_sc_hd__a21oi_1 U23806 ( .A1(n20053), .A2(n19544), .B1(n19543), .Y(
        n19545) );
  sky130_fd_sc_hd__o21a_1 U23807 ( .A1(n19546), .A2(n19917), .B1(n19545), .X(
        n19548) );
  sky130_fd_sc_hd__o211ai_1 U23808 ( .A1(n21138), .A2(n20067), .B1(n19548), 
        .C1(n19547), .Y(n25352) );
  sky130_fd_sc_hd__nor2_1 U23809 ( .A(n19623), .B(n19549), .Y(n19554) );
  sky130_fd_sc_hd__nor2_1 U23810 ( .A(n19554), .B(n19596), .Y(n19694) );
  sky130_fd_sc_hd__a21oi_1 U23811 ( .A1(n19553), .A2(n19552), .B1(n19551), .Y(
        n19698) );
  sky130_fd_sc_hd__nand2_1 U23812 ( .A(n19596), .B(n19554), .Y(n19695) );
  sky130_fd_sc_hd__o21ai_1 U23813 ( .A1(n19694), .A2(n19698), .B1(n19695), .Y(
        n19938) );
  sky130_fd_sc_hd__nor2_1 U23814 ( .A(n19623), .B(n19555), .Y(n19556) );
  sky130_fd_sc_hd__nand2_1 U23815 ( .A(n19596), .B(n19556), .Y(n19936) );
  sky130_fd_sc_hd__a21oi_1 U23816 ( .A1(n19938), .A2(n19937), .B1(n19557), .Y(
        n19590) );
  sky130_fd_sc_hd__nor2_1 U23817 ( .A(n19623), .B(n19558), .Y(n19559) );
  sky130_fd_sc_hd__nor2_1 U23818 ( .A(n19559), .B(n19596), .Y(n19591) );
  sky130_fd_sc_hd__nand2_1 U23819 ( .A(n19596), .B(n19559), .Y(n19589) );
  sky130_fd_sc_hd__nand2_1 U23820 ( .A(n19560), .B(n19589), .Y(n19561) );
  sky130_fd_sc_hd__xor2_1 U23821 ( .A(n19590), .B(n19561), .X(n19562) );
  sky130_fd_sc_hd__nand2_1 U23822 ( .A(n19562), .B(n20030), .Y(n19564) );
  sky130_fd_sc_hd__a22oi_1 U23823 ( .A1(j202_soc_core_j22_cpu_ml_mach[26]), 
        .A2(n20032), .B1(n21692), .B2(n20025), .Y(n19563) );
  sky130_fd_sc_hd__nand2_1 U23824 ( .A(n19564), .B(n19563), .Y(n22199) );
  sky130_fd_sc_hd__nand2_1 U23825 ( .A(n22199), .B(n22125), .Y(n19571) );
  sky130_fd_sc_hd__nand2_1 U23826 ( .A(n19566), .B(n20040), .Y(n19569) );
  sky130_fd_sc_hd__a22oi_1 U23827 ( .A1(j202_soc_core_j22_cpu_ml_bufa[26]), 
        .A2(n22225), .B1(n19953), .B2(j202_soc_core_j22_cpu_ml_macl[26]), .Y(
        n19568) );
  sky130_fd_sc_hd__nand2_1 U23828 ( .A(n21797), .B(n19959), .Y(n19567) );
  sky130_fd_sc_hd__nand3_1 U23829 ( .A(n19569), .B(n19568), .C(n19567), .Y(
        n22220) );
  sky130_fd_sc_hd__a22oi_1 U23830 ( .A1(n19963), .A2(
        j202_soc_core_j22_cpu_ml_bufa[26]), .B1(n22220), .B2(
        j202_soc_core_j22_cpu_macop_MAC_[0]), .Y(n19570) );
  sky130_fd_sc_hd__nand2_1 U23831 ( .A(n19571), .B(n19570), .Y(n20828) );
  sky130_fd_sc_hd__nand2_1 U23832 ( .A(n20828), .B(n20019), .Y(n19585) );
  sky130_fd_sc_hd__nand2_1 U23833 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[26]), .Y(n19574) );
  sky130_fd_sc_hd__nand2_1 U23834 ( .A(n20056), .B(
        j202_soc_core_j22_cpu_rf_pr[26]), .Y(n19573) );
  sky130_fd_sc_hd__nand2_1 U23835 ( .A(n20055), .B(
        j202_soc_core_j22_cpu_rf_gbr[26]), .Y(n19572) );
  sky130_fd_sc_hd__nand3_1 U23836 ( .A(n19574), .B(n19573), .C(n19572), .Y(
        n19580) );
  sky130_fd_sc_hd__nand2_1 U23837 ( .A(n19575), .B(n20053), .Y(n19579) );
  sky130_fd_sc_hd__a2bb2oi_1 U23838 ( .B1(j202_soc_core_j22_cpu_pc[26]), .B2(
        n20046), .A1_N(n19576), .A2_N(n19908), .Y(n19578) );
  sky130_fd_sc_hd__a22oi_1 U23839 ( .A1(n20047), .A2(
        j202_soc_core_j22_cpu_rf_tmp[26]), .B1(n20048), .B2(
        j202_soc_core_j22_cpu_rf_gpr[506]), .Y(n19577) );
  sky130_fd_sc_hd__nand4b_1 U23840 ( .A_N(n19580), .B(n19579), .C(n19578), .D(
        n19577), .Y(n19581) );
  sky130_fd_sc_hd__a21oi_1 U23841 ( .A1(n19582), .A2(n21222), .B1(n19581), .Y(
        n19583) );
  sky130_fd_sc_hd__nand3_1 U23842 ( .A(n19585), .B(n19584), .C(n19583), .Y(
        n25356) );
  sky130_fd_sc_hd__nor2_1 U23843 ( .A(n19623), .B(n19586), .Y(n19587) );
  sky130_fd_sc_hd__or2_0 U23844 ( .A(n19587), .B(n19596), .X(n19627) );
  sky130_fd_sc_hd__nand2_1 U23845 ( .A(n19596), .B(n19587), .Y(n19625) );
  sky130_fd_sc_hd__nand2_1 U23846 ( .A(n19627), .B(n19625), .Y(n19597) );
  sky130_fd_sc_hd__nor2_1 U23847 ( .A(n19623), .B(n19588), .Y(n19595) );
  sky130_fd_sc_hd__nor2_1 U23848 ( .A(n19595), .B(n19596), .Y(n19769) );
  sky130_fd_sc_hd__o21ai_1 U23849 ( .A1(n19591), .A2(n19590), .B1(n19589), .Y(
        n19805) );
  sky130_fd_sc_hd__nor2_1 U23850 ( .A(n19623), .B(n19592), .Y(n19593) );
  sky130_fd_sc_hd__or2_0 U23851 ( .A(n19593), .B(n19596), .X(n19804) );
  sky130_fd_sc_hd__nand2_1 U23852 ( .A(n19596), .B(n19593), .Y(n19803) );
  sky130_fd_sc_hd__a21oi_1 U23853 ( .A1(n19805), .A2(n19804), .B1(n19594), .Y(
        n19773) );
  sky130_fd_sc_hd__nand2_1 U23854 ( .A(n19596), .B(n19595), .Y(n19770) );
  sky130_fd_sc_hd__o21ai_1 U23855 ( .A1(n19769), .A2(n19773), .B1(n19770), .Y(
        n19628) );
  sky130_fd_sc_hd__xnor2_1 U23856 ( .A(n19597), .B(n19628), .Y(n19598) );
  sky130_fd_sc_hd__nand2_1 U23857 ( .A(n19598), .B(n20030), .Y(n19600) );
  sky130_fd_sc_hd__a22oi_1 U23858 ( .A1(j202_soc_core_j22_cpu_ml_mach[29]), 
        .A2(n20032), .B1(n21696), .B2(n20025), .Y(n19599) );
  sky130_fd_sc_hd__nand2_1 U23859 ( .A(n19600), .B(n19599), .Y(n21742) );
  sky130_fd_sc_hd__nand2_1 U23860 ( .A(n21742), .B(n22125), .Y(n19606) );
  sky130_fd_sc_hd__nand2_1 U23861 ( .A(n19601), .B(n20040), .Y(n19603) );
  sky130_fd_sc_hd__a22oi_1 U23862 ( .A1(j202_soc_core_j22_cpu_ml_macl[29]), 
        .A2(n19953), .B1(n22230), .B2(n19959), .Y(n19602) );
  sky130_fd_sc_hd__nand2_1 U23863 ( .A(n19603), .B(n19602), .Y(n21745) );
  sky130_fd_sc_hd__nand2_1 U23864 ( .A(n21745), .B(
        j202_soc_core_j22_cpu_macop_MAC_[0]), .Y(n19605) );
  sky130_fd_sc_hd__nand2_1 U23865 ( .A(n19931), .B(
        j202_soc_core_j22_cpu_ml_bufa[29]), .Y(n19604) );
  sky130_fd_sc_hd__nand3_1 U23866 ( .A(n19606), .B(n19605), .C(n19604), .Y(
        n20402) );
  sky130_fd_sc_hd__nand2_1 U23867 ( .A(n20402), .B(n20019), .Y(n19620) );
  sky130_fd_sc_hd__nand2_1 U23868 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[29]), .Y(n19609) );
  sky130_fd_sc_hd__nand2_1 U23869 ( .A(n20056), .B(
        j202_soc_core_j22_cpu_rf_pr[29]), .Y(n19608) );
  sky130_fd_sc_hd__nand2_1 U23870 ( .A(n20055), .B(
        j202_soc_core_j22_cpu_rf_gbr[29]), .Y(n19607) );
  sky130_fd_sc_hd__nand3_1 U23871 ( .A(n19609), .B(n19608), .C(n19607), .Y(
        n19615) );
  sky130_fd_sc_hd__nand2_1 U23872 ( .A(n19610), .B(n20053), .Y(n19614) );
  sky130_fd_sc_hd__a2bb2oi_1 U23873 ( .B1(j202_soc_core_j22_cpu_pc[29]), .B2(
        n20046), .A1_N(n19611), .A2_N(n19908), .Y(n19613) );
  sky130_fd_sc_hd__a22oi_1 U23874 ( .A1(n20047), .A2(
        j202_soc_core_j22_cpu_rf_tmp[29]), .B1(n20048), .B2(
        j202_soc_core_j22_cpu_rf_gpr[509]), .Y(n19612) );
  sky130_fd_sc_hd__nand4b_1 U23875 ( .A_N(n19615), .B(n19614), .C(n19613), .D(
        n19612), .Y(n19616) );
  sky130_fd_sc_hd__a21oi_1 U23876 ( .A1(n19617), .A2(n21222), .B1(n19616), .Y(
        n19618) );
  sky130_fd_sc_hd__nand3_1 U23877 ( .A(n19620), .B(n19619), .C(n19618), .Y(
        n25359) );
  sky130_fd_sc_hd__or2_0 U23878 ( .A(n19621), .B(n19623), .X(n19630) );
  sky130_fd_sc_hd__nor2_1 U23879 ( .A(n19623), .B(n19622), .Y(n19624) );
  sky130_fd_sc_hd__xor2_1 U23880 ( .A(n19630), .B(n19624), .X(n19632) );
  sky130_fd_sc_hd__nor2_1 U23881 ( .A(n19629), .B(n19630), .Y(n19743) );
  sky130_fd_sc_hd__a21oi_1 U23882 ( .A1(n19628), .A2(n19627), .B1(n19626), .Y(
        n19747) );
  sky130_fd_sc_hd__nand2_1 U23883 ( .A(n19630), .B(n19629), .Y(n19744) );
  sky130_fd_sc_hd__o21ai_1 U23884 ( .A1(n19743), .A2(n19747), .B1(n19744), .Y(
        n19631) );
  sky130_fd_sc_hd__xor2_1 U23885 ( .A(n19632), .B(n19631), .X(n19633) );
  sky130_fd_sc_hd__nand2_1 U23886 ( .A(n19633), .B(n20030), .Y(n19635) );
  sky130_fd_sc_hd__a22oi_1 U23887 ( .A1(j202_soc_core_j22_cpu_ml_mach[31]), 
        .A2(n20032), .B1(n21695), .B2(n20025), .Y(n19634) );
  sky130_fd_sc_hd__nand2_1 U23888 ( .A(n19635), .B(n19634), .Y(n22194) );
  sky130_fd_sc_hd__nand2_1 U23889 ( .A(n22194), .B(n22125), .Y(n19640) );
  sky130_fd_sc_hd__nand2_1 U23890 ( .A(n21701), .B(n20040), .Y(n19637) );
  sky130_fd_sc_hd__a22oi_1 U23891 ( .A1(j202_soc_core_j22_cpu_ml_macl[31]), 
        .A2(n19953), .B1(n22227), .B2(n19959), .Y(n19636) );
  sky130_fd_sc_hd__nand2_1 U23892 ( .A(n19637), .B(n19636), .Y(n22193) );
  sky130_fd_sc_hd__nand2_1 U23893 ( .A(n22193), .B(
        j202_soc_core_j22_cpu_macop_MAC_[0]), .Y(n19639) );
  sky130_fd_sc_hd__nand2_1 U23894 ( .A(n19931), .B(
        j202_soc_core_j22_cpu_ml_bufa[31]), .Y(n19638) );
  sky130_fd_sc_hd__nand3_1 U23895 ( .A(n19640), .B(n19639), .C(n19638), .Y(
        n21006) );
  sky130_fd_sc_hd__nand2_1 U23896 ( .A(n21006), .B(n20019), .Y(n19652) );
  sky130_fd_sc_hd__a22oi_1 U23897 ( .A1(n20047), .A2(
        j202_soc_core_j22_cpu_rf_tmp[31]), .B1(n20048), .B2(
        j202_soc_core_j22_cpu_rf_gpr[511]), .Y(n19645) );
  sky130_fd_sc_hd__a22oi_1 U23898 ( .A1(n20056), .A2(
        j202_soc_core_j22_cpu_rf_pr[31]), .B1(j202_soc_core_j22_cpu_rf_gbr[31]), .B2(n20055), .Y(n19644) );
  sky130_fd_sc_hd__a2bb2oi_1 U23899 ( .B1(j202_soc_core_j22_cpu_pc[31]), .B2(
        n20046), .A1_N(n19641), .A2_N(n19908), .Y(n19643) );
  sky130_fd_sc_hd__nand2_1 U23900 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[31]), .Y(n19642) );
  sky130_fd_sc_hd__nand4_1 U23901 ( .A(n19645), .B(n19644), .C(n19643), .D(
        n19642), .Y(n19646) );
  sky130_fd_sc_hd__a21oi_1 U23902 ( .A1(n20053), .A2(n19647), .B1(n19646), .Y(
        n19648) );
  sky130_fd_sc_hd__o21a_1 U23903 ( .A1(n19764), .A2(n19649), .B1(n19648), .X(
        n19650) );
  sky130_fd_sc_hd__nand3_1 U23904 ( .A(n19652), .B(n19651), .C(n19650), .Y(
        n25362) );
  sky130_fd_sc_hd__nand2_1 U23905 ( .A(n11186), .B(n19653), .Y(n19655) );
  sky130_fd_sc_hd__xnor2_1 U23906 ( .A(n19655), .B(n19654), .Y(n22273) );
  sky130_fd_sc_hd__nand2_1 U23907 ( .A(n22273), .B(n19729), .Y(n19663) );
  sky130_fd_sc_hd__ha_1 U23908 ( .A(j202_soc_core_j22_cpu_pc[15]), .B(n19656), 
        .COUT(n18486), .SUM(n22277) );
  sky130_fd_sc_hd__nand2_1 U23909 ( .A(n25388), .B(n19737), .Y(n19659) );
  sky130_fd_sc_hd__a22oi_1 U23910 ( .A1(n19657), .A2(n22136), .B1(n19736), 
        .B2(n22154), .Y(n19658) );
  sky130_fd_sc_hd__nand2_1 U23911 ( .A(n19659), .B(n19658), .Y(n19660) );
  sky130_fd_sc_hd__a21oi_1 U23912 ( .A1(n22277), .A2(n19661), .B1(n19660), .Y(
        n19662) );
  sky130_fd_sc_hd__nand2_1 U23913 ( .A(n19663), .B(n19662), .Y(n25261) );
  sky130_fd_sc_hd__nand2_1 U23914 ( .A(n21731), .B(n20030), .Y(n19674) );
  sky130_fd_sc_hd__a22oi_1 U23915 ( .A1(j202_soc_core_j22_cpu_ml_mach[16]), 
        .A2(n20032), .B1(n21702), .B2(n20025), .Y(n19673) );
  sky130_fd_sc_hd__nand2_1 U23916 ( .A(n19674), .B(n19673), .Y(n22201) );
  sky130_fd_sc_hd__nand2_1 U23917 ( .A(n22201), .B(n22125), .Y(n19679) );
  sky130_fd_sc_hd__nand2_1 U23918 ( .A(n19675), .B(n20040), .Y(n19677) );
  sky130_fd_sc_hd__a22oi_1 U23919 ( .A1(j202_soc_core_j22_cpu_ml_macl[16]), 
        .A2(n19953), .B1(n22242), .B2(n19959), .Y(n19676) );
  sky130_fd_sc_hd__nand2_1 U23920 ( .A(n19677), .B(n19676), .Y(n22223) );
  sky130_fd_sc_hd__a22oi_1 U23921 ( .A1(j202_soc_core_j22_cpu_ml_bufa[16]), 
        .A2(n19931), .B1(n22223), .B2(j202_soc_core_j22_cpu_macop_MAC_[0]), 
        .Y(n19678) );
  sky130_fd_sc_hd__nand2_1 U23922 ( .A(n19679), .B(n19678), .Y(n20926) );
  sky130_fd_sc_hd__nand2_1 U23923 ( .A(n20926), .B(n20019), .Y(n19693) );
  sky130_fd_sc_hd__clkinv_1 U23924 ( .A(n19908), .Y(n20045) );
  sky130_fd_sc_hd__nand2_1 U23925 ( .A(n20045), .B(
        j202_soc_core_j22_cpu_rf_vbr[16]), .Y(n19683) );
  sky130_fd_sc_hd__nand2_1 U23926 ( .A(n20046), .B(
        j202_soc_core_j22_cpu_pc[16]), .Y(n19682) );
  sky130_fd_sc_hd__nand2_1 U23927 ( .A(n20047), .B(
        j202_soc_core_j22_cpu_rf_tmp[16]), .Y(n19681) );
  sky130_fd_sc_hd__nand2_1 U23928 ( .A(n20048), .B(
        j202_soc_core_j22_cpu_rf_gpr[496]), .Y(n19680) );
  sky130_fd_sc_hd__nand4_1 U23929 ( .A(n19683), .B(n19682), .C(n19681), .D(
        n19680), .Y(n19688) );
  sky130_fd_sc_hd__nand2_1 U23930 ( .A(n19684), .B(n20053), .Y(n19687) );
  sky130_fd_sc_hd__a22oi_1 U23931 ( .A1(n20056), .A2(
        j202_soc_core_j22_cpu_rf_pr[16]), .B1(j202_soc_core_j22_cpu_rf_gbr[16]), .B2(n20055), .Y(n19686) );
  sky130_fd_sc_hd__nand2_1 U23932 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[16]), .Y(n19685) );
  sky130_fd_sc_hd__nand4b_1 U23933 ( .A_N(n19688), .B(n19687), .C(n19686), .D(
        n19685), .Y(n19689) );
  sky130_fd_sc_hd__a21oi_1 U23934 ( .A1(n19690), .A2(n20064), .B1(n19689), .Y(
        n19692) );
  sky130_fd_sc_hd__nand3_1 U23935 ( .A(n19693), .B(n19692), .C(n19691), .Y(
        n25346) );
  sky130_fd_sc_hd__nand2_1 U23936 ( .A(n19696), .B(n19695), .Y(n19697) );
  sky130_fd_sc_hd__xor2_1 U23937 ( .A(n19698), .B(n19697), .X(n19699) );
  sky130_fd_sc_hd__nand2_1 U23938 ( .A(n19699), .B(n20030), .Y(n19702) );
  sky130_fd_sc_hd__nand2_1 U23939 ( .A(n21717), .B(n20025), .Y(n19701) );
  sky130_fd_sc_hd__nand2b_1 U23940 ( .A_N(n20005), .B(
        j202_soc_core_j22_cpu_ml_mach[24]), .Y(n19700) );
  sky130_fd_sc_hd__nand3_1 U23941 ( .A(n19702), .B(n19701), .C(n19700), .Y(
        n21938) );
  sky130_fd_sc_hd__nand2_1 U23942 ( .A(n21938), .B(n22125), .Y(n19708) );
  sky130_fd_sc_hd__nand2_1 U23943 ( .A(n19703), .B(n20040), .Y(n19706) );
  sky130_fd_sc_hd__a22oi_1 U23944 ( .A1(j202_soc_core_j22_cpu_ml_bufa[24]), 
        .A2(n22225), .B1(n19953), .B2(j202_soc_core_j22_cpu_ml_macl[24]), .Y(
        n19705) );
  sky130_fd_sc_hd__nand2_1 U23945 ( .A(n21920), .B(n19959), .Y(n19704) );
  sky130_fd_sc_hd__nand3_1 U23946 ( .A(n19706), .B(n19705), .C(n19704), .Y(
        n21940) );
  sky130_fd_sc_hd__a22oi_1 U23947 ( .A1(n19963), .A2(
        j202_soc_core_j22_cpu_ml_bufa[24]), .B1(n21940), .B2(
        j202_soc_core_j22_cpu_macop_MAC_[0]), .Y(n19707) );
  sky130_fd_sc_hd__nand2_1 U23948 ( .A(n19708), .B(n19707), .Y(n21105) );
  sky130_fd_sc_hd__nand2_1 U23949 ( .A(n21105), .B(n20019), .Y(n19720) );
  sky130_fd_sc_hd__a22oi_1 U23950 ( .A1(n20047), .A2(
        j202_soc_core_j22_cpu_rf_tmp[24]), .B1(n20048), .B2(
        j202_soc_core_j22_cpu_rf_gpr[504]), .Y(n19713) );
  sky130_fd_sc_hd__a22oi_1 U23951 ( .A1(n20056), .A2(
        j202_soc_core_j22_cpu_rf_pr[24]), .B1(j202_soc_core_j22_cpu_rf_gbr[24]), .B2(n20055), .Y(n19712) );
  sky130_fd_sc_hd__a2bb2oi_1 U23952 ( .B1(j202_soc_core_j22_cpu_pc[24]), .B2(
        n20046), .A1_N(n19709), .A2_N(n19908), .Y(n19711) );
  sky130_fd_sc_hd__nand2_1 U23953 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[24]), .Y(n19710) );
  sky130_fd_sc_hd__nand4_1 U23954 ( .A(n19713), .B(n19712), .C(n19711), .D(
        n19710), .Y(n19714) );
  sky130_fd_sc_hd__a21oi_1 U23955 ( .A1(n20053), .A2(n19715), .B1(n19714), .Y(
        n19716) );
  sky130_fd_sc_hd__o21a_1 U23956 ( .A1(n19717), .A2(n19764), .B1(n19716), .X(
        n19718) );
  sky130_fd_sc_hd__nand3_1 U23957 ( .A(n19720), .B(n19719), .C(n19718), .Y(
        n25354) );
  sky130_fd_sc_hd__nand2_1 U23958 ( .A(n19723), .B(n19722), .Y(n19728) );
  sky130_fd_sc_hd__xnor2_1 U23960 ( .A(n19728), .B(n19727), .Y(n21931) );
  sky130_fd_sc_hd__nand2_1 U23961 ( .A(n21931), .B(n19729), .Y(n19740) );
  sky130_fd_sc_hd__ha_1 U23962 ( .A(j202_soc_core_j22_cpu_pc[8]), .B(n19730), 
        .COUT(n18945), .SUM(n21926) );
  sky130_fd_sc_hd__a2bb2oi_1 U23963 ( .B1(n19732), .B2(n21926), .A1_N(n22558), 
        .A2_N(n19731), .Y(n19733) );
  sky130_fd_sc_hd__a21oi_1 U23965 ( .A1(n19736), .A2(n22171), .B1(n19735), .Y(
        n19739) );
  sky130_fd_sc_hd__nand2_1 U23966 ( .A(n25308), .B(n19737), .Y(n19738) );
  sky130_fd_sc_hd__nand3_1 U23967 ( .A(n19740), .B(n19739), .C(n19738), .Y(
        n25378) );
  sky130_fd_sc_hd__nor3_1 U23968 ( .A(n19742), .B(n19741), .C(n20495), .Y(
        n25404) );
  sky130_fd_sc_hd__nand2_1 U23969 ( .A(n19745), .B(n19744), .Y(n19746) );
  sky130_fd_sc_hd__xor2_1 U23970 ( .A(n19747), .B(n19746), .X(n19748) );
  sky130_fd_sc_hd__nand2_1 U23971 ( .A(n19748), .B(n20030), .Y(n19750) );
  sky130_fd_sc_hd__a22oi_1 U23972 ( .A1(j202_soc_core_j22_cpu_ml_mach[30]), 
        .A2(n20032), .B1(n21699), .B2(n20025), .Y(n19749) );
  sky130_fd_sc_hd__nand2_1 U23973 ( .A(n19750), .B(n19749), .Y(n21884) );
  sky130_fd_sc_hd__nand2_1 U23974 ( .A(n21884), .B(n22125), .Y(n19755) );
  sky130_fd_sc_hd__nand2_1 U23975 ( .A(n19751), .B(n20040), .Y(n19753) );
  sky130_fd_sc_hd__a22oi_1 U23976 ( .A1(j202_soc_core_j22_cpu_ml_macl[30]), 
        .A2(n19953), .B1(n21898), .B2(n19959), .Y(n19752) );
  sky130_fd_sc_hd__nand2_1 U23977 ( .A(n19753), .B(n19752), .Y(n21887) );
  sky130_fd_sc_hd__a22oi_1 U23978 ( .A1(j202_soc_core_j22_cpu_ml_bufa[30]), 
        .A2(n19931), .B1(n21887), .B2(j202_soc_core_j22_cpu_macop_MAC_[0]), 
        .Y(n19754) );
  sky130_fd_sc_hd__nand2_1 U23979 ( .A(n19755), .B(n19754), .Y(n21044) );
  sky130_fd_sc_hd__nand2_1 U23980 ( .A(n21044), .B(n20019), .Y(n19768) );
  sky130_fd_sc_hd__a22oi_1 U23981 ( .A1(n20047), .A2(
        j202_soc_core_j22_cpu_rf_tmp[30]), .B1(n20048), .B2(
        j202_soc_core_j22_cpu_rf_gpr[510]), .Y(n19760) );
  sky130_fd_sc_hd__a22oi_1 U23982 ( .A1(n20056), .A2(
        j202_soc_core_j22_cpu_rf_pr[30]), .B1(j202_soc_core_j22_cpu_rf_gbr[30]), .B2(n20055), .Y(n19759) );
  sky130_fd_sc_hd__a2bb2oi_1 U23983 ( .B1(j202_soc_core_j22_cpu_pc[30]), .B2(
        n20046), .A1_N(n19756), .A2_N(n19908), .Y(n19758) );
  sky130_fd_sc_hd__nand2_1 U23984 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[30]), .Y(n19757) );
  sky130_fd_sc_hd__nand4_1 U23985 ( .A(n19760), .B(n19759), .C(n19758), .D(
        n19757), .Y(n19761) );
  sky130_fd_sc_hd__a21oi_1 U23986 ( .A1(n20053), .A2(n19762), .B1(n19761), .Y(
        n19763) );
  sky130_fd_sc_hd__o21a_1 U23987 ( .A1(n19765), .A2(n19764), .B1(n19763), .X(
        n19766) );
  sky130_fd_sc_hd__nand3_1 U23988 ( .A(n19768), .B(n19767), .C(n19766), .Y(
        n25361) );
  sky130_fd_sc_hd__nand2_1 U23989 ( .A(n19771), .B(n19770), .Y(n19772) );
  sky130_fd_sc_hd__xor2_1 U23990 ( .A(n19773), .B(n19772), .X(n19774) );
  sky130_fd_sc_hd__nand2_1 U23991 ( .A(n19774), .B(n20030), .Y(n19776) );
  sky130_fd_sc_hd__a22oi_1 U23992 ( .A1(j202_soc_core_j22_cpu_ml_mach[28]), 
        .A2(n20032), .B1(n21700), .B2(n20025), .Y(n19775) );
  sky130_fd_sc_hd__nand2_1 U23993 ( .A(n19776), .B(n19775), .Y(n22086) );
  sky130_fd_sc_hd__nand2_1 U23994 ( .A(n22086), .B(n22125), .Y(n19781) );
  sky130_fd_sc_hd__nand2_1 U23995 ( .A(n19777), .B(n20040), .Y(n19779) );
  sky130_fd_sc_hd__a22oi_1 U23996 ( .A1(j202_soc_core_j22_cpu_ml_macl[28]), 
        .A2(n19953), .B1(n22096), .B2(n19959), .Y(n19778) );
  sky130_fd_sc_hd__nand2_1 U23997 ( .A(n19779), .B(n19778), .Y(n22089) );
  sky130_fd_sc_hd__a22oi_1 U23998 ( .A1(j202_soc_core_j22_cpu_ml_bufa[28]), 
        .A2(n19931), .B1(n22089), .B2(j202_soc_core_j22_cpu_macop_MAC_[0]), 
        .Y(n19780) );
  sky130_fd_sc_hd__nand2_1 U23999 ( .A(n19781), .B(n19780), .Y(n20378) );
  sky130_fd_sc_hd__nand2_1 U24000 ( .A(n20378), .B(n20019), .Y(n19795) );
  sky130_fd_sc_hd__nand2_1 U24001 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[28]), .Y(n19784) );
  sky130_fd_sc_hd__nand2_1 U24002 ( .A(n20056), .B(
        j202_soc_core_j22_cpu_rf_pr[28]), .Y(n19783) );
  sky130_fd_sc_hd__nand2_1 U24003 ( .A(n20055), .B(
        j202_soc_core_j22_cpu_rf_gbr[28]), .Y(n19782) );
  sky130_fd_sc_hd__nand3_1 U24004 ( .A(n19784), .B(n19783), .C(n19782), .Y(
        n19790) );
  sky130_fd_sc_hd__nand2_1 U24005 ( .A(n19785), .B(n20053), .Y(n19789) );
  sky130_fd_sc_hd__a2bb2oi_1 U24006 ( .B1(j202_soc_core_j22_cpu_pc[28]), .B2(
        n20046), .A1_N(n19786), .A2_N(n19908), .Y(n19788) );
  sky130_fd_sc_hd__a22oi_1 U24007 ( .A1(n20047), .A2(
        j202_soc_core_j22_cpu_rf_tmp[28]), .B1(n20048), .B2(
        j202_soc_core_j22_cpu_rf_gpr[508]), .Y(n19787) );
  sky130_fd_sc_hd__nand4b_1 U24008 ( .A_N(n19790), .B(n19789), .C(n19788), .D(
        n19787), .Y(n19791) );
  sky130_fd_sc_hd__a21oi_1 U24009 ( .A1(n19792), .A2(n21222), .B1(n19791), .Y(
        n19793) );
  sky130_fd_sc_hd__nand3_1 U24010 ( .A(n19795), .B(n19794), .C(n19793), .Y(
        n25358) );
  sky130_fd_sc_hd__nand2_1 U24011 ( .A(n25271), .B(n19798), .Y(n19834) );
  sky130_fd_sc_hd__nand3_1 U24012 ( .A(n21248), .B(n21245), .C(n19796), .Y(
        n19797) );
  sky130_fd_sc_hd__clkinv_1 U24013 ( .A(j202_soc_core_qspi_wb_wdat[31]), .Y(
        n24062) );
  sky130_fd_sc_hd__nor2_1 U24014 ( .A(j202_soc_core_rst), .B(n24062), .Y(
        n25389) );
  sky130_fd_sc_hd__clkinv_1 U24015 ( .A(j202_soc_core_qspi_wb_wdat[30]), .Y(
        n24053) );
  sky130_fd_sc_hd__nor2_1 U24016 ( .A(j202_soc_core_rst), .B(n24053), .Y(
        n25284) );
  sky130_fd_sc_hd__clkinv_1 U24017 ( .A(j202_soc_core_qspi_wb_wdat[29]), .Y(
        n24046) );
  sky130_fd_sc_hd__nor2_1 U24018 ( .A(j202_soc_core_rst), .B(n24046), .Y(
        n25296) );
  sky130_fd_sc_hd__nand2_1 U24019 ( .A(n25731), .B(
        j202_soc_core_qspi_wb_wdat[28]), .Y(n24399) );
  sky130_fd_sc_hd__clkinv_1 U24020 ( .A(j202_soc_core_qspi_wb_wdat[26]), .Y(
        n24026) );
  sky130_fd_sc_hd__nor2_1 U24021 ( .A(j202_soc_core_rst), .B(n24026), .Y(
        n25282) );
  sky130_fd_sc_hd__nand2_1 U24022 ( .A(n25734), .B(
        j202_soc_core_qspi_wb_wdat[24]), .Y(n24392) );
  sky130_fd_sc_hd__clkinv_1 U24023 ( .A(j202_soc_core_qspi_wb_wdat[23]), .Y(
        n24011) );
  sky130_fd_sc_hd__nor2_1 U24024 ( .A(j202_soc_core_rst), .B(n24011), .Y(
        n25292) );
  sky130_fd_sc_hd__clkinv_1 U24025 ( .A(j202_soc_core_qspi_wb_wdat[22]), .Y(
        n24000) );
  sky130_fd_sc_hd__nor2_1 U24026 ( .A(j202_soc_core_rst), .B(n24000), .Y(
        n25289) );
  sky130_fd_sc_hd__clkinv_1 U24027 ( .A(j202_soc_core_qspi_wb_wdat[21]), .Y(
        n23997) );
  sky130_fd_sc_hd__nor2_1 U24028 ( .A(j202_soc_core_rst), .B(n23997), .Y(
        n25283) );
  sky130_fd_sc_hd__nand2_1 U24029 ( .A(n25734), .B(
        j202_soc_core_qspi_wb_wdat[20]), .Y(n24443) );
  sky130_fd_sc_hd__clkinv_1 U24030 ( .A(j202_soc_core_qspi_wb_wdat[18]), .Y(
        n23974) );
  sky130_fd_sc_hd__nor2_1 U24031 ( .A(j202_soc_core_rst), .B(n23974), .Y(
        n25285) );
  sky130_fd_sc_hd__nand2_1 U24032 ( .A(n25734), .B(
        j202_soc_core_qspi_wb_wdat[16]), .Y(n24434) );
  sky130_fd_sc_hd__nand2_1 U24033 ( .A(n25734), .B(
        j202_soc_core_qspi_wb_wdat[12]), .Y(n24426) );
  sky130_fd_sc_hd__nand2_1 U24034 ( .A(n25734), .B(
        j202_soc_core_qspi_wb_wdat[8]), .Y(n24418) );
  sky130_fd_sc_hd__clkinv_1 U24035 ( .A(j202_soc_core_qspi_wb_wdat[7]), .Y(
        n23909) );
  sky130_fd_sc_hd__clkinv_1 U24036 ( .A(j202_soc_core_qspi_wb_wdat[6]), .Y(
        n23903) );
  sky130_fd_sc_hd__nor2_1 U24037 ( .A(j202_soc_core_rst), .B(n23903), .Y(
        n25298) );
  sky130_fd_sc_hd__clkinv_1 U24038 ( .A(j202_soc_core_qspi_wb_wdat[5]), .Y(
        n23897) );
  sky130_fd_sc_hd__nor2_1 U24039 ( .A(j202_soc_core_rst), .B(n23897), .Y(
        n25294) );
  sky130_fd_sc_hd__nand2_1 U24040 ( .A(n25734), .B(
        j202_soc_core_qspi_wb_wdat[4]), .Y(n24481) );
  sky130_fd_sc_hd__clkinv_1 U24041 ( .A(j202_soc_core_qspi_wb_wdat[2]), .Y(
        n23879) );
  sky130_fd_sc_hd__nor2_1 U24042 ( .A(j202_soc_core_rst), .B(n23879), .Y(
        n25286) );
  sky130_fd_sc_hd__nand2_1 U24043 ( .A(n25734), .B(
        j202_soc_core_qspi_wb_wdat[0]), .Y(n24473) );
  sky130_fd_sc_hd__nor2_1 U24044 ( .A(n19798), .B(n25271), .Y(n19801) );
  sky130_fd_sc_hd__nand3_1 U24045 ( .A(n21248), .B(n21245), .C(n19801), .Y(
        n19800) );
  sky130_fd_sc_hd__nand2_1 U24046 ( .A(n25271), .B(n25272), .Y(n20071) );
  sky130_fd_sc_hd__nor2_1 U24047 ( .A(n20071), .B(n19802), .Y(n25322) );
  sky130_fd_sc_hd__nor2_1 U24048 ( .A(n19835), .B(n19802), .Y(n25320) );
  sky130_fd_sc_hd__nor2_1 U24049 ( .A(n19834), .B(n19802), .Y(n25327) );
  sky130_fd_sc_hd__a22oi_1 U24050 ( .A1(j202_soc_core_j22_cpu_ml_mach[27]), 
        .A2(n20032), .B1(n21721), .B2(n20025), .Y(n19809) );
  sky130_fd_sc_hd__nand2_1 U24051 ( .A(n19804), .B(n19803), .Y(n19806) );
  sky130_fd_sc_hd__xnor2_1 U24052 ( .A(n19806), .B(n19805), .Y(n19807) );
  sky130_fd_sc_hd__nand2_1 U24053 ( .A(n19807), .B(n20030), .Y(n19808) );
  sky130_fd_sc_hd__nand2_1 U24054 ( .A(n19809), .B(n19808), .Y(n21943) );
  sky130_fd_sc_hd__nand2_1 U24055 ( .A(n21943), .B(n22125), .Y(n19817) );
  sky130_fd_sc_hd__nand2_1 U24056 ( .A(n19810), .B(n20040), .Y(n19814) );
  sky130_fd_sc_hd__o2bb2ai_1 U24057 ( .B1(n19811), .B2(n22246), .A1_N(
        j202_soc_core_j22_cpu_ml_macl[27]), .A2_N(n19953), .Y(n19812) );
  sky130_fd_sc_hd__a21oi_1 U24058 ( .A1(n21958), .A2(n19959), .B1(n19812), .Y(
        n19813) );
  sky130_fd_sc_hd__nand2_1 U24059 ( .A(n19814), .B(n19813), .Y(n21945) );
  sky130_fd_sc_hd__nand2_1 U24060 ( .A(n21945), .B(
        j202_soc_core_j22_cpu_macop_MAC_[0]), .Y(n19816) );
  sky130_fd_sc_hd__nand2_1 U24061 ( .A(n19963), .B(
        j202_soc_core_j22_cpu_ml_bufa[27]), .Y(n19815) );
  sky130_fd_sc_hd__nand3_1 U24062 ( .A(n19817), .B(n19816), .C(n19815), .Y(
        n20970) );
  sky130_fd_sc_hd__nand2_1 U24063 ( .A(n20970), .B(n20019), .Y(n19831) );
  sky130_fd_sc_hd__nand2_1 U24064 ( .A(n20045), .B(
        j202_soc_core_j22_cpu_rf_vbr[27]), .Y(n19821) );
  sky130_fd_sc_hd__nand2_1 U24065 ( .A(n20046), .B(
        j202_soc_core_j22_cpu_pc[27]), .Y(n19820) );
  sky130_fd_sc_hd__nand2_1 U24066 ( .A(n20047), .B(
        j202_soc_core_j22_cpu_rf_tmp[27]), .Y(n19819) );
  sky130_fd_sc_hd__nand2_1 U24067 ( .A(n20048), .B(
        j202_soc_core_j22_cpu_rf_gpr[507]), .Y(n19818) );
  sky130_fd_sc_hd__nand4_1 U24068 ( .A(n19821), .B(n19820), .C(n19819), .D(
        n19818), .Y(n19826) );
  sky130_fd_sc_hd__nand2_1 U24069 ( .A(n19822), .B(n20053), .Y(n19825) );
  sky130_fd_sc_hd__a22oi_1 U24070 ( .A1(n20056), .A2(
        j202_soc_core_j22_cpu_rf_pr[27]), .B1(j202_soc_core_j22_cpu_rf_gbr[27]), .B2(n20055), .Y(n19824) );
  sky130_fd_sc_hd__nand2_1 U24071 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[27]), .Y(n19823) );
  sky130_fd_sc_hd__nand4b_1 U24072 ( .A_N(n19826), .B(n19825), .C(n19824), .D(
        n19823), .Y(n19827) );
  sky130_fd_sc_hd__a21oi_1 U24073 ( .A1(n21222), .A2(n19828), .B1(n19827), .Y(
        n19829) );
  sky130_fd_sc_hd__nand3_1 U24074 ( .A(n19831), .B(n19830), .C(n19829), .Y(
        n25357) );
  sky130_fd_sc_hd__clkinv_1 U24075 ( .A(j202_soc_core_qspi_wb_wdat[27]), .Y(
        n24037) );
  sky130_fd_sc_hd__nor2_1 U24076 ( .A(j202_soc_core_rst), .B(n24037), .Y(
        n25291) );
  sky130_fd_sc_hd__nand3_1 U24077 ( .A(n19833), .B(n25273), .C(n25374), .Y(
        n20068) );
  sky130_fd_sc_hd__nor2_1 U24078 ( .A(n19834), .B(n20068), .Y(n25332) );
  sky130_fd_sc_hd__nor2_1 U24079 ( .A(n19835), .B(n20068), .Y(n25331) );
  sky130_fd_sc_hd__nor2_1 U24080 ( .A(n19836), .B(n20068), .Y(n25330) );
  sky130_fd_sc_hd__nor2_1 U24081 ( .A(n19834), .B(n20069), .Y(n25328) );
  sky130_fd_sc_hd__nor2_1 U24082 ( .A(n19835), .B(n20069), .Y(n25325) );
  sky130_fd_sc_hd__nand3_1 U24083 ( .A(n19833), .B(n19832), .C(n25273), .Y(
        n20070) );
  sky130_fd_sc_hd__nor2_1 U24084 ( .A(n19834), .B(n20070), .Y(n25323) );
  sky130_fd_sc_hd__nor2_1 U24085 ( .A(n19835), .B(n20070), .Y(n25317) );
  sky130_fd_sc_hd__nor2_1 U24086 ( .A(n19836), .B(n20070), .Y(n25318) );
  sky130_fd_sc_hd__o22ai_1 U24087 ( .A1(n21653), .A2(n19973), .B1(n19837), 
        .B2(n19971), .Y(n19840) );
  sky130_fd_sc_hd__o22ai_1 U24088 ( .A1(n21647), .A2(n19977), .B1(n19838), 
        .B2(n19975), .Y(n19839) );
  sky130_fd_sc_hd__nor2_1 U24089 ( .A(n19840), .B(n19839), .Y(n19847) );
  sky130_fd_sc_hd__a2bb2oi_1 U24090 ( .B1(j202_soc_core_j22_cpu_rf_vbr[1]), 
        .B2(n19985), .A1_N(n19841), .A2_N(n19986), .Y(n19846) );
  sky130_fd_sc_hd__nand2_1 U24091 ( .A(n19842), .B(
        j202_soc_core_j22_cpu_rf_gpr[1]), .Y(n19845) );
  sky130_fd_sc_hd__nand2_1 U24092 ( .A(n19843), .B(
        j202_soc_core_j22_cpu_rf_tmp[1]), .Y(n19844) );
  sky130_fd_sc_hd__nand4_1 U24093 ( .A(n19847), .B(n19846), .C(n19845), .D(
        n19844), .Y(n19848) );
  sky130_fd_sc_hd__a21oi_1 U24094 ( .A1(n19849), .A2(n19969), .B1(n19848), .Y(
        n19968) );
  sky130_fd_sc_hd__nand2_1 U24095 ( .A(n19852), .B(n19851), .Y(n19853) );
  sky130_fd_sc_hd__xor2_1 U24096 ( .A(n19854), .B(n19853), .X(n21697) );
  sky130_fd_sc_hd__nand2_1 U24097 ( .A(n21697), .B(n20030), .Y(n19863) );
  sky130_fd_sc_hd__nand2_1 U24098 ( .A(n19857), .B(n19856), .Y(n19858) );
  sky130_fd_sc_hd__xor2_1 U24099 ( .A(n19859), .B(n19858), .X(n19928) );
  sky130_fd_sc_hd__o22ai_1 U24100 ( .A1(n20007), .A2(n15666), .B1(n19860), 
        .B2(n20005), .Y(n19861) );
  sky130_fd_sc_hd__a21oi_1 U24101 ( .A1(n19928), .A2(n20025), .B1(n19861), .Y(
        n19862) );
  sky130_fd_sc_hd__nand2_1 U24102 ( .A(n19863), .B(n19862), .Y(n22212) );
  sky130_fd_sc_hd__nand2_1 U24103 ( .A(n22212), .B(n22125), .Y(n19872) );
  sky130_fd_sc_hd__nand2_1 U24104 ( .A(n19866), .B(n19865), .Y(n19868) );
  sky130_fd_sc_hd__xor2_1 U24105 ( .A(n19868), .B(n19867), .X(n22239) );
  sky130_fd_sc_hd__o22ai_1 U24106 ( .A1(n20014), .A2(n15666), .B1(n19869), 
        .B2(n20012), .Y(n19870) );
  sky130_fd_sc_hd__a21oi_1 U24107 ( .A1(n22239), .A2(n20016), .B1(n19870), .Y(
        n19871) );
  sky130_fd_sc_hd__nand2_1 U24108 ( .A(n19872), .B(n19871), .Y(n19873) );
  sky130_fd_sc_hd__nand2_1 U24109 ( .A(n19873), .B(n20019), .Y(n19906) );
  sky130_fd_sc_hd__nand2_1 U24110 ( .A(n19873), .B(n21137), .Y(n19904) );
  sky130_fd_sc_hd__nand2_1 U24111 ( .A(n22750), .B(n21178), .Y(n19888) );
  sky130_fd_sc_hd__a2bb2oi_1 U24112 ( .B1(n23301), .B2(n20716), .A1_N(n22314), 
        .A2_N(n20712), .Y(n19887) );
  sky130_fd_sc_hd__nand2_1 U24113 ( .A(n22754), .B(n20805), .Y(n19874) );
  sky130_fd_sc_hd__nand2_1 U24114 ( .A(n22183), .B(n22141), .Y(n22648) );
  sky130_fd_sc_hd__nand2_1 U24115 ( .A(n19874), .B(n22648), .Y(n22439) );
  sky130_fd_sc_hd__o22ai_1 U24116 ( .A1(n21108), .A2(n22439), .B1(n22487), 
        .B2(n21154), .Y(n19883) );
  sky130_fd_sc_hd__o22ai_1 U24117 ( .A1(n22146), .A2(n21155), .B1(n22565), 
        .B2(n19875), .Y(n19882) );
  sky130_fd_sc_hd__a2bb2oi_1 U24118 ( .B1(n21146), .B2(n22141), .A1_N(n21145), 
        .A2_N(n22183), .Y(n19876) );
  sky130_fd_sc_hd__o21ai_1 U24119 ( .A1(n21150), .A2(n22648), .B1(n19876), .Y(
        n19877) );
  sky130_fd_sc_hd__a21oi_1 U24120 ( .A1(n21156), .A2(n20699), .B1(n19877), .Y(
        n19878) );
  sky130_fd_sc_hd__o21ai_1 U24121 ( .A1(n19880), .A2(n19879), .B1(n19878), .Y(
        n19881) );
  sky130_fd_sc_hd__nor3_1 U24122 ( .A(n19883), .B(n19882), .C(n19881), .Y(
        n19886) );
  sky130_fd_sc_hd__nand2_1 U24123 ( .A(n19884), .B(n22183), .Y(n19885) );
  sky130_fd_sc_hd__nand4_1 U24124 ( .A(n19888), .B(n19887), .C(n19886), .D(
        n19885), .Y(n19898) );
  sky130_fd_sc_hd__o2bb2ai_1 U24125 ( .B1(n19891), .B2(n19890), .A1_N(n19889), 
        .A2_N(n25313), .Y(n19892) );
  sky130_fd_sc_hd__a21oi_1 U24126 ( .A1(n22521), .A2(n19893), .B1(n19892), .Y(
        n19894) );
  sky130_fd_sc_hd__nor2_1 U24127 ( .A(n21174), .B(n22662), .Y(n19897) );
  sky130_fd_sc_hd__nor3_1 U24128 ( .A(n20805), .B(n21091), .C(n22662), .Y(
        n19896) );
  sky130_fd_sc_hd__nor3_1 U24129 ( .A(n19898), .B(n19897), .C(n19896), .Y(
        n19903) );
  sky130_fd_sc_hd__nor2_1 U24130 ( .A(n20805), .B(n22662), .Y(n22494) );
  sky130_fd_sc_hd__o21ai_1 U24131 ( .A1(n22509), .A2(n22494), .B1(n20839), .Y(
        n19899) );
  sky130_fd_sc_hd__nand2_1 U24134 ( .A(n19901), .B(n21139), .Y(n19902) );
  sky130_fd_sc_hd__nand2_1 U24135 ( .A(n22122), .B(n19905), .Y(n19966) );
  sky130_fd_sc_hd__o211ai_1 U24136 ( .A1(n19907), .A2(n19968), .B1(n19906), 
        .C1(n19966), .Y(n25306) );
  sky130_fd_sc_hd__clkinv_1 U24137 ( .A(j202_soc_core_qspi_wb_wdat[1]), .Y(
        n23873) );
  sky130_fd_sc_hd__nor2_1 U24138 ( .A(j202_soc_core_rst), .B(n23873), .Y(
        n25288) );
  sky130_fd_sc_hd__a22oi_1 U24139 ( .A1(n20047), .A2(
        j202_soc_core_j22_cpu_rf_tmp[17]), .B1(n20048), .B2(
        j202_soc_core_j22_cpu_rf_gpr[497]), .Y(n19913) );
  sky130_fd_sc_hd__a22oi_1 U24140 ( .A1(n20056), .A2(
        j202_soc_core_j22_cpu_rf_pr[17]), .B1(j202_soc_core_j22_cpu_rf_gbr[17]), .B2(n20055), .Y(n19912) );
  sky130_fd_sc_hd__a2bb2oi_1 U24141 ( .B1(j202_soc_core_j22_cpu_pc[17]), .B2(
        n20046), .A1_N(n19909), .A2_N(n19908), .Y(n19911) );
  sky130_fd_sc_hd__nand2_1 U24142 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[17]), .Y(n19910) );
  sky130_fd_sc_hd__nand4_1 U24143 ( .A(n19913), .B(n19912), .C(n19911), .D(
        n19910), .Y(n19914) );
  sky130_fd_sc_hd__a21oi_1 U24144 ( .A1(n20053), .A2(n19915), .B1(n19914), .Y(
        n19916) );
  sky130_fd_sc_hd__o21a_1 U24145 ( .A1(n19968), .A2(n19917), .B1(n19916), .X(
        n19935) );
  sky130_fd_sc_hd__a21oi_1 U24146 ( .A1(n19920), .A2(n19919), .B1(n19918), .Y(
        n19924) );
  sky130_fd_sc_hd__nand2_1 U24147 ( .A(n19922), .B(n19921), .Y(n19923) );
  sky130_fd_sc_hd__xor2_1 U24148 ( .A(n19924), .B(n19923), .X(n19925) );
  sky130_fd_sc_hd__nand2_1 U24149 ( .A(n19925), .B(n20030), .Y(n19927) );
  sky130_fd_sc_hd__a22oi_1 U24150 ( .A1(j202_soc_core_j22_cpu_ml_mach[17]), 
        .A2(n20032), .B1(n21697), .B2(n20025), .Y(n19926) );
  sky130_fd_sc_hd__nand2_1 U24151 ( .A(n19927), .B(n19926), .Y(n21726) );
  sky130_fd_sc_hd__nand2_1 U24152 ( .A(n21726), .B(n22125), .Y(n19933) );
  sky130_fd_sc_hd__nand2_1 U24153 ( .A(n19928), .B(n20040), .Y(n19930) );
  sky130_fd_sc_hd__a22oi_1 U24154 ( .A1(j202_soc_core_j22_cpu_ml_macl[17]), 
        .A2(n19953), .B1(n22239), .B2(n19959), .Y(n19929) );
  sky130_fd_sc_hd__nand2_1 U24155 ( .A(n19930), .B(n19929), .Y(n21730) );
  sky130_fd_sc_hd__a22oi_1 U24156 ( .A1(j202_soc_core_j22_cpu_ml_bufa[17]), 
        .A2(n19931), .B1(n21730), .B2(j202_soc_core_j22_cpu_macop_MAC_[0]), 
        .Y(n19932) );
  sky130_fd_sc_hd__nand2_1 U24157 ( .A(n19933), .B(n19932), .Y(n20802) );
  sky130_fd_sc_hd__nand2_1 U24158 ( .A(n20802), .B(n20019), .Y(n19934) );
  sky130_fd_sc_hd__nand3_1 U24159 ( .A(n19966), .B(n19935), .C(n19934), .Y(
        n25347) );
  sky130_fd_sc_hd__clkinv_1 U24160 ( .A(j202_soc_core_qspi_wb_wdat[17]), .Y(
        n23968) );
  sky130_fd_sc_hd__nor2_1 U24161 ( .A(j202_soc_core_rst), .B(n23968), .Y(
        n25293) );
  sky130_fd_sc_hd__nand2_1 U24162 ( .A(n19937), .B(n19936), .Y(n19939) );
  sky130_fd_sc_hd__xnor2_1 U24163 ( .A(n19939), .B(n19938), .Y(n19940) );
  sky130_fd_sc_hd__nand2_1 U24164 ( .A(n19940), .B(n20030), .Y(n19948) );
  sky130_fd_sc_hd__nand2_1 U24165 ( .A(n19943), .B(n19942), .Y(n19944) );
  sky130_fd_sc_hd__xor2_1 U24166 ( .A(n19945), .B(n19944), .X(n21715) );
  sky130_fd_sc_hd__nand2_1 U24167 ( .A(n21715), .B(n20025), .Y(n19947) );
  sky130_fd_sc_hd__nand2b_1 U24168 ( .A_N(n20005), .B(
        j202_soc_core_j22_cpu_ml_mach[25]), .Y(n19946) );
  sky130_fd_sc_hd__nand3_1 U24169 ( .A(n19948), .B(n19947), .C(n19946), .Y(
        n21771) );
  sky130_fd_sc_hd__nand2_1 U24170 ( .A(n21771), .B(n22125), .Y(n19965) );
  sky130_fd_sc_hd__nand2_1 U24171 ( .A(n19950), .B(n19949), .Y(n19952) );
  sky130_fd_sc_hd__xnor2_1 U24172 ( .A(n19952), .B(n19951), .Y(n20009) );
  sky130_fd_sc_hd__nand2_1 U24173 ( .A(n20009), .B(n20040), .Y(n19962) );
  sky130_fd_sc_hd__a22oi_1 U24174 ( .A1(j202_soc_core_j22_cpu_ml_bufa[25]), 
        .A2(n22225), .B1(n19953), .B2(j202_soc_core_j22_cpu_ml_macl[25]), .Y(
        n19961) );
  sky130_fd_sc_hd__nand2_1 U24175 ( .A(n19956), .B(n19955), .Y(n19958) );
  sky130_fd_sc_hd__xor2_1 U24176 ( .A(n19958), .B(n19957), .X(n21815) );
  sky130_fd_sc_hd__nand2_1 U24177 ( .A(n21815), .B(n19959), .Y(n19960) );
  sky130_fd_sc_hd__nand3_1 U24178 ( .A(n19962), .B(n19961), .C(n19960), .Y(
        n21773) );
  sky130_fd_sc_hd__a22oi_1 U24179 ( .A1(n19963), .A2(
        j202_soc_core_j22_cpu_ml_bufa[25]), .B1(n21773), .B2(
        j202_soc_core_j22_cpu_macop_MAC_[0]), .Y(n19964) );
  sky130_fd_sc_hd__nand2_1 U24180 ( .A(n19965), .B(n19964), .Y(n21098) );
  sky130_fd_sc_hd__nand2_1 U24181 ( .A(n21098), .B(n20019), .Y(n20004) );
  sky130_fd_sc_hd__o21a_1 U24182 ( .A1(n19968), .A2(n19967), .B1(n19966), .X(
        n20023) );
  sky130_fd_sc_hd__nand2_1 U24183 ( .A(n19970), .B(n19969), .Y(n19992) );
  sky130_fd_sc_hd__o22ai_1 U24184 ( .A1(n19974), .A2(n19973), .B1(n19972), 
        .B2(n19971), .Y(n19980) );
  sky130_fd_sc_hd__o22ai_1 U24185 ( .A1(n19978), .A2(n19977), .B1(n19976), 
        .B2(n19975), .Y(n19979) );
  sky130_fd_sc_hd__nor2_1 U24186 ( .A(n19980), .B(n19979), .Y(n19991) );
  sky130_fd_sc_hd__o22ai_1 U24187 ( .A1(n19984), .A2(n19983), .B1(n19982), 
        .B2(n19981), .Y(n19989) );
  sky130_fd_sc_hd__o2bb2ai_1 U24188 ( .B1(n19987), .B2(n19986), .A1_N(
        j202_soc_core_j22_cpu_rf_vbr[9]), .A2_N(n19985), .Y(n19988) );
  sky130_fd_sc_hd__nor2_1 U24189 ( .A(n19989), .B(n19988), .Y(n19990) );
  sky130_fd_sc_hd__nand3_1 U24190 ( .A(n19992), .B(n19991), .C(n19990), .Y(
        n20021) );
  sky130_fd_sc_hd__nand2_1 U24191 ( .A(n20045), .B(
        j202_soc_core_j22_cpu_rf_vbr[25]), .Y(n19996) );
  sky130_fd_sc_hd__nand2_1 U24192 ( .A(n20046), .B(
        j202_soc_core_j22_cpu_pc[25]), .Y(n19995) );
  sky130_fd_sc_hd__nand2_1 U24193 ( .A(n20047), .B(
        j202_soc_core_j22_cpu_rf_tmp[25]), .Y(n19994) );
  sky130_fd_sc_hd__nand2_1 U24194 ( .A(n20048), .B(
        j202_soc_core_j22_cpu_rf_gpr[505]), .Y(n19993) );
  sky130_fd_sc_hd__nand4_1 U24195 ( .A(n19996), .B(n19995), .C(n19994), .D(
        n19993), .Y(n20001) );
  sky130_fd_sc_hd__nand2_1 U24196 ( .A(n19997), .B(n20053), .Y(n20000) );
  sky130_fd_sc_hd__a22oi_1 U24197 ( .A1(n20056), .A2(
        j202_soc_core_j22_cpu_rf_pr[25]), .B1(j202_soc_core_j22_cpu_rf_gbr[25]), .B2(n20055), .Y(n19999) );
  sky130_fd_sc_hd__nand2_1 U24198 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[25]), .Y(n19998) );
  sky130_fd_sc_hd__nand4b_1 U24199 ( .A_N(n20001), .B(n20000), .C(n19999), .D(
        n19998), .Y(n20002) );
  sky130_fd_sc_hd__a21oi_1 U24200 ( .A1(n21222), .A2(n20021), .B1(n20002), .Y(
        n20003) );
  sky130_fd_sc_hd__nand3_1 U24201 ( .A(n20004), .B(n20023), .C(n20003), .Y(
        n25355) );
  sky130_fd_sc_hd__clkinv_1 U24202 ( .A(j202_soc_core_qspi_wb_wdat[25]), .Y(
        n24019) );
  sky130_fd_sc_hd__nor2_1 U24203 ( .A(j202_soc_core_rst), .B(n24019), .Y(
        n25290) );
  sky130_fd_sc_hd__nand2_1 U24204 ( .A(n21715), .B(n20030), .Y(n20011) );
  sky130_fd_sc_hd__o22ai_1 U24205 ( .A1(n20007), .A2(n21817), .B1(n20006), 
        .B2(n20005), .Y(n20008) );
  sky130_fd_sc_hd__a21oi_1 U24206 ( .A1(n20009), .A2(n20025), .B1(n20008), .Y(
        n20010) );
  sky130_fd_sc_hd__nand2_1 U24207 ( .A(n20011), .B(n20010), .Y(n21813) );
  sky130_fd_sc_hd__nand2_1 U24208 ( .A(n21813), .B(n22125), .Y(n20018) );
  sky130_fd_sc_hd__o22ai_1 U24209 ( .A1(n20014), .A2(n21817), .B1(n20013), 
        .B2(n20012), .Y(n20015) );
  sky130_fd_sc_hd__a21oi_1 U24210 ( .A1(n21815), .A2(n20016), .B1(n20015), .Y(
        n20017) );
  sky130_fd_sc_hd__nand2_1 U24211 ( .A(n20018), .B(n20017), .Y(n20704) );
  sky130_fd_sc_hd__nand2_1 U24212 ( .A(n20704), .B(n20019), .Y(n20024) );
  sky130_fd_sc_hd__nand2_1 U24213 ( .A(n20021), .B(n20020), .Y(n20022) );
  sky130_fd_sc_hd__nand3_1 U24214 ( .A(n20024), .B(n20023), .C(n20022), .Y(
        n25368) );
  sky130_fd_sc_hd__nand2_1 U24215 ( .A(n25734), .B(
        j202_soc_core_qspi_wb_wdat[9]), .Y(n24420) );
  sky130_fd_sc_hd__clkinv_1 U24216 ( .A(j202_soc_core_qspi_wb_wdat[3]), .Y(
        n23885) );
  sky130_fd_sc_hd__nor2_1 U24217 ( .A(j202_soc_core_rst), .B(n23885), .Y(
        n25287) );
  sky130_fd_sc_hd__nand2_1 U24218 ( .A(n21698), .B(n20025), .Y(n20034) );
  sky130_fd_sc_hd__nand2_1 U24219 ( .A(n20027), .B(n20026), .Y(n20029) );
  sky130_fd_sc_hd__xnor2_1 U24220 ( .A(n20029), .B(n20028), .Y(n20031) );
  sky130_fd_sc_hd__a22oi_1 U24221 ( .A1(j202_soc_core_j22_cpu_ml_mach[19]), 
        .A2(n20032), .B1(n20031), .B2(n20030), .Y(n20033) );
  sky130_fd_sc_hd__nand2_1 U24222 ( .A(n20034), .B(n20033), .Y(n21965) );
  sky130_fd_sc_hd__o22ai_1 U24223 ( .A1(n20038), .A2(n20037), .B1(n20036), 
        .B2(n20035), .Y(n20039) );
  sky130_fd_sc_hd__a21oi_1 U24224 ( .A1(n20041), .A2(n20040), .B1(n20039), .Y(
        n21968) );
  sky130_fd_sc_hd__o22ai_1 U24225 ( .A1(n20043), .A2(n20042), .B1(n22125), 
        .B2(n21968), .Y(n20044) );
  sky130_fd_sc_hd__a21oi_1 U24226 ( .A1(n21965), .A2(n22125), .B1(n20044), .Y(
        n20780) );
  sky130_fd_sc_hd__nand2_1 U24227 ( .A(n20045), .B(
        j202_soc_core_j22_cpu_rf_vbr[19]), .Y(n20052) );
  sky130_fd_sc_hd__nand2_1 U24228 ( .A(n20046), .B(
        j202_soc_core_j22_cpu_pc[19]), .Y(n20051) );
  sky130_fd_sc_hd__nand2_1 U24229 ( .A(n20047), .B(
        j202_soc_core_j22_cpu_rf_tmp[19]), .Y(n20050) );
  sky130_fd_sc_hd__nand2_1 U24230 ( .A(n20048), .B(
        j202_soc_core_j22_cpu_rf_gpr[499]), .Y(n20049) );
  sky130_fd_sc_hd__nand4_1 U24231 ( .A(n20052), .B(n20051), .C(n20050), .D(
        n20049), .Y(n20061) );
  sky130_fd_sc_hd__nand2_1 U24232 ( .A(n20054), .B(n20053), .Y(n20060) );
  sky130_fd_sc_hd__a22oi_1 U24233 ( .A1(n20056), .A2(
        j202_soc_core_j22_cpu_rf_pr[19]), .B1(j202_soc_core_j22_cpu_rf_gbr[19]), .B2(n20055), .Y(n20059) );
  sky130_fd_sc_hd__nand2_1 U24234 ( .A(n20057), .B(
        j202_soc_core_j22_cpu_rf_gpr[19]), .Y(n20058) );
  sky130_fd_sc_hd__nand4b_1 U24235 ( .A_N(n20061), .B(n20060), .C(n20059), .D(
        n20058), .Y(n20062) );
  sky130_fd_sc_hd__a21oi_1 U24236 ( .A1(n20064), .A2(n20063), .B1(n20062), .Y(
        n20066) );
  sky130_fd_sc_hd__o211ai_1 U24237 ( .A1(n20780), .A2(n20067), .B1(n20066), 
        .C1(n20065), .Y(n25349) );
  sky130_fd_sc_hd__clkinv_1 U24238 ( .A(j202_soc_core_qspi_wb_wdat[19]), .Y(
        n23981) );
  sky130_fd_sc_hd__nor2_1 U24239 ( .A(j202_soc_core_rst), .B(n23981), .Y(
        n25295) );
  sky130_fd_sc_hd__nand2_1 U24240 ( .A(n25734), .B(
        j202_soc_core_qspi_wb_wdat[13]), .Y(n24428) );
  sky130_fd_sc_hd__nor2_1 U24241 ( .A(j202_soc_core_uart_BRG_cnt[0]), .B(
        j202_soc_core_uart_BRG_cnt[1]), .Y(n25399) );
  sky130_fd_sc_hd__nand2_1 U24242 ( .A(j202_soc_core_uart_sio_ce), .B(
        j202_soc_core_uart_TOP_shift_en), .Y(n21325) );
  sky130_fd_sc_hd__nor2_1 U24243 ( .A(j202_soc_core_rst), .B(n21325), .Y(
        n25401) );
  sky130_fd_sc_hd__nand2_1 U24244 ( .A(n25734), .B(
        j202_soc_core_qspi_wb_wdat[14]), .Y(n24430) );
  sky130_fd_sc_hd__nand2_1 U24245 ( .A(n25734), .B(
        j202_soc_core_qspi_wb_wdat[11]), .Y(n24424) );
  sky130_fd_sc_hd__nor2_1 U24246 ( .A(n20071), .B(n20068), .Y(n25329) );
  sky130_fd_sc_hd__nor2_1 U24247 ( .A(n20071), .B(n20069), .Y(n25326) );
  sky130_fd_sc_hd__nor2_1 U24248 ( .A(n20071), .B(n20070), .Y(n25319) );
  sky130_fd_sc_hd__nand2_1 U24249 ( .A(j202_soc_core_bldc_core_00_comm[2]), 
        .B(j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld), .Y(n23805) );
  sky130_fd_sc_hd__nor2_1 U24250 ( .A(j202_soc_core_bldc_core_00_comm[1]), .B(
        n23805), .Y(n25397) );
  sky130_fd_sc_hd__clkinv_1 U24251 ( .A(j202_soc_core_bldc_core_00_comm[1]), 
        .Y(n25161) );
  sky130_fd_sc_hd__nand2b_1 U24252 ( .A_N(j202_soc_core_bldc_core_00_comm[2]), 
        .B(j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld), .Y(n23807) );
  sky130_fd_sc_hd__nor2_1 U24253 ( .A(n25161), .B(n23807), .Y(n25398) );
  sky130_fd_sc_hd__clkbuf_1 U24254 ( .A(la_data_out[17]), .X(io_out[37]) );
  sky130_fd_sc_hd__and3_1 U24255 ( .A(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[0]), .C(n20102), .X(io_oeb[12]) );
  sky130_fd_sc_hd__clkbuf_1 U24256 ( .A(la_data_out[16]), .X(io_out[36]) );
  sky130_fd_sc_hd__clkbuf_1 U24257 ( .A(io_oeb[12]), .X(io_oeb[10]) );
  sky130_fd_sc_hd__clkbuf_1 U24258 ( .A(la_data_out[15]), .X(io_out[35]) );
  sky130_fd_sc_hd__clkbuf_1 U24259 ( .A(la_data_out[14]), .X(io_out[34]) );
  sky130_fd_sc_hd__clkbuf_1 U24260 ( .A(la_data_out[13]), .X(io_out[33]) );
  sky130_fd_sc_hd__clkbuf_1 U24261 ( .A(la_data_out[0]), .X(io_out[0]) );
  sky130_fd_sc_hd__clkbuf_1 U24262 ( .A(la_data_out[12]), .X(io_out[32]) );
  sky130_fd_sc_hd__clkbuf_1 U24263 ( .A(la_data_out[11]), .X(io_out[31]) );
  sky130_fd_sc_hd__clkbuf_1 U24264 ( .A(la_data_out[9]), .X(io_out[29]) );
  sky130_fd_sc_hd__clkbuf_1 U24265 ( .A(la_data_out[2]), .X(io_out[2]) );
  sky130_fd_sc_hd__clkbuf_1 U24266 ( .A(la_data_out[8]), .X(io_out[28]) );
  sky130_fd_sc_hd__clkbuf_1 U24267 ( .A(la_data_out[7]), .X(io_out[27]) );
  sky130_fd_sc_hd__clkbuf_1 U24268 ( .A(la_data_out[3]), .X(io_out[3]) );
  sky130_fd_sc_hd__clkbuf_1 U24269 ( .A(la_data_out[6]), .X(io_out[26]) );
  sky130_fd_sc_hd__clkbuf_1 U24270 ( .A(la_data_out[5]), .X(io_out[7]) );
  sky130_fd_sc_hd__clkbuf_1 U24271 ( .A(la_data_out[4]), .X(io_out[4]) );
  sky130_fd_sc_hd__nand2_1 U24272 ( .A(j202_soc_core_uart_TOP_rx_go), .B(
        j202_soc_core_uart_TOP_rx_sio_ce), .Y(n23821) );
  sky130_fd_sc_hd__clkinv_1 U24273 ( .A(n23821), .Y(j202_soc_core_uart_TOP_N95) );
  sky130_fd_sc_hd__clkinv_1 U24274 ( .A(j202_soc_core_uart_TOP_rx_fifo_gb), 
        .Y(n20074) );
  sky130_fd_sc_hd__nor2_1 U24276 ( .A(j202_soc_core_uart_TOP_rx_valid_r), .B(
        n20075), .Y(n25235) );
  sky130_fd_sc_hd__nand2_1 U24277 ( .A(j202_soc_core_uart_TOP_rx_fifo_wp[0]), 
        .B(n25235), .Y(n25231) );
  sky130_fd_sc_hd__nand2_1 U24278 ( .A(n22104), .B(j202_soc_core_aquc_SEL__0_), 
        .Y(n23254) );
  sky130_fd_sc_hd__nand3_1 U24279 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[0]), 
        .B(j202_soc_core_uart_WRTXD1), .C(n23254), .Y(n25200) );
  sky130_fd_sc_hd__nor2_1 U24280 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[1]), 
        .B(n25200), .Y(j202_soc_core_uart_TOP_tx_fifo_N31) );
  sky130_fd_sc_hd__nand2b_1 U24281 ( .A_N(n25403), .B(n25734), .Y(
        j202_soc_core_ahb2apb_00_N127) );
  sky130_fd_sc_hd__nor2_1 U24282 ( .A(j202_soc_core_rst), .B(
        j202_soc_core_qspi_wb_wdat[12]), .Y(n23940) );
  sky130_fd_sc_hd__and3_1 U24283 ( .A(n21224), .B(n20076), .C(
        j202_soc_core_ahb2apb_01_state[1]), .X(n20093) );
  sky130_fd_sc_hd__nor2_1 U24284 ( .A(j202_soc_core_intc_core_00_bs_addr[10]), 
        .B(j202_soc_core_intc_core_00_bs_addr[11]), .Y(n20079) );
  sky130_fd_sc_hd__nand4_1 U24285 ( .A(j202_soc_core_pstrb[5]), .B(
        j202_soc_core_pstrb[4]), .C(j202_soc_core_pstrb[6]), .D(
        j202_soc_core_pstrb[7]), .Y(n20077) );
  sky130_fd_sc_hd__nand2_1 U24286 ( .A(j202_soc_core_pwrite[1]), .B(n20077), 
        .Y(n20078) );
  sky130_fd_sc_hd__nand3_1 U24287 ( .A(n20093), .B(n20079), .C(n20078), .Y(
        n24451) );
  sky130_fd_sc_hd__nor2_1 U24288 ( .A(j202_soc_core_intc_core_00_bs_addr[5]), 
        .B(n24451), .Y(n24461) );
  sky130_fd_sc_hd__clkinv_1 U24289 ( .A(j202_soc_core_intc_core_00_bs_addr[4]), 
        .Y(n24467) );
  sky130_fd_sc_hd__nand2_1 U24290 ( .A(n24467), .B(
        j202_soc_core_intc_core_00_bs_addr[9]), .Y(n20080) );
  sky130_fd_sc_hd__nand2_1 U24291 ( .A(n24468), .B(n24573), .Y(n20095) );
  sky130_fd_sc_hd__nor2_1 U24292 ( .A(n20080), .B(n20095), .Y(n20081) );
  sky130_fd_sc_hd__nand3_1 U24293 ( .A(n24461), .B(n24471), .C(n20081), .Y(
        n24292) );
  sky130_fd_sc_hd__nor2_1 U24294 ( .A(j202_soc_core_intc_core_00_bs_addr[3]), 
        .B(j202_soc_core_intc_core_00_bs_addr[2]), .Y(n24469) );
  sky130_fd_sc_hd__nand3_1 U24295 ( .A(n20083), .B(
        j202_soc_core_intc_core_00_bs_addr[8]), .C(n24469), .Y(n24548) );
  sky130_fd_sc_hd__nand2_1 U24296 ( .A(n20082), .B(j202_soc_core_pwrite[1]), 
        .Y(n24290) );
  sky130_fd_sc_hd__nand2_1 U24297 ( .A(n25734), .B(n24290), .Y(n24291) );
  sky130_fd_sc_hd__o2bb2ai_1 U24298 ( .B1(n23940), .B2(n20115), .A1_N(n24290), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[3]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__nor2_1 U24299 ( .A(j202_soc_core_rst), .B(
        j202_soc_core_qspi_wb_wdat[8]), .Y(n23918) );
  sky130_fd_sc_hd__nor2_1 U24300 ( .A(j202_soc_core_rst), .B(
        j202_soc_core_qspi_wb_wdat[20]), .Y(n23990) );
  sky130_fd_sc_hd__o2bb2ai_1 U24301 ( .B1(n23990), .B2(n20115), .A1_N(n24290), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[5]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__nor2_1 U24302 ( .A(j202_soc_core_rst), .B(
        j202_soc_core_qspi_wb_wdat[28]), .Y(n24043) );
  sky130_fd_sc_hd__o2bb2ai_1 U24303 ( .B1(n24043), .B2(n20115), .A1_N(n24290), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[7]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__nor2_1 U24304 ( .A(j202_soc_core_rst), .B(
        j202_soc_core_qspi_wb_wdat[24]), .Y(n24015) );
  sky130_fd_sc_hd__o2bb2ai_1 U24305 ( .B1(n24015), .B2(n20115), .A1_N(n24290), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[6]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__nor2_1 U24306 ( .A(j202_soc_core_rst), .B(
        j202_soc_core_qspi_wb_wdat[4]), .Y(n23893) );
  sky130_fd_sc_hd__o2bb2ai_1 U24307 ( .B1(n23893), .B2(n20115), .A1_N(n24290), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[1]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__nor2_1 U24308 ( .A(j202_soc_core_rst), .B(
        j202_soc_core_qspi_wb_wdat[0]), .Y(n23868) );
  sky130_fd_sc_hd__o2bb2ai_1 U24309 ( .B1(n23868), .B2(n20115), .A1_N(n24290), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[0]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__nor2_1 U24310 ( .A(j202_soc_core_rst), .B(
        j202_soc_core_qspi_wb_wdat[16]), .Y(n23965) );
  sky130_fd_sc_hd__o2bb2ai_1 U24311 ( .B1(n23965), .B2(n20115), .A1_N(n24290), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[4]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o2bb2ai_1 U24312 ( .B1(n24422), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[66]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o2bb2ai_1 U24313 ( .B1(n24430), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[67]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__clkinv_1 U24314 ( .A(n25389), .Y(n24405) );
  sky130_fd_sc_hd__o2bb2ai_1 U24315 ( .B1(n24405), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[103]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o2bb2ai_1 U24316 ( .B1(n24420), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[34]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o2bb2ai_1 U24317 ( .B1(n24428), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[35]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o2bb2ai_1 U24318 ( .B1(n24432), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[99]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o2bb2ai_1 U24319 ( .B1(n24395), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[70]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o2bb2ai_1 U24320 ( .B1(n24387), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[37]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o2bb2ai_1 U24321 ( .B1(n24402), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[71]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o2bb2ai_1 U24322 ( .B1(n24438), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[68]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o2bb2ai_1 U24323 ( .B1(n24477), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[64]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o2bb2ai_1 U24324 ( .B1(n24479), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[96]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__nor2_1 U24325 ( .A(j202_soc_core_wbqspiflash_00_state[2]), 
        .B(n25070), .Y(n23542) );
  sky130_fd_sc_hd__nand2_1 U24326 ( .A(j202_soc_core_wbqspiflash_00_state[4]), 
        .B(n23542), .Y(n23356) );
  sky130_fd_sc_hd__nor2_1 U24327 ( .A(n23395), .B(n22847), .Y(n23535) );
  sky130_fd_sc_hd__nor2_1 U24328 ( .A(n23356), .B(n23433), .Y(n25044) );
  sky130_fd_sc_hd__nor2_1 U24329 ( .A(j202_soc_core_rst), .B(n25044), .Y(
        n23585) );
  sky130_fd_sc_hd__o2bb2ai_1 U24330 ( .B1(n24393), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[38]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o2bb2ai_1 U24331 ( .B1(n24397), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[102]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o2bb2ai_1 U24332 ( .B1(n24390), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[101]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__nor2_1 U24333 ( .A(j202_soc_core_intc_core_00_bs_addr[2]), 
        .B(n24453), .Y(n24452) );
  sky130_fd_sc_hd__nand3_1 U24334 ( .A(n20083), .B(
        j202_soc_core_intc_core_00_bs_addr[8]), .C(n24452), .Y(n24498) );
  sky130_fd_sc_hd__nand2_1 U24335 ( .A(n20084), .B(j202_soc_core_pwrite[1]), 
        .Y(n20475) );
  sky130_fd_sc_hd__o2bb2ai_1 U24336 ( .B1(n23918), .B2(n20473), .A1_N(n20475), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[18]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o2bb2ai_1 U24337 ( .B1(n23868), .B2(n20473), .A1_N(n20475), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[16]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__nand2_1 U24338 ( .A(n20087), .B(n20086), .Y(n20088) );
  sky130_fd_sc_hd__nand2_1 U24339 ( .A(n20089), .B(n21664), .Y(n22187) );
  sky130_fd_sc_hd__nand2_1 U24340 ( .A(n23345), .B(n22153), .Y(n22149) );
  sky130_fd_sc_hd__o31ai_1 U24341 ( .A1(j202_soc_core_j22_cpu_macop_MAC_[4]), 
        .A2(n20101), .A3(n21669), .B1(n22186), .Y(n20090) );
  sky130_fd_sc_hd__nand2_1 U24342 ( .A(j202_soc_core_intc_core_00_bs_addr[2]), 
        .B(j202_soc_core_intc_core_00_bs_addr[8]), .Y(n20091) );
  sky130_fd_sc_hd__nand2_1 U24343 ( .A(n24579), .B(
        j202_soc_core_intc_core_00_bs_addr[3]), .Y(n24492) );
  sky130_fd_sc_hd__nand2_1 U24344 ( .A(n20092), .B(j202_soc_core_pwrite[1]), 
        .Y(n20477) );
  sky130_fd_sc_hd__o2bb2ai_1 U24345 ( .B1(n20474), .B2(n23918), .A1_N(n20477), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[26]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o2bb2ai_1 U24346 ( .B1(n20474), .B2(n23940), .A1_N(n20477), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[27]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o2bb2ai_1 U24347 ( .B1(n23868), .B2(n20474), .A1_N(n20477), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[24]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o2bb2ai_1 U24348 ( .B1(n24422), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[82]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o2bb2ai_1 U24349 ( .B1(n24475), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[48]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o2bb2ai_1 U24350 ( .B1(n24479), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[112]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o2bb2ai_1 U24351 ( .B1(n24428), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[51]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o2bb2ai_1 U24352 ( .B1(n24477), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[80]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o2bb2ai_1 U24353 ( .B1(n24483), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[49]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__nand2b_1 U24354 ( .A_N(n20093), .B(n25734), .Y(n25531) );
  sky130_fd_sc_hd__o2bb2ai_1 U24355 ( .B1(n20477), .B2(n24483), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[57]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o2bb2ai_1 U24356 ( .B1(n20477), .B2(n24420), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[58]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o2bb2ai_1 U24357 ( .B1(n20477), .B2(n24422), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[90]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o2bb2ai_1 U24358 ( .B1(n20477), .B2(n24432), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[123]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o2bb2ai_1 U24359 ( .B1(n20477), .B2(n24428), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[59]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o2bb2ai_1 U24360 ( .B1(n20477), .B2(n24479), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[120]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__nor3_1 U24361 ( .A(j202_soc_core_intc_core_00_bs_addr[4]), 
        .B(j202_soc_core_intc_core_00_bs_addr[9]), .C(n24448), .Y(n20094) );
  sky130_fd_sc_hd__nand4_1 U24362 ( .A(n24461), .B(n24471), .C(n20094), .D(
        n24469), .Y(n24495) );
  sky130_fd_sc_hd__nand2_1 U24363 ( .A(n20096), .B(j202_soc_core_pwrite[1]), 
        .Y(n24442) );
  sky130_fd_sc_hd__nand2_1 U24364 ( .A(n25734), .B(n24442), .Y(n24444) );
  sky130_fd_sc_hd__o2bb2ai_1 U24365 ( .B1(n24397), .B2(n24442), .A1_N(
        j202_soc_core_intc_core_00_rg_ie[27]), .A2_N(n20114), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o2bb2ai_1 U24366 ( .B1(n24389), .B2(n24442), .A1_N(
        j202_soc_core_intc_core_00_rg_ie[22]), .A2_N(n20114), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o2bb2ai_1 U24367 ( .B1(n24399), .B2(n24442), .A1_N(
        j202_soc_core_intc_core_00_rg_ie[28]), .A2_N(n20114), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o2bb2ai_1 U24368 ( .B1(n24402), .B2(n24442), .A1_N(
        j202_soc_core_intc_core_00_rg_ie[30]), .A2_N(n20114), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o2bb2ai_1 U24369 ( .B1(n24390), .B2(n24442), .A1_N(
        j202_soc_core_intc_core_00_rg_ie[23]), .A2_N(n20114), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o2bb2ai_1 U24370 ( .B1(n24395), .B2(n24442), .A1_N(
        j202_soc_core_intc_core_00_rg_ie[26]), .A2_N(n20114), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o2bb2ai_1 U24371 ( .B1(n24392), .B2(n24442), .A1_N(
        j202_soc_core_intc_core_00_rg_ie[24]), .A2_N(n20114), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o2bb2ai_1 U24372 ( .B1(n24387), .B2(n24442), .A1_N(
        j202_soc_core_intc_core_00_rg_ie[21]), .A2_N(n20114), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o2bb2ai_1 U24373 ( .B1(n23965), .B2(n20473), .A1_N(n20475), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[20]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o2bb2ai_1 U24374 ( .B1(n20474), .B2(n23965), .A1_N(n20477), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[28]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o2bb2ai_1 U24375 ( .B1(n20477), .B2(n24430), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[91]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o2bb2ai_1 U24376 ( .B1(n20477), .B2(n24393), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[62]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o2bb2ai_1 U24377 ( .B1(n20477), .B2(n24387), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[61]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o2bb2ai_1 U24378 ( .B1(n20477), .B2(n24395), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[94]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o2bb2ai_1 U24379 ( .B1(n20477), .B2(n24436), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[60]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o2bb2ai_1 U24380 ( .B1(n20477), .B2(n24389), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[93]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o2bb2ai_1 U24381 ( .B1(n20477), .B2(n24402), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[95]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o2bb2ai_1 U24382 ( .B1(n20477), .B2(n24438), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[92]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o2bb2ai_1 U24383 ( .B1(n20477), .B2(n24390), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[125]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__nand2_1 U24384 ( .A(n20098), .B(n20097), .Y(n22135) );
  sky130_fd_sc_hd__nor3_1 U24385 ( .A(n20099), .B(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .C(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]), .Y(n21681) );
  sky130_fd_sc_hd__o31ai_1 U24386 ( .A1(n21675), .A2(
        j202_soc_core_j22_cpu_macop_MAC_[4]), .A3(n20101), .B1(n22143), .Y(
        j202_soc_core_j22_cpu_ml_N323) );
  sky130_fd_sc_hd__o2bb2ai_1 U24387 ( .B1(n24395), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[86]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o2bb2ai_1 U24388 ( .B1(n24389), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[85]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o2bb2ai_1 U24389 ( .B1(n24436), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[52]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o2bb2ai_1 U24390 ( .B1(n24430), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[83]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o2bb2ai_1 U24391 ( .B1(n24402), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[87]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o2bb2ai_1 U24392 ( .B1(n24387), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[53]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o2bb2ai_1 U24393 ( .B1(n24397), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[118]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o2bb2ai_1 U24394 ( .B1(n24438), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[84]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o2bb2ai_1 U24395 ( .B1(n24390), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[117]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o2bb2ai_1 U24396 ( .B1(n20477), .B2(n24440), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[124]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o2bb2ai_1 U24397 ( .B1(n24440), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[100]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__clkinv_1 U24398 ( .A(gpio_en_o[0]), .Y(io_oeb[0]) );
  sky130_fd_sc_hd__clkinv_1 U24399 ( .A(gpio_en_o[4]), .Y(io_oeb[4]) );
  sky130_fd_sc_hd__clkinv_1 U24400 ( .A(gpio_en_o[16]), .Y(io_oeb[36]) );
  sky130_fd_sc_hd__clkinv_1 U24401 ( .A(gpio_en_o[8]), .Y(io_oeb[28]) );
  sky130_fd_sc_hd__a22oi_1 U24402 ( .A1(
        j202_soc_core_wbqspiflash_00_spif_override), .A2(
        j202_soc_core_wbqspiflash_00_alt_cmd), .B1(n20102), .B2(
        j202_soc_core_wbqspiflash_00_w_qspi_cs_n), .Y(n23534) );
  sky130_fd_sc_hd__nor2_1 U24403 ( .A(j202_soc_core_wbqspiflash_00_state[4]), 
        .B(n24899), .Y(n23526) );
  sky130_fd_sc_hd__nand2_1 U24404 ( .A(n22847), .B(
        j202_soc_core_wbqspiflash_00_state[3]), .Y(n23435) );
  sky130_fd_sc_hd__nor2_1 U24405 ( .A(n23435), .B(n25070), .Y(n23450) );
  sky130_fd_sc_hd__nor2_1 U24406 ( .A(n23526), .B(n23366), .Y(n23455) );
  sky130_fd_sc_hd__nand2_1 U24407 ( .A(n25070), .B(n24899), .Y(n23398) );
  sky130_fd_sc_hd__nand3_1 U24408 ( .A(j202_soc_core_wbqspiflash_00_state[3]), 
        .B(n25001), .C(n22847), .Y(n25011) );
  sky130_fd_sc_hd__nand2_1 U24409 ( .A(j202_soc_core_wbqspiflash_00_state[3]), 
        .B(n23542), .Y(n22852) );
  sky130_fd_sc_hd__nand2_1 U24410 ( .A(n25011), .B(n22852), .Y(n23578) );
  sky130_fd_sc_hd__nor2_1 U24411 ( .A(n23455), .B(n23578), .Y(n23483) );
  sky130_fd_sc_hd__nor2_1 U24412 ( .A(j202_soc_core_wbqspiflash_00_spi_busy), 
        .B(n23534), .Y(n22838) );
  sky130_fd_sc_hd__clkinv_1 U24413 ( .A(n22838), .Y(n23511) );
  sky130_fd_sc_hd__nand2_1 U24414 ( .A(n23395), .B(
        j202_soc_core_wbqspiflash_00_state[1]), .Y(n23500) );
  sky130_fd_sc_hd__nor3_1 U24415 ( .A(n23513), .B(n23500), .C(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n23457) );
  sky130_fd_sc_hd__nor2_1 U24416 ( .A(n23511), .B(n23442), .Y(n22854) );
  sky130_fd_sc_hd__o21ai_1 U24417 ( .A1(j202_soc_core_wbqspiflash_00_spif_cmd), 
        .A2(n24903), .B1(j202_soc_core_wbqspiflash_00_spif_ctrl), .Y(n24995)
         );
  sky130_fd_sc_hd__nand2_1 U24418 ( .A(n23513), .B(n25027), .Y(n23528) );
  sky130_fd_sc_hd__nor2_1 U24419 ( .A(n23528), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n23462) );
  sky130_fd_sc_hd__nand2_1 U24420 ( .A(j202_soc_core_qspi_wb_addr[24]), .B(
        j202_soc_core_ahb2wbqspi_00_stb_o), .Y(n23359) );
  sky130_fd_sc_hd__nor2_1 U24421 ( .A(n23494), .B(n23359), .Y(n23403) );
  sky130_fd_sc_hd__nand2_1 U24422 ( .A(n23409), .B(n25053), .Y(n23564) );
  sky130_fd_sc_hd__nand2_1 U24423 ( .A(j202_soc_core_qspi_wb_addr[3]), .B(
        j202_soc_core_qspi_wb_addr[2]), .Y(n22833) );
  sky130_fd_sc_hd__nor2_1 U24424 ( .A(j202_soc_core_qspi_wb_we), .B(n23359), 
        .Y(n23425) );
  sky130_fd_sc_hd__nand3_1 U24425 ( .A(n25111), .B(
        j202_soc_core_wbqspiflash_00_write_in_progress), .C(n20103), .Y(n23431) );
  sky130_fd_sc_hd__clkinv_1 U24426 ( .A(n23431), .Y(n23463) );
  sky130_fd_sc_hd__a211oi_1 U24427 ( .A1(n22775), .A2(n22833), .B1(n23425), 
        .C1(n23463), .Y(n23477) );
  sky130_fd_sc_hd__clkinv_1 U24428 ( .A(n23477), .Y(n20105) );
  sky130_fd_sc_hd__clkinv_1 U24429 ( .A(
        j202_soc_core_wbqspiflash_00_write_in_progress), .Y(n23495) );
  sky130_fd_sc_hd__nor2_1 U24430 ( .A(
        j202_soc_core_wbqspiflash_00_write_in_progress), .B(n23564), .Y(n23428) );
  sky130_fd_sc_hd__nor2_1 U24431 ( .A(j202_soc_core_qspi_wb_addr[24]), .B(
        n20103), .Y(n20217) );
  sky130_fd_sc_hd__nand2_1 U24432 ( .A(n20217), .B(n23494), .Y(n23422) );
  sky130_fd_sc_hd__clkinv_1 U24433 ( .A(n23422), .Y(n23382) );
  sky130_fd_sc_hd__clkinv_1 U24434 ( .A(
        j202_soc_core_wbqspiflash_00_write_protect), .Y(n23758) );
  sky130_fd_sc_hd__nand2_1 U24435 ( .A(n23403), .B(
        j202_soc_core_qspi_wb_wdat[31]), .Y(n23407) );
  sky130_fd_sc_hd__nor2_1 U24436 ( .A(j202_soc_core_qspi_wb_addr[2]), .B(
        n23407), .Y(n23519) );
  sky130_fd_sc_hd__o22ai_1 U24437 ( .A1(n23382), .A2(n23758), .B1(n20217), 
        .B2(n23519), .Y(n20104) );
  sky130_fd_sc_hd__o21ai_1 U24438 ( .A1(n23477), .A2(n23428), .B1(n20104), .Y(
        n23518) );
  sky130_fd_sc_hd__nor2_1 U24440 ( .A(n24899), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n23541) );
  sky130_fd_sc_hd__nand2_1 U24441 ( .A(n25027), .B(n23541), .Y(n23468) );
  sky130_fd_sc_hd__a21oi_1 U24443 ( .A1(n22854), .A2(n24995), .B1(n20106), .Y(
        n23392) );
  sky130_fd_sc_hd__nand2_1 U24444 ( .A(n23395), .B(n22847), .Y(n23529) );
  sky130_fd_sc_hd__nor2_1 U24445 ( .A(j202_soc_core_wbqspiflash_00_spi_wr), 
        .B(j202_soc_core_wbqspiflash_00_spi_busy), .Y(n25100) );
  sky130_fd_sc_hd__nand2_1 U24446 ( .A(n25100), .B(io_out[8]), .Y(n23515) );
  sky130_fd_sc_hd__nor2_1 U24447 ( .A(n24899), .B(n23515), .Y(n22770) );
  sky130_fd_sc_hd__nand2_1 U24448 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .Y(n22839) );
  sky130_fd_sc_hd__nand2_1 U24449 ( .A(n24903), .B(n24901), .Y(n23757) );
  sky130_fd_sc_hd__nand2_1 U24450 ( .A(n22839), .B(n23757), .Y(n23447) );
  sky130_fd_sc_hd__nand2_1 U24452 ( .A(j202_soc_core_wbqspiflash_00_spif_cmd), 
        .B(j202_soc_core_wbqspiflash_00_spif_ctrl), .Y(n23562) );
  sky130_fd_sc_hd__a21oi_1 U24453 ( .A1(n23447), .A2(n23402), .B1(n23562), .Y(
        n23498) );
  sky130_fd_sc_hd__clkinv_1 U24454 ( .A(j202_soc_core_wbqspiflash_00_spif_ctrl), .Y(n25015) );
  sky130_fd_sc_hd__nor3_1 U24455 ( .A(n23760), .B(
        j202_soc_core_wbqspiflash_00_spif_cmd), .C(n25015), .Y(n23481) );
  sky130_fd_sc_hd__nor2_1 U24456 ( .A(n23498), .B(n23481), .Y(n20107) );
  sky130_fd_sc_hd__nand2_1 U24457 ( .A(n25015), .B(
        j202_soc_core_wbqspiflash_00_spif_cmd), .Y(n25031) );
  sky130_fd_sc_hd__clkinv_1 U24458 ( .A(n25031), .Y(n24998) );
  sky130_fd_sc_hd__nand3_1 U24459 ( .A(n24998), .B(n23495), .C(n23758), .Y(
        n23401) );
  sky130_fd_sc_hd__nand2_1 U24460 ( .A(n20107), .B(n23401), .Y(n23377) );
  sky130_fd_sc_hd__nand2_1 U24461 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(n23788), .Y(n23478) );
  sky130_fd_sc_hd__nor3_1 U24462 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[2]), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[0]), .C(
        j202_soc_core_wbqspiflash_00_reset_counter[1]), .Y(n23767) );
  sky130_fd_sc_hd__clkinv_1 U24463 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[3]), .Y(n23802) );
  sky130_fd_sc_hd__nand2_1 U24464 ( .A(n23767), .B(n23802), .Y(n23771) );
  sky130_fd_sc_hd__nor2_1 U24465 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[4]), .B(n23771), .Y(n23773)
         );
  sky130_fd_sc_hd__nand2b_1 U24466 ( .A_N(
        j202_soc_core_wbqspiflash_00_reset_counter[5]), .B(n23773), .Y(n23776)
         );
  sky130_fd_sc_hd__nor2_1 U24467 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[6]), .B(n23776), .Y(n23778)
         );
  sky130_fd_sc_hd__nand2b_1 U24468 ( .A_N(
        j202_soc_core_wbqspiflash_00_reset_counter[7]), .B(n23778), .Y(n23781)
         );
  sky130_fd_sc_hd__nor2_1 U24469 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[8]), .B(n23781), .Y(n23783)
         );
  sky130_fd_sc_hd__clkinv_1 U24470 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[9]), .Y(n23801) );
  sky130_fd_sc_hd__nand2_1 U24471 ( .A(n23783), .B(n23801), .Y(n23785) );
  sky130_fd_sc_hd__nand2_1 U24472 ( .A(j202_soc_core_wbqspiflash_00_state[2]), 
        .B(n25064), .Y(n25068) );
  sky130_fd_sc_hd__nor2_1 U24473 ( .A(n25070), .B(n25068), .Y(n25085) );
  sky130_fd_sc_hd__clkinv_1 U24474 ( .A(n23564), .Y(n20109) );
  sky130_fd_sc_hd__nand2_1 U24475 ( .A(n23494), .B(
        j202_soc_core_qspi_wb_addr[24]), .Y(n22834) );
  sky130_fd_sc_hd__clkinv_1 U24476 ( .A(n22834), .Y(n20108) );
  sky130_fd_sc_hd__nand2_1 U24477 ( .A(n20109), .B(n20108), .Y(n20119) );
  sky130_fd_sc_hd__nor2_1 U24478 ( .A(j202_soc_core_wbqspiflash_00_state[4]), 
        .B(j202_soc_core_wbqspiflash_00_state[2]), .Y(n25005) );
  sky130_fd_sc_hd__nand2_1 U24479 ( .A(n25005), .B(n25027), .Y(n23756) );
  sky130_fd_sc_hd__nand2_1 U24480 ( .A(j202_soc_core_ahb2wbqspi_00_stb_o), .B(
        n23762), .Y(n25118) );
  sky130_fd_sc_hd__clkinv_1 U24481 ( .A(n25118), .Y(n20110) );
  sky130_fd_sc_hd__nand2_1 U24482 ( .A(n20110), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n20118) );
  sky130_fd_sc_hd__clkinv_1 U24483 ( .A(n20118), .Y(n20111) );
  sky130_fd_sc_hd__nor2_1 U24484 ( .A(n25085), .B(n23525), .Y(n23375) );
  sky130_fd_sc_hd__nor2_1 U24485 ( .A(n23513), .B(n23529), .Y(n25000) );
  sky130_fd_sc_hd__nor2_1 U24486 ( .A(j202_soc_core_wbqspiflash_00_spi_busy), 
        .B(n23491), .Y(n23372) );
  sky130_fd_sc_hd__nor2_1 U24487 ( .A(n25005), .B(n23478), .Y(n22858) );
  sky130_fd_sc_hd__nor3_1 U24488 ( .A(n24898), .B(n23372), .C(n22858), .Y(
        n20112) );
  sky130_fd_sc_hd__o211ai_1 U24489 ( .A1(n23478), .A2(n23785), .B1(n23375), 
        .C1(n20112), .Y(n20113) );
  sky130_fd_sc_hd__a31oi_1 U24490 ( .A1(n23788), .A2(n22770), .A3(n23377), 
        .B1(n20113), .Y(n22850) );
  sky130_fd_sc_hd__a31oi_1 U24491 ( .A1(n23483), .A2(n23392), .A3(n22850), 
        .B1(j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N752) );
  sky130_fd_sc_hd__nor2b_1 U24492 ( .B_N(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[0]), .A(
        j202_soc_core_wbqspiflash_00_spif_override), .Y(io_out[10]) );
  sky130_fd_sc_hd__nor2b_1 U24493 ( .B_N(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[1]), .A(
        j202_soc_core_wbqspiflash_00_spif_override), .Y(io_out[11]) );
  sky130_fd_sc_hd__o2bb2ai_1 U24494 ( .B1(n24400), .B2(n24442), .A1_N(
        j202_soc_core_intc_core_00_rg_ie[29]), .A2_N(n20114), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o2bb2ai_1 U24495 ( .B1(n24400), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[55]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o2bb2ai_1 U24496 ( .B1(n24400), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[39]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o2bb2ai_1 U24497 ( .B1(n20477), .B2(n24488), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[121]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o2bb2ai_1 U24498 ( .B1(n20477), .B2(n24485), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[89]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o2bb2ai_1 U24499 ( .B1(n24488), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[113]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o2bb2ai_1 U24500 ( .B1(n24485), .B2(n20475), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[81]), .A2_N(n20473), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o2bb2ai_1 U24501 ( .B1(n24488), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[97]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o2bb2ai_1 U24502 ( .B1(n24485), .B2(n24290), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[65]), .A2_N(n20115), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__nand2_1 U24503 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_state[1]), .B(n20116), .Y(n23597) );
  sky130_fd_sc_hd__nand2_1 U24504 ( .A(n25734), .B(n23597), .Y(n23589) );
  sky130_fd_sc_hd__nor2_1 U24505 ( .A(n21324), .B(n23589), .Y(n23599) );
  sky130_fd_sc_hd__nand2_1 U24506 ( .A(n23599), .B(n23587), .Y(n23750) );
  sky130_fd_sc_hd__nor2_1 U24507 ( .A(n20116), .B(j202_soc_core_rst), .Y(
        n20117) );
  sky130_fd_sc_hd__nand3_1 U24508 ( .A(n23750), .B(n22886), .C(n20117), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N311) );
  sky130_fd_sc_hd__nand2_1 U24509 ( .A(n25027), .B(n25070), .Y(n22843) );
  sky130_fd_sc_hd__nor2_1 U24510 ( .A(n23451), .B(n22843), .Y(n23364) );
  sky130_fd_sc_hd__nand2_1 U24511 ( .A(n23364), .B(n23425), .Y(n25065) );
  sky130_fd_sc_hd__nor2_1 U24512 ( .A(n20119), .B(n20118), .Y(n22779) );
  sky130_fd_sc_hd__nor2_1 U24513 ( .A(j202_soc_core_wbqspiflash_00_spi_len[0]), 
        .B(j202_soc_core_wbqspiflash_00_spi_len[1]), .Y(n23510) );
  sky130_fd_sc_hd__nand2_1 U24514 ( .A(n23526), .B(n25070), .Y(n25018) );
  sky130_fd_sc_hd__nand2_1 U24515 ( .A(n23384), .B(n23479), .Y(n23509) );
  sky130_fd_sc_hd__nand2_1 U24516 ( .A(n23526), .B(n23450), .Y(n25108) );
  sky130_fd_sc_hd__a21oi_1 U24517 ( .A1(n23510), .A2(n20120), .B1(n23787), .Y(
        n20121) );
  sky130_fd_sc_hd__nor2_1 U24518 ( .A(n23363), .B(
        j202_soc_core_wbqspiflash_00_spi_in[31]), .Y(n23292) );
  sky130_fd_sc_hd__nor2_1 U24519 ( .A(n25070), .B(n23451), .Y(n23536) );
  sky130_fd_sc_hd__nand2_1 U24520 ( .A(n23384), .B(n23536), .Y(n25107) );
  sky130_fd_sc_hd__o22ai_1 U24521 ( .A1(n20121), .A2(n23363), .B1(n25109), 
        .B2(n25107), .Y(n22771) );
  sky130_fd_sc_hd__a211oi_1 U24522 ( .A1(n23428), .A2(n25047), .B1(n22779), 
        .C1(n22771), .Y(n20122) );
  sky130_fd_sc_hd__nor2_1 U24523 ( .A(n25018), .B(n23433), .Y(n23754) );
  sky130_fd_sc_hd__nand2_1 U24524 ( .A(j202_soc_core_wbqspiflash_00_spi_valid), 
        .B(n23754), .Y(n23368) );
  sky130_fd_sc_hd__clkbuf_1 U24525 ( .A(j202_soc_core_wbqspiflash_00_N755), 
        .X(n25536) );
  sky130_fd_sc_hd__nand3_1 U24526 ( .A(n21218), .B(
        j202_soc_core_ahb2apb_02_state[1]), .C(n20123), .Y(n24069) );
  sky130_fd_sc_hd__and3_1 U24527 ( .A(j202_soc_core_pwrite[2]), .B(
        j202_soc_core_pstrb[2]), .C(j202_soc_core_pstrb[0]), .X(n20124) );
  sky130_fd_sc_hd__nand4_1 U24528 ( .A(n20125), .B(j202_soc_core_pstrb[3]), 
        .C(j202_soc_core_pstrb[1]), .D(n20124), .Y(n23867) );
  sky130_fd_sc_hd__clkinv_1 U24529 ( .A(j202_soc_core_gpio_core_00_reg_addr[2]), .Y(n20126) );
  sky130_fd_sc_hd__nor2_1 U24530 ( .A(j202_soc_core_gpio_core_00_reg_addr[7]), 
        .B(n20126), .Y(n20127) );
  sky130_fd_sc_hd__nor2_1 U24531 ( .A(j202_soc_core_gpio_core_00_reg_addr[1]), 
        .B(j202_soc_core_gpio_core_00_reg_addr[0]), .Y(n20133) );
  sky130_fd_sc_hd__nor2_1 U24532 ( .A(j202_soc_core_gpio_core_00_reg_addr[6]), 
        .B(j202_soc_core_gpio_core_00_reg_addr[5]), .Y(n20131) );
  sky130_fd_sc_hd__nand3_1 U24533 ( .A(n20127), .B(n20133), .C(n20131), .Y(
        n24073) );
  sky130_fd_sc_hd__nor2_1 U24534 ( .A(j202_soc_core_gpio_core_00_reg_addr[4]), 
        .B(j202_soc_core_gpio_core_00_reg_addr[3]), .Y(n24070) );
  sky130_fd_sc_hd__nand2_1 U24535 ( .A(n20130), .B(n24070), .Y(n20128) );
  sky130_fd_sc_hd__o21ai_2 U24536 ( .A1(n23867), .A2(n20128), .B1(n25730), .Y(
        n10673) );
  sky130_fd_sc_hd__nor2b_1 U24537 ( .B_N(
        j202_soc_core_gpio_core_00_reg_addr[4]), .A(
        j202_soc_core_gpio_core_00_reg_addr[3]), .Y(n23866) );
  sky130_fd_sc_hd__nand2_1 U24538 ( .A(n20130), .B(n23866), .Y(n24077) );
  sky130_fd_sc_hd__o21ai_1 U24539 ( .A1(n23867), .A2(n24077), .B1(n25734), .Y(
        n10670) );
  sky130_fd_sc_hd__clkbuf_1 U24540 ( .A(n10670), .X(n25534) );
  sky130_fd_sc_hd__clkinv_1 U24541 ( .A(j202_soc_core_gpio_core_00_reg_addr[3]), .Y(n20129) );
  sky130_fd_sc_hd__nor2_1 U24542 ( .A(j202_soc_core_gpio_core_00_reg_addr[4]), 
        .B(n20129), .Y(n20134) );
  sky130_fd_sc_hd__nand2_1 U24543 ( .A(n20130), .B(n20134), .Y(n24076) );
  sky130_fd_sc_hd__o21ai_1 U24544 ( .A1(n23867), .A2(n24076), .B1(n25734), .Y(
        n10671) );
  sky130_fd_sc_hd__nor2_1 U24545 ( .A(j202_soc_core_gpio_core_00_reg_addr[2]), 
        .B(j202_soc_core_gpio_core_00_reg_addr[7]), .Y(n20132) );
  sky130_fd_sc_hd__and3_1 U24546 ( .A(n20133), .B(n20132), .C(n20131), .X(
        n24071) );
  sky130_fd_sc_hd__nand2_1 U24547 ( .A(n24071), .B(n20134), .Y(n24078) );
  sky130_fd_sc_hd__o21ai_1 U24548 ( .A1(n23867), .A2(n24078), .B1(n25734), .Y(
        n10672) );
  sky130_fd_sc_hd__nand2_1 U24549 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(n25027), .Y(n23476) );
  sky130_fd_sc_hd__nor2_1 U24550 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]), .B(n25067), .Y(n20137)
         );
  sky130_fd_sc_hd__nor2_1 U24551 ( .A(j202_soc_core_qspi_wb_addr[21]), .B(
        n25069), .Y(n20135) );
  sky130_fd_sc_hd__nor2_1 U24552 ( .A(n20137), .B(n20135), .Y(n20138) );
  sky130_fd_sc_hd__nor2_1 U24553 ( .A(n22839), .B(n24905), .Y(n20144) );
  sky130_fd_sc_hd__nand2_1 U24554 ( .A(n20144), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[5]), .Y(n20163) );
  sky130_fd_sc_hd__nor2_1 U24555 ( .A(n20163), .B(n24909), .Y(n20162) );
  sky130_fd_sc_hd__nand2_1 U24556 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[7]), .B(n20162), .Y(n20161)
         );
  sky130_fd_sc_hd__nor2_1 U24557 ( .A(n24940), .B(n20161), .Y(n20146) );
  sky130_fd_sc_hd__nand2_1 U24558 ( .A(n20146), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[9]), .Y(n20154) );
  sky130_fd_sc_hd__nor3_1 U24559 ( .A(n20154), .B(n24925), .C(n24922), .Y(
        n20152) );
  sky130_fd_sc_hd__nand2_1 U24560 ( .A(n20152), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[12]), .Y(n20151) );
  sky130_fd_sc_hd__nand2_1 U24561 ( .A(n20187), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[13]), .Y(n20186) );
  sky130_fd_sc_hd__nand2b_1 U24562 ( .A_N(n20186), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]), .Y(n20179) );
  sky130_fd_sc_hd__nor3_1 U24563 ( .A(n20179), .B(n24944), .C(n24987), .Y(
        n23380) );
  sky130_fd_sc_hd__nor2b_1 U24564 ( .B_N(n23380), .A(n25019), .Y(n20195) );
  sky130_fd_sc_hd__nand2_1 U24565 ( .A(n20195), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .Y(n20196) );
  sky130_fd_sc_hd__nor2_1 U24566 ( .A(n20196), .B(n23567), .Y(n20206) );
  sky130_fd_sc_hd__xnor2_1 U24567 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .B(
        j202_soc_core_qspi_wb_addr[22]), .Y(n20208) );
  sky130_fd_sc_hd__o22ai_1 U24569 ( .A1(n20138), .A2(n20207), .B1(n20137), 
        .B2(n20136), .Y(n20216) );
  sky130_fd_sc_hd__nor2_1 U24570 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[10]), .B(n20139), .Y(n20155)
         );
  sky130_fd_sc_hd__xnor2_1 U24571 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[11]), .B(
        j202_soc_core_qspi_wb_addr[11]), .Y(n20171) );
  sky130_fd_sc_hd__xnor2_1 U24572 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[8]), .B(
        j202_soc_core_qspi_wb_addr[8]), .Y(n20218) );
  sky130_fd_sc_hd__nand2_1 U24573 ( .A(n20218), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[7]), .Y(n20140) );
  sky130_fd_sc_hd__o21ai_1 U24574 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[7]), .A2(n20162), .B1(n20161), 
        .Y(n20156) );
  sky130_fd_sc_hd__a21oi_1 U24575 ( .A1(n20140), .A2(n20156), .B1(
        j202_soc_core_qspi_wb_addr[7]), .Y(n20141) );
  sky130_fd_sc_hd__a31oi_1 U24576 ( .A1(n20143), .A2(n20142), .A3(n20171), 
        .B1(n20141), .Y(n20194) );
  sky130_fd_sc_hd__xor2_1 U24578 ( .A(j202_soc_core_qspi_wb_addr[5]), .B(
        n20145), .X(n20178) );
  sky130_fd_sc_hd__xnor2_1 U24579 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[4]), .B(
        j202_soc_core_qspi_wb_addr[4]), .Y(n20173) );
  sky130_fd_sc_hd__o21ai_1 U24580 ( .A1(n20146), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[9]), .B1(n20154), .Y(n20147)
         );
  sky130_fd_sc_hd__xnor2_1 U24581 ( .A(j202_soc_core_qspi_wb_addr[9]), .B(
        n20147), .Y(n20148) );
  sky130_fd_sc_hd__a31oi_1 U24582 ( .A1(n23757), .A2(n23409), .A3(n20173), 
        .B1(n20148), .Y(n20177) );
  sky130_fd_sc_hd__nor2_1 U24583 ( .A(j202_soc_core_qspi_wb_addr[15]), .B(
        n24987), .Y(n20150) );
  sky130_fd_sc_hd__xnor2_1 U24584 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]), .B(
        j202_soc_core_qspi_wb_addr[16]), .Y(n20181) );
  sky130_fd_sc_hd__xnor2_1 U24585 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .B(n25053), .Y(n20149)
         );
  sky130_fd_sc_hd__o21ai_1 U24586 ( .A1(n20150), .A2(n20181), .B1(n20149), .Y(
        n20160) );
  sky130_fd_sc_hd__xor2_1 U24588 ( .A(j202_soc_core_qspi_wb_addr[12]), .B(
        n20153), .X(n20159) );
  sky130_fd_sc_hd__nor2_1 U24589 ( .A(j202_soc_core_qspi_wb_addr[10]), .B(
        n24922), .Y(n20172) );
  sky130_fd_sc_hd__nand2_1 U24591 ( .A(n20156), .B(
        j202_soc_core_qspi_wb_addr[7]), .Y(n20157) );
  sky130_fd_sc_hd__nand4b_1 U24592 ( .A_N(n20160), .B(n20159), .C(n20158), .D(
        n20157), .Y(n20170) );
  sky130_fd_sc_hd__xnor2_1 U24593 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[15]), .B(
        j202_soc_core_qspi_wb_addr[15]), .Y(n20182) );
  sky130_fd_sc_hd__xnor2_1 U24594 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]), .B(
        j202_soc_core_qspi_wb_addr[23]), .Y(n20209) );
  sky130_fd_sc_hd__o22ai_1 U24595 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]), .A2(n20182), .B1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .B2(n20209), .Y(n20169)
         );
  sky130_fd_sc_hd__a21oi_1 U24596 ( .A1(n24909), .A2(n20163), .B1(n20162), .Y(
        n20164) );
  sky130_fd_sc_hd__xnor2_1 U24597 ( .A(j202_soc_core_qspi_wb_addr[6]), .B(
        n20164), .Y(n20166) );
  sky130_fd_sc_hd__nand2_1 U24598 ( .A(n23447), .B(
        j202_soc_core_qspi_wb_addr[3]), .Y(n20165) );
  sky130_fd_sc_hd__o211ai_1 U24599 ( .A1(n20167), .A2(n20218), .B1(n20166), 
        .C1(n20165), .Y(n20168) );
  sky130_fd_sc_hd__nor3_1 U24600 ( .A(n20170), .B(n20169), .C(n20168), .Y(
        n20176) );
  sky130_fd_sc_hd__o22ai_1 U24601 ( .A1(n20174), .A2(n20173), .B1(n20172), 
        .B2(n20171), .Y(n20175) );
  sky130_fd_sc_hd__and4b_1 U24602 ( .B(n20178), .C(n20177), .D(n20176), .A_N(
        n20175), .X(n20193) );
  sky130_fd_sc_hd__xor2_1 U24603 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]), .B(
        j202_soc_core_qspi_wb_addr[14]), .X(n20185) );
  sky130_fd_sc_hd__nor2_1 U24604 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[15]), .B(n24986), .Y(n20180)
         );
  sky130_fd_sc_hd__nor3b_1 U24605 ( .C_N(n20181), .A(n20180), .B(n20179), .Y(
        n20184) );
  sky130_fd_sc_hd__a21oi_1 U24606 ( .A1(n20182), .A2(n20186), .B1(n20185), .Y(
        n20183) );
  sky130_fd_sc_hd__a211oi_1 U24607 ( .A1(n20185), .A2(n20186), .B1(n20184), 
        .C1(n20183), .Y(n20192) );
  sky130_fd_sc_hd__xor2_1 U24608 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .B(
        j202_soc_core_qspi_wb_addr[19]), .X(n20190) );
  sky130_fd_sc_hd__xnor2_1 U24610 ( .A(j202_soc_core_qspi_wb_addr[13]), .B(
        n20188), .Y(n20189) );
  sky130_fd_sc_hd__a21oi_1 U24611 ( .A1(n20196), .A2(n20190), .B1(n20189), .Y(
        n20191) );
  sky130_fd_sc_hd__nand4_1 U24612 ( .A(n20194), .B(n20193), .C(n20192), .D(
        n20191), .Y(n20215) );
  sky130_fd_sc_hd__xor2_1 U24613 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]), .B(
        j202_soc_core_qspi_wb_addr[20]), .X(n20198) );
  sky130_fd_sc_hd__nor2_1 U24614 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .B(n20195), .Y(n20199)
         );
  sky130_fd_sc_hd__nand2_1 U24615 ( .A(n20199), .B(
        j202_soc_core_qspi_wb_addr[18]), .Y(n20204) );
  sky130_fd_sc_hd__a21oi_1 U24616 ( .A1(j202_soc_core_qspi_wb_addr[19]), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .B1(
        j202_soc_core_qspi_wb_addr[18]), .Y(n20197) );
  sky130_fd_sc_hd__o21ai_1 U24617 ( .A1(j202_soc_core_qspi_wb_addr[19]), .A2(
        n20198), .B1(n20197), .Y(n20201) );
  sky130_fd_sc_hd__nor3_1 U24618 ( .A(j202_soc_core_qspi_wb_addr[18]), .B(
        n20199), .C(n20202), .Y(n20200) );
  sky130_fd_sc_hd__a21oi_1 U24619 ( .A1(n20202), .A2(n20201), .B1(n20200), .Y(
        n20203) );
  sky130_fd_sc_hd__o211ai_1 U24620 ( .A1(n20206), .A2(n20205), .B1(n20204), 
        .C1(n20203), .Y(n20214) );
  sky130_fd_sc_hd__nand2_1 U24621 ( .A(n20207), .B(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]), .Y(n20212) );
  sky130_fd_sc_hd__o21ai_1 U24622 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[23]), .A2(n25088), .B1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .Y(n20211) );
  sky130_fd_sc_hd__a21bo_2 U24623 ( .A1(n20209), .A2(n20208), .B1_N(n20212), 
        .X(n20210) );
  sky130_fd_sc_hd__nor4_1 U24625 ( .A(n20216), .B(n20215), .C(n20214), .D(
        n20213), .Y(n23383) );
  sky130_fd_sc_hd__xor2_1 U24626 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[17]), .B(
        j202_soc_core_qspi_wb_addr[17]), .X(n23381) );
  sky130_fd_sc_hd__nor2_1 U24627 ( .A(n23380), .B(n23381), .Y(n23379) );
  sky130_fd_sc_hd__nand4_1 U24628 ( .A(n23383), .B(n23379), .C(n23404), .D(
        n20218), .Y(n23291) );
  sky130_fd_sc_hd__nor2_1 U24629 ( .A(j202_soc_core_wbqspiflash_00_spi_wr), 
        .B(n23291), .Y(n23550) );
  sky130_fd_sc_hd__nand2_1 U24630 ( .A(j202_soc_core_qspi_wb_cyc), .B(n23550), 
        .Y(n23506) );
  sky130_fd_sc_hd__nor2_1 U24631 ( .A(n23476), .B(n23506), .Y(n25117) );
  sky130_fd_sc_hd__nand2_1 U24632 ( .A(n24899), .B(
        j202_soc_core_wbqspiflash_00_state[4]), .Y(n23412) );
  sky130_fd_sc_hd__nor2_1 U24633 ( .A(n23526), .B(n22856), .Y(n25102) );
  sky130_fd_sc_hd__nor2_1 U24635 ( .A(j202_soc_core_rst), .B(n23360), .Y(
        n25492) );
  sky130_fd_sc_hd__nor2_1 U24636 ( .A(n20220), .B(n22798), .Y(n20224) );
  sky130_fd_sc_hd__nor2_1 U24637 ( .A(n20225), .B(j202_soc_core_j22_cpu_rte4), 
        .Y(n20222) );
  sky130_fd_sc_hd__and3_1 U24638 ( .A(n22800), .B(n20222), .C(n20221), .X(
        n20223) );
  sky130_fd_sc_hd__nand2_1 U24639 ( .A(n20224), .B(n20223), .Y(n21618) );
  sky130_fd_sc_hd__nand2_1 U24640 ( .A(n25734), .B(n20225), .Y(n22374) );
  sky130_fd_sc_hd__nor2_1 U24641 ( .A(n20225), .B(j202_soc_core_rst), .Y(
        n21617) );
  sky130_fd_sc_hd__nand3_1 U24642 ( .A(n23239), .B(
        j202_soc_core_j22_cpu_regop_We__1_), .C(n20478), .Y(n20483) );
  sky130_fd_sc_hd__nand2b_1 U24643 ( .A_N(n20483), .B(n20237), .Y(n20227) );
  sky130_fd_sc_hd__nand3_1 U24644 ( .A(n23239), .B(
        j202_soc_core_j22_cpu_regop_We__2_), .C(n20226), .Y(n21997) );
  sky130_fd_sc_hd__nand2_1 U24645 ( .A(n20227), .B(n21997), .Y(n21619) );
  sky130_fd_sc_hd__o22ai_1 U24646 ( .A1(n21672), .A2(n22374), .B1(n20228), 
        .B2(n21619), .Y(n20229) );
  sky130_fd_sc_hd__nand2_1 U24647 ( .A(n20235), .B(n20230), .Y(n23236) );
  sky130_fd_sc_hd__nand2_1 U24648 ( .A(n21672), .B(n20232), .Y(n20481) );
  sky130_fd_sc_hd__nor2_1 U24649 ( .A(j202_soc_core_j22_cpu_regop_We__1_), .B(
        j202_soc_core_j22_cpu_regop_We__2_), .Y(n20233) );
  sky130_fd_sc_hd__nor2_1 U24650 ( .A(n20234), .B(n21657), .Y(n20264) );
  sky130_fd_sc_hd__nand3_1 U24651 ( .A(n20264), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__3_), .C(
        j202_soc_core_j22_cpu_regop_M_Rn__2_), .Y(n20324) );
  sky130_fd_sc_hd__nand2_1 U24652 ( .A(j202_soc_core_j22_cpu_regop_M_Rn__1_), 
        .B(j202_soc_core_j22_cpu_regop_M_Rn__0_), .Y(n20320) );
  sky130_fd_sc_hd__nand3_1 U24653 ( .A(n20236), .B(
        j202_soc_core_j22_cpu_regop_M_Wm__2_), .C(n20235), .Y(n20244) );
  sky130_fd_sc_hd__nand3_1 U24654 ( .A(n20237), .B(
        j202_soc_core_j22_cpu_regop_We__2_), .C(
        j202_soc_core_j22_cpu_regop_We__1_), .Y(n20242) );
  sky130_fd_sc_hd__nand2_1 U24655 ( .A(n20256), .B(n20238), .Y(n20240) );
  sky130_fd_sc_hd__o211ai_2 U24656 ( .A1(n20324), .A2(n20320), .B1(n20244), 
        .C1(n21188), .Y(j202_soc_core_j22_cpu_rf_N3264) );
  sky130_fd_sc_hd__nand2_1 U24657 ( .A(n20264), .B(n20246), .Y(n20322) );
  sky130_fd_sc_hd__nand2_1 U24658 ( .A(n21672), .B(n20247), .Y(n20254) );
  sky130_fd_sc_hd__a21o_1 U24659 ( .A1(n20249), .A2(
        j202_soc_core_j22_cpu_regop_We__1_), .B1(n20248), .X(n20252) );
  sky130_fd_sc_hd__nand2_1 U24660 ( .A(n20256), .B(n20250), .Y(n20251) );
  sky130_fd_sc_hd__nand2_1 U24661 ( .A(n20252), .B(n20251), .Y(n20253) );
  sky130_fd_sc_hd__o211ai_2 U24662 ( .A1(n20268), .A2(n20322), .B1(n20254), 
        .C1(n21190), .Y(j202_soc_core_j22_cpu_rf_N2709) );
  sky130_fd_sc_hd__nand3_1 U24663 ( .A(n20264), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__3_), .C(n20255), .Y(n20319) );
  sky130_fd_sc_hd__a22oi_1 U24664 ( .A1(n20306), .A2(n20258), .B1(n20271), 
        .B2(n20257), .Y(n20259) );
  sky130_fd_sc_hd__o21ai_2 U24665 ( .A1(n20268), .A2(n20319), .B1(n21193), .Y(
        j202_soc_core_j22_cpu_rf_N3005) );
  sky130_fd_sc_hd__a22oi_1 U24666 ( .A1(n20306), .A2(n20261), .B1(n20271), 
        .B2(n20260), .Y(n20262) );
  sky130_fd_sc_hd__nand3_1 U24667 ( .A(n20264), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__2_), .C(n20263), .Y(n20321) );
  sky130_fd_sc_hd__a22oi_1 U24668 ( .A1(n20306), .A2(n20266), .B1(n20271), 
        .B2(n20265), .Y(n20267) );
  sky130_fd_sc_hd__o21ai_2 U24669 ( .A1(n20268), .A2(n20321), .B1(n21194), .Y(
        j202_soc_core_j22_cpu_rf_N2857) );
  sky130_fd_sc_hd__nand2_1 U24670 ( .A(n20269), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__1_), .Y(n20325) );
  sky130_fd_sc_hd__a22oi_1 U24671 ( .A1(n20306), .A2(n20272), .B1(n20271), 
        .B2(n20270), .Y(n20273) );
  sky130_fd_sc_hd__nand3_1 U24672 ( .A(n23239), .B(n20276), .C(n20275), .Y(
        n22372) );
  sky130_fd_sc_hd__nand2_1 U24673 ( .A(n20306), .B(n20280), .Y(n20281) );
  sky130_fd_sc_hd__o211ai_2 U24674 ( .A1(n20309), .A2(n20282), .B1(n20281), 
        .C1(n20307), .Y(n21068) );
  sky130_fd_sc_hd__nand2_1 U24675 ( .A(n20306), .B(n20283), .Y(n20284) );
  sky130_fd_sc_hd__nand2_1 U24676 ( .A(n20306), .B(n20286), .Y(n20287) );
  sky130_fd_sc_hd__o211ai_2 U24677 ( .A1(n20309), .A2(n20288), .B1(n20287), 
        .C1(n20307), .Y(n21134) );
  sky130_fd_sc_hd__nand2_1 U24678 ( .A(n20306), .B(n20289), .Y(n20290) );
  sky130_fd_sc_hd__o211ai_2 U24679 ( .A1(n20309), .A2(n11183), .B1(n20290), 
        .C1(n20307), .Y(n21073) );
  sky130_fd_sc_hd__nand2_1 U24680 ( .A(n20306), .B(n20291), .Y(n20292) );
  sky130_fd_sc_hd__o211ai_2 U24681 ( .A1(n20309), .A2(n20293), .B1(n20292), 
        .C1(n20307), .Y(n21202) );
  sky130_fd_sc_hd__nand2_1 U24682 ( .A(n20306), .B(n20294), .Y(n20295) );
  sky130_fd_sc_hd__o211ai_2 U24683 ( .A1(n20309), .A2(n20296), .B1(n20295), 
        .C1(n20307), .Y(n21072) );
  sky130_fd_sc_hd__nand2_1 U24684 ( .A(n20306), .B(n20297), .Y(n20298) );
  sky130_fd_sc_hd__o211ai_2 U24685 ( .A1(n20309), .A2(n11191), .B1(n20298), 
        .C1(n20307), .Y(n21132) );
  sky130_fd_sc_hd__nand2_1 U24686 ( .A(n20306), .B(n20299), .Y(n20300) );
  sky130_fd_sc_hd__o211ai_2 U24687 ( .A1(n20309), .A2(n20301), .B1(n20300), 
        .C1(n20307), .Y(n21133) );
  sky130_fd_sc_hd__nand2_1 U24688 ( .A(n20306), .B(n20302), .Y(n20303) );
  sky130_fd_sc_hd__o211ai_2 U24689 ( .A1(n20309), .A2(n20304), .B1(n20303), 
        .C1(n20307), .Y(n21200) );
  sky130_fd_sc_hd__nand2_1 U24690 ( .A(n20306), .B(n20305), .Y(n20308) );
  sky130_fd_sc_hd__o211ai_2 U24691 ( .A1(n20309), .A2(n11193), .B1(n20308), 
        .C1(n20307), .Y(n21205) );
  sky130_fd_sc_hd__nor2_1 U24692 ( .A(n20310), .B(n21253), .Y(n20311) );
  sky130_fd_sc_hd__buf_4 U24693 ( .A(n20311), .X(n25523) );
  sky130_fd_sc_hd__nor2_1 U24694 ( .A(n20312), .B(n21253), .Y(n20313) );
  sky130_fd_sc_hd__buf_4 U24695 ( .A(n20313), .X(n25500) );
  sky130_fd_sc_hd__nor2_1 U24696 ( .A(n20314), .B(n21253), .Y(n20315) );
  sky130_fd_sc_hd__nand2_1 U24698 ( .A(n20318), .B(
        j202_soc_core_j22_cpu_regop_M_Rn__0_), .Y(n20323) );
  sky130_fd_sc_hd__o21ai_2 U24699 ( .A1(n20319), .A2(n20323), .B1(n21102), .Y(
        j202_soc_core_j22_cpu_rf_N3042) );
  sky130_fd_sc_hd__o21ai_2 U24700 ( .A1(n20321), .A2(n20323), .B1(n21200), .Y(
        j202_soc_core_j22_cpu_rf_N2894) );
  sky130_fd_sc_hd__o21ai_2 U24701 ( .A1(n20322), .A2(n20320), .B1(n21072), .Y(
        j202_soc_core_j22_cpu_rf_N2820) );
  sky130_fd_sc_hd__o21ai_2 U24702 ( .A1(n20321), .A2(n20320), .B1(n21133), .Y(
        j202_soc_core_j22_cpu_rf_N2968) );
  sky130_fd_sc_hd__o21ai_2 U24703 ( .A1(n20321), .A2(n20325), .B1(n21132), .Y(
        j202_soc_core_j22_cpu_rf_N2931) );
  sky130_fd_sc_hd__o21ai_2 U24704 ( .A1(n20322), .A2(n20323), .B1(n21202), .Y(
        j202_soc_core_j22_cpu_rf_N2746) );
  sky130_fd_sc_hd__o21ai_2 U24705 ( .A1(n20325), .A2(n20324), .B1(n21073), .Y(
        j202_soc_core_j22_cpu_rf_N3227) );
  sky130_fd_sc_hd__nand2_1 U24706 ( .A(n20339), .B(n20979), .Y(n22412) );
  sky130_fd_sc_hd__nor2_1 U24707 ( .A(n20327), .B(n20326), .Y(n20739) );
  sky130_fd_sc_hd__nand4_1 U24708 ( .A(n24872), .B(n25303), .C(n25315), .D(
        n25304), .Y(n20746) );
  sky130_fd_sc_hd__nand3_1 U24709 ( .A(n22342), .B(n24869), .C(n21424), .Y(
        n22413) );
  sky130_fd_sc_hd__nand3b_1 U24710 ( .A_N(n20739), .B(n20746), .C(n22413), .Y(
        n21532) );
  sky130_fd_sc_hd__nor2b_1 U24711 ( .B_N(n22412), .A(n21532), .Y(n21800) );
  sky130_fd_sc_hd__nand2_1 U24712 ( .A(n22342), .B(n21336), .Y(n22419) );
  sky130_fd_sc_hd__nor4_1 U24713 ( .A(n20328), .B(n21575), .C(n25377), .D(
        n20335), .Y(n20329) );
  sky130_fd_sc_hd__nor2_1 U24715 ( .A(n21420), .B(n25377), .Y(n20767) );
  sky130_fd_sc_hd__o21ai_1 U24716 ( .A1(n21575), .A2(n20767), .B1(n21563), .Y(
        n22740) );
  sky130_fd_sc_hd__nand2_1 U24717 ( .A(n20741), .B(n25377), .Y(n22384) );
  sky130_fd_sc_hd__nor2_1 U24718 ( .A(n22390), .B(n22384), .Y(n20994) );
  sky130_fd_sc_hd__nand2b_1 U24719 ( .A_N(n21734), .B(n25303), .Y(n21801) );
  sky130_fd_sc_hd__nand2_1 U24720 ( .A(n25304), .B(n21735), .Y(n21413) );
  sky130_fd_sc_hd__nor4b_1 U24721 ( .D_N(n22740), .A(n20994), .B(n22306), .C(
        n21492), .Y(n20345) );
  sky130_fd_sc_hd__nor2_1 U24722 ( .A(n21586), .B(n20340), .Y(n21332) );
  sky130_fd_sc_hd__nor2_1 U24723 ( .A(n21486), .B(n22387), .Y(n20333) );
  sky130_fd_sc_hd__nand2_1 U24724 ( .A(n20736), .B(n20333), .Y(n21556) );
  sky130_fd_sc_hd__nand2_1 U24725 ( .A(n22330), .B(n20766), .Y(n20987) );
  sky130_fd_sc_hd__nor2_1 U24726 ( .A(n21569), .B(n20987), .Y(n21608) );
  sky130_fd_sc_hd__nand3_1 U24727 ( .A(n20761), .B(n20981), .C(n25387), .Y(
        n21522) );
  sky130_fd_sc_hd__nor2_1 U24728 ( .A(n22342), .B(n21522), .Y(n24830) );
  sky130_fd_sc_hd__nor2_1 U24729 ( .A(n22333), .B(n22385), .Y(n21412) );
  sky130_fd_sc_hd__nor2_1 U24730 ( .A(n21505), .B(n21456), .Y(n24854) );
  sky130_fd_sc_hd__nand2_1 U24731 ( .A(n25381), .B(n20986), .Y(n22386) );
  sky130_fd_sc_hd__nor2_1 U24732 ( .A(n25380), .B(n22386), .Y(n20332) );
  sky130_fd_sc_hd__nand2_1 U24733 ( .A(n20332), .B(n21403), .Y(n23220) );
  sky130_fd_sc_hd__nor2_1 U24734 ( .A(n22386), .B(n21420), .Y(n24871) );
  sky130_fd_sc_hd__nand2_1 U24735 ( .A(n20737), .B(n24871), .Y(n24849) );
  sky130_fd_sc_hd__nand2_1 U24736 ( .A(n21403), .B(n21412), .Y(n24838) );
  sky130_fd_sc_hd__nor2_1 U24737 ( .A(n21505), .B(n20988), .Y(n24828) );
  sky130_fd_sc_hd__nor2b_1 U24738 ( .B_N(n24838), .A(n24828), .Y(n24846) );
  sky130_fd_sc_hd__nand3_1 U24739 ( .A(n23220), .B(n24849), .C(n24846), .Y(
        n20749) );
  sky130_fd_sc_hd__nor2_1 U24740 ( .A(n24854), .B(n20749), .Y(n21504) );
  sky130_fd_sc_hd__nand2_1 U24741 ( .A(n21640), .B(n20333), .Y(n21473) );
  sky130_fd_sc_hd__nand2_1 U24742 ( .A(n21504), .B(n21473), .Y(n21411) );
  sky130_fd_sc_hd__nor4b_1 U24743 ( .D_N(n21556), .A(n21608), .B(n24830), .C(
        n21411), .Y(n20338) );
  sky130_fd_sc_hd__nor3_1 U24744 ( .A(n25380), .B(n21569), .C(n20742), .Y(
        n20764) );
  sky130_fd_sc_hd__o22ai_1 U24745 ( .A1(n21480), .A2(n22409), .B1(n21569), 
        .B2(n21474), .Y(n20334) );
  sky130_fd_sc_hd__a211oi_1 U24746 ( .A1(n21564), .A2(n21330), .B1(n20764), 
        .C1(n20334), .Y(n21507) );
  sky130_fd_sc_hd__nor3_1 U24747 ( .A(n20986), .B(n20983), .C(n22407), .Y(
        n20751) );
  sky130_fd_sc_hd__nor2_1 U24748 ( .A(n20335), .B(n20992), .Y(n21406) );
  sky130_fd_sc_hd__nor3_1 U24749 ( .A(n20751), .B(n21464), .C(n21406), .Y(
        n21594) );
  sky130_fd_sc_hd__nand2_1 U24750 ( .A(n22330), .B(n20336), .Y(n20975) );
  sky130_fd_sc_hd__nor2_1 U24751 ( .A(n21505), .B(n20975), .Y(n21510) );
  sky130_fd_sc_hd__a21oi_1 U24752 ( .A1(n24826), .A2(n24825), .B1(n21510), .Y(
        n21414) );
  sky130_fd_sc_hd__and3_1 U24753 ( .A(n21507), .B(n21594), .C(n21414), .X(
        n20337) );
  sky130_fd_sc_hd__nand2_1 U24754 ( .A(n20338), .B(n20337), .Y(n21543) );
  sky130_fd_sc_hd__nand3_1 U24755 ( .A(n22762), .B(n20761), .C(n20339), .Y(
        n20993) );
  sky130_fd_sc_hd__nand2_1 U24756 ( .A(n25387), .B(n20342), .Y(n21431) );
  sky130_fd_sc_hd__a21oi_1 U24757 ( .A1(n21522), .A2(n21431), .B1(n25369), .Y(
        n21426) );
  sky130_fd_sc_hd__o22ai_1 U24758 ( .A1(n24872), .A2(n20340), .B1(n21536), 
        .B2(n25387), .Y(n21438) );
  sky130_fd_sc_hd__nor2_1 U24759 ( .A(n21426), .B(n21438), .Y(n21447) );
  sky130_fd_sc_hd__nand2_1 U24760 ( .A(n20750), .B(n21447), .Y(n21643) );
  sky130_fd_sc_hd__nand3_1 U24761 ( .A(n24826), .B(n25369), .C(n25387), .Y(
        n20977) );
  sky130_fd_sc_hd__o21ai_1 U24762 ( .A1(n24869), .A2(n22419), .B1(n20977), .Y(
        n21494) );
  sky130_fd_sc_hd__nand3_1 U24763 ( .A(n22762), .B(n20761), .C(n24825), .Y(
        n21417) );
  sky130_fd_sc_hd__nor2_1 U24764 ( .A(n21734), .B(n20341), .Y(n21519) );
  sky130_fd_sc_hd__a21oi_1 U24765 ( .A1(n20342), .A2(n25369), .B1(n21519), .Y(
        n21432) );
  sky130_fd_sc_hd__nor4_1 U24767 ( .A(n21543), .B(n21643), .C(n21494), .D(
        n24832), .Y(n20344) );
  sky130_fd_sc_hd__nand4_1 U24768 ( .A(n21800), .B(n21580), .C(n20345), .D(
        n20344), .Y(n20346) );
  sky130_fd_sc_hd__nand2_1 U24769 ( .A(n20346), .B(n24858), .Y(n20351) );
  sky130_fd_sc_hd__nand2_1 U24770 ( .A(n24879), .B(n24897), .Y(n24844) );
  sky130_fd_sc_hd__nor3_1 U24771 ( .A(j202_soc_core_j22_cpu_opst[1]), .B(
        j202_soc_core_j22_cpu_opst[4]), .C(n20773), .Y(n20501) );
  sky130_fd_sc_hd__nand2_1 U24772 ( .A(n21604), .B(n20501), .Y(n21339) );
  sky130_fd_sc_hd__nand2_1 U24773 ( .A(n24879), .B(n20347), .Y(n24874) );
  sky130_fd_sc_hd__nand2_1 U24774 ( .A(j202_soc_core_j22_cpu_opst[0]), .B(
        n20348), .Y(n21395) );
  sky130_fd_sc_hd__nor2_1 U24775 ( .A(n21441), .B(n21395), .Y(n21527) );
  sky130_fd_sc_hd__nand2_1 U24776 ( .A(n24879), .B(n21527), .Y(n22339) );
  sky130_fd_sc_hd__nand2_1 U24777 ( .A(n24874), .B(n22339), .Y(n24835) );
  sky130_fd_sc_hd__nor3_1 U24778 ( .A(n24888), .B(n24863), .C(n24835), .Y(
        n20349) );
  sky130_fd_sc_hd__nor2_1 U24779 ( .A(n22551), .B(n22525), .Y(n20356) );
  sky130_fd_sc_hd__nand2b_1 U24780 ( .A_N(n20353), .B(n20352), .Y(n20354) );
  sky130_fd_sc_hd__nand2_1 U24781 ( .A(n22073), .B(n21178), .Y(n20381) );
  sky130_fd_sc_hd__o21a_1 U24782 ( .A1(n21150), .A2(n22074), .B1(n20905), .X(
        n20358) );
  sky130_fd_sc_hd__nand2_1 U24783 ( .A(n23335), .B(n20904), .Y(n20357) );
  sky130_fd_sc_hd__o211ai_1 U24784 ( .A1(n21091), .A2(n23335), .B1(n20358), 
        .C1(n20357), .Y(n20377) );
  sky130_fd_sc_hd__nand2_1 U24785 ( .A(n20955), .B(n20904), .Y(n20359) );
  sky130_fd_sc_hd__a21o_1 U24786 ( .A1(n21010), .A2(n20359), .B1(n23335), .X(
        n20375) );
  sky130_fd_sc_hd__o22ai_1 U24787 ( .A1(n21145), .A2(n23333), .B1(n22610), 
        .B2(n21155), .Y(n20363) );
  sky130_fd_sc_hd__nand2_1 U24788 ( .A(n22592), .B(n22705), .Y(n21116) );
  sky130_fd_sc_hd__o22ai_1 U24789 ( .A1(n22641), .A2(n21116), .B1(n21048), 
        .B2(n21154), .Y(n20362) );
  sky130_fd_sc_hd__nand2_1 U24790 ( .A(n20360), .B(n22592), .Y(n21158) );
  sky130_fd_sc_hd__xor2_1 U24791 ( .A(n22631), .B(n22074), .X(n22449) );
  sky130_fd_sc_hd__o22ai_1 U24792 ( .A1(n22560), .A2(n21158), .B1(n21108), 
        .B2(n22449), .Y(n20361) );
  sky130_fd_sc_hd__nor3_1 U24793 ( .A(n20363), .B(n20362), .C(n20361), .Y(
        n20374) );
  sky130_fd_sc_hd__nand2_1 U24794 ( .A(n20364), .B(n21017), .Y(n20838) );
  sky130_fd_sc_hd__nand2_1 U24795 ( .A(n20838), .B(n21139), .Y(n21167) );
  sky130_fd_sc_hd__nor2_1 U24796 ( .A(n22064), .B(n21167), .Y(n20369) );
  sky130_fd_sc_hd__nand2_1 U24797 ( .A(n21164), .B(n22573), .Y(n20367) );
  sky130_fd_sc_hd__nand4_1 U24798 ( .A(n20649), .B(n22141), .C(n22704), .D(
        n21019), .Y(n20531) );
  sky130_fd_sc_hd__nand3_1 U24799 ( .A(n20365), .B(n22154), .C(n22141), .Y(
        n20366) );
  sky130_fd_sc_hd__nand2_1 U24800 ( .A(n20531), .B(n20366), .Y(n20833) );
  sky130_fd_sc_hd__nand2_1 U24801 ( .A(n20833), .B(n21139), .Y(n21166) );
  sky130_fd_sc_hd__o211ai_1 U24802 ( .A1(n22604), .A2(n21163), .B1(n20367), 
        .C1(n21166), .Y(n20368) );
  sky130_fd_sc_hd__nor2_1 U24803 ( .A(n20369), .B(n20368), .Y(n20373) );
  sky130_fd_sc_hd__nand2_1 U24804 ( .A(n20371), .B(n20370), .Y(n20834) );
  sky130_fd_sc_hd__nand2_1 U24805 ( .A(n20834), .B(n21139), .Y(n21085) );
  sky130_fd_sc_hd__nand2_1 U24806 ( .A(n21144), .B(n23333), .Y(n20372) );
  sky130_fd_sc_hd__nand4_1 U24807 ( .A(n20375), .B(n20374), .C(n20373), .D(
        n20372), .Y(n20376) );
  sky130_fd_sc_hd__a21oi_1 U24808 ( .A1(n20377), .A2(n22631), .B1(n20376), .Y(
        n20380) );
  sky130_fd_sc_hd__nand2_1 U24809 ( .A(n20378), .B(n21137), .Y(n20379) );
  sky130_fd_sc_hd__nand2_1 U24810 ( .A(n21984), .B(n21178), .Y(n20405) );
  sky130_fd_sc_hd__nor2_1 U24811 ( .A(n21048), .B(n23338), .Y(n20396) );
  sky130_fd_sc_hd__nand2_1 U24812 ( .A(n20383), .B(n21139), .Y(n20384) );
  sky130_fd_sc_hd__nand2_1 U24813 ( .A(n20384), .B(n21141), .Y(n20401) );
  sky130_fd_sc_hd__a21oi_1 U24814 ( .A1(n23338), .A2(n21048), .B1(n21143), .Y(
        n20400) );
  sky130_fd_sc_hd__nand2_1 U24815 ( .A(n21118), .B(n22591), .Y(n20391) );
  sky130_fd_sc_hd__nand2b_1 U24816 ( .A_N(n21985), .B(n22575), .Y(n22633) );
  sky130_fd_sc_hd__a22oi_1 U24817 ( .A1(n22575), .A2(n21146), .B1(n21985), 
        .B2(n20385), .Y(n20387) );
  sky130_fd_sc_hd__nand2_1 U24818 ( .A(n21048), .B(n21985), .Y(n22452) );
  sky130_fd_sc_hd__nand3_1 U24819 ( .A(n22633), .B(n22452), .C(n21147), .Y(
        n20386) );
  sky130_fd_sc_hd__o211ai_1 U24820 ( .A1(n21150), .A2(n22633), .B1(n20387), 
        .C1(n20386), .Y(n20389) );
  sky130_fd_sc_hd__o22ai_1 U24821 ( .A1(n20955), .A2(n21155), .B1(n22604), 
        .B2(n21154), .Y(n20388) );
  sky130_fd_sc_hd__nor2_1 U24822 ( .A(n20389), .B(n20388), .Y(n20390) );
  sky130_fd_sc_hd__o211ai_1 U24823 ( .A1(n21985), .A2(n21085), .B1(n20391), 
        .C1(n20390), .Y(n20395) );
  sky130_fd_sc_hd__o22ai_1 U24824 ( .A1(n22600), .A2(n21116), .B1(n22561), 
        .B2(n21158), .Y(n20392) );
  sky130_fd_sc_hd__a21oi_1 U24825 ( .A1(n21164), .A2(n22576), .B1(n20392), .Y(
        n20393) );
  sky130_fd_sc_hd__o211ai_1 U24826 ( .A1(n22300), .A2(n21167), .B1(n21166), 
        .C1(n20393), .Y(n20394) );
  sky130_fd_sc_hd__nor2_1 U24827 ( .A(n20395), .B(n20394), .Y(n20398) );
  sky130_fd_sc_hd__nand2_1 U24828 ( .A(n20396), .B(n21170), .Y(n20397) );
  sky130_fd_sc_hd__o211ai_1 U24829 ( .A1(n23338), .A2(n21174), .B1(n20398), 
        .C1(n20397), .Y(n20399) );
  sky130_fd_sc_hd__a21oi_1 U24830 ( .A1(n20401), .A2(n20400), .B1(n20399), .Y(
        n20404) );
  sky130_fd_sc_hd__nand2_1 U24831 ( .A(n20402), .B(n21137), .Y(n20403) );
  sky130_fd_sc_hd__nand2_1 U24832 ( .A(n20407), .B(n21137), .Y(n20428) );
  sky130_fd_sc_hd__a21oi_1 U24833 ( .A1(n23312), .A2(n22641), .B1(n21143), .Y(
        n20425) );
  sky130_fd_sc_hd__nand2_1 U24835 ( .A(n20408), .B(n21141), .Y(n20424) );
  sky130_fd_sc_hd__xnor2_1 U24836 ( .A(n22577), .B(n23310), .Y(n22466) );
  sky130_fd_sc_hd__clkinv_1 U24837 ( .A(n22466), .Y(n20411) );
  sky130_fd_sc_hd__o22ai_1 U24838 ( .A1(n21145), .A2(n23310), .B1(n22643), 
        .B2(n21155), .Y(n20410) );
  sky130_fd_sc_hd__a21oi_1 U24839 ( .A1(n20411), .A2(n21147), .B1(n20410), .Y(
        n20415) );
  sky130_fd_sc_hd__o22ai_1 U24840 ( .A1(n22560), .A2(n21116), .B1(n22647), 
        .B2(n21158), .Y(n20413) );
  sky130_fd_sc_hd__o2bb2ai_1 U24841 ( .B1(n22600), .B2(n21154), .A1_N(n21156), 
        .A2_N(n22631), .Y(n20412) );
  sky130_fd_sc_hd__nor2_1 U24842 ( .A(n20413), .B(n20412), .Y(n20414) );
  sky130_fd_sc_hd__o211ai_1 U24843 ( .A1(n22640), .A2(n21085), .B1(n20415), 
        .C1(n20414), .Y(n20418) );
  sky130_fd_sc_hd__a2bb2oi_1 U24844 ( .B1(n21775), .B2(n21164), .A1_N(n22567), 
        .A2_N(n21163), .Y(n20416) );
  sky130_fd_sc_hd__o211ai_1 U24845 ( .A1(n22646), .A2(n21167), .B1(n21166), 
        .C1(n20416), .Y(n20417) );
  sky130_fd_sc_hd__nor2_1 U24846 ( .A(n20418), .B(n20417), .Y(n20422) );
  sky130_fd_sc_hd__a21oi_1 U24847 ( .A1(n23310), .A2(n21089), .B1(n21146), .Y(
        n20419) );
  sky130_fd_sc_hd__nand2_1 U24849 ( .A(n20420), .B(n22577), .Y(n20421) );
  sky130_fd_sc_hd__o211ai_1 U24850 ( .A1(n23312), .A2(n21174), .B1(n20422), 
        .C1(n20421), .Y(n20423) );
  sky130_fd_sc_hd__a21oi_1 U24851 ( .A1(n20425), .A2(n20424), .B1(n20423), .Y(
        n20427) );
  sky130_fd_sc_hd__nand2_1 U24852 ( .A(n22020), .B(n21178), .Y(n20426) );
  sky130_fd_sc_hd__nand2_1 U24853 ( .A(j202_soc_core_uart_TOP_load), .B(
        j202_soc_core_uart_sio_ce), .Y(n25122) );
  sky130_fd_sc_hd__nor2_1 U24854 ( .A(n25123), .B(n25122), .Y(n25121) );
  sky130_fd_sc_hd__o2bb2ai_1 U24855 ( .B1(n23831), .B2(n25121), .A1_N(n23831), 
        .A2_N(n25121), .Y(n22) );
  sky130_fd_sc_hd__clkinv_1 U24856 ( .A(n23254), .Y(j202_soc_core_uart_N5) );
  sky130_fd_sc_hd__clkinv_1 U24857 ( .A(n25406), .Y(n25244) );
  sky130_fd_sc_hd__o2bb2ai_1 U24858 ( .B1(n25244), .B2(n20429), .A1_N(n25244), 
        .A2_N(j202_soc_core_bldc_core_00_hall_value[1]), .Y(n136) );
  sky130_fd_sc_hd__and3b_1 U24859 ( .B(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[1]), .C(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_addr_1[2]), .A_N(
        j202_soc_core_bldc_core_00_bldc_wb_slave_00_state[0]), .X(n25164) );
  sky130_fd_sc_hd__nand2_1 U24860 ( .A(n20430), .B(n25164), .Y(n25158) );
  sky130_fd_sc_hd__clkinv_1 U24861 ( .A(j202_soc_core_bldc_core_00_wdata[0]), 
        .Y(n25171) );
  sky130_fd_sc_hd__o2bb2ai_1 U24862 ( .B1(n25158), .B2(n25171), .A1_N(n25158), 
        .A2_N(j202_soc_core_bldc_core_00_pwm_en), .Y(n48) );
  sky130_fd_sc_hd__nand3_1 U24863 ( .A(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[1]), .B(
        j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen_2), .C(n20431), .Y(n23103) );
  sky130_fd_sc_hd__or4_1 U24864 ( .A(j202_soc_core_cmt_core_00_reg_addr[1]), 
        .B(j202_soc_core_cmt_core_00_reg_addr[0]), .C(
        j202_soc_core_cmt_core_00_reg_addr[6]), .D(
        j202_soc_core_cmt_core_00_reg_addr[7]), .X(n20432) );
  sky130_fd_sc_hd__nor2_1 U24865 ( .A(j202_soc_core_cmt_core_00_reg_addr[5]), 
        .B(n20432), .Y(n22968) );
  sky130_fd_sc_hd__clkinv_1 U24866 ( .A(j202_soc_core_cmt_core_00_reg_addr[4]), 
        .Y(n22967) );
  sky130_fd_sc_hd__nand2_1 U24867 ( .A(n22968), .B(n22967), .Y(n20433) );
  sky130_fd_sc_hd__nor2_1 U24868 ( .A(n23103), .B(n20433), .Y(n20436) );
  sky130_fd_sc_hd__clkinv_1 U24869 ( .A(n20436), .Y(n20435) );
  sky130_fd_sc_hd__nand2b_1 U24870 ( .A_N(
        j202_soc_core_cmt_core_00_reg_addr[3]), .B(
        j202_soc_core_cmt_core_00_reg_addr[2]), .Y(n22971) );
  sky130_fd_sc_hd__nor2_1 U24871 ( .A(n20435), .B(n22971), .Y(n25240) );
  sky130_fd_sc_hd__clkinv_1 U24872 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[3]), .Y(n25220) );
  sky130_fd_sc_hd__o2bb2ai_1 U24873 ( .B1(n25239), .B2(n25220), .A1_N(n25239), 
        .A2_N(j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[3]), .Y(n112) );
  sky130_fd_sc_hd__clkinv_1 U24874 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[5]), .Y(n25210) );
  sky130_fd_sc_hd__o2bb2ai_1 U24875 ( .B1(n25239), .B2(n25210), .A1_N(n25239), 
        .A2_N(j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[5]), .Y(n99) );
  sky130_fd_sc_hd__clkinv_1 U24876 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[2]), .Y(n25195) );
  sky130_fd_sc_hd__o2bb2ai_1 U24877 ( .B1(n25239), .B2(n25195), .A1_N(n25239), 
        .A2_N(j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[2]), .Y(n75) );
  sky130_fd_sc_hd__clkinv_1 U24878 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[1]), .Y(n25154) );
  sky130_fd_sc_hd__o2bb2ai_1 U24879 ( .B1(n25239), .B2(n25154), .A1_N(n25239), 
        .A2_N(j202_soc_core_cmt_core_00_cks0[1]), .Y(n33) );
  sky130_fd_sc_hd__clkinv_1 U24880 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[4]), .Y(n25207) );
  sky130_fd_sc_hd__o2bb2ai_1 U24881 ( .B1(n25239), .B2(n25207), .A1_N(n25239), 
        .A2_N(j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[4]), .Y(n95) );
  sky130_fd_sc_hd__clkinv_1 U24882 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[0]), .Y(n25198) );
  sky130_fd_sc_hd__o2bb2ai_1 U24883 ( .B1(n25239), .B2(n25198), .A1_N(n25239), 
        .A2_N(j202_soc_core_cmt_core_00_cks0[0]), .Y(n81) );
  sky130_fd_sc_hd__or3_1 U24884 ( .A(j202_soc_core_cmt_core_00_reg_addr[3]), 
        .B(j202_soc_core_cmt_core_00_reg_addr[2]), .C(n20435), .X(n20434) );
  sky130_fd_sc_hd__o2bb2ai_1 U24885 ( .B1(n20434), .B2(n25154), .A1_N(n20434), 
        .A2_N(j202_soc_core_cmt_core_00_str1), .Y(n32) );
  sky130_fd_sc_hd__o2bb2ai_1 U24886 ( .B1(n20434), .B2(n25198), .A1_N(n20434), 
        .A2_N(j202_soc_core_cmt_core_00_str0), .Y(n80) );
  sky130_fd_sc_hd__nand2b_1 U24887 ( .A_N(
        j202_soc_core_cmt_core_00_reg_addr[2]), .B(
        j202_soc_core_cmt_core_00_reg_addr[3]), .Y(n22975) );
  sky130_fd_sc_hd__nor2_1 U24888 ( .A(n20435), .B(n22975), .Y(n25213) );
  sky130_fd_sc_hd__o2bb2ai_1 U24889 ( .B1(n25212), .B2(n25210), .A1_N(n25212), 
        .A2_N(j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[5]), .Y(n100) );
  sky130_fd_sc_hd__o2bb2ai_1 U24890 ( .B1(n25212), .B2(n25207), .A1_N(n25212), 
        .A2_N(j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[4]), .Y(n96) );
  sky130_fd_sc_hd__o2bb2ai_1 U24891 ( .B1(n25212), .B2(n25195), .A1_N(n25212), 
        .A2_N(j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[2]), .Y(n76) );
  sky130_fd_sc_hd__o2bb2ai_1 U24892 ( .B1(n25212), .B2(n25220), .A1_N(n25212), 
        .A2_N(j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[3]), .Y(n113) );
  sky130_fd_sc_hd__o2bb2ai_1 U24893 ( .B1(n25212), .B2(n25154), .A1_N(n25212), 
        .A2_N(j202_soc_core_cmt_core_00_cks1[1]), .Y(n34) );
  sky130_fd_sc_hd__clkinv_1 U24894 ( .A(j202_soc_core_cmt_core_00_cnt0[11]), 
        .Y(n20468) );
  sky130_fd_sc_hd__clkinv_1 U24895 ( .A(j202_soc_core_cmt_core_00_cnt0[9]), 
        .Y(n23079) );
  sky130_fd_sc_hd__nand3_1 U24896 ( .A(n20436), .B(
        j202_soc_core_cmt_core_00_reg_addr[3]), .C(
        j202_soc_core_cmt_core_00_reg_addr[2]), .Y(n23101) );
  sky130_fd_sc_hd__clkinv_1 U24897 ( .A(j202_soc_core_cmt_core_00_cnt0[13]), 
        .Y(n20438) );
  sky130_fd_sc_hd__clkinv_1 U24898 ( .A(j202_soc_core_cmt_core_00_cnt0[7]), 
        .Y(n23067) );
  sky130_fd_sc_hd__o22ai_1 U24899 ( .A1(n20438), .A2(
        j202_soc_core_cmt_core_00_const0[13]), .B1(n23067), .B2(
        j202_soc_core_cmt_core_00_const0[7]), .Y(n20437) );
  sky130_fd_sc_hd__a221oi_1 U24900 ( .A1(n20438), .A2(
        j202_soc_core_cmt_core_00_const0[13]), .B1(
        j202_soc_core_cmt_core_00_const0[7]), .B2(n23067), .C1(n20437), .Y(
        n20458) );
  sky130_fd_sc_hd__clkinv_1 U24901 ( .A(j202_soc_core_cmt_core_00_cnt0[14]), 
        .Y(n23095) );
  sky130_fd_sc_hd__o22ai_1 U24902 ( .A1(n20468), .A2(
        j202_soc_core_cmt_core_00_const0[11]), .B1(n23095), .B2(
        j202_soc_core_cmt_core_00_const0[14]), .Y(n20439) );
  sky130_fd_sc_hd__a221oi_1 U24903 ( .A1(n20468), .A2(
        j202_soc_core_cmt_core_00_const0[11]), .B1(
        j202_soc_core_cmt_core_00_const0[14]), .B2(n23095), .C1(n20439), .Y(
        n20457) );
  sky130_fd_sc_hd__clkinv_1 U24904 ( .A(j202_soc_core_cmt_core_00_cnt0[3]), 
        .Y(n20493) );
  sky130_fd_sc_hd__clkinv_1 U24905 ( .A(j202_soc_core_cmt_core_00_const0[3]), 
        .Y(n25219) );
  sky130_fd_sc_hd__o22ai_1 U24906 ( .A1(j202_soc_core_cmt_core_00_const0[3]), 
        .A2(n20493), .B1(n25219), .B2(j202_soc_core_cmt_core_00_cnt0[3]), .Y(
        n20455) );
  sky130_fd_sc_hd__clkinv_1 U24907 ( .A(j202_soc_core_cmt_core_00_cnt0[6]), 
        .Y(n23063) );
  sky130_fd_sc_hd__clkinv_1 U24908 ( .A(j202_soc_core_cmt_core_00_const0[6]), 
        .Y(n25214) );
  sky130_fd_sc_hd__clkinv_1 U24909 ( .A(j202_soc_core_cmt_core_00_const0[8]), 
        .Y(n25222) );
  sky130_fd_sc_hd__clkinv_1 U24910 ( .A(j202_soc_core_cmt_core_00_const0[4]), 
        .Y(n25208) );
  sky130_fd_sc_hd__o22ai_1 U24911 ( .A1(n25222), .A2(
        j202_soc_core_cmt_core_00_cnt0[8]), .B1(n25208), .B2(
        j202_soc_core_cmt_core_00_cnt0[4]), .Y(n20440) );
  sky130_fd_sc_hd__a221oi_1 U24912 ( .A1(n25222), .A2(
        j202_soc_core_cmt_core_00_cnt0[8]), .B1(
        j202_soc_core_cmt_core_00_cnt0[4]), .B2(n25208), .C1(n20440), .Y(
        n20441) );
  sky130_fd_sc_hd__o221ai_1 U24913 ( .A1(j202_soc_core_cmt_core_00_const0[6]), 
        .A2(n23063), .B1(n25214), .B2(j202_soc_core_cmt_core_00_cnt0[6]), .C1(
        n20441), .Y(n20454) );
  sky130_fd_sc_hd__clkinv_1 U24914 ( .A(j202_soc_core_cmt_core_00_cnt0[12]), 
        .Y(n23084) );
  sky130_fd_sc_hd__clkinv_1 U24915 ( .A(j202_soc_core_cmt_core_00_cnt0[2]), 
        .Y(n23057) );
  sky130_fd_sc_hd__o22ai_1 U24916 ( .A1(n23084), .A2(
        j202_soc_core_cmt_core_00_const0[12]), .B1(n23057), .B2(
        j202_soc_core_cmt_core_00_const0[2]), .Y(n20442) );
  sky130_fd_sc_hd__a221oi_1 U24917 ( .A1(n23084), .A2(
        j202_soc_core_cmt_core_00_const0[12]), .B1(
        j202_soc_core_cmt_core_00_const0[2]), .B2(n23057), .C1(n20442), .Y(
        n20452) );
  sky130_fd_sc_hd__clkinv_1 U24918 ( .A(j202_soc_core_cmt_core_00_cnt0[15]), 
        .Y(n20444) );
  sky130_fd_sc_hd__clkinv_1 U24919 ( .A(j202_soc_core_cmt_core_00_const0[0]), 
        .Y(n25197) );
  sky130_fd_sc_hd__o22ai_1 U24920 ( .A1(n20444), .A2(
        j202_soc_core_cmt_core_00_const0[15]), .B1(n25197), .B2(
        j202_soc_core_cmt_core_00_cnt0[0]), .Y(n20443) );
  sky130_fd_sc_hd__a221oi_1 U24921 ( .A1(n20444), .A2(
        j202_soc_core_cmt_core_00_const0[15]), .B1(
        j202_soc_core_cmt_core_00_cnt0[0]), .B2(n25197), .C1(n20443), .Y(
        n20451) );
  sky130_fd_sc_hd__clkinv_1 U24922 ( .A(j202_soc_core_cmt_core_00_cnt0[10]), 
        .Y(n20447) );
  sky130_fd_sc_hd__clkinv_1 U24923 ( .A(j202_soc_core_cmt_core_00_cnt0[1]), 
        .Y(n20446) );
  sky130_fd_sc_hd__o22ai_1 U24924 ( .A1(n20447), .A2(
        j202_soc_core_cmt_core_00_const0[10]), .B1(n20446), .B2(
        j202_soc_core_cmt_core_00_const0[1]), .Y(n20445) );
  sky130_fd_sc_hd__a221oi_1 U24925 ( .A1(n20447), .A2(
        j202_soc_core_cmt_core_00_const0[10]), .B1(
        j202_soc_core_cmt_core_00_const0[1]), .B2(n20446), .C1(n20445), .Y(
        n20450) );
  sky130_fd_sc_hd__clkinv_1 U24926 ( .A(j202_soc_core_cmt_core_00_const0[5]), 
        .Y(n25209) );
  sky130_fd_sc_hd__o22ai_1 U24927 ( .A1(n23079), .A2(
        j202_soc_core_cmt_core_00_const0[9]), .B1(n25209), .B2(
        j202_soc_core_cmt_core_00_cnt0[5]), .Y(n20448) );
  sky130_fd_sc_hd__a221oi_1 U24928 ( .A1(n23079), .A2(
        j202_soc_core_cmt_core_00_const0[9]), .B1(
        j202_soc_core_cmt_core_00_cnt0[5]), .B2(n25209), .C1(n20448), .Y(
        n20449) );
  sky130_fd_sc_hd__nand4_1 U24929 ( .A(n20452), .B(n20451), .C(n20450), .D(
        n20449), .Y(n20453) );
  sky130_fd_sc_hd__nor3_1 U24930 ( .A(n20455), .B(n20454), .C(n20453), .Y(
        n20456) );
  sky130_fd_sc_hd__nand3_1 U24931 ( .A(n20458), .B(n20457), .C(n20456), .Y(
        n23049) );
  sky130_fd_sc_hd__nand2_1 U24932 ( .A(n23101), .B(n23049), .Y(n20471) );
  sky130_fd_sc_hd__clkinv_1 U24933 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[9]), .Y(n23045) );
  sky130_fd_sc_hd__clkinv_1 U24934 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[7]), .Y(n23040) );
  sky130_fd_sc_hd__nor3_1 U24935 ( .A(j202_soc_core_cmt_core_00_cks0[1]), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[5]), .C(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[3]), .Y(n20459) );
  sky130_fd_sc_hd__a31oi_1 U24936 ( .A1(j202_soc_core_cmt_core_00_cks0[1]), 
        .A2(n23045), .A3(n23040), .B1(n20459), .Y(n20466) );
  sky130_fd_sc_hd__nor4_1 U24937 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[8]), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[2]), .C(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[0]), .D(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[1]), .Y(n20465) );
  sky130_fd_sc_hd__clkinv_1 U24938 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[5]), .Y(n23036) );
  sky130_fd_sc_hd__a21oi_1 U24939 ( .A1(j202_soc_core_cmt_core_00_cks0[0]), 
        .A2(n23045), .B1(n23036), .Y(n20463) );
  sky130_fd_sc_hd__a21oi_1 U24940 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[7]), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[3]), .B1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[9]), .Y(n20461) );
  sky130_fd_sc_hd__nor4_1 U24943 ( .A(n20463), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[4]), .C(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[6]), .D(n20462), .Y(
        n20464) );
  sky130_fd_sc_hd__nand3_1 U24944 ( .A(n20466), .B(n20465), .C(n20464), .Y(
        n20470) );
  sky130_fd_sc_hd__nor2_1 U24945 ( .A(n20471), .B(n20470), .Y(n23046) );
  sky130_fd_sc_hd__clkinv_1 U24946 ( .A(j202_soc_core_cmt_core_00_cnt0[8]), 
        .Y(n23077) );
  sky130_fd_sc_hd__nand2_1 U24947 ( .A(j202_soc_core_cmt_core_00_cnt0[0]), .B(
        j202_soc_core_cmt_core_00_cnt0[1]), .Y(n23054) );
  sky130_fd_sc_hd__nor2_1 U24948 ( .A(n23057), .B(n23054), .Y(n23053) );
  sky130_fd_sc_hd__and3_1 U24949 ( .A(j202_soc_core_cmt_core_00_cnt0[6]), .B(
        j202_soc_core_cmt_core_00_cnt0[4]), .C(
        j202_soc_core_cmt_core_00_cnt0[5]), .X(n20467) );
  sky130_fd_sc_hd__nand4_1 U24950 ( .A(j202_soc_core_cmt_core_00_cnt0[7]), .B(
        j202_soc_core_cmt_core_00_cnt0[3]), .C(n23053), .D(n20467), .Y(n23072)
         );
  sky130_fd_sc_hd__nor2_1 U24951 ( .A(n23077), .B(n23072), .Y(n23071) );
  sky130_fd_sc_hd__nand2_1 U24952 ( .A(n23046), .B(n23071), .Y(n23078) );
  sky130_fd_sc_hd__nor2_1 U24953 ( .A(n23079), .B(n23078), .Y(n23081) );
  sky130_fd_sc_hd__nand2_1 U24954 ( .A(j202_soc_core_cmt_core_00_cnt0[10]), 
        .B(n23081), .Y(n20469) );
  sky130_fd_sc_hd__nor2_1 U24955 ( .A(n20468), .B(n20469), .Y(n23085) );
  sky130_fd_sc_hd__clkinv_1 U24956 ( .A(n20469), .Y(n23083) );
  sky130_fd_sc_hd__nand2_1 U24957 ( .A(n23101), .B(n20470), .Y(n23076) );
  sky130_fd_sc_hd__nand2_1 U24958 ( .A(n20471), .B(n23076), .Y(n23086) );
  sky130_fd_sc_hd__o21ai_1 U24959 ( .A1(j202_soc_core_cmt_core_00_cnt0[11]), 
        .A2(n23083), .B1(n23086), .Y(n20472) );
  sky130_fd_sc_hd__clkinv_1 U24960 ( .A(n23101), .Y(n23074) );
  sky130_fd_sc_hd__o2bb2ai_1 U24961 ( .B1(n23085), .B2(n20472), .A1_N(n23074), 
        .A2_N(j202_soc_core_cmt_core_00_wdata_cnt0[11]), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[11]) );
  sky130_fd_sc_hd__nand2_1 U24962 ( .A(j202_soc_core_cmt_core_00_reg_addr[4]), 
        .B(n22968), .Y(n22972) );
  sky130_fd_sc_hd__nor3_1 U24963 ( .A(n23103), .B(n22972), .C(n22971), .Y(
        n25230) );
  sky130_fd_sc_hd__o2bb2ai_1 U24964 ( .B1(n25229), .B2(n25195), .A1_N(n25229), 
        .A2_N(j202_soc_core_cmt_core_00_const0[2]), .Y(n77) );
  sky130_fd_sc_hd__clkinv_1 U24965 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[13]), .Y(n23091) );
  sky130_fd_sc_hd__o2bb2ai_1 U24966 ( .B1(n25229), .B2(n23091), .A1_N(n25229), 
        .A2_N(j202_soc_core_cmt_core_00_const0[13]), .Y(n128) );
  sky130_fd_sc_hd__clkinv_1 U24967 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[9]), .Y(n25150) );
  sky130_fd_sc_hd__o2bb2ai_1 U24968 ( .B1(n25229), .B2(n25150), .A1_N(n25229), 
        .A2_N(j202_soc_core_cmt_core_00_const0[9]), .Y(n28) );
  sky130_fd_sc_hd__clkinv_1 U24969 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[15]), .Y(n23218) );
  sky130_fd_sc_hd__o2bb2ai_1 U24970 ( .B1(n25229), .B2(n23218), .A1_N(n25229), 
        .A2_N(j202_soc_core_cmt_core_00_const0[15]), .Y(n124) );
  sky130_fd_sc_hd__clkinv_1 U24971 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[12]), .Y(n23200) );
  sky130_fd_sc_hd__o2bb2ai_1 U24972 ( .B1(n25229), .B2(n23200), .A1_N(n25229), 
        .A2_N(j202_soc_core_cmt_core_00_const0[12]), .Y(n127) );
  sky130_fd_sc_hd__o2bb2ai_1 U24973 ( .B1(n25229), .B2(n25154), .A1_N(n25229), 
        .A2_N(j202_soc_core_cmt_core_00_const0[1]), .Y(n35) );
  sky130_fd_sc_hd__clkinv_1 U24974 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[10]), .Y(n25225) );
  sky130_fd_sc_hd__o2bb2ai_1 U24975 ( .B1(n25229), .B2(n25225), .A1_N(n25229), 
        .A2_N(j202_soc_core_cmt_core_00_const0[10]), .Y(n125) );
  sky130_fd_sc_hd__clkinv_1 U24976 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[14]), .Y(n23094) );
  sky130_fd_sc_hd__o2bb2ai_1 U24977 ( .B1(n25229), .B2(n23094), .A1_N(n25229), 
        .A2_N(j202_soc_core_cmt_core_00_const0[14]), .Y(n129) );
  sky130_fd_sc_hd__clkinv_1 U24978 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[7]), .Y(n25217) );
  sky130_fd_sc_hd__o2bb2ai_1 U24979 ( .B1(n25229), .B2(n25217), .A1_N(n25229), 
        .A2_N(j202_soc_core_cmt_core_00_const0[7]), .Y(n106) );
  sky130_fd_sc_hd__nor3_1 U24980 ( .A(n23103), .B(n22972), .C(n22975), .Y(
        n25228) );
  sky130_fd_sc_hd__o2bb2ai_1 U24981 ( .B1(n25227), .B2(n25207), .A1_N(n25227), 
        .A2_N(j202_soc_core_cmt_core_00_const1[4]), .Y(n98) );
  sky130_fd_sc_hd__o2bb2ai_1 U24982 ( .B1(n25227), .B2(n23200), .A1_N(n25227), 
        .A2_N(j202_soc_core_cmt_core_00_const1[12]), .Y(n121) );
  sky130_fd_sc_hd__o2bb2ai_1 U24983 ( .B1(n25227), .B2(n23091), .A1_N(n25227), 
        .A2_N(j202_soc_core_cmt_core_00_const1[13]), .Y(n122) );
  sky130_fd_sc_hd__o2bb2ai_1 U24984 ( .B1(n25227), .B2(n23094), .A1_N(n25227), 
        .A2_N(j202_soc_core_cmt_core_00_const1[14]), .Y(n123) );
  sky130_fd_sc_hd__o2bb2ai_1 U24985 ( .B1(n25227), .B2(n23218), .A1_N(n25227), 
        .A2_N(j202_soc_core_cmt_core_00_const1[15]), .Y(n118) );
  sky130_fd_sc_hd__o2bb2ai_1 U24986 ( .B1(n23990), .B2(n20473), .A1_N(n20475), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[21]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o2bb2ai_1 U24987 ( .B1(n23893), .B2(n20473), .A1_N(n20475), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[17]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o2bb2ai_1 U24988 ( .B1(n20474), .B2(n23990), .A1_N(n20477), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[29]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o2bb2ai_1 U24989 ( .B1(n20474), .B2(n24015), .A1_N(n20477), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[30]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o2bb2ai_1 U24990 ( .B1(n20474), .B2(n23893), .A1_N(n20477), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[25]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__nand2_1 U24991 ( .A(n24579), .B(n24453), .Y(n24496) );
  sky130_fd_sc_hd__nor2_1 U24992 ( .A(n24447), .B(n24496), .Y(n24289) );
  sky130_fd_sc_hd__nor2_1 U24993 ( .A(j202_soc_core_rst), .B(n24289), .Y(
        n24288) );
  sky130_fd_sc_hd__o2bb2ai_1 U24994 ( .B1(n23990), .B2(n24288), .A1_N(n20497), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[13]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o2bb2ai_1 U24995 ( .B1(n23940), .B2(n24288), .A1_N(n20497), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[11]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o2bb2ai_1 U24996 ( .B1(n23893), .B2(n24288), .A1_N(n20497), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[9]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o2bb2ai_1 U24997 ( .B1(n24015), .B2(n24288), .A1_N(n20497), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[14]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o2bb2ai_1 U24998 ( .B1(n23918), .B2(n24288), .A1_N(n20497), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[10]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o2bb2ai_1 U24999 ( .B1(n23965), .B2(n24288), .A1_N(n20497), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[12]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o2bb2ai_1 U25000 ( .B1(n24043), .B2(n24288), .A1_N(n20497), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[15]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o2bb2ai_1 U25001 ( .B1(n23868), .B2(n24288), .A1_N(n20497), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[8]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o2bb2ai_1 U25002 ( .B1(n24387), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[45]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o2bb2ai_1 U25003 ( .B1(n24430), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[75]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o2bb2ai_1 U25004 ( .B1(n24477), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[72]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o2bb2ai_1 U25005 ( .B1(n24428), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[43]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o2bb2ai_1 U25006 ( .B1(n24436), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[44]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o2bb2ai_1 U25007 ( .B1(n24405), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[111]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__o2bb2ai_1 U25008 ( .B1(n24479), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[104]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o2bb2ai_1 U25009 ( .B1(n24422), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[74]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o2bb2ai_1 U25010 ( .B1(n24475), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[40]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o2bb2ai_1 U25011 ( .B1(n24395), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[78]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o2bb2ai_1 U25012 ( .B1(n24438), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[76]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o2bb2ai_1 U25013 ( .B1(n24432), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[107]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o2bb2ai_1 U25014 ( .B1(n24483), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[41]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o2bb2ai_1 U25015 ( .B1(n24420), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[42]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o2bb2ai_1 U25016 ( .B1(n24402), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[79]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o2bb2ai_1 U25017 ( .B1(n24393), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[46]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o2bb2ai_1 U25018 ( .B1(n24397), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[110]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o2bb2ai_1 U25019 ( .B1(n24389), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[77]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o2bb2ai_1 U25020 ( .B1(n24390), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[109]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o2bb2ai_1 U25021 ( .B1(n24015), .B2(n20473), .A1_N(n20475), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[22]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o2bb2ai_1 U25022 ( .B1(n24043), .B2(n20473), .A1_N(n20475), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[23]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_2__rg_itgt_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o2bb2ai_1 U25023 ( .B1(n20474), .B2(n24043), .A1_N(n20477), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[31]), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__clkinv_1 U25024 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[29]), .Y(n23693) );
  sky130_fd_sc_hd__nand2_1 U25025 ( .A(n23740), .B(
        j202_soc_core_wbqspiflash_00_spi_spd), .Y(n23738) );
  sky130_fd_sc_hd__o2bb2ai_1 U25026 ( .B1(n23693), .B2(n23738), .A1_N(n23732), 
        .A2_N(j202_soc_core_wbqspiflash_00_lldriver_r_word[29]), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N317) );
  sky130_fd_sc_hd__nand2_1 U25027 ( .A(n21324), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd), .Y(n23588) );
  sky130_fd_sc_hd__clkinv_1 U25028 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_dir), .Y(n20476) );
  sky130_fd_sc_hd__o2bb2ai_1 U25029 ( .B1(n23588), .B2(n20476), .A1_N(n23689), 
        .A2_N(j202_soc_core_wbqspiflash_00_spi_dir), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N355) );
  sky130_fd_sc_hd__o2bb2ai_1 U25030 ( .B1(n20477), .B2(n24400), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[63]), .A2_N(n20474), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_3__rg_itgt_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o2bb2ai_1 U25031 ( .B1(n24400), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[47]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__nand2_1 U25032 ( .A(n20478), .B(
        j202_soc_core_j22_cpu_regop_We__0_), .Y(n20480) );
  sky130_fd_sc_hd__nor2_1 U25033 ( .A(n20480), .B(n20479), .Y(n22722) );
  sky130_fd_sc_hd__nand2_1 U25034 ( .A(n23239), .B(n22722), .Y(n22721) );
  sky130_fd_sc_hd__o21ai_1 U25035 ( .A1(n20482), .A2(n20481), .B1(n22721), .Y(
        j202_soc_core_j22_cpu_rf_N2627) );
  sky130_fd_sc_hd__nand2_1 U25036 ( .A(n20485), .B(n20484), .Y(n20486) );
  sky130_fd_sc_hd__nor3_1 U25037 ( .A(n20487), .B(n20486), .C(n21657), .Y(
        n21217) );
  sky130_fd_sc_hd__nand2_1 U25038 ( .A(n20488), .B(n25731), .Y(n10559) );
  sky130_fd_sc_hd__nor2_1 U25039 ( .A(n20489), .B(n11036), .Y(n20490) );
  sky130_fd_sc_hd__buf_4 U25040 ( .A(n20490), .X(n25506) );
  sky130_fd_sc_hd__o2bb2ai_1 U25043 ( .B1(n21191), .B2(n23312), .A1_N(n21191), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N2700) );
  sky130_fd_sc_hd__o2bb2ai_1 U25044 ( .B1(n23312), .B2(n21197), .A1_N(n21216), 
        .A2_N(n22017), .Y(j202_soc_core_j22_cpu_rf_N3331) );
  sky130_fd_sc_hd__nand2_1 U25045 ( .A(n23046), .B(n23053), .Y(n20492) );
  sky130_fd_sc_hd__nor2_1 U25046 ( .A(n20493), .B(n20492), .Y(n23058) );
  sky130_fd_sc_hd__a21oi_1 U25047 ( .A1(n20493), .A2(n20492), .B1(n23058), .Y(
        n20494) );
  sky130_fd_sc_hd__o2bb2ai_1 U25048 ( .B1(n23101), .B2(n25220), .A1_N(n20494), 
        .A2_N(n23086), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[3])
         );
  sky130_fd_sc_hd__o2bb2ai_1 U25049 ( .B1(n25193), .B2(n25128), .A1_N(n25193), 
        .A2_N(j202_soc_core_bldc_core_00_wdata[12]), .Y(n60) );
  sky130_fd_sc_hd__o2bb2ai_1 U25050 ( .B1(n25193), .B2(n25135), .A1_N(n25193), 
        .A2_N(j202_soc_core_bldc_core_00_wdata[17]), .Y(n31) );
  sky130_fd_sc_hd__o2bb2ai_1 U25051 ( .B1(n25193), .B2(n25139), .A1_N(n25193), 
        .A2_N(j202_soc_core_bldc_core_00_wdata[21]), .Y(n67) );
  sky130_fd_sc_hd__o2bb2ai_1 U25052 ( .B1(n25193), .B2(n25136), .A1_N(n25193), 
        .A2_N(j202_soc_core_bldc_core_00_wdata[18]), .Y(n65) );
  sky130_fd_sc_hd__nor2b_1 U25053 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[23]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N26) );
  sky130_fd_sc_hd__nor2b_1 U25054 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[30]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N33) );
  sky130_fd_sc_hd__nor2b_1 U25055 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[27]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N30) );
  sky130_fd_sc_hd__o2bb2ai_1 U25056 ( .B1(n24440), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[108]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__nor2b_1 U25057 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[31]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N34) );
  sky130_fd_sc_hd__o2bb2ai_1 U25058 ( .B1(n24488), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[105]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o2bb2ai_1 U25059 ( .B1(n24485), .B2(n20497), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[73]), .A2_N(n24288), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__clkinv_1 U25060 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[0]), 
        .Y(n23816) );
  sky130_fd_sc_hd__nor2_1 U25061 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[1]), 
        .B(n23816), .Y(n23815) );
  sky130_fd_sc_hd__nor2b_1 U25062 ( .B_N(j202_soc_core_uart_TOP_rx_bit_cnt[3]), 
        .A(j202_soc_core_uart_TOP_rx_bit_cnt[2]), .Y(n23219) );
  sky130_fd_sc_hd__and2_0 U25063 ( .A(n23815), .B(n23219), .X(n10908) );
  sky130_fd_sc_hd__and2_0 U25064 ( .A(n23853), .B(
        j202_soc_core_uart_TOP_hold_reg[1]), .X(j202_soc_core_uart_TOP_N25) );
  sky130_fd_sc_hd__nand2_1 U25065 ( .A(n25107), .B(n23509), .Y(n23761) );
  sky130_fd_sc_hd__and2_0 U25066 ( .A(j202_soc_core_wbqspiflash_00_spi_out[11]), .B(n23761), .X(j202_soc_core_wbqspiflash_00_N678) );
  sky130_fd_sc_hd__and2_0 U25067 ( .A(j202_soc_core_wbqspiflash_00_spi_out[22]), .B(n23761), .X(j202_soc_core_wbqspiflash_00_N689) );
  sky130_fd_sc_hd__and2_0 U25068 ( .A(j202_soc_core_wbqspiflash_00_spi_out[8]), 
        .B(n23761), .X(j202_soc_core_wbqspiflash_00_N675) );
  sky130_fd_sc_hd__and2_0 U25069 ( .A(j202_soc_core_wbqspiflash_00_spi_out[9]), 
        .B(n23761), .X(j202_soc_core_wbqspiflash_00_N676) );
  sky130_fd_sc_hd__and2_0 U25070 ( .A(j202_soc_core_wbqspiflash_00_spi_out[26]), .B(n23761), .X(j202_soc_core_wbqspiflash_00_N693) );
  sky130_fd_sc_hd__and2_0 U25071 ( .A(j202_soc_core_wbqspiflash_00_spi_out[12]), .B(n23761), .X(j202_soc_core_wbqspiflash_00_N679) );
  sky130_fd_sc_hd__and2_0 U25072 ( .A(j202_soc_core_wbqspiflash_00_spi_out[13]), .B(n23761), .X(j202_soc_core_wbqspiflash_00_N680) );
  sky130_fd_sc_hd__and2_0 U25073 ( .A(j202_soc_core_wbqspiflash_00_spi_out[10]), .B(n23761), .X(j202_soc_core_wbqspiflash_00_N677) );
  sky130_fd_sc_hd__and2_0 U25074 ( .A(j202_soc_core_wbqspiflash_00_spi_out[25]), .B(n23761), .X(j202_soc_core_wbqspiflash_00_N692) );
  sky130_fd_sc_hd__and2_0 U25075 ( .A(j202_soc_core_wbqspiflash_00_spi_out[23]), .B(n23761), .X(j202_soc_core_wbqspiflash_00_N690) );
  sky130_fd_sc_hd__and2_0 U25076 ( .A(j202_soc_core_wbqspiflash_00_spi_out[24]), .B(n23761), .X(j202_soc_core_wbqspiflash_00_N691) );
  sky130_fd_sc_hd__nand2_1 U25077 ( .A(n25005), .B(n23788), .Y(n23784) );
  sky130_fd_sc_hd__o21bai_1 U25078 ( .A1(n25070), .A2(n23785), .B1_N(n23784), 
        .Y(n23361) );
  sky130_fd_sc_hd__nor2_1 U25079 ( .A(j202_soc_core_rst), .B(n23361), .Y(
        j202_soc_core_wbqspiflash_00_N751) );
  sky130_fd_sc_hd__nand2_1 U25080 ( .A(n24894), .B(n25731), .Y(n10562) );
  sky130_fd_sc_hd__nand2_1 U25081 ( .A(n20499), .B(n21599), .Y(n10560) );
  sky130_fd_sc_hd__nor2_1 U25082 ( .A(n21329), .B(n22417), .Y(n21465) );
  sky130_fd_sc_hd__nor3b_1 U25083 ( .C_N(n21339), .A(n24897), .B(n21465), .Y(
        n21528) );
  sky130_fd_sc_hd__nor2_1 U25084 ( .A(n20500), .B(n21527), .Y(n21499) );
  sky130_fd_sc_hd__nand2_1 U25085 ( .A(n21328), .B(n20501), .Y(n21467) );
  sky130_fd_sc_hd__nand3_1 U25086 ( .A(n21528), .B(n21499), .C(n21467), .Y(
        n21003) );
  sky130_fd_sc_hd__nand3_1 U25087 ( .A(j202_soc_core_j22_cpu_opst[3]), .B(
        n20774), .C(n21328), .Y(n23249) );
  sky130_fd_sc_hd__clkinv_1 U25088 ( .A(n23249), .Y(n24895) );
  sky130_fd_sc_hd__a21oi_1 U25089 ( .A1(n24878), .A2(n21441), .B1(n24895), .Y(
        n21002) );
  sky130_fd_sc_hd__nand3_1 U25090 ( .A(n21002), .B(n21408), .C(n22803), .Y(
        n20502) );
  sky130_fd_sc_hd__nor2_1 U25091 ( .A(n21003), .B(n20502), .Y(n21440) );
  sky130_fd_sc_hd__nand2_1 U25092 ( .A(n21440), .B(n21395), .Y(n20503) );
  sky130_fd_sc_hd__a31oi_1 U25093 ( .A1(n21604), .A2(
        j202_soc_core_j22_cpu_opst[1]), .A3(n20773), .B1(n20503), .Y(n20504)
         );
  sky130_fd_sc_hd__o21ai_1 U25094 ( .A1(n20504), .A2(n21592), .B1(n21607), .Y(
        n10568) );
  sky130_fd_sc_hd__o22ai_1 U25095 ( .A1(n20506), .A2(n21997), .B1(n21236), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N2645) );
  sky130_fd_sc_hd__o22ai_1 U25096 ( .A1(n22486), .A2(n21189), .B1(n21188), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N3235) );
  sky130_fd_sc_hd__o22ai_1 U25097 ( .A1(n22486), .A2(n21191), .B1(n21190), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N2680) );
  sky130_fd_sc_hd__o22ai_1 U25098 ( .A1(n22486), .A2(n21070), .B1(n21194), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N2828) );
  sky130_fd_sc_hd__o22ai_1 U25099 ( .A1(n22486), .A2(n21103), .B1(n21192), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N2754) );
  sky130_fd_sc_hd__o22ai_1 U25100 ( .A1(n22486), .A2(n21069), .B1(n21193), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N2976) );
  sky130_fd_sc_hd__o22ai_1 U25101 ( .A1(n22486), .A2(n21071), .B1(n21195), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N3124) );
  sky130_fd_sc_hd__o22ai_1 U25102 ( .A1(n22519), .A2(n21191), .B1(n21190), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N2681) );
  sky130_fd_sc_hd__o22ai_1 U25103 ( .A1(n22519), .A2(n21189), .B1(n21188), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N3236) );
  sky130_fd_sc_hd__o22ai_1 U25104 ( .A1(n22519), .A2(n21069), .B1(n21193), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N2977) );
  sky130_fd_sc_hd__o22ai_1 U25105 ( .A1(n22519), .A2(n21103), .B1(n21192), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N2755) );
  sky130_fd_sc_hd__o22ai_1 U25106 ( .A1(n22519), .A2(n21070), .B1(n21194), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N2829) );
  sky130_fd_sc_hd__o22ai_1 U25107 ( .A1(n22519), .A2(n21071), .B1(n21195), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N3125) );
  sky130_fd_sc_hd__o22ai_1 U25108 ( .A1(n22486), .A2(n21197), .B1(n21196), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N3311) );
  sky130_fd_sc_hd__o22ai_1 U25109 ( .A1(n22486), .A2(n21187), .B1(n21073), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N3198) );
  sky130_fd_sc_hd__o22ai_1 U25110 ( .A1(n22519), .A2(n21197), .B1(n21196), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N3313) );
  sky130_fd_sc_hd__o22ai_1 U25111 ( .A1(n22519), .A2(n21187), .B1(n21073), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N3199) );
  sky130_fd_sc_hd__o22ai_1 U25112 ( .A1(n22519), .A2(n21182), .B1(n21072), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N2792) );
  sky130_fd_sc_hd__o22ai_1 U25113 ( .A1(n22519), .A2(n21184), .B1(n21068), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N3088) );
  sky130_fd_sc_hd__nor2_1 U25114 ( .A(j202_soc_core_j22_cpu_intack), .B(n22721), .Y(n20664) );
  sky130_fd_sc_hd__nand2_1 U25115 ( .A(n22033), .B(n20664), .Y(n20510) );
  sky130_fd_sc_hd__nand2_1 U25116 ( .A(n23239), .B(
        j202_soc_core_j22_cpu_intack), .Y(n21398) );
  sky130_fd_sc_hd__nand2_1 U25117 ( .A(n20666), .B(
        j202_soc_core_intr_level__4_), .Y(n20507) );
  sky130_fd_sc_hd__a21oi_1 U25119 ( .A1(j202_soc_core_intr_level__1_), .A2(
        n20666), .B1(n20665), .Y(n20509) );
  sky130_fd_sc_hd__nor2_1 U25120 ( .A(n22124), .B(n20666), .Y(n20667) );
  sky130_fd_sc_hd__nand2_1 U25121 ( .A(n22555), .B(n20667), .Y(n20508) );
  sky130_fd_sc_hd__nand3_1 U25122 ( .A(n20510), .B(n20509), .C(n20508), .Y(
        j202_soc_core_j22_cpu_rf_N3388) );
  sky130_fd_sc_hd__nand2_1 U25123 ( .A(n21850), .B(n20664), .Y(n20513) );
  sky130_fd_sc_hd__a21oi_1 U25124 ( .A1(j202_soc_core_intr_level__2_), .A2(
        n20666), .B1(n20665), .Y(n20512) );
  sky130_fd_sc_hd__nand2_1 U25125 ( .A(n22045), .B(n20667), .Y(n20511) );
  sky130_fd_sc_hd__nand3_1 U25126 ( .A(n20513), .B(n20512), .C(n20511), .Y(
        j202_soc_core_j22_cpu_rf_N3390) );
  sky130_fd_sc_hd__o22ai_1 U25127 ( .A1(n22723), .A2(n21191), .B1(n21190), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N2678) );
  sky130_fd_sc_hd__o22ai_1 U25128 ( .A1(n22723), .A2(n21189), .B1(n21188), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N3233) );
  sky130_fd_sc_hd__o22ai_1 U25129 ( .A1(n22723), .A2(n21070), .B1(n21194), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N2826) );
  sky130_fd_sc_hd__o22ai_1 U25130 ( .A1(n22723), .A2(n21071), .B1(n21195), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N3122) );
  sky130_fd_sc_hd__o22ai_1 U25131 ( .A1(n22723), .A2(n21069), .B1(n21193), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N2974) );
  sky130_fd_sc_hd__o22ai_1 U25132 ( .A1(n22723), .A2(n21103), .B1(n21192), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N2752) );
  sky130_fd_sc_hd__o22ai_1 U25133 ( .A1(n22723), .A2(n21197), .B1(n21196), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N3307) );
  sky130_fd_sc_hd__o22ai_1 U25134 ( .A1(n22723), .A2(n21187), .B1(n21073), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N3196) );
  sky130_fd_sc_hd__o22ai_1 U25135 ( .A1(n22723), .A2(n21199), .B1(n21198), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N3011) );
  sky130_fd_sc_hd__o22ai_1 U25136 ( .A1(n22723), .A2(n21184), .B1(n21068), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N3085) );
  sky130_fd_sc_hd__o22ai_1 U25137 ( .A1(n22723), .A2(n21201), .B1(n21200), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N2863) );
  sky130_fd_sc_hd__o22ai_1 U25138 ( .A1(n22723), .A2(n21185), .B1(n21132), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N2900) );
  sky130_fd_sc_hd__o22ai_1 U25139 ( .A1(n22723), .A2(n21186), .B1(n21134), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N3159) );
  sky130_fd_sc_hd__o22ai_1 U25140 ( .A1(n22723), .A2(n21183), .B1(n21133), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N2937) );
  sky130_fd_sc_hd__o22ai_1 U25141 ( .A1(n22723), .A2(n21203), .B1(n21202), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N2715) );
  sky130_fd_sc_hd__o22ai_1 U25142 ( .A1(n22723), .A2(n21206), .B1(n21205), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N3048) );
  sky130_fd_sc_hd__o22ai_1 U25143 ( .A1(n22492), .A2(n21189), .B1(n21188), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N3238) );
  sky130_fd_sc_hd__o22ai_1 U25144 ( .A1(n22492), .A2(n21191), .B1(n21190), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N2683) );
  sky130_fd_sc_hd__o22ai_1 U25145 ( .A1(n22492), .A2(n21070), .B1(n21194), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N2831) );
  sky130_fd_sc_hd__o22ai_1 U25146 ( .A1(n22492), .A2(n21069), .B1(n21193), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N2979) );
  sky130_fd_sc_hd__o22ai_1 U25147 ( .A1(n22492), .A2(n21071), .B1(n21195), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N3127) );
  sky130_fd_sc_hd__o22ai_1 U25148 ( .A1(n22492), .A2(n21103), .B1(n21192), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N2757) );
  sky130_fd_sc_hd__o22ai_1 U25149 ( .A1(n22492), .A2(n21197), .B1(n21196), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N3315) );
  sky130_fd_sc_hd__o22ai_1 U25150 ( .A1(n22492), .A2(n21184), .B1(n21068), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N3090) );
  sky130_fd_sc_hd__o22ai_1 U25151 ( .A1(n22492), .A2(n21201), .B1(n21200), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N2868) );
  sky130_fd_sc_hd__o22ai_1 U25152 ( .A1(n22492), .A2(n21187), .B1(n21073), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N3201) );
  sky130_fd_sc_hd__o22ai_1 U25153 ( .A1(n22492), .A2(n21185), .B1(n21132), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N2905) );
  sky130_fd_sc_hd__o22ai_1 U25154 ( .A1(n22492), .A2(n21186), .B1(n21134), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N3164) );
  sky130_fd_sc_hd__o22ai_1 U25155 ( .A1(n22492), .A2(n21183), .B1(n21133), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N2942) );
  sky130_fd_sc_hd__o22ai_1 U25156 ( .A1(n22492), .A2(n21182), .B1(n21072), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N2794) );
  sky130_fd_sc_hd__o22ai_1 U25157 ( .A1(n22492), .A2(n21203), .B1(n21202), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N2720) );
  sky130_fd_sc_hd__o22ai_1 U25158 ( .A1(n22492), .A2(n21199), .B1(n21198), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N3016) );
  sky130_fd_sc_hd__o22ai_1 U25159 ( .A1(n22492), .A2(n21206), .B1(n21205), 
        .B2(n20514), .Y(j202_soc_core_j22_cpu_rf_N3053) );
  sky130_fd_sc_hd__o22ai_1 U25160 ( .A1(n22520), .A2(n21189), .B1(n21188), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N3239) );
  sky130_fd_sc_hd__o22ai_1 U25161 ( .A1(n22520), .A2(n21191), .B1(n21190), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N2684) );
  sky130_fd_sc_hd__o22ai_1 U25162 ( .A1(n22520), .A2(n21103), .B1(n21192), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N2758) );
  sky130_fd_sc_hd__o22ai_1 U25163 ( .A1(n22520), .A2(n21069), .B1(n21193), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N2980) );
  sky130_fd_sc_hd__o22ai_1 U25164 ( .A1(n22520), .A2(n21070), .B1(n21194), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N2832) );
  sky130_fd_sc_hd__o22ai_1 U25165 ( .A1(n22520), .A2(n21071), .B1(n21195), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N3128) );
  sky130_fd_sc_hd__o22ai_1 U25166 ( .A1(n22520), .A2(n21197), .B1(n21196), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N3316) );
  sky130_fd_sc_hd__o22ai_1 U25167 ( .A1(n22520), .A2(n21187), .B1(n21073), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N3202) );
  sky130_fd_sc_hd__o22ai_1 U25168 ( .A1(n22520), .A2(n21201), .B1(n21200), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N2869) );
  sky130_fd_sc_hd__o22ai_1 U25169 ( .A1(n22520), .A2(n21199), .B1(n21198), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N3017) );
  sky130_fd_sc_hd__o22ai_1 U25170 ( .A1(n22520), .A2(n21184), .B1(n21068), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N3091) );
  sky130_fd_sc_hd__o22ai_1 U25171 ( .A1(n22520), .A2(n21203), .B1(n21202), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N2721) );
  sky130_fd_sc_hd__o22ai_1 U25172 ( .A1(n22520), .A2(n21183), .B1(n21133), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N2943) );
  sky130_fd_sc_hd__o22ai_1 U25173 ( .A1(n22520), .A2(n21185), .B1(n21132), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N2906) );
  sky130_fd_sc_hd__o22ai_1 U25174 ( .A1(n22520), .A2(n21186), .B1(n21134), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N3165) );
  sky130_fd_sc_hd__o22ai_1 U25175 ( .A1(n22520), .A2(n21182), .B1(n21072), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N2795) );
  sky130_fd_sc_hd__o22ai_1 U25176 ( .A1(n22520), .A2(n21206), .B1(n21205), 
        .B2(n20515), .Y(j202_soc_core_j22_cpu_rf_N3054) );
  sky130_fd_sc_hd__nand2_1 U25177 ( .A(n22286), .B(n20664), .Y(n20518) );
  sky130_fd_sc_hd__a21oi_1 U25178 ( .A1(j202_soc_core_intr_level__3_), .A2(
        n20666), .B1(n20665), .Y(n20517) );
  sky130_fd_sc_hd__nand2_1 U25179 ( .A(n22495), .B(n20667), .Y(n20516) );
  sky130_fd_sc_hd__nand3_1 U25180 ( .A(n20518), .B(n20517), .C(n20516), .Y(
        j202_soc_core_j22_cpu_rf_N3392) );
  sky130_fd_sc_hd__o22ai_1 U25181 ( .A1(n22486), .A2(n21201), .B1(n21200), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N2865) );
  sky130_fd_sc_hd__o22ai_1 U25182 ( .A1(n22486), .A2(n21199), .B1(n21102), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N3013) );
  sky130_fd_sc_hd__o22ai_1 U25183 ( .A1(n22486), .A2(n21185), .B1(n21132), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N2902) );
  sky130_fd_sc_hd__o22ai_1 U25184 ( .A1(n22723), .A2(n21182), .B1(n21072), 
        .B2(n22720), .Y(j202_soc_core_j22_cpu_rf_N2789) );
  sky130_fd_sc_hd__o22ai_1 U25185 ( .A1(n22486), .A2(n21184), .B1(n21068), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N3087) );
  sky130_fd_sc_hd__o22ai_1 U25186 ( .A1(n22486), .A2(n21183), .B1(n21133), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N2939) );
  sky130_fd_sc_hd__o22ai_1 U25187 ( .A1(n22486), .A2(n21206), .B1(n21205), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N3050) );
  sky130_fd_sc_hd__o22ai_1 U25188 ( .A1(n22519), .A2(n21201), .B1(n21200), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N2866) );
  sky130_fd_sc_hd__o22ai_1 U25189 ( .A1(n22519), .A2(n21183), .B1(n21133), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N2940) );
  sky130_fd_sc_hd__o22ai_1 U25190 ( .A1(n22519), .A2(n21199), .B1(n21102), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N3014) );
  sky130_fd_sc_hd__o22ai_1 U25191 ( .A1(n22519), .A2(n21185), .B1(n21132), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N2903) );
  sky130_fd_sc_hd__o22ai_1 U25192 ( .A1(n22519), .A2(n21206), .B1(n21205), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N3051) );
  sky130_fd_sc_hd__o22ai_1 U25193 ( .A1(n22486), .A2(n21182), .B1(n21072), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N2791) );
  sky130_fd_sc_hd__o22ai_1 U25194 ( .A1(n22486), .A2(n21186), .B1(n21134), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N3161) );
  sky130_fd_sc_hd__o22ai_1 U25195 ( .A1(n22519), .A2(n21186), .B1(n21134), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N3162) );
  sky130_fd_sc_hd__o22ai_1 U25196 ( .A1(n22519), .A2(n21203), .B1(n21202), 
        .B2(n20519), .Y(j202_soc_core_j22_cpu_rf_N2718) );
  sky130_fd_sc_hd__o22ai_1 U25197 ( .A1(n22486), .A2(n21203), .B1(n21202), 
        .B2(n20520), .Y(j202_soc_core_j22_cpu_rf_N2717) );
  sky130_fd_sc_hd__a22oi_1 U25198 ( .A1(n20707), .A2(n22524), .B1(n25308), 
        .B2(n20706), .Y(n22549) );
  sky130_fd_sc_hd__nand2_1 U25199 ( .A(n20708), .B(n22549), .Y(n21925) );
  sky130_fd_sc_hd__nand2_1 U25200 ( .A(n20521), .B(n21137), .Y(n20543) );
  sky130_fd_sc_hd__nand2_1 U25201 ( .A(n21925), .B(n21170), .Y(n20522) );
  sky130_fd_sc_hd__o211ai_1 U25202 ( .A1(n20908), .A2(n21925), .B1(n20905), 
        .C1(n20522), .Y(n20540) );
  sky130_fd_sc_hd__o21ai_1 U25203 ( .A1(n20908), .A2(n20721), .B1(n21010), .Y(
        n20523) );
  sky130_fd_sc_hd__nand2_1 U25204 ( .A(n21925), .B(n20523), .Y(n20538) );
  sky130_fd_sc_hd__nand2_1 U25205 ( .A(n20524), .B(n21139), .Y(n20651) );
  sky130_fd_sc_hd__a2bb2oi_1 U25206 ( .B1(n21935), .B2(n20711), .A1_N(n21627), 
        .A2_N(n20712), .Y(n20525) );
  sky130_fd_sc_hd__o21ai_1 U25207 ( .A1(n21929), .A2(n20651), .B1(n20525), .Y(
        n20536) );
  sky130_fd_sc_hd__nand2_1 U25208 ( .A(n21153), .B(n22584), .Y(n20528) );
  sky130_fd_sc_hd__nand2_1 U25209 ( .A(n22171), .B(n20721), .Y(n22621) );
  sky130_fd_sc_hd__nand2_1 U25210 ( .A(n21929), .B(n22558), .Y(n22473) );
  sky130_fd_sc_hd__o22ai_1 U25211 ( .A1(n22171), .A2(n21145), .B1(n21150), 
        .B2(n22621), .Y(n20526) );
  sky130_fd_sc_hd__a31oi_1 U25212 ( .A1(n21147), .A2(n22621), .A3(n22473), 
        .B1(n20526), .Y(n20527) );
  sky130_fd_sc_hd__o211ai_1 U25213 ( .A1(n22559), .A2(n21154), .B1(n20528), 
        .C1(n20527), .Y(n20529) );
  sky130_fd_sc_hd__a21oi_1 U25214 ( .A1(n20716), .A2(n23322), .B1(n20529), .Y(
        n20534) );
  sky130_fd_sc_hd__a2bb2oi_1 U25215 ( .B1(n21156), .B2(n22133), .A1_N(n22645), 
        .A2_N(n21155), .Y(n20533) );
  sky130_fd_sc_hd__a2bb2oi_1 U25216 ( .B1(n20530), .B2(n21164), .A1_N(n22557), 
        .A2_N(n21163), .Y(n20532) );
  sky130_fd_sc_hd__nand2b_1 U25217 ( .A_N(n20531), .B(n21139), .Y(n20723) );
  sky130_fd_sc_hd__nand4_1 U25218 ( .A(n20534), .B(n20533), .C(n20532), .D(
        n20723), .Y(n20535) );
  sky130_fd_sc_hd__nor2_1 U25219 ( .A(n20536), .B(n20535), .Y(n20537) );
  sky130_fd_sc_hd__nand2_1 U25220 ( .A(n20538), .B(n20537), .Y(n20539) );
  sky130_fd_sc_hd__a21oi_1 U25221 ( .A1(n20540), .A2(n20721), .B1(n20539), .Y(
        n20542) );
  sky130_fd_sc_hd__nand2_1 U25222 ( .A(n21931), .B(n21178), .Y(n20541) );
  sky130_fd_sc_hd__o22ai_1 U25223 ( .A1(n21199), .A2(n22173), .B1(n21102), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N3020) );
  sky130_fd_sc_hd__o22ai_1 U25224 ( .A1(n21184), .A2(n22173), .B1(n21068), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N3094) );
  sky130_fd_sc_hd__o22ai_1 U25225 ( .A1(n21185), .A2(n22173), .B1(n21132), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N2909) );
  sky130_fd_sc_hd__o22ai_1 U25226 ( .A1(n21186), .A2(n22173), .B1(n21134), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N3168) );
  sky130_fd_sc_hd__o22ai_1 U25227 ( .A1(n21203), .A2(n22173), .B1(n21202), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N2724) );
  sky130_fd_sc_hd__o22ai_1 U25228 ( .A1(n21206), .A2(n22173), .B1(n21205), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N3057) );
  sky130_fd_sc_hd__o22ai_1 U25229 ( .A1(n21201), .A2(n22173), .B1(n21200), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N2872) );
  sky130_fd_sc_hd__o22ai_1 U25230 ( .A1(n21183), .A2(n22173), .B1(n21133), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N2946) );
  sky130_fd_sc_hd__o22ai_1 U25231 ( .A1(n21189), .A2(n22173), .B1(n21188), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N3242) );
  sky130_fd_sc_hd__o22ai_1 U25232 ( .A1(n21191), .A2(n22173), .B1(n21190), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N2687) );
  sky130_fd_sc_hd__o22ai_1 U25233 ( .A1(n21071), .A2(n22173), .B1(n21195), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N3131) );
  sky130_fd_sc_hd__o22ai_1 U25234 ( .A1(n21103), .A2(n22173), .B1(n21192), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N2761) );
  sky130_fd_sc_hd__o22ai_1 U25235 ( .A1(n21069), .A2(n22173), .B1(n21193), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N2983) );
  sky130_fd_sc_hd__o22ai_1 U25236 ( .A1(n21070), .A2(n22173), .B1(n21194), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N2835) );
  sky130_fd_sc_hd__o22ai_1 U25237 ( .A1(n22173), .A2(n21197), .B1(n21196), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N3318) );
  sky130_fd_sc_hd__o22ai_1 U25238 ( .A1(n21187), .A2(n22173), .B1(n21073), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N3205) );
  sky130_fd_sc_hd__o22ai_1 U25239 ( .A1(n21182), .A2(n22173), .B1(n21072), 
        .B2(n20544), .Y(j202_soc_core_j22_cpu_rf_N2798) );
  sky130_fd_sc_hd__o22ai_1 U25240 ( .A1(n22290), .A2(n21203), .B1(n21202), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N2723) );
  sky130_fd_sc_hd__o22ai_1 U25241 ( .A1(n22290), .A2(n21201), .B1(n21200), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N2871) );
  sky130_fd_sc_hd__o22ai_1 U25242 ( .A1(n22290), .A2(n21206), .B1(n21205), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N3056) );
  sky130_fd_sc_hd__o22ai_1 U25243 ( .A1(n22290), .A2(n21185), .B1(n21132), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N2908) );
  sky130_fd_sc_hd__o22ai_1 U25244 ( .A1(n22290), .A2(n21187), .B1(n21073), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N3204) );
  sky130_fd_sc_hd__o22ai_1 U25245 ( .A1(n22290), .A2(n21186), .B1(n21134), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N3167) );
  sky130_fd_sc_hd__o22ai_1 U25246 ( .A1(n22290), .A2(n21199), .B1(n21102), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N3019) );
  sky130_fd_sc_hd__o22ai_1 U25247 ( .A1(n22290), .A2(n21183), .B1(n21133), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N2945) );
  sky130_fd_sc_hd__o22ai_1 U25248 ( .A1(n22290), .A2(n21184), .B1(n21068), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N3093) );
  sky130_fd_sc_hd__o22ai_1 U25249 ( .A1(n22290), .A2(n21191), .B1(n21190), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N2686) );
  sky130_fd_sc_hd__o22ai_1 U25250 ( .A1(n22290), .A2(n21189), .B1(n21188), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N3241) );
  sky130_fd_sc_hd__o22ai_1 U25251 ( .A1(n22290), .A2(n21071), .B1(n21195), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N3130) );
  sky130_fd_sc_hd__o22ai_1 U25252 ( .A1(n22290), .A2(n21103), .B1(n21192), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N2760) );
  sky130_fd_sc_hd__o22ai_1 U25253 ( .A1(n22290), .A2(n21069), .B1(n21193), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N2982) );
  sky130_fd_sc_hd__o22ai_1 U25254 ( .A1(n22290), .A2(n21070), .B1(n21194), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N2834) );
  sky130_fd_sc_hd__o22ai_1 U25255 ( .A1(n22290), .A2(n21197), .B1(n21196), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N3317) );
  sky130_fd_sc_hd__o22ai_1 U25256 ( .A1(n22290), .A2(n21182), .B1(n21072), 
        .B2(n20545), .Y(j202_soc_core_j22_cpu_rf_N2797) );
  sky130_fd_sc_hd__nand2_1 U25257 ( .A(n25309), .B(n20706), .Y(n20548) );
  sky130_fd_sc_hd__nand2_1 U25258 ( .A(n20546), .B(n20707), .Y(n20547) );
  sky130_fd_sc_hd__nand3_1 U25259 ( .A(n20708), .B(n20548), .C(n20547), .Y(
        n22554) );
  sky130_fd_sc_hd__o21ai_1 U25260 ( .A1(n20908), .A2(n22554), .B1(n20905), .Y(
        n20549) );
  sky130_fd_sc_hd__nand2_1 U25261 ( .A(n20549), .B(n20648), .Y(n20565) );
  sky130_fd_sc_hd__o2bb2ai_1 U25262 ( .B1(n22037), .B2(n20712), .A1_N(n22575), 
        .A2_N(n20711), .Y(n20550) );
  sky130_fd_sc_hd__a21oi_1 U25263 ( .A1(n20714), .A2(n22159), .B1(n20550), .Y(
        n20564) );
  sky130_fd_sc_hd__nand2b_1 U25264 ( .A_N(n22300), .B(n20648), .Y(n22626) );
  sky130_fd_sc_hd__nand2_1 U25265 ( .A(n22561), .B(n22300), .Y(n22470) );
  sky130_fd_sc_hd__o22ai_1 U25266 ( .A1(n21145), .A2(n22159), .B1(n21150), 
        .B2(n22626), .Y(n20551) );
  sky130_fd_sc_hd__a31oi_1 U25267 ( .A1(n21147), .A2(n22626), .A3(n22470), 
        .B1(n20551), .Y(n20554) );
  sky130_fd_sc_hd__nand2_1 U25268 ( .A(n20716), .B(n23336), .Y(n20553) );
  sky130_fd_sc_hd__a2bb2oi_1 U25269 ( .B1(n21156), .B2(n22578), .A1_N(n22560), 
        .A2_N(n21155), .Y(n20552) );
  sky130_fd_sc_hd__nand3_1 U25270 ( .A(n20554), .B(n20553), .C(n20552), .Y(
        n20559) );
  sky130_fd_sc_hd__nand2_1 U25271 ( .A(n21118), .B(n22136), .Y(n20557) );
  sky130_fd_sc_hd__o22a_1 U25272 ( .A1(n22580), .A2(n21116), .B1(n22562), .B2(
        n21154), .X(n20556) );
  sky130_fd_sc_hd__nand2_1 U25273 ( .A(n21164), .B(n20689), .Y(n20555) );
  sky130_fd_sc_hd__nand4_1 U25274 ( .A(n20557), .B(n20556), .C(n20723), .D(
        n20555), .Y(n20558) );
  sky130_fd_sc_hd__nor2_1 U25275 ( .A(n20559), .B(n20558), .Y(n20563) );
  sky130_fd_sc_hd__nand2_1 U25276 ( .A(n20648), .B(n21170), .Y(n20560) );
  sky130_fd_sc_hd__o211ai_1 U25277 ( .A1(n20908), .A2(n20648), .B1(n21010), 
        .C1(n20560), .Y(n20561) );
  sky130_fd_sc_hd__nand2_1 U25278 ( .A(n22554), .B(n20561), .Y(n20562) );
  sky130_fd_sc_hd__nand4_1 U25279 ( .A(n20565), .B(n20564), .C(n20563), .D(
        n20562), .Y(n20566) );
  sky130_fd_sc_hd__a21oi_1 U25280 ( .A1(n22302), .A2(n21178), .B1(n20566), .Y(
        n20567) );
  sky130_fd_sc_hd__nor2_1 U25281 ( .A(n21236), .B(n22297), .Y(
        j202_soc_core_j22_cpu_rf_N2656) );
  sky130_fd_sc_hd__nand2_1 U25282 ( .A(n25310), .B(n20706), .Y(n20570) );
  sky130_fd_sc_hd__nand2_1 U25283 ( .A(n22517), .B(n20707), .Y(n20569) );
  sky130_fd_sc_hd__nand3_1 U25284 ( .A(n20708), .B(n20570), .C(n20569), .Y(
        n22514) );
  sky130_fd_sc_hd__nand2_1 U25285 ( .A(n20571), .B(n21137), .Y(n20590) );
  sky130_fd_sc_hd__nand2_1 U25286 ( .A(n22514), .B(n21170), .Y(n20572) );
  sky130_fd_sc_hd__o211ai_1 U25287 ( .A1(n20908), .A2(n22514), .B1(n20905), 
        .C1(n20572), .Y(n20587) );
  sky130_fd_sc_hd__nand2_1 U25289 ( .A(n21156), .B(n21867), .Y(n20573) );
  sky130_fd_sc_hd__o211ai_1 U25290 ( .A1(n22612), .A2(n21116), .B1(n20573), 
        .C1(n20723), .Y(n20575) );
  sky130_fd_sc_hd__o2bb2ai_1 U25291 ( .B1(n22563), .B2(n21163), .A1_N(n21164), 
        .A2_N(n20720), .Y(n20574) );
  sky130_fd_sc_hd__nor2_1 U25292 ( .A(n20575), .B(n20574), .Y(n20583) );
  sky130_fd_sc_hd__o2bb2ai_1 U25293 ( .B1(n22611), .B2(n20712), .A1_N(n22579), 
        .A2_N(n20711), .Y(n20576) );
  sky130_fd_sc_hd__a21oi_1 U25294 ( .A1(n20714), .A2(n22156), .B1(n20576), .Y(
        n20582) );
  sky130_fd_sc_hd__nor2_1 U25295 ( .A(n21152), .B(n22156), .Y(n22475) );
  sky130_fd_sc_hd__nand2_1 U25296 ( .A(n22156), .B(n21152), .Y(n22627) );
  sky130_fd_sc_hd__clkinv_1 U25297 ( .A(n22627), .Y(n22474) );
  sky130_fd_sc_hd__nor3_1 U25298 ( .A(n21108), .B(n22475), .C(n22474), .Y(
        n20579) );
  sky130_fd_sc_hd__o22ai_1 U25299 ( .A1(n22156), .A2(n21145), .B1(n21150), 
        .B2(n22627), .Y(n20578) );
  sky130_fd_sc_hd__o22ai_1 U25300 ( .A1(n22561), .A2(n21155), .B1(n22556), 
        .B2(n21154), .Y(n20577) );
  sky130_fd_sc_hd__nor3_1 U25301 ( .A(n20579), .B(n20578), .C(n20577), .Y(
        n20581) );
  sky130_fd_sc_hd__nand2_1 U25302 ( .A(n20716), .B(n23340), .Y(n20580) );
  sky130_fd_sc_hd__nand4_1 U25303 ( .A(n20583), .B(n20582), .C(n20581), .D(
        n20580), .Y(n20584) );
  sky130_fd_sc_hd__a21oi_1 U25304 ( .A1(n22514), .A2(n20585), .B1(n20584), .Y(
        n20586) );
  sky130_fd_sc_hd__nand2_1 U25305 ( .A(n21861), .B(n21178), .Y(n20588) );
  sky130_fd_sc_hd__nand3_1 U25306 ( .A(n20590), .B(n20589), .C(n20588), .Y(
        n21858) );
  sky130_fd_sc_hd__o22ai_1 U25307 ( .A1(n22158), .A2(n21206), .B1(n21205), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N3064) );
  sky130_fd_sc_hd__o22ai_1 U25308 ( .A1(n22158), .A2(n21203), .B1(n21202), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N2731) );
  sky130_fd_sc_hd__o22ai_1 U25309 ( .A1(n22158), .A2(n21183), .B1(n21133), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N2953) );
  sky130_fd_sc_hd__o22ai_1 U25310 ( .A1(n22158), .A2(n21186), .B1(n21134), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N3175) );
  sky130_fd_sc_hd__o22ai_1 U25311 ( .A1(n22158), .A2(n21184), .B1(n21068), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N3101) );
  sky130_fd_sc_hd__o22ai_1 U25312 ( .A1(n22158), .A2(n21201), .B1(n21200), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N2879) );
  sky130_fd_sc_hd__o22ai_1 U25313 ( .A1(n22158), .A2(n21185), .B1(n21132), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N2916) );
  sky130_fd_sc_hd__o22ai_1 U25314 ( .A1(n22158), .A2(n21182), .B1(n21072), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N2805) );
  sky130_fd_sc_hd__o22ai_1 U25315 ( .A1(n22158), .A2(n21187), .B1(n21073), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N3212) );
  sky130_fd_sc_hd__o22ai_1 U25316 ( .A1(n22158), .A2(n21199), .B1(n21102), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N3027) );
  sky130_fd_sc_hd__o22ai_1 U25317 ( .A1(n22158), .A2(n21189), .B1(n21188), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N3249) );
  sky130_fd_sc_hd__o22ai_1 U25318 ( .A1(n22158), .A2(n21191), .B1(n21190), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N2694) );
  sky130_fd_sc_hd__o22ai_1 U25319 ( .A1(n22158), .A2(n21069), .B1(n21193), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N2990) );
  sky130_fd_sc_hd__o22ai_1 U25320 ( .A1(n22158), .A2(n21103), .B1(n21192), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N2768) );
  sky130_fd_sc_hd__o22ai_1 U25321 ( .A1(n22158), .A2(n21071), .B1(n21195), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N3138) );
  sky130_fd_sc_hd__o22ai_1 U25322 ( .A1(n22158), .A2(n21070), .B1(n21194), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N2842) );
  sky130_fd_sc_hd__o22ai_1 U25323 ( .A1(n22158), .A2(n21197), .B1(n21196), 
        .B2(n20591), .Y(j202_soc_core_j22_cpu_rf_N3325) );
  sky130_fd_sc_hd__nand2b_1 U25324 ( .A_N(n22538), .B(n20707), .Y(n20593) );
  sky130_fd_sc_hd__nand2_1 U25325 ( .A(n25311), .B(n20706), .Y(n20592) );
  sky130_fd_sc_hd__nand3_1 U25326 ( .A(n20708), .B(n20593), .C(n20592), .Y(
        n22515) );
  sky130_fd_sc_hd__nand2_1 U25327 ( .A(n20594), .B(n21137), .Y(n20614) );
  sky130_fd_sc_hd__nand2_1 U25328 ( .A(n22515), .B(n21170), .Y(n20595) );
  sky130_fd_sc_hd__o211ai_1 U25329 ( .A1(n20908), .A2(n22515), .B1(n20905), 
        .C1(n20595), .Y(n20611) );
  sky130_fd_sc_hd__o21ai_1 U25330 ( .A1(n20908), .A2(n20689), .B1(n21010), .Y(
        n20596) );
  sky130_fd_sc_hd__nand2_1 U25331 ( .A(n22515), .B(n20596), .Y(n20609) );
  sky130_fd_sc_hd__o2bb2ai_1 U25332 ( .B1(n22711), .B2(n20712), .A1_N(n22576), 
        .A2_N(n20711), .Y(n20597) );
  sky130_fd_sc_hd__a21oi_1 U25333 ( .A1(n20714), .A2(n22164), .B1(n20597), .Y(
        n20608) );
  sky130_fd_sc_hd__nand2b_1 U25334 ( .A_N(n22351), .B(n20689), .Y(n22629) );
  sky130_fd_sc_hd__nand2_1 U25335 ( .A(n22564), .B(n22351), .Y(n22478) );
  sky130_fd_sc_hd__o22ai_1 U25336 ( .A1(n21145), .A2(n22164), .B1(n21150), 
        .B2(n22629), .Y(n20598) );
  sky130_fd_sc_hd__a31oi_1 U25337 ( .A1(n21147), .A2(n22629), .A3(n22478), 
        .B1(n20598), .Y(n20601) );
  sky130_fd_sc_hd__nand2_1 U25338 ( .A(n20716), .B(n23330), .Y(n20600) );
  sky130_fd_sc_hd__a2bb2oi_1 U25339 ( .B1(n21963), .B2(n21156), .A1_N(n22488), 
        .A2_N(n21116), .Y(n20599) );
  sky130_fd_sc_hd__nand3_1 U25340 ( .A(n20601), .B(n20600), .C(n20599), .Y(
        n20606) );
  sky130_fd_sc_hd__nand2_1 U25341 ( .A(n21118), .B(n20648), .Y(n20604) );
  sky130_fd_sc_hd__o22a_1 U25342 ( .A1(n22557), .A2(n21155), .B1(n22560), .B2(
        n21154), .X(n20603) );
  sky130_fd_sc_hd__nand2_1 U25343 ( .A(n21164), .B(n20699), .Y(n20602) );
  sky130_fd_sc_hd__nand4_1 U25344 ( .A(n20604), .B(n20603), .C(n20723), .D(
        n20602), .Y(n20605) );
  sky130_fd_sc_hd__nor2_1 U25345 ( .A(n20606), .B(n20605), .Y(n20607) );
  sky130_fd_sc_hd__nand3_1 U25346 ( .A(n20609), .B(n20608), .C(n20607), .Y(
        n20610) );
  sky130_fd_sc_hd__a21oi_1 U25347 ( .A1(n20611), .A2(n20689), .B1(n20610), .Y(
        n20613) );
  sky130_fd_sc_hd__nand2_1 U25348 ( .A(n22353), .B(n21178), .Y(n20612) );
  sky130_fd_sc_hd__nand3_1 U25349 ( .A(n20614), .B(n20613), .C(n20612), .Y(
        n22346) );
  sky130_fd_sc_hd__o22ai_1 U25350 ( .A1(n22350), .A2(n21203), .B1(n21202), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N2727) );
  sky130_fd_sc_hd__o22ai_1 U25351 ( .A1(n22350), .A2(n21199), .B1(n21102), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N3023) );
  sky130_fd_sc_hd__o22ai_1 U25352 ( .A1(n22350), .A2(n21185), .B1(n21132), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N2912) );
  sky130_fd_sc_hd__o22ai_1 U25353 ( .A1(n22350), .A2(n21187), .B1(n21073), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N3208) );
  sky130_fd_sc_hd__o22ai_1 U25354 ( .A1(n22350), .A2(n21186), .B1(n21134), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N3171) );
  sky130_fd_sc_hd__o22ai_1 U25355 ( .A1(n22350), .A2(n21182), .B1(n21072), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N2801) );
  sky130_fd_sc_hd__o22ai_1 U25356 ( .A1(n22350), .A2(n21206), .B1(n21205), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N3060) );
  sky130_fd_sc_hd__o22ai_1 U25357 ( .A1(n22350), .A2(n21201), .B1(n21200), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N2875) );
  sky130_fd_sc_hd__o22ai_1 U25358 ( .A1(n22350), .A2(n21183), .B1(n21133), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N2949) );
  sky130_fd_sc_hd__o22ai_1 U25359 ( .A1(n22350), .A2(n21184), .B1(n21068), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N3097) );
  sky130_fd_sc_hd__o22ai_1 U25360 ( .A1(n22350), .A2(n21189), .B1(n21188), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N3245) );
  sky130_fd_sc_hd__o22ai_1 U25361 ( .A1(n22350), .A2(n21191), .B1(n21190), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N2690) );
  sky130_fd_sc_hd__o22ai_1 U25362 ( .A1(n22350), .A2(n21103), .B1(n21192), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N2764) );
  sky130_fd_sc_hd__o22ai_1 U25363 ( .A1(n22350), .A2(n21070), .B1(n21194), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N2838) );
  sky130_fd_sc_hd__o22ai_1 U25364 ( .A1(n22350), .A2(n21069), .B1(n21193), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N2986) );
  sky130_fd_sc_hd__o22ai_1 U25365 ( .A1(n22350), .A2(n21071), .B1(n21195), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N3134) );
  sky130_fd_sc_hd__o22ai_1 U25366 ( .A1(n22350), .A2(n21197), .B1(n21196), 
        .B2(n20615), .Y(j202_soc_core_j22_cpu_rf_N3322) );
  sky130_fd_sc_hd__o2bb2ai_1 U25367 ( .B1(n22525), .B2(n20616), .A1_N(n25312), 
        .A2_N(n20706), .Y(n22528) );
  sky130_fd_sc_hd__nand2_1 U25368 ( .A(n20708), .B(n20617), .Y(n22093) );
  sky130_fd_sc_hd__nand2_1 U25369 ( .A(n22093), .B(n21170), .Y(n20618) );
  sky130_fd_sc_hd__o211ai_1 U25370 ( .A1(n20908), .A2(n22093), .B1(n20905), 
        .C1(n20618), .Y(n20619) );
  sky130_fd_sc_hd__nand2_1 U25371 ( .A(n20619), .B(n20720), .Y(n20634) );
  sky130_fd_sc_hd__o2bb2ai_1 U25372 ( .B1(n22646), .B2(n20712), .A1_N(n22631), 
        .A2_N(n20711), .Y(n20620) );
  sky130_fd_sc_hd__a21oi_1 U25373 ( .A1(n20714), .A2(n22161), .B1(n20620), .Y(
        n20633) );
  sky130_fd_sc_hd__nand2b_1 U25374 ( .A_N(n22064), .B(n20720), .Y(n22628) );
  sky130_fd_sc_hd__nand2_1 U25375 ( .A(n22560), .B(n22064), .Y(n22477) );
  sky130_fd_sc_hd__o22ai_1 U25376 ( .A1(n21145), .A2(n22161), .B1(n21150), 
        .B2(n22628), .Y(n20621) );
  sky130_fd_sc_hd__a31oi_1 U25377 ( .A1(n21147), .A2(n22628), .A3(n22477), 
        .B1(n20621), .Y(n20624) );
  sky130_fd_sc_hd__nand2_1 U25378 ( .A(n20716), .B(n23333), .Y(n20623) );
  sky130_fd_sc_hd__a2bb2oi_1 U25379 ( .B1(n21156), .B2(n22577), .A1_N(n22561), 
        .A2_N(n21154), .Y(n20622) );
  sky130_fd_sc_hd__nand3_1 U25380 ( .A(n20624), .B(n20623), .C(n20622), .Y(
        n20629) );
  sky130_fd_sc_hd__nand2_1 U25381 ( .A(n21118), .B(n21152), .Y(n20627) );
  sky130_fd_sc_hd__o22a_1 U25382 ( .A1(n22647), .A2(n21116), .B1(n22564), .B2(
        n21155), .X(n20626) );
  sky130_fd_sc_hd__nand2_1 U25383 ( .A(n21164), .B(n20935), .Y(n20625) );
  sky130_fd_sc_hd__nand4_1 U25384 ( .A(n20627), .B(n20626), .C(n20723), .D(
        n20625), .Y(n20628) );
  sky130_fd_sc_hd__nor2_1 U25385 ( .A(n20629), .B(n20628), .Y(n20632) );
  sky130_fd_sc_hd__nand2_1 U25387 ( .A(n22093), .B(n20630), .Y(n20631) );
  sky130_fd_sc_hd__nand4_1 U25388 ( .A(n20634), .B(n20633), .C(n20632), .D(
        n20631), .Y(n20635) );
  sky130_fd_sc_hd__a21oi_1 U25389 ( .A1(n22066), .A2(n21178), .B1(n20635), .Y(
        n20636) );
  sky130_fd_sc_hd__nor2_1 U25390 ( .A(n21236), .B(n22072), .Y(
        j202_soc_core_j22_cpu_rf_N2655) );
  sky130_fd_sc_hd__o22ai_1 U25391 ( .A1(n22299), .A2(n21191), .B1(n21190), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N2692) );
  sky130_fd_sc_hd__o22ai_1 U25392 ( .A1(n22299), .A2(n21189), .B1(n21188), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N3247) );
  sky130_fd_sc_hd__o22ai_1 U25393 ( .A1(n22299), .A2(n21071), .B1(n21195), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N3136) );
  sky130_fd_sc_hd__o22ai_1 U25394 ( .A1(n22299), .A2(n21070), .B1(n21194), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N2840) );
  sky130_fd_sc_hd__o22ai_1 U25395 ( .A1(n22299), .A2(n21103), .B1(n21192), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N2766) );
  sky130_fd_sc_hd__o22ai_1 U25396 ( .A1(n22299), .A2(n21069), .B1(n21193), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N2988) );
  sky130_fd_sc_hd__o22ai_1 U25397 ( .A1(n22299), .A2(n21197), .B1(n21196), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N3324) );
  sky130_fd_sc_hd__o22ai_1 U25398 ( .A1(n22299), .A2(n21199), .B1(n21198), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N3025) );
  sky130_fd_sc_hd__o22ai_1 U25399 ( .A1(n22299), .A2(n21186), .B1(n21134), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N3173) );
  sky130_fd_sc_hd__o22ai_1 U25400 ( .A1(n22299), .A2(n21183), .B1(n21133), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N2951) );
  sky130_fd_sc_hd__o22ai_1 U25401 ( .A1(n22299), .A2(n21185), .B1(n21132), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N2914) );
  sky130_fd_sc_hd__o22ai_1 U25402 ( .A1(n22299), .A2(n21182), .B1(n21072), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N2803) );
  sky130_fd_sc_hd__o22ai_1 U25403 ( .A1(n22299), .A2(n21187), .B1(n21073), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N3210) );
  sky130_fd_sc_hd__o22ai_1 U25404 ( .A1(n22299), .A2(n21184), .B1(n21068), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N3099) );
  sky130_fd_sc_hd__o22ai_1 U25405 ( .A1(n22299), .A2(n21201), .B1(n21200), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N2877) );
  sky130_fd_sc_hd__o22ai_1 U25406 ( .A1(n22299), .A2(n21203), .B1(n21202), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N2729) );
  sky130_fd_sc_hd__o22ai_1 U25407 ( .A1(n22299), .A2(n21206), .B1(n21205), 
        .B2(n22297), .Y(j202_soc_core_j22_cpu_rf_N3062) );
  sky130_fd_sc_hd__o22ai_1 U25408 ( .A1(n21189), .A2(n22163), .B1(n21188), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N3246) );
  sky130_fd_sc_hd__o22ai_1 U25409 ( .A1(n21191), .A2(n22163), .B1(n21190), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N2691) );
  sky130_fd_sc_hd__o22ai_1 U25410 ( .A1(n21070), .A2(n22163), .B1(n21194), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N2839) );
  sky130_fd_sc_hd__o22ai_1 U25411 ( .A1(n21069), .A2(n22163), .B1(n21193), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N2987) );
  sky130_fd_sc_hd__o22ai_1 U25412 ( .A1(n21103), .A2(n22163), .B1(n21192), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N2765) );
  sky130_fd_sc_hd__o22ai_1 U25413 ( .A1(n21071), .A2(n22163), .B1(n21195), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N3135) );
  sky130_fd_sc_hd__o22ai_1 U25414 ( .A1(n22163), .A2(n21197), .B1(n21196), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N3323) );
  sky130_fd_sc_hd__o22ai_1 U25415 ( .A1(n21185), .A2(n22163), .B1(n21132), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N2913) );
  sky130_fd_sc_hd__o22ai_1 U25416 ( .A1(n21184), .A2(n22163), .B1(n21068), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N3098) );
  sky130_fd_sc_hd__o22ai_1 U25417 ( .A1(n21187), .A2(n22163), .B1(n21073), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N3209) );
  sky130_fd_sc_hd__o22ai_1 U25418 ( .A1(n21186), .A2(n22163), .B1(n21134), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N3172) );
  sky130_fd_sc_hd__o22ai_1 U25419 ( .A1(n21203), .A2(n22163), .B1(n21202), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N2728) );
  sky130_fd_sc_hd__o22ai_1 U25420 ( .A1(n21183), .A2(n22163), .B1(n21133), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N2950) );
  sky130_fd_sc_hd__o22ai_1 U25421 ( .A1(n21199), .A2(n22163), .B1(n21198), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N3024) );
  sky130_fd_sc_hd__o22ai_1 U25422 ( .A1(n21182), .A2(n22163), .B1(n21072), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N2802) );
  sky130_fd_sc_hd__o22ai_1 U25423 ( .A1(n21201), .A2(n22163), .B1(n21200), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N2876) );
  sky130_fd_sc_hd__o22ai_1 U25424 ( .A1(n21206), .A2(n22163), .B1(n21205), 
        .B2(n22072), .Y(j202_soc_core_j22_cpu_rf_N3061) );
  sky130_fd_sc_hd__nand2_1 U25425 ( .A(n20640), .B(n21137), .Y(n20663) );
  sky130_fd_sc_hd__a21oi_1 U25426 ( .A1(n22274), .A2(n20904), .B1(n20641), .Y(
        n20660) );
  sky130_fd_sc_hd__nand2_1 U25427 ( .A(n22136), .B(n21170), .Y(n20642) );
  sky130_fd_sc_hd__o211ai_1 U25428 ( .A1(n20908), .A2(n22136), .B1(n21010), 
        .C1(n20642), .Y(n20658) );
  sky130_fd_sc_hd__a2bb2oi_1 U25429 ( .B1(n21828), .B2(n21156), .A1_N(n22645), 
        .A2_N(n21116), .Y(n20645) );
  sky130_fd_sc_hd__nand2_1 U25430 ( .A(n22154), .B(n22136), .Y(n22622) );
  sky130_fd_sc_hd__nand2_1 U25431 ( .A(n22275), .B(n22556), .Y(n22472) );
  sky130_fd_sc_hd__o22ai_1 U25432 ( .A1(n22154), .A2(n21145), .B1(n21150), 
        .B2(n22622), .Y(n20643) );
  sky130_fd_sc_hd__a31oi_1 U25433 ( .A1(n21147), .A2(n22622), .A3(n22472), 
        .B1(n20643), .Y(n20644) );
  sky130_fd_sc_hd__nand2_1 U25434 ( .A(n20645), .B(n20644), .Y(n20646) );
  sky130_fd_sc_hd__a21oi_1 U25435 ( .A1(n20716), .A2(n23344), .B1(n20646), .Y(
        n20656) );
  sky130_fd_sc_hd__o22ai_1 U25436 ( .A1(n22562), .A2(n21155), .B1(n22563), 
        .B2(n21154), .Y(n20647) );
  sky130_fd_sc_hd__a21oi_1 U25437 ( .A1(n21164), .A2(n20648), .B1(n20647), .Y(
        n20655) );
  sky130_fd_sc_hd__nand3_1 U25438 ( .A(n20649), .B(n21139), .C(n22141), .Y(
        n20650) );
  sky130_fd_sc_hd__nand2_1 U25439 ( .A(n20712), .B(n20650), .Y(n20652) );
  sky130_fd_sc_hd__a2bb2oi_1 U25440 ( .B1(n22704), .B2(n20652), .A1_N(n22275), 
        .A2_N(n20651), .Y(n20654) );
  sky130_fd_sc_hd__a2bb2oi_1 U25441 ( .B1(n22591), .B2(n20711), .A1_N(n22565), 
        .A2_N(n21163), .Y(n20653) );
  sky130_fd_sc_hd__nand4_1 U25442 ( .A(n20656), .B(n20655), .C(n20654), .D(
        n20653), .Y(n20657) );
  sky130_fd_sc_hd__a21oi_1 U25443 ( .A1(n22270), .A2(n20658), .B1(n20657), .Y(
        n20659) );
  sky130_fd_sc_hd__o21a_1 U25444 ( .A1(n22556), .A2(n20660), .B1(n20659), .X(
        n20662) );
  sky130_fd_sc_hd__nand2_1 U25445 ( .A(n22273), .B(n21178), .Y(n20661) );
  sky130_fd_sc_hd__o22ai_1 U25446 ( .A1(n21187), .A2(n22274), .B1(n21073), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N3213) );
  sky130_fd_sc_hd__o22ai_1 U25447 ( .A1(n21183), .A2(n22274), .B1(n21133), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N2954) );
  sky130_fd_sc_hd__o22ai_1 U25448 ( .A1(n21206), .A2(n22274), .B1(n21205), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N3065) );
  sky130_fd_sc_hd__o22ai_1 U25449 ( .A1(n21182), .A2(n22274), .B1(n21072), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N2806) );
  sky130_fd_sc_hd__o22ai_1 U25450 ( .A1(n21199), .A2(n22274), .B1(n21198), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N3028) );
  sky130_fd_sc_hd__o22ai_1 U25451 ( .A1(n21201), .A2(n22274), .B1(n21200), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N2880) );
  sky130_fd_sc_hd__o22ai_1 U25452 ( .A1(n21184), .A2(n22274), .B1(n21068), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N3102) );
  sky130_fd_sc_hd__o22ai_1 U25453 ( .A1(n21185), .A2(n22274), .B1(n21132), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N2917) );
  sky130_fd_sc_hd__o22ai_1 U25454 ( .A1(n21186), .A2(n22274), .B1(n21134), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N3176) );
  sky130_fd_sc_hd__o22ai_1 U25455 ( .A1(n21203), .A2(n22274), .B1(n21202), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N2732) );
  sky130_fd_sc_hd__nand2_1 U25456 ( .A(n22057), .B(n20664), .Y(n20670) );
  sky130_fd_sc_hd__a21oi_1 U25457 ( .A1(j202_soc_core_intr_level__0_), .A2(
        n20666), .B1(n20665), .Y(n20669) );
  sky130_fd_sc_hd__nand2_1 U25458 ( .A(n22484), .B(n20667), .Y(n20668) );
  sky130_fd_sc_hd__nand3_1 U25459 ( .A(n20670), .B(n20669), .C(n20668), .Y(
        j202_soc_core_j22_cpu_rf_N3386) );
  sky130_fd_sc_hd__o22ai_1 U25460 ( .A1(n21069), .A2(n22274), .B1(n21193), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N2991) );
  sky130_fd_sc_hd__o22ai_1 U25461 ( .A1(n21071), .A2(n22274), .B1(n21195), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N3139) );
  sky130_fd_sc_hd__o22ai_1 U25462 ( .A1(n21103), .A2(n22274), .B1(n21192), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N2769) );
  sky130_fd_sc_hd__o22ai_1 U25463 ( .A1(n21070), .A2(n22274), .B1(n21194), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N2843) );
  sky130_fd_sc_hd__o22ai_1 U25464 ( .A1(n21191), .A2(n22274), .B1(n21190), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N2695) );
  sky130_fd_sc_hd__o22ai_1 U25465 ( .A1(n21189), .A2(n22274), .B1(n21188), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N3250) );
  sky130_fd_sc_hd__o22ai_1 U25466 ( .A1(n22274), .A2(n21197), .B1(n21196), 
        .B2(n20671), .Y(j202_soc_core_j22_cpu_rf_N3326) );
  sky130_fd_sc_hd__nor2_1 U25467 ( .A(n22700), .B(n22594), .Y(n22501) );
  sky130_fd_sc_hd__nand2_1 U25468 ( .A(n22501), .B(n22693), .Y(n22698) );
  sky130_fd_sc_hd__nand2_1 U25469 ( .A(n21925), .B(n22721), .Y(n20672) );
  sky130_fd_sc_hd__nand2_1 U25470 ( .A(n23239), .B(n20681), .Y(n21934) );
  sky130_fd_sc_hd__nand2_1 U25471 ( .A(n20672), .B(n21934), .Y(n20673) );
  sky130_fd_sc_hd__a21oi_1 U25472 ( .A1(n21924), .A2(n22124), .B1(n20673), .Y(
        n20680) );
  sky130_fd_sc_hd__fah_1 U25473 ( .A(n22424), .B(n22423), .CI(n20674), .COUT(
        n22511), .SUM(n22426) );
  sky130_fd_sc_hd__xor2_1 U25474 ( .A(j202_soc_core_j22_cpu_rfuo_sr__q_), .B(
        n22591), .X(n20675) );
  sky130_fd_sc_hd__xnor2_1 U25475 ( .A(n22511), .B(n20675), .Y(n22427) );
  sky130_fd_sc_hd__nand2_1 U25476 ( .A(n22501), .B(n22510), .Y(n22596) );
  sky130_fd_sc_hd__o21ai_1 U25477 ( .A1(n22608), .A2(n22596), .B1(n23239), .Y(
        n20676) );
  sky130_fd_sc_hd__a21oi_1 U25478 ( .A1(n22427), .A2(n20677), .B1(n20676), .Y(
        n20678) );
  sky130_fd_sc_hd__o22ai_1 U25479 ( .A1(n20681), .A2(n20680), .B1(n20679), 
        .B2(n20678), .Y(j202_soc_core_j22_cpu_rf_N2638) );
  sky130_fd_sc_hd__nand2_1 U25480 ( .A(n22316), .B(n21178), .Y(n20702) );
  sky130_fd_sc_hd__a22oi_1 U25481 ( .A1(n20707), .A2(n22541), .B1(n25313), 
        .B2(n20706), .Y(n22533) );
  sky130_fd_sc_hd__nand2_1 U25482 ( .A(n20708), .B(n22533), .Y(n22322) );
  sky130_fd_sc_hd__nand2_1 U25483 ( .A(n22322), .B(n21170), .Y(n20682) );
  sky130_fd_sc_hd__o211ai_1 U25484 ( .A1(n20908), .A2(n22322), .B1(n20905), 
        .C1(n20682), .Y(n20700) );
  sky130_fd_sc_hd__o21ai_1 U25485 ( .A1(n20908), .A2(n20699), .B1(n21010), .Y(
        n20683) );
  sky130_fd_sc_hd__nand2_1 U25486 ( .A(n22322), .B(n20683), .Y(n20697) );
  sky130_fd_sc_hd__o2bb2ai_1 U25487 ( .B1(n22754), .B2(n20712), .A1_N(n22574), 
        .A2_N(n20711), .Y(n20684) );
  sky130_fd_sc_hd__a21oi_1 U25488 ( .A1(n20714), .A2(n22169), .B1(n20684), .Y(
        n20696) );
  sky130_fd_sc_hd__nand2b_1 U25489 ( .A_N(n22314), .B(n20699), .Y(n22625) );
  sky130_fd_sc_hd__nand2_1 U25490 ( .A(n22559), .B(n22314), .Y(n22471) );
  sky130_fd_sc_hd__o22ai_1 U25491 ( .A1(n21145), .A2(n22169), .B1(n21150), 
        .B2(n22625), .Y(n20685) );
  sky130_fd_sc_hd__a31oi_1 U25492 ( .A1(n21147), .A2(n22625), .A3(n22471), 
        .B1(n20685), .Y(n20688) );
  sky130_fd_sc_hd__nand2_1 U25493 ( .A(n20716), .B(n23324), .Y(n20687) );
  sky130_fd_sc_hd__o22a_1 U25494 ( .A1(n20805), .A2(n21116), .B1(n22558), .B2(
        n21155), .X(n20686) );
  sky130_fd_sc_hd__nand3_1 U25495 ( .A(n20688), .B(n20687), .C(n20686), .Y(
        n20694) );
  sky130_fd_sc_hd__nand2_1 U25496 ( .A(n21118), .B(n20689), .Y(n20692) );
  sky130_fd_sc_hd__a2bb2oi_1 U25497 ( .B1(n21156), .B2(n21683), .A1_N(n22557), 
        .A2_N(n21154), .Y(n20691) );
  sky130_fd_sc_hd__nand2_1 U25498 ( .A(n21164), .B(n22496), .Y(n20690) );
  sky130_fd_sc_hd__nand4_1 U25499 ( .A(n20692), .B(n20691), .C(n20723), .D(
        n20690), .Y(n20693) );
  sky130_fd_sc_hd__nor2_1 U25500 ( .A(n20694), .B(n20693), .Y(n20695) );
  sky130_fd_sc_hd__nand3_1 U25501 ( .A(n20697), .B(n20696), .C(n20695), .Y(
        n20698) );
  sky130_fd_sc_hd__a21oi_1 U25502 ( .A1(n20700), .A2(n20699), .B1(n20698), .Y(
        n20701) );
  sky130_fd_sc_hd__nand2_1 U25503 ( .A(n20702), .B(n20701), .Y(n20703) );
  sky130_fd_sc_hd__nor2_1 U25504 ( .A(n21236), .B(n22319), .Y(
        j202_soc_core_j22_cpu_rf_N2652) );
  sky130_fd_sc_hd__o22ai_1 U25505 ( .A1(n21189), .A2(n20705), .B1(n21188), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N3243) );
  sky130_fd_sc_hd__o22ai_1 U25506 ( .A1(n21191), .A2(n20705), .B1(n21190), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N2688) );
  sky130_fd_sc_hd__o22ai_1 U25507 ( .A1(n21070), .A2(n20705), .B1(n21194), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N2836) );
  sky130_fd_sc_hd__o22ai_1 U25508 ( .A1(n21103), .A2(n20705), .B1(n21192), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N2762) );
  sky130_fd_sc_hd__o22ai_1 U25509 ( .A1(n21069), .A2(n20705), .B1(n21193), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N2984) );
  sky130_fd_sc_hd__o22ai_1 U25510 ( .A1(n21071), .A2(n20705), .B1(n21195), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N3132) );
  sky130_fd_sc_hd__o22ai_1 U25511 ( .A1(n20705), .A2(n21197), .B1(n21196), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N3319) );
  sky130_fd_sc_hd__o22ai_1 U25512 ( .A1(n21201), .A2(n20705), .B1(n21200), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N2873) );
  sky130_fd_sc_hd__o22ai_1 U25513 ( .A1(n21184), .A2(n20705), .B1(n21068), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N3095) );
  sky130_fd_sc_hd__o22ai_1 U25514 ( .A1(n21199), .A2(n20705), .B1(n21198), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N3021) );
  sky130_fd_sc_hd__o22ai_1 U25515 ( .A1(n21185), .A2(n20705), .B1(n21132), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N2910) );
  sky130_fd_sc_hd__o22ai_1 U25516 ( .A1(n21187), .A2(n20705), .B1(n21073), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N3206) );
  sky130_fd_sc_hd__o22ai_1 U25517 ( .A1(n21183), .A2(n20705), .B1(n21133), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N2947) );
  sky130_fd_sc_hd__o22ai_1 U25518 ( .A1(n21186), .A2(n20705), .B1(n21134), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N3169) );
  sky130_fd_sc_hd__o22ai_1 U25519 ( .A1(n21182), .A2(n20705), .B1(n21072), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N2799) );
  sky130_fd_sc_hd__o22ai_1 U25520 ( .A1(n21203), .A2(n20705), .B1(n21202), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N2725) );
  sky130_fd_sc_hd__o22ai_1 U25521 ( .A1(n21206), .A2(n20705), .B1(n21205), 
        .B2(n22319), .Y(j202_soc_core_j22_cpu_rf_N3058) );
  sky130_fd_sc_hd__a22oi_1 U25522 ( .A1(n20707), .A2(n20825), .B1(n25314), 
        .B2(n20706), .Y(n22534) );
  sky130_fd_sc_hd__nand2_1 U25523 ( .A(n20708), .B(n22534), .Y(n21803) );
  sky130_fd_sc_hd__nand2_1 U25524 ( .A(n21803), .B(n21170), .Y(n20709) );
  sky130_fd_sc_hd__o211ai_1 U25525 ( .A1(n20908), .A2(n21803), .B1(n20905), 
        .C1(n20709), .Y(n20710) );
  sky130_fd_sc_hd__nand2_1 U25526 ( .A(n20710), .B(n20935), .Y(n20732) );
  sky130_fd_sc_hd__o2bb2ai_1 U25527 ( .B1(n22264), .B2(n20712), .A1_N(n22573), 
        .A2_N(n20711), .Y(n20713) );
  sky130_fd_sc_hd__a21oi_1 U25528 ( .A1(n20714), .A2(n22166), .B1(n20713), .Y(
        n20731) );
  sky130_fd_sc_hd__nand2b_1 U25529 ( .A_N(n21807), .B(n20935), .Y(n22630) );
  sky130_fd_sc_hd__nand2b_1 U25530 ( .A_N(n20935), .B(n21807), .Y(n22476) );
  sky130_fd_sc_hd__o22ai_1 U25531 ( .A1(n21145), .A2(n22166), .B1(n21150), 
        .B2(n22630), .Y(n20715) );
  sky130_fd_sc_hd__a31oi_1 U25532 ( .A1(n21147), .A2(n22630), .A3(n22476), 
        .B1(n20715), .Y(n20719) );
  sky130_fd_sc_hd__nand2_1 U25533 ( .A(n20716), .B(n23327), .Y(n20718) );
  sky130_fd_sc_hd__a2bb2oi_1 U25534 ( .B1(n21156), .B2(n21775), .A1_N(n22559), 
        .A2_N(n21155), .Y(n20717) );
  sky130_fd_sc_hd__nand3_1 U25535 ( .A(n20719), .B(n20718), .C(n20717), .Y(
        n20727) );
  sky130_fd_sc_hd__nand2_1 U25536 ( .A(n21118), .B(n20720), .Y(n20725) );
  sky130_fd_sc_hd__o22a_1 U25537 ( .A1(n22487), .A2(n21116), .B1(n22564), .B2(
        n21154), .X(n20724) );
  sky130_fd_sc_hd__nand2_1 U25538 ( .A(n21164), .B(n20721), .Y(n20722) );
  sky130_fd_sc_hd__nand4_1 U25539 ( .A(n20725), .B(n20724), .C(n20723), .D(
        n20722), .Y(n20726) );
  sky130_fd_sc_hd__nor2_1 U25540 ( .A(n20727), .B(n20726), .Y(n20730) );
  sky130_fd_sc_hd__nand2_1 U25542 ( .A(n21803), .B(n20728), .Y(n20729) );
  sky130_fd_sc_hd__nand4_1 U25543 ( .A(n20732), .B(n20731), .C(n20730), .D(
        n20729), .Y(n20733) );
  sky130_fd_sc_hd__a21oi_1 U25544 ( .A1(n21809), .A2(n21178), .B1(n20733), .Y(
        n20734) );
  sky130_fd_sc_hd__nor2_1 U25545 ( .A(n21236), .B(n21805), .Y(
        j202_soc_core_j22_cpu_rf_N2653) );
  sky130_fd_sc_hd__o22ai_1 U25546 ( .A1(n21187), .A2(n22168), .B1(n21073), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N3207) );
  sky130_fd_sc_hd__o22ai_1 U25547 ( .A1(n21201), .A2(n22168), .B1(n21200), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N2874) );
  sky130_fd_sc_hd__o22ai_1 U25548 ( .A1(n21203), .A2(n22168), .B1(n21202), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N2726) );
  sky130_fd_sc_hd__o22ai_1 U25549 ( .A1(n21199), .A2(n22168), .B1(n21102), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N3022) );
  sky130_fd_sc_hd__o22ai_1 U25550 ( .A1(n21206), .A2(n22168), .B1(n21205), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N3059) );
  sky130_fd_sc_hd__o22ai_1 U25551 ( .A1(n21189), .A2(n22168), .B1(n21188), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N3244) );
  sky130_fd_sc_hd__o22ai_1 U25552 ( .A1(n21071), .A2(n22168), .B1(n21195), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N3133) );
  sky130_fd_sc_hd__o22ai_1 U25553 ( .A1(n21103), .A2(n22168), .B1(n21192), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N2763) );
  sky130_fd_sc_hd__o22ai_1 U25554 ( .A1(n22168), .A2(n21197), .B1(n21196), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N3321) );
  sky130_fd_sc_hd__o22ai_1 U25555 ( .A1(n21185), .A2(n22168), .B1(n21132), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N2911) );
  sky130_fd_sc_hd__nand2_1 U25556 ( .A(n20737), .B(n20736), .Y(n20976) );
  sky130_fd_sc_hd__nor2_1 U25557 ( .A(n20975), .B(n20976), .Y(n20740) );
  sky130_fd_sc_hd__nand2b_1 U25558 ( .A_N(n20998), .B(n22328), .Y(n21410) );
  sky130_fd_sc_hd__nor2_1 U25559 ( .A(n24827), .B(n20752), .Y(n21582) );
  sky130_fd_sc_hd__nand2_1 U25560 ( .A(n21640), .B(n20737), .Y(n20760) );
  sky130_fd_sc_hd__and3_1 U25561 ( .A(n22328), .B(n21547), .C(n21416), .X(
        n21553) );
  sky130_fd_sc_hd__a31oi_1 U25562 ( .A1(n21548), .A2(n20737), .A3(n21582), 
        .B1(n21553), .Y(n21523) );
  sky130_fd_sc_hd__nor3_1 U25564 ( .A(n20740), .B(n20739), .C(n20738), .Y(
        n20763) );
  sky130_fd_sc_hd__nor2_1 U25565 ( .A(n22386), .B(n20998), .Y(n22732) );
  sky130_fd_sc_hd__nand2_1 U25566 ( .A(n20741), .B(n21435), .Y(n22738) );
  sky130_fd_sc_hd__nand2b_1 U25567 ( .A_N(n22738), .B(n21547), .Y(n20974) );
  sky130_fd_sc_hd__nand2_1 U25568 ( .A(n20974), .B(n22740), .Y(n21489) );
  sky130_fd_sc_hd__nand2_1 U25569 ( .A(n21635), .B(n20741), .Y(n21485) );
  sky130_fd_sc_hd__nand2_1 U25570 ( .A(n20742), .B(n22735), .Y(n20743) );
  sky130_fd_sc_hd__nand3_1 U25571 ( .A(n21635), .B(n21454), .C(n25372), .Y(
        n22388) );
  sky130_fd_sc_hd__a31oi_1 U25573 ( .A1(n20744), .A2(n25381), .A3(n22743), 
        .B1(n20765), .Y(n20745) );
  sky130_fd_sc_hd__nor2_1 U25575 ( .A(n21608), .B(n20984), .Y(n20747) );
  sky130_fd_sc_hd__nand4_1 U25576 ( .A(n20747), .B(n22741), .C(n20746), .D(
        n22797), .Y(n21513) );
  sky130_fd_sc_hd__nor4_1 U25577 ( .A(n22732), .B(n20994), .C(n21489), .D(
        n21513), .Y(n20748) );
  sky130_fd_sc_hd__nand3b_1 U25578 ( .A_N(n20749), .B(n20763), .C(n20748), .Y(
        n21589) );
  sky130_fd_sc_hd__nand2_1 U25579 ( .A(n20750), .B(n21632), .Y(n21459) );
  sky130_fd_sc_hd__nor2_1 U25580 ( .A(n20751), .B(n21459), .Y(n21039) );
  sky130_fd_sc_hd__nor3_1 U25581 ( .A(n20752), .B(n21455), .C(n22409), .Y(
        n21562) );
  sky130_fd_sc_hd__nor2_1 U25582 ( .A(n24854), .B(n21562), .Y(n21633) );
  sky130_fd_sc_hd__nand2b_1 U25583 ( .A_N(n21505), .B(n21564), .Y(n21401) );
  sky130_fd_sc_hd__nand4_1 U25584 ( .A(n21039), .B(n21633), .C(n20753), .D(
        n21401), .Y(n21476) );
  sky130_fd_sc_hd__o22ai_1 U25585 ( .A1(n21505), .A2(n21474), .B1(n20976), 
        .B2(n20759), .Y(n20754) );
  sky130_fd_sc_hd__nor4_1 U25586 ( .A(n21589), .B(n21476), .C(n21494), .D(
        n20754), .Y(n20756) );
  sky130_fd_sc_hd__a21oi_1 U25587 ( .A1(n22306), .A2(n25315), .B1(n23229), .Y(
        n20755) );
  sky130_fd_sc_hd__a21oi_1 U25588 ( .A1(n20756), .A2(n20755), .B1(n21607), .Y(
        n10575) );
  sky130_fd_sc_hd__o22ai_1 U25589 ( .A1(n22662), .A2(n21187), .B1(n21073), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N3197) );
  sky130_fd_sc_hd__o22ai_1 U25590 ( .A1(n22662), .A2(n21191), .B1(n21190), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N2679) );
  sky130_fd_sc_hd__o22ai_1 U25591 ( .A1(n22662), .A2(n21189), .B1(n21188), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N3234) );
  sky130_fd_sc_hd__o22ai_1 U25592 ( .A1(n22662), .A2(n21070), .B1(n21194), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N2827) );
  sky130_fd_sc_hd__o22ai_1 U25593 ( .A1(n22662), .A2(n21103), .B1(n21192), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N2753) );
  sky130_fd_sc_hd__o22ai_1 U25594 ( .A1(n22662), .A2(n21071), .B1(n21195), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N3123) );
  sky130_fd_sc_hd__o22ai_1 U25595 ( .A1(n22662), .A2(n21069), .B1(n21193), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N2975) );
  sky130_fd_sc_hd__o22ai_1 U25596 ( .A1(n22662), .A2(n21197), .B1(n21196), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N3309) );
  sky130_fd_sc_hd__o22ai_1 U25597 ( .A1(n22662), .A2(n21185), .B1(n21132), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N2901) );
  sky130_fd_sc_hd__o22ai_1 U25598 ( .A1(n22662), .A2(n21201), .B1(n21200), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N2864) );
  sky130_fd_sc_hd__o22ai_1 U25599 ( .A1(n22662), .A2(n21182), .B1(n21072), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N2790) );
  sky130_fd_sc_hd__o22ai_1 U25600 ( .A1(n22662), .A2(n21199), .B1(n21198), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N3012) );
  sky130_fd_sc_hd__o22ai_1 U25601 ( .A1(n22662), .A2(n21184), .B1(n21068), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N3086) );
  sky130_fd_sc_hd__o22ai_1 U25602 ( .A1(n22662), .A2(n21203), .B1(n21202), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N2716) );
  sky130_fd_sc_hd__o22ai_1 U25603 ( .A1(n22662), .A2(n21183), .B1(n21133), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N2938) );
  sky130_fd_sc_hd__o22ai_1 U25604 ( .A1(n22662), .A2(n21186), .B1(n21134), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N3160) );
  sky130_fd_sc_hd__o22ai_1 U25605 ( .A1(n22662), .A2(n21206), .B1(n21205), 
        .B2(n20757), .Y(j202_soc_core_j22_cpu_rf_N3049) );
  sky130_fd_sc_hd__nand2_1 U25606 ( .A(n24869), .B(n20768), .Y(n20758) );
  sky130_fd_sc_hd__nand2_1 U25607 ( .A(n22413), .B(n20758), .Y(n21498) );
  sky130_fd_sc_hd__a21o_1 U25608 ( .A1(n20976), .A2(n20760), .B1(n20759), .X(
        n21506) );
  sky130_fd_sc_hd__nand2_1 U25609 ( .A(n20761), .B(n25387), .Y(n20762) );
  sky130_fd_sc_hd__nand3b_1 U25611 ( .A_N(n21562), .B(n20763), .C(n24860), .Y(
        n22396) );
  sky130_fd_sc_hd__nor2_1 U25612 ( .A(n20764), .B(n22396), .Y(n22415) );
  sky130_fd_sc_hd__nor4_1 U25614 ( .A(n21519), .B(n20994), .C(n20765), .D(
        n22744), .Y(n20769) );
  sky130_fd_sc_hd__nand3_1 U25615 ( .A(n22330), .B(n20766), .C(n22735), .Y(
        n21566) );
  sky130_fd_sc_hd__nand2_1 U25616 ( .A(n20767), .B(n20995), .Y(n20990) );
  sky130_fd_sc_hd__nand2_1 U25617 ( .A(n20768), .B(n25387), .Y(n22736) );
  sky130_fd_sc_hd__nand4_1 U25618 ( .A(n20769), .B(n21566), .C(n20990), .D(
        n22736), .Y(n20770) );
  sky130_fd_sc_hd__nor4_1 U25619 ( .A(n21498), .B(n20772), .C(n20771), .D(
        n20770), .Y(n20777) );
  sky130_fd_sc_hd__nand3_1 U25620 ( .A(j202_soc_core_j22_cpu_opst[2]), .B(
        n20774), .C(n20773), .Y(n20775) );
  sky130_fd_sc_hd__nand2_1 U25621 ( .A(n21467), .B(n20775), .Y(n21526) );
  sky130_fd_sc_hd__nand2_1 U25622 ( .A(n24879), .B(n21526), .Y(n21583) );
  sky130_fd_sc_hd__nand2_1 U25623 ( .A(n20776), .B(n22418), .Y(n22748) );
  sky130_fd_sc_hd__nand2_1 U25624 ( .A(n24879), .B(n21465), .Y(n21490) );
  sky130_fd_sc_hd__o211ai_1 U25625 ( .A1(n24882), .A2(n20777), .B1(n22748), 
        .C1(n21490), .Y(n10593) );
  sky130_fd_sc_hd__nand2_1 U25626 ( .A(n21007), .B(n20778), .Y(n20779) );
  sky130_fd_sc_hd__nand2b_1 U25627 ( .A_N(n20780), .B(n21137), .Y(n20798) );
  sky130_fd_sc_hd__nand2_1 U25628 ( .A(n23309), .B(n20904), .Y(n20781) );
  sky130_fd_sc_hd__o211ai_1 U25629 ( .A1(n22642), .A2(n21150), .B1(n20905), 
        .C1(n20781), .Y(n20795) );
  sky130_fd_sc_hd__nand2_1 U25630 ( .A(n21963), .B(n21170), .Y(n20782) );
  sky130_fd_sc_hd__o211a_2 U25631 ( .A1(n20908), .A2(n21963), .B1(n21010), 
        .C1(n20782), .X(n20793) );
  sky130_fd_sc_hd__xnor2_1 U25632 ( .A(n21963), .B(n23307), .Y(n22456) );
  sky130_fd_sc_hd__clkinv_1 U25633 ( .A(n22456), .Y(n20784) );
  sky130_fd_sc_hd__o22ai_1 U25634 ( .A1(n23307), .A2(n21145), .B1(n22566), 
        .B2(n21155), .Y(n20783) );
  sky130_fd_sc_hd__a21oi_1 U25635 ( .A1(n20784), .A2(n21147), .B1(n20783), .Y(
        n20788) );
  sky130_fd_sc_hd__o22ai_1 U25636 ( .A1(n22564), .A2(n21116), .B1(n22488), 
        .B2(n21158), .Y(n20786) );
  sky130_fd_sc_hd__o2bb2ai_1 U25637 ( .B1(n22641), .B2(n21154), .A1_N(n21156), 
        .A2_N(n22576), .Y(n20785) );
  sky130_fd_sc_hd__nor2_1 U25638 ( .A(n20786), .B(n20785), .Y(n20787) );
  sky130_fd_sc_hd__o211ai_1 U25639 ( .A1(n22642), .A2(n21085), .B1(n20788), 
        .C1(n20787), .Y(n20791) );
  sky130_fd_sc_hd__a2bb2oi_1 U25640 ( .B1(n21683), .B2(n21164), .A1_N(n22600), 
        .A2_N(n21163), .Y(n20789) );
  sky130_fd_sc_hd__o211ai_1 U25641 ( .A1(n22711), .A2(n21167), .B1(n21166), 
        .C1(n20789), .Y(n20790) );
  sky130_fd_sc_hd__nor2_1 U25642 ( .A(n20791), .B(n20790), .Y(n20792) );
  sky130_fd_sc_hd__a21oi_1 U25644 ( .A1(n21963), .A2(n20795), .B1(n20794), .Y(
        n20797) );
  sky130_fd_sc_hd__nand2_1 U25645 ( .A(n21756), .B(n21178), .Y(n20796) );
  sky130_fd_sc_hd__o22ai_1 U25646 ( .A1(n21186), .A2(n23309), .B1(n21134), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N3180) );
  sky130_fd_sc_hd__o22ai_1 U25647 ( .A1(n21184), .A2(n23309), .B1(n21068), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N3106) );
  sky130_fd_sc_hd__o22ai_1 U25648 ( .A1(n21203), .A2(n23309), .B1(n21202), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N2736) );
  sky130_fd_sc_hd__o22ai_1 U25649 ( .A1(n21183), .A2(n23309), .B1(n21133), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N2958) );
  sky130_fd_sc_hd__o22ai_1 U25650 ( .A1(n21206), .A2(n23309), .B1(n21205), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N3069) );
  sky130_fd_sc_hd__o22ai_1 U25651 ( .A1(n21185), .A2(n23309), .B1(n21132), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N2921) );
  sky130_fd_sc_hd__o22ai_1 U25652 ( .A1(n21199), .A2(n23309), .B1(n21102), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N3032) );
  sky130_fd_sc_hd__o22ai_1 U25653 ( .A1(n21201), .A2(n23309), .B1(n21200), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N2884) );
  sky130_fd_sc_hd__o22ai_1 U25654 ( .A1(n21189), .A2(n23309), .B1(n21188), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N3254) );
  sky130_fd_sc_hd__o22ai_1 U25655 ( .A1(n21191), .A2(n23309), .B1(n21190), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N2699) );
  sky130_fd_sc_hd__o22ai_1 U25656 ( .A1(n21071), .A2(n23309), .B1(n21195), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N3143) );
  sky130_fd_sc_hd__o22ai_1 U25657 ( .A1(n21070), .A2(n23309), .B1(n21194), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N2847) );
  sky130_fd_sc_hd__o22ai_1 U25658 ( .A1(n21103), .A2(n23309), .B1(n21192), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N2773) );
  sky130_fd_sc_hd__o22ai_1 U25659 ( .A1(n21069), .A2(n23309), .B1(n21193), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N2995) );
  sky130_fd_sc_hd__o22ai_1 U25660 ( .A1(n21197), .A2(n23309), .B1(n21196), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N3330) );
  sky130_fd_sc_hd__o22ai_1 U25661 ( .A1(n21182), .A2(n23309), .B1(n21072), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N2810) );
  sky130_fd_sc_hd__o22ai_1 U25662 ( .A1(n21187), .A2(n23309), .B1(n21073), 
        .B2(n20799), .Y(j202_soc_core_j22_cpu_rf_N3217) );
  sky130_fd_sc_hd__nand2_1 U25663 ( .A(n21007), .B(n20800), .Y(n20801) );
  sky130_fd_sc_hd__nand2_1 U25664 ( .A(n20802), .B(n21137), .Y(n20823) );
  sky130_fd_sc_hd__nand2_1 U25665 ( .A(n23303), .B(n20904), .Y(n20803) );
  sky130_fd_sc_hd__nand2_1 U25666 ( .A(n20803), .B(n20905), .Y(n20820) );
  sky130_fd_sc_hd__nand2_1 U25667 ( .A(n21683), .B(n21170), .Y(n20804) );
  sky130_fd_sc_hd__o211a_2 U25668 ( .A1(n20908), .A2(n21683), .B1(n21010), 
        .C1(n20804), .X(n20818) );
  sky130_fd_sc_hd__o22ai_1 U25669 ( .A1(n22559), .A2(n21116), .B1(n20805), 
        .B2(n21158), .Y(n20807) );
  sky130_fd_sc_hd__o2bb2ai_1 U25670 ( .B1(n22566), .B2(n21154), .A1_N(n21156), 
        .A2_N(n22574), .Y(n20806) );
  sky130_fd_sc_hd__nor2_1 U25671 ( .A(n20807), .B(n20806), .Y(n20813) );
  sky130_fd_sc_hd__nand2_1 U25672 ( .A(n21144), .B(n23301), .Y(n20812) );
  sky130_fd_sc_hd__nand2_1 U25673 ( .A(n23301), .B(n21683), .Y(n22623) );
  sky130_fd_sc_hd__nand2_1 U25674 ( .A(n22116), .B(n22565), .Y(n22461) );
  sky130_fd_sc_hd__o22ai_1 U25675 ( .A1(n23301), .A2(n21145), .B1(n21150), 
        .B2(n22623), .Y(n20808) );
  sky130_fd_sc_hd__a31oi_1 U25676 ( .A1(n21147), .A2(n22623), .A3(n22461), 
        .B1(n20808), .Y(n20811) );
  sky130_fd_sc_hd__nand2_1 U25677 ( .A(n20809), .B(n22133), .Y(n20810) );
  sky130_fd_sc_hd__nand4_1 U25678 ( .A(n20813), .B(n20812), .C(n20811), .D(
        n20810), .Y(n20816) );
  sky130_fd_sc_hd__a2bb2oi_1 U25679 ( .B1(n22136), .B2(n21164), .A1_N(n22643), 
        .A2_N(n21163), .Y(n20814) );
  sky130_fd_sc_hd__o211ai_1 U25680 ( .A1(n22754), .A2(n21167), .B1(n21166), 
        .C1(n20814), .Y(n20815) );
  sky130_fd_sc_hd__nor2_1 U25681 ( .A(n20816), .B(n20815), .Y(n20817) );
  sky130_fd_sc_hd__o21ai_1 U25682 ( .A1(n20818), .A2(n23303), .B1(n20817), .Y(
        n20819) );
  sky130_fd_sc_hd__a21oi_1 U25683 ( .A1(n21683), .A2(n20820), .B1(n20819), .Y(
        n20822) );
  sky130_fd_sc_hd__nand2_1 U25684 ( .A(n22115), .B(n21178), .Y(n20821) );
  sky130_fd_sc_hd__nand3_1 U25685 ( .A(n20823), .B(n20822), .C(n20821), .Y(
        n22111) );
  sky130_fd_sc_hd__o22ai_1 U25686 ( .A1(n21182), .A2(n23303), .B1(n21072), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N2808) );
  sky130_fd_sc_hd__o22ai_1 U25687 ( .A1(n21187), .A2(n23303), .B1(n21073), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N3215) );
  sky130_fd_sc_hd__o22ai_1 U25688 ( .A1(n21189), .A2(n23303), .B1(n21188), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N3252) );
  sky130_fd_sc_hd__o22ai_1 U25689 ( .A1(n21191), .A2(n23303), .B1(n21190), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N2697) );
  sky130_fd_sc_hd__o22ai_1 U25690 ( .A1(n21070), .A2(n23303), .B1(n21194), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N2845) );
  sky130_fd_sc_hd__o22ai_1 U25691 ( .A1(n21103), .A2(n23303), .B1(n21192), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N2771) );
  sky130_fd_sc_hd__o22ai_1 U25692 ( .A1(n21069), .A2(n23303), .B1(n21193), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N2993) );
  sky130_fd_sc_hd__o22ai_1 U25693 ( .A1(n21071), .A2(n23303), .B1(n21195), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N3141) );
  sky130_fd_sc_hd__o22ai_1 U25694 ( .A1(n21197), .A2(n23303), .B1(n21196), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N3328) );
  sky130_fd_sc_hd__o22ai_1 U25695 ( .A1(n21183), .A2(n23303), .B1(n21133), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N2956) );
  sky130_fd_sc_hd__o22ai_1 U25696 ( .A1(n21184), .A2(n23303), .B1(n21068), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N3104) );
  sky130_fd_sc_hd__o22ai_1 U25697 ( .A1(n21199), .A2(n23303), .B1(n21198), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N3030) );
  sky130_fd_sc_hd__o22ai_1 U25698 ( .A1(n21201), .A2(n23303), .B1(n21200), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N2882) );
  sky130_fd_sc_hd__o22ai_1 U25699 ( .A1(n21185), .A2(n23303), .B1(n21132), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N2919) );
  sky130_fd_sc_hd__o22ai_1 U25700 ( .A1(n21186), .A2(n23303), .B1(n21134), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N3178) );
  sky130_fd_sc_hd__o22ai_1 U25701 ( .A1(n21203), .A2(n23303), .B1(n21202), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N2734) );
  sky130_fd_sc_hd__o22ai_1 U25702 ( .A1(n21206), .A2(n23303), .B1(n21205), 
        .B2(n20824), .Y(j202_soc_core_j22_cpu_rf_N3067) );
  sky130_fd_sc_hd__nand2_1 U25703 ( .A(n21007), .B(n20826), .Y(n20827) );
  sky130_fd_sc_hd__nand2_1 U25704 ( .A(n20828), .B(n21137), .Y(n20855) );
  sky130_fd_sc_hd__nand2_1 U25705 ( .A(n22252), .B(n21178), .Y(n20854) );
  sky130_fd_sc_hd__nand2_1 U25706 ( .A(n23329), .B(n21063), .Y(n20830) );
  sky130_fd_sc_hd__o211ai_1 U25707 ( .A1(n22602), .A2(n20831), .B1(n22691), 
        .C1(n20830), .Y(n20832) );
  sky130_fd_sc_hd__nand2_1 U25708 ( .A(n20832), .B(n22573), .Y(n20844) );
  sky130_fd_sc_hd__a21oi_1 U25709 ( .A1(n20834), .A2(n23327), .B1(n20833), .Y(
        n20843) );
  sky130_fd_sc_hd__xor2_1 U25710 ( .A(n22573), .B(n22602), .X(n22453) );
  sky130_fd_sc_hd__o22ai_1 U25711 ( .A1(n20836), .A2(n23327), .B1(n20835), 
        .B2(n22453), .Y(n20837) );
  sky130_fd_sc_hd__a21oi_1 U25712 ( .A1(n22166), .A2(n20838), .B1(n20837), .Y(
        n20842) );
  sky130_fd_sc_hd__o211ai_1 U25713 ( .A1(n22601), .A2(n20840), .B1(n21063), 
        .C1(n22512), .Y(n20841) );
  sky130_fd_sc_hd__nand4_1 U25714 ( .A(n20844), .B(n20843), .C(n20842), .D(
        n20841), .Y(n20852) );
  sky130_fd_sc_hd__a21oi_1 U25715 ( .A1(n22573), .A2(n21170), .B1(n20845), .Y(
        n20850) );
  sky130_fd_sc_hd__o22ai_1 U25716 ( .A1(n22606), .A2(n21155), .B1(n22610), 
        .B2(n21154), .Y(n20848) );
  sky130_fd_sc_hd__o22ai_1 U25717 ( .A1(n22566), .A2(n21116), .B1(n22557), 
        .B2(n21158), .Y(n20847) );
  sky130_fd_sc_hd__o2bb2ai_1 U25718 ( .B1(n20955), .B2(n21163), .A1_N(n21164), 
        .A2_N(n21935), .Y(n20846) );
  sky130_fd_sc_hd__nor3_1 U25719 ( .A(n20848), .B(n20847), .C(n20846), .Y(
        n20849) );
  sky130_fd_sc_hd__a21oi_1 U25721 ( .A1(n20852), .A2(n21139), .B1(n20851), .Y(
        n20853) );
  sky130_fd_sc_hd__nand3_1 U25722 ( .A(n20855), .B(n20854), .C(n20853), .Y(
        n22248) );
  sky130_fd_sc_hd__o22ai_1 U25723 ( .A1(n21187), .A2(n23329), .B1(n21073), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N3225) );
  sky130_fd_sc_hd__o22ai_1 U25724 ( .A1(n21182), .A2(n23329), .B1(n21072), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N2818) );
  sky130_fd_sc_hd__o22ai_1 U25725 ( .A1(n21103), .A2(n23329), .B1(n21192), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N2781) );
  sky130_fd_sc_hd__o22ai_1 U25726 ( .A1(n21069), .A2(n23329), .B1(n21193), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N3003) );
  sky130_fd_sc_hd__o22ai_1 U25727 ( .A1(n21071), .A2(n23329), .B1(n21195), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N3151) );
  sky130_fd_sc_hd__o22ai_1 U25728 ( .A1(n21070), .A2(n23329), .B1(n21194), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N2855) );
  sky130_fd_sc_hd__o22ai_1 U25729 ( .A1(n21191), .A2(n23329), .B1(n21190), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N2707) );
  sky130_fd_sc_hd__o22ai_1 U25730 ( .A1(n21189), .A2(n23329), .B1(n21188), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N3262) );
  sky130_fd_sc_hd__o22ai_1 U25731 ( .A1(n21183), .A2(n23329), .B1(n21133), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N2966) );
  sky130_fd_sc_hd__o22ai_1 U25732 ( .A1(n21185), .A2(n23329), .B1(n21132), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N2929) );
  sky130_fd_sc_hd__o22ai_1 U25733 ( .A1(n21199), .A2(n23329), .B1(n21198), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N3040) );
  sky130_fd_sc_hd__o22ai_1 U25734 ( .A1(n21201), .A2(n23329), .B1(n21200), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N2892) );
  sky130_fd_sc_hd__o22ai_1 U25735 ( .A1(n21184), .A2(n23329), .B1(n21068), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N3114) );
  sky130_fd_sc_hd__o22ai_1 U25736 ( .A1(n21203), .A2(n23329), .B1(n21202), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N2744) );
  sky130_fd_sc_hd__o22ai_1 U25737 ( .A1(n21186), .A2(n23329), .B1(n21134), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N3188) );
  sky130_fd_sc_hd__o22ai_1 U25738 ( .A1(n21206), .A2(n23329), .B1(n21205), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N3077) );
  sky130_fd_sc_hd__o22ai_1 U25739 ( .A1(n23329), .A2(n21197), .B1(n21196), 
        .B2(n22251), .Y(j202_soc_core_j22_cpu_rf_N3338) );
  sky130_fd_sc_hd__o22ai_1 U25740 ( .A1(n21191), .A2(n22168), .B1(n21190), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N2689) );
  sky130_fd_sc_hd__o22ai_1 U25741 ( .A1(n21070), .A2(n22168), .B1(n21194), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N2837) );
  sky130_fd_sc_hd__o22ai_1 U25742 ( .A1(n21069), .A2(n22168), .B1(n21193), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N2985) );
  sky130_fd_sc_hd__nor2_1 U25743 ( .A(n22551), .B(n22526), .Y(n20856) );
  sky130_fd_sc_hd__nand2b_1 U25744 ( .A_N(n20857), .B(n21137), .Y(n20877) );
  sky130_fd_sc_hd__a21oi_1 U25745 ( .A1(n23315), .A2(n22600), .B1(n21143), .Y(
        n20874) );
  sky130_fd_sc_hd__o21ai_0 U25746 ( .A1(n22600), .A2(n23315), .B1(n21139), .Y(
        n20858) );
  sky130_fd_sc_hd__nand2_1 U25747 ( .A(n20858), .B(n21141), .Y(n20873) );
  sky130_fd_sc_hd__xnor2_1 U25748 ( .A(n22578), .B(n23313), .Y(n22467) );
  sky130_fd_sc_hd__clkinv_1 U25749 ( .A(n22467), .Y(n20860) );
  sky130_fd_sc_hd__o22ai_1 U25750 ( .A1(n23313), .A2(n21145), .B1(n22641), 
        .B2(n21155), .Y(n20859) );
  sky130_fd_sc_hd__a21oi_1 U25751 ( .A1(n20860), .A2(n21147), .B1(n20859), .Y(
        n20864) );
  sky130_fd_sc_hd__o22ai_1 U25752 ( .A1(n22561), .A2(n21116), .B1(n22580), 
        .B2(n21158), .Y(n20862) );
  sky130_fd_sc_hd__o2bb2ai_1 U25753 ( .B1(n22567), .B2(n21154), .A1_N(n21156), 
        .A2_N(n22575), .Y(n20861) );
  sky130_fd_sc_hd__nor2_1 U25754 ( .A(n20862), .B(n20861), .Y(n20863) );
  sky130_fd_sc_hd__o211ai_1 U25755 ( .A1(n22599), .A2(n21085), .B1(n20864), 
        .C1(n20863), .Y(n20867) );
  sky130_fd_sc_hd__a2bb2oi_1 U25756 ( .B1(n21963), .B2(n21164), .A1_N(n22614), 
        .A2_N(n21163), .Y(n20865) );
  sky130_fd_sc_hd__o211ai_1 U25757 ( .A1(n22037), .A2(n21167), .B1(n21166), 
        .C1(n20865), .Y(n20866) );
  sky130_fd_sc_hd__nor2_1 U25758 ( .A(n20867), .B(n20866), .Y(n20871) );
  sky130_fd_sc_hd__a21oi_1 U25759 ( .A1(n23313), .A2(n21089), .B1(n21146), .Y(
        n20868) );
  sky130_fd_sc_hd__nand2_1 U25761 ( .A(n20869), .B(n22578), .Y(n20870) );
  sky130_fd_sc_hd__o211ai_1 U25762 ( .A1(n23315), .A2(n21174), .B1(n20871), 
        .C1(n20870), .Y(n20872) );
  sky130_fd_sc_hd__a21oi_1 U25763 ( .A1(n20874), .A2(n20873), .B1(n20872), .Y(
        n20876) );
  sky130_fd_sc_hd__nand2_1 U25764 ( .A(n21974), .B(n21178), .Y(n20875) );
  sky130_fd_sc_hd__nand3_1 U25765 ( .A(n20877), .B(n20876), .C(n20875), .Y(
        n21970) );
  sky130_fd_sc_hd__o22ai_1 U25766 ( .A1(n21184), .A2(n23315), .B1(n21068), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N3109) );
  sky130_fd_sc_hd__o22ai_1 U25767 ( .A1(n21185), .A2(n23315), .B1(n21132), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N2924) );
  sky130_fd_sc_hd__o22ai_1 U25768 ( .A1(n21199), .A2(n23315), .B1(n21102), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N3035) );
  sky130_fd_sc_hd__o22ai_1 U25769 ( .A1(n21206), .A2(n23315), .B1(n21205), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N3072) );
  sky130_fd_sc_hd__o22ai_1 U25770 ( .A1(n21201), .A2(n23315), .B1(n21200), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N2887) );
  sky130_fd_sc_hd__o22ai_1 U25771 ( .A1(n21183), .A2(n23315), .B1(n21133), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N2961) );
  sky130_fd_sc_hd__o22ai_1 U25772 ( .A1(n21203), .A2(n23315), .B1(n21202), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N2739) );
  sky130_fd_sc_hd__o22ai_1 U25773 ( .A1(n21186), .A2(n23315), .B1(n21134), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N3183) );
  sky130_fd_sc_hd__o22ai_1 U25774 ( .A1(n21189), .A2(n23315), .B1(n21188), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N3257) );
  sky130_fd_sc_hd__o22ai_1 U25775 ( .A1(n21191), .A2(n23315), .B1(n21190), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N2702) );
  sky130_fd_sc_hd__o22ai_1 U25776 ( .A1(n21071), .A2(n23315), .B1(n21195), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N3146) );
  sky130_fd_sc_hd__o22ai_1 U25777 ( .A1(n21070), .A2(n23315), .B1(n21194), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N2850) );
  sky130_fd_sc_hd__o22ai_1 U25778 ( .A1(n21103), .A2(n23315), .B1(n21192), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N2776) );
  sky130_fd_sc_hd__o22ai_1 U25779 ( .A1(n21069), .A2(n23315), .B1(n21193), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N2998) );
  sky130_fd_sc_hd__o22ai_1 U25780 ( .A1(n21184), .A2(n22168), .B1(n21068), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N3096) );
  sky130_fd_sc_hd__o22ai_1 U25781 ( .A1(n21183), .A2(n22168), .B1(n21133), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N2948) );
  sky130_fd_sc_hd__o22ai_1 U25782 ( .A1(n21182), .A2(n22168), .B1(n21072), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N2800) );
  sky130_fd_sc_hd__o22ai_1 U25783 ( .A1(n21186), .A2(n22168), .B1(n21134), 
        .B2(n21805), .Y(j202_soc_core_j22_cpu_rf_N3170) );
  sky130_fd_sc_hd__o22ai_1 U25784 ( .A1(n23315), .A2(n21197), .B1(n21196), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N3333) );
  sky130_fd_sc_hd__o22ai_1 U25785 ( .A1(n21182), .A2(n23315), .B1(n21072), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N2813) );
  sky130_fd_sc_hd__o22ai_1 U25786 ( .A1(n21187), .A2(n23315), .B1(n21073), 
        .B2(n20878), .Y(j202_soc_core_j22_cpu_rf_N3220) );
  sky130_fd_sc_hd__nand2_1 U25787 ( .A(n21007), .B(n20879), .Y(n20880) );
  sky130_fd_sc_hd__nand2b_1 U25788 ( .A_N(n20881), .B(n21137), .Y(n20901) );
  sky130_fd_sc_hd__a21oi_1 U25789 ( .A1(n23321), .A2(n22614), .B1(n21143), .Y(
        n20898) );
  sky130_fd_sc_hd__o21ai_1 U25790 ( .A1(n22614), .A2(n23321), .B1(n21139), .Y(
        n20882) );
  sky130_fd_sc_hd__nand2_1 U25791 ( .A(n20882), .B(n21141), .Y(n20897) );
  sky130_fd_sc_hd__xnor2_1 U25792 ( .A(n21828), .B(n23319), .Y(n22457) );
  sky130_fd_sc_hd__clkinv_1 U25793 ( .A(n22457), .Y(n20884) );
  sky130_fd_sc_hd__o22ai_1 U25794 ( .A1(n23319), .A2(n21145), .B1(n22567), 
        .B2(n21155), .Y(n20883) );
  sky130_fd_sc_hd__a21oi_1 U25795 ( .A1(n20884), .A2(n21147), .B1(n20883), .Y(
        n20888) );
  sky130_fd_sc_hd__o22ai_1 U25796 ( .A1(n22556), .A2(n21116), .B1(n22645), 
        .B2(n21158), .Y(n20886) );
  sky130_fd_sc_hd__o2bb2ai_1 U25797 ( .B1(n22568), .B2(n21154), .A1_N(n21156), 
        .A2_N(n22591), .Y(n20885) );
  sky130_fd_sc_hd__nor2_1 U25798 ( .A(n20886), .B(n20885), .Y(n20887) );
  sky130_fd_sc_hd__o211ai_1 U25799 ( .A1(n22613), .A2(n21085), .B1(n20888), 
        .C1(n20887), .Y(n20891) );
  sky130_fd_sc_hd__a2bb2oi_1 U25800 ( .B1(n22578), .B2(n21164), .A1_N(n22606), 
        .A2_N(n21163), .Y(n20889) );
  sky130_fd_sc_hd__o211ai_1 U25801 ( .A1(n22644), .A2(n21167), .B1(n21166), 
        .C1(n20889), .Y(n20890) );
  sky130_fd_sc_hd__nor2_1 U25802 ( .A(n20891), .B(n20890), .Y(n20895) );
  sky130_fd_sc_hd__a21oi_1 U25803 ( .A1(n23319), .A2(n21089), .B1(n21146), .Y(
        n20892) );
  sky130_fd_sc_hd__o21ai_1 U25804 ( .A1(n21091), .A2(n23321), .B1(n20892), .Y(
        n20893) );
  sky130_fd_sc_hd__nand2_1 U25805 ( .A(n20893), .B(n21828), .Y(n20894) );
  sky130_fd_sc_hd__o211ai_1 U25806 ( .A1(n23321), .A2(n21174), .B1(n20895), 
        .C1(n20894), .Y(n20896) );
  sky130_fd_sc_hd__a21oi_1 U25807 ( .A1(n20898), .A2(n20897), .B1(n20896), .Y(
        n20900) );
  sky130_fd_sc_hd__nand2_1 U25808 ( .A(n21823), .B(n21178), .Y(n20899) );
  sky130_fd_sc_hd__nand3_1 U25809 ( .A(n20901), .B(n20900), .C(n20899), .Y(
        n21819) );
  sky130_fd_sc_hd__o22ai_1 U25810 ( .A1(n21182), .A2(n23321), .B1(n21072), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N2815) );
  sky130_fd_sc_hd__o22ai_1 U25811 ( .A1(n21189), .A2(n23321), .B1(n21188), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N3259) );
  sky130_fd_sc_hd__o22ai_1 U25812 ( .A1(n21191), .A2(n23321), .B1(n21190), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N2704) );
  sky130_fd_sc_hd__o22ai_1 U25813 ( .A1(n21069), .A2(n23321), .B1(n21193), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N3000) );
  sky130_fd_sc_hd__o22ai_1 U25814 ( .A1(n21103), .A2(n23321), .B1(n21192), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N2778) );
  sky130_fd_sc_hd__o22ai_1 U25815 ( .A1(n21071), .A2(n23321), .B1(n21195), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N3148) );
  sky130_fd_sc_hd__o22ai_1 U25816 ( .A1(n21070), .A2(n23321), .B1(n21194), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N2852) );
  sky130_fd_sc_hd__nand2_1 U25817 ( .A(n22373), .B(n21178), .Y(n20924) );
  sky130_fd_sc_hd__nand2_1 U25818 ( .A(n21007), .B(n20902), .Y(n20903) );
  sky130_fd_sc_hd__nand2_1 U25819 ( .A(n23300), .B(n20904), .Y(n20906) );
  sky130_fd_sc_hd__a21oi_1 U25820 ( .A1(n20906), .A2(n20905), .B1(n22563), .Y(
        n20922) );
  sky130_fd_sc_hd__nand2_1 U25821 ( .A(n22133), .B(n21170), .Y(n20907) );
  sky130_fd_sc_hd__o211ai_1 U25822 ( .A1(n20908), .A2(n22133), .B1(n21010), 
        .C1(n20907), .Y(n20909) );
  sky130_fd_sc_hd__nand2_1 U25823 ( .A(n22368), .B(n20909), .Y(n20920) );
  sky130_fd_sc_hd__o2bb2ai_1 U25824 ( .B1(n22556), .B2(n21155), .A1_N(n21156), 
        .A2_N(n21935), .Y(n20914) );
  sky130_fd_sc_hd__o22ai_1 U25825 ( .A1(n22558), .A2(n21116), .B1(n22146), 
        .B2(n21158), .Y(n20913) );
  sky130_fd_sc_hd__nand2_1 U25826 ( .A(n23298), .B(n22133), .Y(n22624) );
  sky130_fd_sc_hd__nand2_1 U25827 ( .A(n22375), .B(n22563), .Y(n22459) );
  sky130_fd_sc_hd__o22ai_1 U25828 ( .A1(n23298), .A2(n21145), .B1(n21150), 
        .B2(n22624), .Y(n20910) );
  sky130_fd_sc_hd__a31oi_1 U25829 ( .A1(n21147), .A2(n22624), .A3(n22459), 
        .B1(n20910), .Y(n20911) );
  sky130_fd_sc_hd__o21ai_1 U25830 ( .A1(n22565), .A2(n21154), .B1(n20911), .Y(
        n20912) );
  sky130_fd_sc_hd__nor3_1 U25831 ( .A(n20914), .B(n20913), .C(n20912), .Y(
        n20919) );
  sky130_fd_sc_hd__nand2_1 U25832 ( .A(n21164), .B(n21152), .Y(n20915) );
  sky130_fd_sc_hd__o211ai_1 U25833 ( .A1(n22566), .A2(n21163), .B1(n20915), 
        .C1(n21166), .Y(n20916) );
  sky130_fd_sc_hd__a21oi_1 U25834 ( .A1(n21053), .A2(n22185), .B1(n20916), .Y(
        n20918) );
  sky130_fd_sc_hd__nand2_1 U25835 ( .A(n21144), .B(n23298), .Y(n20917) );
  sky130_fd_sc_hd__nand4_1 U25836 ( .A(n20920), .B(n20919), .C(n20918), .D(
        n20917), .Y(n20921) );
  sky130_fd_sc_hd__nor2_1 U25837 ( .A(n20922), .B(n20921), .Y(n20923) );
  sky130_fd_sc_hd__nand2_1 U25838 ( .A(n20924), .B(n20923), .Y(n20925) );
  sky130_fd_sc_hd__nor2_1 U25839 ( .A(n21236), .B(n22371), .Y(
        j202_soc_core_j22_cpu_rf_N2660) );
  sky130_fd_sc_hd__o22ai_1 U25840 ( .A1(n21197), .A2(n23321), .B1(n21196), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N3335) );
  sky130_fd_sc_hd__o22ai_1 U25841 ( .A1(n21183), .A2(n23321), .B1(n21133), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N2963) );
  sky130_fd_sc_hd__o22ai_1 U25842 ( .A1(n21185), .A2(n23321), .B1(n21132), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N2926) );
  sky130_fd_sc_hd__o22ai_1 U25843 ( .A1(n21184), .A2(n23321), .B1(n21068), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N3111) );
  sky130_fd_sc_hd__o22ai_1 U25844 ( .A1(n21201), .A2(n23321), .B1(n21200), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N2889) );
  sky130_fd_sc_hd__o22ai_1 U25845 ( .A1(n21199), .A2(n23321), .B1(n21198), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N3037) );
  sky130_fd_sc_hd__o22ai_1 U25846 ( .A1(n21203), .A2(n23321), .B1(n21202), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N2741) );
  sky130_fd_sc_hd__o22ai_1 U25847 ( .A1(n21186), .A2(n23321), .B1(n21134), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N3185) );
  sky130_fd_sc_hd__o22ai_1 U25848 ( .A1(n21187), .A2(n23321), .B1(n21073), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N3222) );
  sky130_fd_sc_hd__o22ai_1 U25849 ( .A1(n21206), .A2(n23321), .B1(n21205), 
        .B2(n20927), .Y(j202_soc_core_j22_cpu_rf_N3074) );
  sky130_fd_sc_hd__nand2_1 U25850 ( .A(n21007), .B(n20928), .Y(n20929) );
  sky130_fd_sc_hd__nand2b_1 U25851 ( .A_N(n20930), .B(n21137), .Y(n20951) );
  sky130_fd_sc_hd__nor2_1 U25852 ( .A(n22566), .B(n23306), .Y(n20943) );
  sky130_fd_sc_hd__nand2_1 U25854 ( .A(n23306), .B(n22566), .Y(n20947) );
  sky130_fd_sc_hd__nand2_1 U25855 ( .A(n23304), .B(n21775), .Y(n22650) );
  sky130_fd_sc_hd__a2bb2oi_1 U25856 ( .B1(n21146), .B2(n21775), .A1_N(n21145), 
        .A2_N(n23304), .Y(n20933) );
  sky130_fd_sc_hd__nand2_1 U25857 ( .A(n21787), .B(n22566), .Y(n22460) );
  sky130_fd_sc_hd__nand3_1 U25858 ( .A(n22460), .B(n21147), .C(n22650), .Y(
        n20932) );
  sky130_fd_sc_hd__o211ai_1 U25859 ( .A1(n21150), .A2(n22650), .B1(n20933), 
        .C1(n20932), .Y(n20934) );
  sky130_fd_sc_hd__a21oi_1 U25860 ( .A1(n21153), .A2(n20935), .B1(n20934), .Y(
        n20939) );
  sky130_fd_sc_hd__o2bb2ai_1 U25861 ( .B1(n22643), .B2(n21154), .A1_N(n21156), 
        .A2_N(n22573), .Y(n20937) );
  sky130_fd_sc_hd__o22ai_1 U25862 ( .A1(n22565), .A2(n21155), .B1(n22487), 
        .B2(n21158), .Y(n20936) );
  sky130_fd_sc_hd__nor2_1 U25863 ( .A(n20937), .B(n20936), .Y(n20938) );
  sky130_fd_sc_hd__o211ai_1 U25864 ( .A1(n21787), .A2(n21085), .B1(n20939), 
        .C1(n20938), .Y(n20942) );
  sky130_fd_sc_hd__a2bb2oi_1 U25865 ( .B1(n22133), .B2(n21164), .A1_N(n22641), 
        .A2_N(n21163), .Y(n20940) );
  sky130_fd_sc_hd__o211ai_1 U25866 ( .A1(n22264), .A2(n21167), .B1(n21166), 
        .C1(n20940), .Y(n20941) );
  sky130_fd_sc_hd__nor2_1 U25867 ( .A(n20942), .B(n20941), .Y(n20945) );
  sky130_fd_sc_hd__nand2_1 U25868 ( .A(n20943), .B(n21170), .Y(n20944) );
  sky130_fd_sc_hd__o211ai_1 U25869 ( .A1(n23306), .A2(n21174), .B1(n20945), 
        .C1(n20944), .Y(n20946) );
  sky130_fd_sc_hd__a31oi_1 U25870 ( .A1(n20948), .A2(n21063), .A3(n20947), 
        .B1(n20946), .Y(n20950) );
  sky130_fd_sc_hd__nand2_1 U25871 ( .A(n21786), .B(n21178), .Y(n20949) );
  sky130_fd_sc_hd__nand3_1 U25872 ( .A(n20951), .B(n20950), .C(n20949), .Y(
        n21782) );
  sky130_fd_sc_hd__o22ai_1 U25873 ( .A1(n21206), .A2(n23306), .B1(n21205), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N3068) );
  sky130_fd_sc_hd__o22ai_1 U25874 ( .A1(n21184), .A2(n23306), .B1(n21068), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N3105) );
  sky130_fd_sc_hd__o22ai_1 U25875 ( .A1(n21183), .A2(n23306), .B1(n21133), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N2957) );
  sky130_fd_sc_hd__o22ai_1 U25876 ( .A1(n21185), .A2(n23306), .B1(n21132), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N2920) );
  sky130_fd_sc_hd__o22ai_1 U25877 ( .A1(n21199), .A2(n23306), .B1(n21102), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N3031) );
  sky130_fd_sc_hd__o22ai_1 U25878 ( .A1(n21201), .A2(n23306), .B1(n21200), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N2883) );
  sky130_fd_sc_hd__o22ai_1 U25879 ( .A1(n21203), .A2(n23306), .B1(n21202), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N2735) );
  sky130_fd_sc_hd__o22ai_1 U25880 ( .A1(n21186), .A2(n23306), .B1(n21134), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N3179) );
  sky130_fd_sc_hd__o22ai_1 U25881 ( .A1(n21189), .A2(n23306), .B1(n21188), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N3253) );
  sky130_fd_sc_hd__o22ai_1 U25882 ( .A1(n21191), .A2(n23306), .B1(n21190), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N2698) );
  sky130_fd_sc_hd__o22ai_1 U25883 ( .A1(n21103), .A2(n23306), .B1(n21192), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N2772) );
  sky130_fd_sc_hd__o22ai_1 U25884 ( .A1(n21069), .A2(n23306), .B1(n21193), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N2994) );
  sky130_fd_sc_hd__o22ai_1 U25885 ( .A1(n21071), .A2(n23306), .B1(n21195), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N3142) );
  sky130_fd_sc_hd__o22ai_1 U25886 ( .A1(n21070), .A2(n23306), .B1(n21194), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N2846) );
  sky130_fd_sc_hd__o22ai_1 U25887 ( .A1(n21197), .A2(n23306), .B1(n21196), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N3329) );
  sky130_fd_sc_hd__o22ai_1 U25888 ( .A1(n21182), .A2(n23306), .B1(n21072), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N2809) );
  sky130_fd_sc_hd__o22ai_1 U25889 ( .A1(n21187), .A2(n23306), .B1(n21073), 
        .B2(n20952), .Y(j202_soc_core_j22_cpu_rf_N3216) );
  sky130_fd_sc_hd__nand2_1 U25890 ( .A(n21007), .B(n22538), .Y(n20953) );
  sky130_fd_sc_hd__nand2_1 U25891 ( .A(n21952), .B(n21178), .Y(n20973) );
  sky130_fd_sc_hd__a21oi_1 U25892 ( .A1(n23332), .A2(n22610), .B1(n21143), .Y(
        n20969) );
  sky130_fd_sc_hd__nand2_1 U25894 ( .A(n20954), .B(n21141), .Y(n20968) );
  sky130_fd_sc_hd__xnor2_1 U25895 ( .A(n22576), .B(n23330), .Y(n22447) );
  sky130_fd_sc_hd__o22a_1 U25896 ( .A1(n22643), .A2(n21116), .B1(n21108), .B2(
        n22447), .X(n20959) );
  sky130_fd_sc_hd__o22ai_1 U25897 ( .A1(n23330), .A2(n21145), .B1(n22601), 
        .B2(n21155), .Y(n20957) );
  sky130_fd_sc_hd__o22ai_1 U25898 ( .A1(n20955), .A2(n21154), .B1(n22564), 
        .B2(n21158), .Y(n20956) );
  sky130_fd_sc_hd__nor2_1 U25899 ( .A(n20957), .B(n20956), .Y(n20958) );
  sky130_fd_sc_hd__o211ai_1 U25900 ( .A1(n22609), .A2(n21085), .B1(n20959), 
        .C1(n20958), .Y(n20962) );
  sky130_fd_sc_hd__a2bb2oi_1 U25901 ( .B1(n22574), .B2(n21164), .A1_N(n21048), 
        .A2_N(n21163), .Y(n20960) );
  sky130_fd_sc_hd__o211ai_1 U25902 ( .A1(n22351), .A2(n21167), .B1(n21166), 
        .C1(n20960), .Y(n20961) );
  sky130_fd_sc_hd__nor2_1 U25903 ( .A(n20962), .B(n20961), .Y(n20966) );
  sky130_fd_sc_hd__a21oi_1 U25904 ( .A1(n23330), .A2(n21089), .B1(n21146), .Y(
        n20963) );
  sky130_fd_sc_hd__nand2_1 U25906 ( .A(n20964), .B(n22576), .Y(n20965) );
  sky130_fd_sc_hd__o211ai_1 U25907 ( .A1(n23332), .A2(n21174), .B1(n20966), 
        .C1(n20965), .Y(n20967) );
  sky130_fd_sc_hd__a21oi_1 U25908 ( .A1(n20969), .A2(n20968), .B1(n20967), .Y(
        n20972) );
  sky130_fd_sc_hd__nand2_1 U25909 ( .A(n20970), .B(n21137), .Y(n20971) );
  sky130_fd_sc_hd__nand3_1 U25910 ( .A(n20973), .B(n20972), .C(n20971), .Y(
        n21947) );
  sky130_fd_sc_hd__o22ai_1 U25911 ( .A1(n21182), .A2(n23332), .B1(n21072), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N2819) );
  sky130_fd_sc_hd__o22ai_1 U25912 ( .A1(n21187), .A2(n23332), .B1(n21073), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N3226) );
  sky130_fd_sc_hd__o22ai_1 U25913 ( .A1(n21191), .A2(n23332), .B1(n21190), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N2708) );
  sky130_fd_sc_hd__o22ai_1 U25914 ( .A1(n21189), .A2(n23332), .B1(n21188), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N3263) );
  sky130_fd_sc_hd__o22ai_1 U25915 ( .A1(n21103), .A2(n23332), .B1(n21192), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N2782) );
  sky130_fd_sc_hd__o22ai_1 U25916 ( .A1(n21069), .A2(n23332), .B1(n21193), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N3004) );
  sky130_fd_sc_hd__o22ai_1 U25917 ( .A1(n21070), .A2(n23332), .B1(n21194), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N2856) );
  sky130_fd_sc_hd__o22ai_1 U25918 ( .A1(n21071), .A2(n23332), .B1(n21195), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N3152) );
  sky130_fd_sc_hd__o22ai_1 U25919 ( .A1(n21197), .A2(n23332), .B1(n21196), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N3339) );
  sky130_fd_sc_hd__o22ai_1 U25920 ( .A1(n21199), .A2(n23332), .B1(n21198), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N3041) );
  sky130_fd_sc_hd__o22ai_1 U25921 ( .A1(n21185), .A2(n23332), .B1(n21132), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N2930) );
  sky130_fd_sc_hd__o22ai_1 U25922 ( .A1(n21184), .A2(n23332), .B1(n21068), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N3115) );
  sky130_fd_sc_hd__o22ai_1 U25923 ( .A1(n21201), .A2(n23332), .B1(n21200), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N2893) );
  sky130_fd_sc_hd__o22ai_1 U25924 ( .A1(n21183), .A2(n23332), .B1(n21133), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N2967) );
  sky130_fd_sc_hd__o22ai_1 U25925 ( .A1(n21203), .A2(n23332), .B1(n21202), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N2745) );
  sky130_fd_sc_hd__o22ai_1 U25926 ( .A1(n21186), .A2(n23332), .B1(n21134), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N3189) );
  sky130_fd_sc_hd__o22ai_1 U25927 ( .A1(n21206), .A2(n23332), .B1(n21205), 
        .B2(n21951), .Y(j202_soc_core_j22_cpu_rf_N3078) );
  sky130_fd_sc_hd__o21ai_1 U25929 ( .A1(n24872), .A2(n21413), .B1(n20977), .Y(
        n21565) );
  sky130_fd_sc_hd__nor2_1 U25930 ( .A(n21546), .B(n21565), .Y(n21515) );
  sky130_fd_sc_hd__nand2_1 U25932 ( .A(n20980), .B(n21522), .Y(n22282) );
  sky130_fd_sc_hd__nand4_1 U25933 ( .A(n21523), .B(n21515), .C(n21430), .D(
        n21506), .Y(n21001) );
  sky130_fd_sc_hd__a21oi_1 U25934 ( .A1(n22309), .A2(n20981), .B1(n24867), .Y(
        n20982) );
  sky130_fd_sc_hd__nand3_1 U25935 ( .A(n20982), .B(n21556), .C(n21473), .Y(
        n21524) );
  sky130_fd_sc_hd__nand2b_1 U25936 ( .A_N(n21524), .B(n24861), .Y(n21497) );
  sky130_fd_sc_hd__nor3_1 U25937 ( .A(n20986), .B(n20983), .C(n21455), .Y(
        n21554) );
  sky130_fd_sc_hd__a211oi_1 U25938 ( .A1(n24872), .A2(n21492), .B1(n21554), 
        .C1(n20984), .Y(n21000) );
  sky130_fd_sc_hd__nor2_1 U25939 ( .A(n20988), .B(n22407), .Y(n22746) );
  sky130_fd_sc_hd__nor2_1 U25940 ( .A(n21455), .B(n20985), .Y(n21422) );
  sky130_fd_sc_hd__nor2_1 U25941 ( .A(n20986), .B(n21409), .Y(n24841) );
  sky130_fd_sc_hd__a21oi_1 U25942 ( .A1(n22743), .A2(n20987), .B1(n22742), .Y(
        n22411) );
  sky130_fd_sc_hd__o22ai_1 U25943 ( .A1(n20988), .A2(n21455), .B1(n22407), 
        .B2(n21474), .Y(n24847) );
  sky130_fd_sc_hd__nor4_1 U25944 ( .A(n22746), .B(n24841), .C(n22411), .D(
        n24847), .Y(n20991) );
  sky130_fd_sc_hd__nand2_1 U25945 ( .A(n22734), .B(n20989), .Y(n24850) );
  sky130_fd_sc_hd__nand3_1 U25946 ( .A(n20991), .B(n24850), .C(n20990), .Y(
        n21590) );
  sky130_fd_sc_hd__nand3_1 U25947 ( .A(n21454), .B(n22735), .C(n25372), .Y(
        n21636) );
  sky130_fd_sc_hd__nand2_1 U25950 ( .A(n20996), .B(n20995), .Y(n21404) );
  sky130_fd_sc_hd__nand2_1 U25951 ( .A(n21431), .B(n21404), .Y(n20997) );
  sky130_fd_sc_hd__nor4_1 U25952 ( .A(n21590), .B(n24848), .C(n21496), .D(
        n20997), .Y(n20999) );
  sky130_fd_sc_hd__nand4_1 U25953 ( .A(n21000), .B(n20999), .C(n20998), .D(
        n21402), .Y(n21593) );
  sky130_fd_sc_hd__o31ai_1 U25954 ( .A1(n21001), .A2(n21497), .A3(n21593), 
        .B1(n24858), .Y(n21005) );
  sky130_fd_sc_hd__nand2_1 U25956 ( .A(n24879), .B(n21003), .Y(n21452) );
  sky130_fd_sc_hd__nand3_1 U25957 ( .A(n21005), .B(n21004), .C(n21452), .Y(
        n10578) );
  sky130_fd_sc_hd__nand2_1 U25958 ( .A(n21006), .B(n21137), .Y(n21037) );
  sky130_fd_sc_hd__nand2_1 U25959 ( .A(n21007), .B(n22542), .Y(n21008) );
  sky130_fd_sc_hd__nor2_1 U25961 ( .A(n21011), .B(n22619), .Y(n22590) );
  sky130_fd_sc_hd__o211ai_1 U25963 ( .A1(n22590), .A2(n22176), .B1(n22181), 
        .C1(n21012), .Y(n21016) );
  sky130_fd_sc_hd__o22ai_1 U25964 ( .A1(n23344), .A2(n21145), .B1(n22604), 
        .B2(n21155), .Y(n21014) );
  sky130_fd_sc_hd__o22ai_1 U25965 ( .A1(n22614), .A2(n21116), .B1(n22556), 
        .B2(n21158), .Y(n21013) );
  sky130_fd_sc_hd__nor2_1 U25966 ( .A(n21014), .B(n21013), .Y(n21015) );
  sky130_fd_sc_hd__o211ai_1 U25967 ( .A1(n22607), .A2(n21085), .B1(n21016), 
        .C1(n21015), .Y(n21024) );
  sky130_fd_sc_hd__xnor2_1 U25968 ( .A(n22591), .B(n23344), .Y(n22595) );
  sky130_fd_sc_hd__nand3_1 U25970 ( .A(n21020), .B(n21139), .C(n22154), .Y(
        n21021) );
  sky130_fd_sc_hd__a21oi_1 U25972 ( .A1(n21164), .A2(n22575), .B1(n21022), .Y(
        n21023) );
  sky130_fd_sc_hd__nand3b_1 U25973 ( .A_N(n21024), .B(n21023), .C(n21166), .Y(
        n21025) );
  sky130_fd_sc_hd__a21oi_1 U25974 ( .A1(n22358), .A2(n21026), .B1(n21025), .Y(
        n21036) );
  sky130_fd_sc_hd__nand2_1 U25975 ( .A(n22358), .B(n21170), .Y(n21033) );
  sky130_fd_sc_hd__a21oi_1 U25976 ( .A1(n23344), .A2(n21089), .B1(n21146), .Y(
        n21032) );
  sky130_fd_sc_hd__nand2_1 U25977 ( .A(n23348), .B(n21028), .Y(n21031) );
  sky130_fd_sc_hd__nand3_1 U25978 ( .A(n21029), .B(n22264), .C(n22176), .Y(
        n21030) );
  sky130_fd_sc_hd__nand4_1 U25979 ( .A(n21033), .B(n21032), .C(n21031), .D(
        n21030), .Y(n21034) );
  sky130_fd_sc_hd__nand2_1 U25980 ( .A(n21034), .B(n22591), .Y(n21035) );
  sky130_fd_sc_hd__nand3_1 U25981 ( .A(n21037), .B(n21036), .C(n21035), .Y(
        n21038) );
  sky130_fd_sc_hd__nor2_1 U25982 ( .A(n21236), .B(n11201), .Y(
        j202_soc_core_j22_cpu_rf_N2676) );
  sky130_fd_sc_hd__nor2_1 U25983 ( .A(n22282), .B(n21532), .Y(n21043) );
  sky130_fd_sc_hd__nand2_1 U25984 ( .A(n25383), .B(n24858), .Y(n22308) );
  sky130_fd_sc_hd__a21oi_1 U25985 ( .A1(n21492), .A2(n25316), .B1(n24826), .Y(
        n22307) );
  sky130_fd_sc_hd__nand3_1 U25986 ( .A(n22280), .B(n24858), .C(n25384), .Y(
        n21042) );
  sky130_fd_sc_hd__nand3_1 U25987 ( .A(n24861), .B(n21039), .C(n21599), .Y(
        n21041) );
  sky130_fd_sc_hd__o211ai_1 U25988 ( .A1(n21043), .A2(n22308), .B1(n21042), 
        .C1(n22283), .Y(n10492) );
  sky130_fd_sc_hd__o22ai_1 U25989 ( .A1(n21182), .A2(n23300), .B1(n21072), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N2807) );
  sky130_fd_sc_hd__o22ai_1 U25990 ( .A1(n21187), .A2(n23300), .B1(n21073), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N3214) );
  sky130_fd_sc_hd__o22ai_1 U25991 ( .A1(n21191), .A2(n23300), .B1(n21190), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N2696) );
  sky130_fd_sc_hd__o22ai_1 U25992 ( .A1(n21189), .A2(n23300), .B1(n21188), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N3251) );
  sky130_fd_sc_hd__o22ai_1 U25993 ( .A1(n21070), .A2(n23300), .B1(n21194), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N2844) );
  sky130_fd_sc_hd__o22ai_1 U25994 ( .A1(n21103), .A2(n23300), .B1(n21192), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N2770) );
  sky130_fd_sc_hd__o22ai_1 U25995 ( .A1(n21069), .A2(n23300), .B1(n21193), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N2992) );
  sky130_fd_sc_hd__o22ai_1 U25996 ( .A1(n21071), .A2(n23300), .B1(n21195), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N3140) );
  sky130_fd_sc_hd__nand2_1 U25997 ( .A(n21044), .B(n21137), .Y(n21066) );
  sky130_fd_sc_hd__nor2_1 U25998 ( .A(n22551), .B(n21045), .Y(n21046) );
  sky130_fd_sc_hd__a21oi_1 U25999 ( .A1(n23340), .A2(n21089), .B1(n21146), .Y(
        n21047) );
  sky130_fd_sc_hd__o22ai_1 U26001 ( .A1(n21145), .A2(n23340), .B1(n21048), 
        .B2(n21155), .Y(n21051) );
  sky130_fd_sc_hd__o22ai_1 U26002 ( .A1(n22567), .A2(n21116), .B1(n22608), 
        .B2(n21154), .Y(n21050) );
  sky130_fd_sc_hd__nor3_1 U26003 ( .A(n21051), .B(n21050), .C(n21049), .Y(
        n21057) );
  sky130_fd_sc_hd__xnor2_1 U26004 ( .A(n22579), .B(n23340), .Y(n22448) );
  sky130_fd_sc_hd__o22ai_1 U26005 ( .A1(n22562), .A2(n21158), .B1(n21108), 
        .B2(n22448), .Y(n21052) );
  sky130_fd_sc_hd__a21oi_1 U26006 ( .A1(n21164), .A2(n22631), .B1(n21052), .Y(
        n21056) );
  sky130_fd_sc_hd__nand2_1 U26007 ( .A(n21144), .B(n23340), .Y(n21055) );
  sky130_fd_sc_hd__nand2_1 U26008 ( .A(n21053), .B(n22156), .Y(n21054) );
  sky130_fd_sc_hd__nand4_1 U26009 ( .A(n21057), .B(n21056), .C(n21055), .D(
        n21054), .Y(n21058) );
  sky130_fd_sc_hd__o21bai_1 U26010 ( .A1(n21174), .A2(n23342), .B1_N(n21058), 
        .Y(n21059) );
  sky130_fd_sc_hd__a21oi_1 U26011 ( .A1(n21060), .A2(n22579), .B1(n21059), .Y(
        n21065) );
  sky130_fd_sc_hd__o21ai_1 U26012 ( .A1(n22604), .A2(n23342), .B1(n21139), .Y(
        n21061) );
  sky130_fd_sc_hd__nand2_1 U26013 ( .A(n21061), .B(n21141), .Y(n21062) );
  sky130_fd_sc_hd__o211ai_1 U26014 ( .A1(n22579), .A2(n21890), .B1(n21063), 
        .C1(n21062), .Y(n21064) );
  sky130_fd_sc_hd__nand3_1 U26015 ( .A(n21066), .B(n21065), .C(n21064), .Y(
        n21067) );
  sky130_fd_sc_hd__nor2_1 U26016 ( .A(n21236), .B(n11199), .Y(
        j202_soc_core_j22_cpu_rf_N2675) );
  sky130_fd_sc_hd__o22ai_1 U26017 ( .A1(n21197), .A2(n23300), .B1(n21196), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N3327) );
  sky130_fd_sc_hd__o22ai_1 U26018 ( .A1(n21199), .A2(n23300), .B1(n21198), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N3029) );
  sky130_fd_sc_hd__o22ai_1 U26019 ( .A1(n21185), .A2(n23300), .B1(n21132), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N2918) );
  sky130_fd_sc_hd__o22ai_1 U26020 ( .A1(n21184), .A2(n23300), .B1(n21068), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N3103) );
  sky130_fd_sc_hd__o22ai_1 U26021 ( .A1(n21201), .A2(n23300), .B1(n21200), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N2881) );
  sky130_fd_sc_hd__o22ai_1 U26022 ( .A1(n21183), .A2(n23300), .B1(n21133), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N2955) );
  sky130_fd_sc_hd__o22ai_1 U26023 ( .A1(n21186), .A2(n23300), .B1(n21134), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N3177) );
  sky130_fd_sc_hd__o22ai_1 U26024 ( .A1(n21203), .A2(n23300), .B1(n21202), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N2733) );
  sky130_fd_sc_hd__o22ai_1 U26025 ( .A1(n21206), .A2(n23300), .B1(n21205), 
        .B2(n22371), .Y(j202_soc_core_j22_cpu_rf_N3066) );
  sky130_fd_sc_hd__o22ai_1 U26026 ( .A1(n21201), .A2(n23348), .B1(n21200), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N2898) );
  sky130_fd_sc_hd__o22ai_1 U26027 ( .A1(n21184), .A2(n23348), .B1(n21068), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N3120) );
  sky130_fd_sc_hd__o22ai_1 U26028 ( .A1(n21199), .A2(n23348), .B1(n21102), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N3046) );
  sky130_fd_sc_hd__o22ai_1 U26029 ( .A1(n21206), .A2(n23348), .B1(n21205), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N3083) );
  sky130_fd_sc_hd__o22ai_1 U26030 ( .A1(n21182), .A2(n23348), .B1(n21072), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N2824) );
  sky130_fd_sc_hd__o22ai_1 U26031 ( .A1(n21185), .A2(n23348), .B1(n21132), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N2935) );
  sky130_fd_sc_hd__o22ai_1 U26032 ( .A1(n21183), .A2(n23348), .B1(n21133), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N2972) );
  sky130_fd_sc_hd__o22ai_1 U26033 ( .A1(n21203), .A2(n23348), .B1(n21202), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N2750) );
  sky130_fd_sc_hd__o22ai_1 U26034 ( .A1(n21186), .A2(n23348), .B1(n21134), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N3194) );
  sky130_fd_sc_hd__o22ai_1 U26035 ( .A1(n21191), .A2(n23348), .B1(n21190), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N2713) );
  sky130_fd_sc_hd__o22ai_1 U26036 ( .A1(n21189), .A2(n23348), .B1(n21188), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N3268) );
  sky130_fd_sc_hd__o22ai_1 U26037 ( .A1(n21071), .A2(n23348), .B1(n21195), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N3157) );
  sky130_fd_sc_hd__o22ai_1 U26038 ( .A1(n21070), .A2(n23348), .B1(n21194), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N2861) );
  sky130_fd_sc_hd__o22ai_1 U26039 ( .A1(n21103), .A2(n23348), .B1(n21192), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N2787) );
  sky130_fd_sc_hd__o22ai_1 U26040 ( .A1(n21069), .A2(n23348), .B1(n21193), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N3009) );
  sky130_fd_sc_hd__o22ai_1 U26041 ( .A1(n23348), .A2(n21197), .B1(n21196), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N3343) );
  sky130_fd_sc_hd__o22ai_1 U26042 ( .A1(n21187), .A2(n23348), .B1(n21073), 
        .B2(n11201), .Y(j202_soc_core_j22_cpu_rf_N3231) );
  sky130_fd_sc_hd__o22ai_1 U26043 ( .A1(n21183), .A2(n23342), .B1(n21133), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N2971) );
  sky130_fd_sc_hd__o22ai_1 U26044 ( .A1(n21184), .A2(n23342), .B1(n21068), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N3119) );
  sky130_fd_sc_hd__o22ai_1 U26045 ( .A1(n21199), .A2(n23342), .B1(n21102), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N3045) );
  sky130_fd_sc_hd__o22ai_1 U26046 ( .A1(n21185), .A2(n23342), .B1(n21132), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N2934) );
  sky130_fd_sc_hd__o22ai_1 U26047 ( .A1(n21206), .A2(n23342), .B1(n21205), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N3082) );
  sky130_fd_sc_hd__o22ai_1 U26048 ( .A1(n21201), .A2(n23342), .B1(n21200), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N2897) );
  sky130_fd_sc_hd__o22ai_1 U26049 ( .A1(n21203), .A2(n23342), .B1(n21202), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N2749) );
  sky130_fd_sc_hd__o22ai_1 U26050 ( .A1(n21186), .A2(n23342), .B1(n21134), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N3193) );
  sky130_fd_sc_hd__o22ai_1 U26051 ( .A1(n21189), .A2(n23342), .B1(n21188), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N3267) );
  sky130_fd_sc_hd__o22ai_1 U26052 ( .A1(n21191), .A2(n23342), .B1(n21190), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N2712) );
  sky130_fd_sc_hd__o22ai_1 U26053 ( .A1(n21103), .A2(n23342), .B1(n21192), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N2786) );
  sky130_fd_sc_hd__o22ai_1 U26054 ( .A1(n21070), .A2(n23342), .B1(n21194), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N2860) );
  sky130_fd_sc_hd__o22ai_1 U26055 ( .A1(n21071), .A2(n23342), .B1(n21195), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N3156) );
  sky130_fd_sc_hd__o22ai_1 U26056 ( .A1(n21069), .A2(n23342), .B1(n21193), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N3008) );
  sky130_fd_sc_hd__o22ai_1 U26057 ( .A1(n23342), .A2(n21197), .B1(n21196), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N3342) );
  sky130_fd_sc_hd__o22ai_1 U26058 ( .A1(n21182), .A2(n23342), .B1(n21072), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N2823) );
  sky130_fd_sc_hd__o22ai_1 U26059 ( .A1(n21187), .A2(n23342), .B1(n21073), 
        .B2(n11199), .Y(j202_soc_core_j22_cpu_rf_N3230) );
  sky130_fd_sc_hd__nand3_1 U26060 ( .A(n21075), .B(n25543), .C(n21074), .Y(
        n21077) );
  sky130_fd_sc_hd__nor2_1 U26061 ( .A(n21077), .B(n21076), .Y(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_N487) );
  sky130_fd_sc_hd__nand2_1 U26062 ( .A(n21765), .B(n21178), .Y(n21101) );
  sky130_fd_sc_hd__a21oi_1 U26063 ( .A1(n23326), .A2(n22606), .B1(n21143), .Y(
        n21097) );
  sky130_fd_sc_hd__nand2_1 U26065 ( .A(n21080), .B(n21141), .Y(n21096) );
  sky130_fd_sc_hd__xnor2_1 U26066 ( .A(n22574), .B(n23324), .Y(n22446) );
  sky130_fd_sc_hd__o22a_1 U26067 ( .A1(n21108), .A2(n22446), .B1(n22559), .B2(
        n21158), .X(n21084) );
  sky130_fd_sc_hd__o22ai_1 U26068 ( .A1(n23324), .A2(n21145), .B1(n22568), 
        .B2(n21155), .Y(n21082) );
  sky130_fd_sc_hd__o22ai_1 U26069 ( .A1(n22565), .A2(n21116), .B1(n22601), 
        .B2(n21154), .Y(n21081) );
  sky130_fd_sc_hd__nor2_1 U26070 ( .A(n21082), .B(n21081), .Y(n21083) );
  sky130_fd_sc_hd__o211ai_1 U26071 ( .A1(n22605), .A2(n21085), .B1(n21084), 
        .C1(n21083), .Y(n21088) );
  sky130_fd_sc_hd__a2bb2oi_1 U26072 ( .B1(n21828), .B2(n21164), .A1_N(n22610), 
        .A2_N(n21163), .Y(n21086) );
  sky130_fd_sc_hd__o211ai_1 U26073 ( .A1(n22314), .A2(n21167), .B1(n21166), 
        .C1(n21086), .Y(n21087) );
  sky130_fd_sc_hd__nor2_1 U26074 ( .A(n21088), .B(n21087), .Y(n21094) );
  sky130_fd_sc_hd__a21oi_1 U26075 ( .A1(n23324), .A2(n21089), .B1(n21146), .Y(
        n21090) );
  sky130_fd_sc_hd__nand2_1 U26077 ( .A(n21092), .B(n22574), .Y(n21093) );
  sky130_fd_sc_hd__o211ai_1 U26078 ( .A1(n23326), .A2(n21174), .B1(n21094), 
        .C1(n21093), .Y(n21095) );
  sky130_fd_sc_hd__a21oi_1 U26079 ( .A1(n21097), .A2(n21096), .B1(n21095), .Y(
        n21100) );
  sky130_fd_sc_hd__nand2_1 U26080 ( .A(n21098), .B(n21137), .Y(n21099) );
  sky130_fd_sc_hd__nand3_1 U26081 ( .A(n21101), .B(n21100), .C(n21099), .Y(
        n21761) );
  sky130_fd_sc_hd__o22ai_1 U26082 ( .A1(n21184), .A2(n23326), .B1(n21068), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N3113) );
  sky130_fd_sc_hd__o22ai_1 U26083 ( .A1(n21199), .A2(n23326), .B1(n21102), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N3039) );
  sky130_fd_sc_hd__o22ai_1 U26084 ( .A1(n21185), .A2(n23326), .B1(n21132), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N2928) );
  sky130_fd_sc_hd__o22ai_1 U26085 ( .A1(n21206), .A2(n23326), .B1(n21205), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N3076) );
  sky130_fd_sc_hd__o22ai_1 U26086 ( .A1(n21201), .A2(n23326), .B1(n21200), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N2891) );
  sky130_fd_sc_hd__o22ai_1 U26087 ( .A1(n21183), .A2(n23326), .B1(n21133), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N2965) );
  sky130_fd_sc_hd__o22ai_1 U26088 ( .A1(n21182), .A2(n23326), .B1(n21072), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N2817) );
  sky130_fd_sc_hd__o22ai_1 U26089 ( .A1(n21187), .A2(n23326), .B1(n21073), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N3224) );
  sky130_fd_sc_hd__o22ai_1 U26090 ( .A1(n21186), .A2(n23326), .B1(n21134), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N3187) );
  sky130_fd_sc_hd__o22ai_1 U26091 ( .A1(n21203), .A2(n23326), .B1(n21202), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N2743) );
  sky130_fd_sc_hd__o22ai_1 U26092 ( .A1(n21191), .A2(n23326), .B1(n21190), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N2706) );
  sky130_fd_sc_hd__o22ai_1 U26093 ( .A1(n21189), .A2(n23326), .B1(n21188), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N3261) );
  sky130_fd_sc_hd__o22ai_1 U26094 ( .A1(n21069), .A2(n23326), .B1(n21193), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N3002) );
  sky130_fd_sc_hd__o22ai_1 U26095 ( .A1(n21103), .A2(n23326), .B1(n21192), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N2780) );
  sky130_fd_sc_hd__o22ai_1 U26096 ( .A1(n21071), .A2(n23326), .B1(n21195), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N3150) );
  sky130_fd_sc_hd__o22ai_1 U26097 ( .A1(n21070), .A2(n23326), .B1(n21194), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N2854) );
  sky130_fd_sc_hd__o22ai_1 U26098 ( .A1(n23326), .A2(n21197), .B1(n21196), 
        .B2(n21764), .Y(j202_soc_core_j22_cpu_rf_N3337) );
  sky130_fd_sc_hd__nand2_1 U26099 ( .A(n21105), .B(n21137), .Y(n21130) );
  sky130_fd_sc_hd__nand2_1 U26100 ( .A(n21839), .B(n21178), .Y(n21129) );
  sky130_fd_sc_hd__nor2_1 U26101 ( .A(n22568), .B(n21937), .Y(n21122) );
  sky130_fd_sc_hd__nand2_1 U26102 ( .A(n21106), .B(n21139), .Y(n21107) );
  sky130_fd_sc_hd__nand2_1 U26103 ( .A(n21107), .B(n21141), .Y(n21127) );
  sky130_fd_sc_hd__a21oi_1 U26104 ( .A1(n21937), .A2(n22568), .B1(n21143), .Y(
        n21126) );
  sky130_fd_sc_hd__nand2_1 U26105 ( .A(n21144), .B(n23322), .Y(n21115) );
  sky130_fd_sc_hd__nor2_1 U26106 ( .A(n21935), .B(n23322), .Y(n22451) );
  sky130_fd_sc_hd__nor2_1 U26107 ( .A(n21108), .B(n22451), .Y(n21111) );
  sky130_fd_sc_hd__nand2_1 U26108 ( .A(n23322), .B(n21935), .Y(n22632) );
  sky130_fd_sc_hd__a2bb2oi_1 U26109 ( .B1(n21146), .B2(n21935), .A1_N(n21145), 
        .A2_N(n23322), .Y(n21109) );
  sky130_fd_sc_hd__a21oi_1 U26111 ( .A1(n21111), .A2(n22632), .B1(n21110), .Y(
        n21114) );
  sky130_fd_sc_hd__o22a_1 U26112 ( .A1(n22614), .A2(n21155), .B1(n22606), .B2(
        n21154), .X(n21113) );
  sky130_fd_sc_hd__nand2_1 U26113 ( .A(n21164), .B(n21867), .Y(n21112) );
  sky130_fd_sc_hd__nand4_1 U26114 ( .A(n21115), .B(n21114), .C(n21113), .D(
        n21112), .Y(n21121) );
  sky130_fd_sc_hd__o22ai_1 U26115 ( .A1(n22563), .A2(n21116), .B1(n22558), 
        .B2(n21158), .Y(n21117) );
  sky130_fd_sc_hd__a21oi_1 U26116 ( .A1(n21118), .A2(n22573), .B1(n21117), .Y(
        n21119) );
  sky130_fd_sc_hd__o211ai_1 U26117 ( .A1(n21929), .A2(n21167), .B1(n21166), 
        .C1(n21119), .Y(n21120) );
  sky130_fd_sc_hd__nor2_1 U26118 ( .A(n21121), .B(n21120), .Y(n21124) );
  sky130_fd_sc_hd__nand2_1 U26119 ( .A(n21122), .B(n21170), .Y(n21123) );
  sky130_fd_sc_hd__o211ai_1 U26120 ( .A1(n21937), .A2(n21174), .B1(n21124), 
        .C1(n21123), .Y(n21125) );
  sky130_fd_sc_hd__a21oi_1 U26121 ( .A1(n21127), .A2(n21126), .B1(n21125), .Y(
        n21128) );
  sky130_fd_sc_hd__nand3_1 U26122 ( .A(n21130), .B(n21129), .C(n21128), .Y(
        n21834) );
  sky130_fd_sc_hd__o22ai_1 U26123 ( .A1(n21184), .A2(n21937), .B1(n21068), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N3112) );
  sky130_fd_sc_hd__o22ai_1 U26124 ( .A1(n21182), .A2(n21937), .B1(n21072), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N2816) );
  sky130_fd_sc_hd__o22ai_1 U26125 ( .A1(n21187), .A2(n21937), .B1(n21073), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N3223) );
  sky130_fd_sc_hd__o22ai_1 U26126 ( .A1(n21189), .A2(n21937), .B1(n21188), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N3260) );
  sky130_fd_sc_hd__o22ai_1 U26127 ( .A1(n21191), .A2(n21937), .B1(n21190), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N2705) );
  sky130_fd_sc_hd__o22ai_1 U26128 ( .A1(n21071), .A2(n21937), .B1(n21195), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N3149) );
  sky130_fd_sc_hd__o22ai_1 U26129 ( .A1(n21103), .A2(n21937), .B1(n21192), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N2779) );
  sky130_fd_sc_hd__o22ai_1 U26130 ( .A1(n21069), .A2(n21937), .B1(n21193), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N3001) );
  sky130_fd_sc_hd__o22ai_1 U26131 ( .A1(n21070), .A2(n21937), .B1(n21194), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N2853) );
  sky130_fd_sc_hd__nand2_1 U26132 ( .A(n22829), .B(n22827), .Y(n21131) );
  sky130_fd_sc_hd__nand3_1 U26133 ( .A(n21904), .B(n21208), .C(n21131), .Y(
        j202_soc_core_ahb2aqu_00_N128) );
  sky130_fd_sc_hd__o22ai_1 U26134 ( .A1(n21937), .A2(n21197), .B1(n21196), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N3336) );
  sky130_fd_sc_hd__o22ai_1 U26135 ( .A1(n21185), .A2(n21937), .B1(n21132), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N2927) );
  sky130_fd_sc_hd__o22ai_1 U26136 ( .A1(n21199), .A2(n21937), .B1(n21198), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N3038) );
  sky130_fd_sc_hd__o22ai_1 U26137 ( .A1(n21201), .A2(n21937), .B1(n21200), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N2890) );
  sky130_fd_sc_hd__o22ai_1 U26138 ( .A1(n21183), .A2(n21937), .B1(n21133), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N2964) );
  sky130_fd_sc_hd__o22ai_1 U26139 ( .A1(n21186), .A2(n21937), .B1(n21134), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N3186) );
  sky130_fd_sc_hd__o22ai_1 U26140 ( .A1(n21203), .A2(n21937), .B1(n21202), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N2742) );
  sky130_fd_sc_hd__o22ai_1 U26141 ( .A1(n21206), .A2(n21937), .B1(n21205), 
        .B2(n21838), .Y(j202_soc_core_j22_cpu_rf_N3075) );
  sky130_fd_sc_hd__nand2b_1 U26142 ( .A_N(n21138), .B(n21137), .Y(n21181) );
  sky130_fd_sc_hd__nor2_1 U26143 ( .A(n22567), .B(n23318), .Y(n21171) );
  sky130_fd_sc_hd__nand2_1 U26144 ( .A(n21140), .B(n21139), .Y(n21142) );
  sky130_fd_sc_hd__nand2_1 U26145 ( .A(n21142), .B(n21141), .Y(n21177) );
  sky130_fd_sc_hd__a21oi_1 U26146 ( .A1(n23318), .A2(n22567), .B1(n21143), .Y(
        n21176) );
  sky130_fd_sc_hd__nand2_1 U26147 ( .A(n21144), .B(n23316), .Y(n21162) );
  sky130_fd_sc_hd__nand2_1 U26148 ( .A(n23316), .B(n21867), .Y(n22634) );
  sky130_fd_sc_hd__a2bb2oi_1 U26149 ( .B1(n21146), .B2(n21867), .A1_N(n21145), 
        .A2_N(n23316), .Y(n21149) );
  sky130_fd_sc_hd__nand2_1 U26150 ( .A(n21878), .B(n22567), .Y(n22458) );
  sky130_fd_sc_hd__nand3_1 U26151 ( .A(n22458), .B(n21147), .C(n22634), .Y(
        n21148) );
  sky130_fd_sc_hd__o211ai_1 U26152 ( .A1(n21150), .A2(n22634), .B1(n21149), 
        .C1(n21148), .Y(n21151) );
  sky130_fd_sc_hd__a21oi_1 U26153 ( .A1(n21153), .A2(n21152), .B1(n21151), .Y(
        n21161) );
  sky130_fd_sc_hd__o22a_1 U26154 ( .A1(n22600), .A2(n21155), .B1(n22614), .B2(
        n21154), .X(n21160) );
  sky130_fd_sc_hd__o22a_1 U26155 ( .A1(n22612), .A2(n21158), .B1(n22604), .B2(
        n21157), .X(n21159) );
  sky130_fd_sc_hd__nand4_1 U26156 ( .A(n21162), .B(n21161), .C(n21160), .D(
        n21159), .Y(n21169) );
  sky130_fd_sc_hd__a2bb2oi_1 U26157 ( .B1(n22577), .B2(n21164), .A1_N(n22568), 
        .A2_N(n21163), .Y(n21165) );
  sky130_fd_sc_hd__o211ai_1 U26158 ( .A1(n22611), .A2(n21167), .B1(n21166), 
        .C1(n21165), .Y(n21168) );
  sky130_fd_sc_hd__nor2_1 U26159 ( .A(n21169), .B(n21168), .Y(n21173) );
  sky130_fd_sc_hd__nand2_1 U26160 ( .A(n21171), .B(n21170), .Y(n21172) );
  sky130_fd_sc_hd__o211ai_1 U26161 ( .A1(n23318), .A2(n21174), .B1(n21173), 
        .C1(n21172), .Y(n21175) );
  sky130_fd_sc_hd__a21oi_1 U26162 ( .A1(n21177), .A2(n21176), .B1(n21175), .Y(
        n21180) );
  sky130_fd_sc_hd__nand2_1 U26163 ( .A(n21877), .B(n21178), .Y(n21179) );
  sky130_fd_sc_hd__o22ai_1 U26164 ( .A1(n23318), .A2(n21182), .B1(n21072), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N2814) );
  sky130_fd_sc_hd__o22ai_1 U26165 ( .A1(n23318), .A2(n21183), .B1(n21133), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N2962) );
  sky130_fd_sc_hd__o22ai_1 U26166 ( .A1(n23318), .A2(n21184), .B1(n21068), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N3110) );
  sky130_fd_sc_hd__o22ai_1 U26167 ( .A1(n23318), .A2(n21185), .B1(n21132), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N2925) );
  sky130_fd_sc_hd__o22ai_1 U26168 ( .A1(n23318), .A2(n21186), .B1(n21134), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N3184) );
  sky130_fd_sc_hd__o22ai_1 U26169 ( .A1(n23318), .A2(n21187), .B1(n21073), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N3221) );
  sky130_fd_sc_hd__o22ai_1 U26170 ( .A1(n23318), .A2(n21189), .B1(n21188), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N3258) );
  sky130_fd_sc_hd__o22ai_1 U26171 ( .A1(n23318), .A2(n21191), .B1(n21190), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N2703) );
  sky130_fd_sc_hd__o22ai_1 U26172 ( .A1(n23318), .A2(n21103), .B1(n21192), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N2777) );
  sky130_fd_sc_hd__o22ai_1 U26173 ( .A1(n23318), .A2(n21069), .B1(n21193), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N2999) );
  sky130_fd_sc_hd__o22ai_1 U26174 ( .A1(n23318), .A2(n21070), .B1(n21194), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N2851) );
  sky130_fd_sc_hd__o22ai_1 U26175 ( .A1(n23318), .A2(n21071), .B1(n21195), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N3147) );
  sky130_fd_sc_hd__o22ai_1 U26176 ( .A1(n23318), .A2(n21197), .B1(n21196), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N3334) );
  sky130_fd_sc_hd__o22ai_1 U26177 ( .A1(n23318), .A2(n21199), .B1(n21198), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N3036) );
  sky130_fd_sc_hd__o22ai_1 U26178 ( .A1(n23318), .A2(n21201), .B1(n21200), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N2888) );
  sky130_fd_sc_hd__o22ai_1 U26179 ( .A1(n23318), .A2(n21203), .B1(n21202), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N2740) );
  sky130_fd_sc_hd__o22ai_1 U26180 ( .A1(n23318), .A2(n21206), .B1(n21205), 
        .B2(n21204), .Y(j202_soc_core_j22_cpu_rf_N3073) );
  sky130_fd_sc_hd__nor2_1 U26181 ( .A(n23250), .B(n21207), .Y(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_N497) );
  sky130_fd_sc_hd__nand2_1 U26182 ( .A(n21208), .B(n22403), .Y(n21209) );
  sky130_fd_sc_hd__nor2_1 U26183 ( .A(n22825), .B(n21210), .Y(
        j202_soc_core_ahb2aqu_00_N131) );
  sky130_fd_sc_hd__nor2_1 U26184 ( .A(n22816), .B(n21210), .Y(
        j202_soc_core_ahb2aqu_00_N130) );
  sky130_fd_sc_hd__nor2_1 U26185 ( .A(n22817), .B(n21210), .Y(
        j202_soc_core_ahb2aqu_00_N129) );
  sky130_fd_sc_hd__nor2_1 U26186 ( .A(n22819), .B(n21210), .Y(
        j202_soc_core_ahb2aqu_00_N136) );
  sky130_fd_sc_hd__nor2_1 U26187 ( .A(n22820), .B(n21210), .Y(
        j202_soc_core_ahb2aqu_00_N134) );
  sky130_fd_sc_hd__nor2_1 U26188 ( .A(n22818), .B(n21210), .Y(
        j202_soc_core_ahb2aqu_00_N135) );
  sky130_fd_sc_hd__nor2_1 U26189 ( .A(n22823), .B(n21210), .Y(
        j202_soc_core_ahb2aqu_00_N132) );
  sky130_fd_sc_hd__nor2_1 U26190 ( .A(n22822), .B(n21210), .Y(
        j202_soc_core_ahb2aqu_00_N133) );
  sky130_fd_sc_hd__nand3_1 U26191 ( .A(n21213), .B(n21212), .C(n21211), .Y(
        n21214) );
  sky130_fd_sc_hd__a21o_1 U26192 ( .A1(n22816), .A2(n21215), .B1(n21214), .X(
        n21906) );
  sky130_fd_sc_hd__or3_1 U26193 ( .A(j202_soc_core_rst), .B(n21217), .C(n21216), .X(n25433) );
  sky130_fd_sc_hd__and3_1 U26194 ( .A(n25339), .B(n21219), .C(n21218), .X(
        n25436) );
  sky130_fd_sc_hd__nand2_1 U26195 ( .A(n23242), .B(
        j202_soc_core_j22_cpu_memop_MEM__2_), .Y(n21221) );
  sky130_fd_sc_hd__nor2_1 U26196 ( .A(n21221), .B(n21220), .Y(n21223) );
  sky130_fd_sc_hd__nor2_1 U26197 ( .A(n21223), .B(n21222), .Y(n21250) );
  sky130_fd_sc_hd__and3_1 U26199 ( .A(n25340), .B(n21225), .C(n21224), .X(
        n25463) );
  sky130_fd_sc_hd__nand2_1 U26200 ( .A(n22860), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd), .Y(n23600) );
  sky130_fd_sc_hd__nand2_1 U26201 ( .A(n25392), .B(
        j202_soc_core_wbqspiflash_00_spi_spd), .Y(n21226) );
  sky130_fd_sc_hd__and3_1 U26202 ( .A(n23600), .B(n21226), .C(n23588), .X(
        n25482) );
  sky130_fd_sc_hd__and3_1 U26203 ( .A(n21228), .B(n21227), .C(
        j202_soc_core_aquc_WE_), .X(n25483) );
  sky130_fd_sc_hd__nor2_1 U26204 ( .A(j202_soc_core_ahb2apb_01_state[2]), .B(
        j202_soc_core_rst), .Y(n21230) );
  sky130_fd_sc_hd__and3_1 U26205 ( .A(n21230), .B(
        j202_soc_core_ahb2apb_01_state[0]), .C(n21229), .X(n25484) );
  sky130_fd_sc_hd__and3_1 U26206 ( .A(n21230), .B(
        j202_soc_core_ahb2apb_01_state[1]), .C(
        j202_soc_core_ahb2apb_01_state[0]), .X(n25485) );
  sky130_fd_sc_hd__nor2_1 U26207 ( .A(j202_soc_core_ahb2apb_02_state[2]), .B(
        j202_soc_core_rst), .Y(n21232) );
  sky130_fd_sc_hd__and3_1 U26208 ( .A(n21232), .B(
        j202_soc_core_ahb2apb_02_state[0]), .C(n21231), .X(n25486) );
  sky130_fd_sc_hd__and3_1 U26209 ( .A(n21232), .B(
        j202_soc_core_ahb2apb_02_state[1]), .C(
        j202_soc_core_ahb2apb_02_state[0]), .X(n25487) );
  sky130_fd_sc_hd__nand2_1 U26210 ( .A(n23747), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[1]), .Y(n22863) );
  sky130_fd_sc_hd__nand2_1 U26211 ( .A(n23747), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[0]), .Y(n22867) );
  sky130_fd_sc_hd__nand2_1 U26212 ( .A(n25392), .B(n23735), .Y(n22861) );
  sky130_fd_sc_hd__clkinv_1 U26213 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd), .Y(n21233) );
  sky130_fd_sc_hd__nand2_1 U26214 ( .A(n22860), .B(n21233), .Y(n23602) );
  sky130_fd_sc_hd__o211ai_1 U26215 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd), .A2(n21234), .B1(n22861), 
        .C1(n23602), .Y(n22868) );
  sky130_fd_sc_hd__nand2_1 U26216 ( .A(n22867), .B(n22868), .Y(n22866) );
  sky130_fd_sc_hd__nand2_1 U26217 ( .A(n22863), .B(n21235), .Y(
        DP_OP_1501J1_126_8405_n4) );
  sky130_fd_sc_hd__nand3_1 U26218 ( .A(n21236), .B(n25734), .C(n21997), .Y(
        n25489) );
  sky130_fd_sc_hd__nor2_1 U26219 ( .A(n21237), .B(n22816), .Y(n21907) );
  sky130_fd_sc_hd__nand2b_1 U26220 ( .A_N(n21253), .B(n21238), .Y(n21242) );
  sky130_fd_sc_hd__nor2_1 U26221 ( .A(n21241), .B(n25379), .Y(n21321) );
  sky130_fd_sc_hd__nand3_1 U26222 ( .A(n21246), .B(n21245), .C(n21244), .Y(
        n21913) );
  sky130_fd_sc_hd__o22ai_1 U26223 ( .A1(n21908), .A2(n21252), .B1(n21251), 
        .B2(n22816), .Y(n22828) );
  sky130_fd_sc_hd__a21oi_1 U26224 ( .A1(n25391), .A2(n25379), .B1(n22828), .Y(
        n21254) );
  sky130_fd_sc_hd__nor2_1 U26225 ( .A(n25109), .B(n25107), .Y(n21256) );
  sky130_fd_sc_hd__nand2_1 U26226 ( .A(j202_soc_core_wbqspiflash_00_spi_wr), 
        .B(n21256), .Y(n25119) );
  sky130_fd_sc_hd__o21ai_1 U26227 ( .A1(j202_soc_core_rst), .A2(n25119), .B1(
        n20219), .Y(n25494) );
  sky130_fd_sc_hd__buf_4 U26228 ( .A(n21300), .X(n25515) );
  sky130_fd_sc_hd__or2b_4 U26229 ( .A(n11036), .B_N(n25488), .X(n10539) );
  sky130_fd_sc_hd__a21oi_1 U26230 ( .A1(n21321), .A2(n25391), .B1(n22828), .Y(
        n21322) );
  sky130_fd_sc_hd__nand2_1 U26231 ( .A(n21324), .B(n23587), .Y(n23608) );
  sky130_fd_sc_hd__nand4_1 U26232 ( .A(n23731), .B(n22862), .C(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .D(n23608), .Y(n25527) );
  sky130_fd_sc_hd__nand2_1 U26233 ( .A(n25734), .B(n23731), .Y(n25528) );
  sky130_fd_sc_hd__nand2_1 U26234 ( .A(n25734), .B(n23699), .Y(n25529) );
  sky130_fd_sc_hd__nand2_1 U26235 ( .A(n21325), .B(n25122), .Y(
        j202_soc_core_uart_TOP_N24) );
  sky130_fd_sc_hd__nand2_1 U26236 ( .A(n25734), .B(n24069), .Y(n25530) );
  sky130_fd_sc_hd__nand2_1 U26237 ( .A(n24867), .B(n25387), .Y(n23223) );
  sky130_fd_sc_hd__nand4_1 U26238 ( .A(n24861), .B(n24860), .C(n24884), .D(
        n23223), .Y(n21326) );
  sky130_fd_sc_hd__nor3_1 U26240 ( .A(n21329), .B(n22336), .C(n22802), .Y(
        n23232) );
  sky130_fd_sc_hd__nand2_1 U26241 ( .A(n21331), .B(n21330), .Y(n21549) );
  sky130_fd_sc_hd__o21ai_1 U26242 ( .A1(n25369), .A2(n22412), .B1(n21549), .Y(
        n21335) );
  sky130_fd_sc_hd__nand2_1 U26243 ( .A(n21582), .B(n21332), .Y(n22739) );
  sky130_fd_sc_hd__nor4b_1 U26245 ( .D_N(n23220), .A(n24828), .B(n21335), .C(
        n21334), .Y(n24868) );
  sky130_fd_sc_hd__a21oi_1 U26246 ( .A1(n21336), .A2(n24825), .B1(n21482), .Y(
        n21337) );
  sky130_fd_sc_hd__a31oi_1 U26247 ( .A1(n24868), .A2(n21337), .A3(n22797), 
        .B1(n24882), .Y(n22787) );
  sky130_fd_sc_hd__nor2_1 U26248 ( .A(j202_soc_core_rst), .B(n23229), .Y(
        n24893) );
  sky130_fd_sc_hd__nor3_1 U26249 ( .A(n23232), .B(n22787), .C(n23238), .Y(
        n21340) );
  sky130_fd_sc_hd__a21o_1 U26250 ( .A1(n21339), .A2(n21338), .B1(n22401), .X(
        n23221) );
  sky130_fd_sc_hd__nand4_1 U26251 ( .A(n21341), .B(n21340), .C(n23221), .D(
        n21644), .Y(n10566) );
  sky130_fd_sc_hd__nand2_1 U26252 ( .A(n21388), .B(n25731), .Y(n22785) );
  sky130_fd_sc_hd__o22ai_1 U26253 ( .A1(n21365), .A2(n21381), .B1(n21385), 
        .B2(n21377), .Y(n21342) );
  sky130_fd_sc_hd__a22o_1 U26254 ( .A1(n25390), .A2(n21366), .B1(n21393), .B2(
        n21342), .X(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N5) );
  sky130_fd_sc_hd__o21ai_0 U26255 ( .A1(n21365), .A2(n22785), .B1(n21344), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N6) );
  sky130_fd_sc_hd__o22ai_1 U26256 ( .A1(n21347), .A2(n21346), .B1(n21379), 
        .B2(n21345), .Y(n21352) );
  sky130_fd_sc_hd__o2bb2ai_1 U26257 ( .B1(n21350), .B2(n21349), .A1_N(n21350), 
        .A2_N(n21348), .Y(n21351) );
  sky130_fd_sc_hd__o22ai_1 U26258 ( .A1(n21353), .A2(n21352), .B1(n21381), 
        .B2(n21351), .Y(n21364) );
  sky130_fd_sc_hd__a22o_1 U26259 ( .A1(n21356), .A2(n21378), .B1(n21355), .B2(
        n21354), .X(n21362) );
  sky130_fd_sc_hd__o2bb2ai_1 U26260 ( .B1(n21359), .B2(n21358), .A1_N(n21359), 
        .A2_N(n21357), .Y(n21360) );
  sky130_fd_sc_hd__o22ai_1 U26261 ( .A1(n21377), .A2(n21362), .B1(n21361), 
        .B2(n21360), .Y(n21363) );
  sky130_fd_sc_hd__o22ai_1 U26262 ( .A1(n21365), .A2(n21364), .B1(n21385), 
        .B2(n21363), .Y(n21374) );
  sky130_fd_sc_hd__nand2_1 U26263 ( .A(n21367), .B(n25731), .Y(n21389) );
  sky130_fd_sc_hd__nand2_1 U26264 ( .A(n21387), .B(n21369), .Y(n21370) );
  sky130_fd_sc_hd__nor3_1 U26266 ( .A(n21389), .B(n21372), .C(n21388), .Y(
        n21373) );
  sky130_fd_sc_hd__a211o_1 U26267 ( .A1(n21393), .A2(n21374), .B1(n25370), 
        .C1(n21373), .X(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N3) );
  sky130_fd_sc_hd__nand2_1 U26268 ( .A(n21377), .B(n21375), .Y(n21376) );
  sky130_fd_sc_hd__o21ai_1 U26269 ( .A1(n21378), .A2(n21377), .B1(n21376), .Y(
        n21386) );
  sky130_fd_sc_hd__nand2_1 U26270 ( .A(n21379), .B(n21381), .Y(n21380) );
  sky130_fd_sc_hd__nand2_1 U26272 ( .A(n21383), .B(n21385), .Y(n21384) );
  sky130_fd_sc_hd__o21ai_1 U26273 ( .A1(n21386), .A2(n21385), .B1(n21384), .Y(
        n21392) );
  sky130_fd_sc_hd__nor3_1 U26274 ( .A(n21390), .B(n21389), .C(n21388), .Y(
        n21391) );
  sky130_fd_sc_hd__a211o_1 U26275 ( .A1(n21393), .A2(n21392), .B1(n25370), 
        .C1(n21391), .X(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_vec_N4) );
  sky130_fd_sc_hd__or3_1 U26276 ( .A(j202_soc_core_intr_vec__4_), .B(
        j202_soc_core_intr_vec__0_), .C(j202_soc_core_intr_vec__6_), .X(n21394) );
  sky130_fd_sc_hd__nor3_1 U26277 ( .A(j202_soc_core_intr_vec__2_), .B(
        j202_soc_core_intr_vec__3_), .C(n21394), .Y(n23228) );
  sky130_fd_sc_hd__clkinv_1 U26278 ( .A(n21395), .Y(n21396) );
  sky130_fd_sc_hd__nand2_1 U26279 ( .A(n24879), .B(n21396), .Y(n24885) );
  sky130_fd_sc_hd__a31oi_1 U26280 ( .A1(j202_soc_core_j22_cpu_opst[1]), .A2(
        n23228), .A3(n22899), .B1(n24885), .Y(
        j202_soc_core_j22_cpu_id_idec_N822) );
  sky130_fd_sc_hd__nand2_1 U26281 ( .A(n21398), .B(n25731), .Y(n22906) );
  sky130_fd_sc_hd__a211oi_1 U26282 ( .A1(n21400), .A2(n21399), .B1(
        j202_soc_core_intc_core_00_cp_intack_all_0_), .C1(n22906), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_intr_req_N3) );
  sky130_fd_sc_hd__o21ai_1 U26283 ( .A1(n22330), .A2(n21402), .B1(n21401), .Y(
        n21421) );
  sky130_fd_sc_hd__nand2_1 U26284 ( .A(n21403), .B(n21564), .Y(n21425) );
  sky130_fd_sc_hd__nand3_1 U26285 ( .A(n21504), .B(n21425), .C(n21404), .Y(
        n21405) );
  sky130_fd_sc_hd__o31ai_1 U26286 ( .A1(n21406), .A2(n21421), .A3(n21405), 
        .B1(n24858), .Y(n21407) );
  sky130_fd_sc_hd__o21ai_1 U26287 ( .A1(n21408), .A2(n22401), .B1(n21407), .Y(
        n10501) );
  sky130_fd_sc_hd__nand2_1 U26288 ( .A(n21410), .B(n21409), .Y(n21434) );
  sky130_fd_sc_hd__a21oi_1 U26289 ( .A1(n21412), .A2(n21563), .B1(n21411), .Y(
        n22331) );
  sky130_fd_sc_hd__nand3_1 U26290 ( .A(n21414), .B(n22331), .C(n21413), .Y(
        n21415) );
  sky130_fd_sc_hd__a21oi_1 U26291 ( .A1(n21416), .A2(n21434), .B1(n21415), .Y(
        n21451) );
  sky130_fd_sc_hd__nor3_1 U26292 ( .A(n24872), .B(n21418), .C(n21417), .Y(
        n21419) );
  sky130_fd_sc_hd__a31oi_1 U26293 ( .A1(n21420), .A2(n21563), .A3(n22733), 
        .B1(n21419), .Y(n21463) );
  sky130_fd_sc_hd__a21oi_1 U26294 ( .A1(n22733), .A2(n21422), .B1(n21421), .Y(
        n21429) );
  sky130_fd_sc_hd__nand2_1 U26295 ( .A(n21506), .B(n21801), .Y(n21423) );
  sky130_fd_sc_hd__a21oi_1 U26296 ( .A1(n21424), .A2(n25387), .B1(n21423), .Y(
        n21516) );
  sky130_fd_sc_hd__nand3_1 U26297 ( .A(n21516), .B(n21556), .C(n21425), .Y(
        n21477) );
  sky130_fd_sc_hd__nor4_1 U26298 ( .A(n21427), .B(n24867), .C(n21477), .D(
        n21426), .Y(n21428) );
  sky130_fd_sc_hd__nand4_1 U26299 ( .A(n21451), .B(n21463), .C(n21429), .D(
        n21428), .Y(n21446) );
  sky130_fd_sc_hd__nand2_1 U26300 ( .A(n21431), .B(n21430), .Y(n22107) );
  sky130_fd_sc_hd__o21a_1 U26301 ( .A1(n22390), .A2(n21568), .B1(n22797), .X(
        n21596) );
  sky130_fd_sc_hd__o21ai_1 U26302 ( .A1(n22332), .A2(n21432), .B1(n21596), .Y(
        n21433) );
  sky130_fd_sc_hd__a211oi_1 U26303 ( .A1(n21435), .A2(n21434), .B1(n24830), 
        .C1(n21433), .Y(n21450) );
  sky130_fd_sc_hd__nand2_1 U26304 ( .A(n21436), .B(n21450), .Y(n21437) );
  sky130_fd_sc_hd__o31ai_1 U26305 ( .A1(n21446), .A2(n21438), .A3(n21437), 
        .B1(n24858), .Y(n21439) );
  sky130_fd_sc_hd__o21ai_1 U26306 ( .A1(n21440), .A2(n22401), .B1(n21439), .Y(
        n10570) );
  sky130_fd_sc_hd__nand2_1 U26307 ( .A(n24878), .B(n21441), .Y(n21442) );
  sky130_fd_sc_hd__nand2_1 U26309 ( .A(n24879), .B(n21444), .Y(n21471) );
  sky130_fd_sc_hd__o21ai_1 U26310 ( .A1(j202_soc_core_j22_cpu_opst[0]), .A2(
        n21471), .B1(n24844), .Y(n21445) );
  sky130_fd_sc_hd__a211o_1 U26311 ( .A1(n21446), .A2(n24858), .B1(n24835), 
        .C1(n21445), .X(j202_soc_core_j22_cpu_id_idec_N937) );
  sky130_fd_sc_hd__a21oi_1 U26312 ( .A1(n24884), .A2(n21447), .B1(n24882), .Y(
        n21448) );
  sky130_fd_sc_hd__nor2_1 U26313 ( .A(n25371), .B(n21448), .Y(n21449) );
  sky130_fd_sc_hd__a21o_1 U26315 ( .A1(n21451), .A2(n21450), .B1(n24882), .X(
        n21453) );
  sky130_fd_sc_hd__nand2_1 U26316 ( .A(n21453), .B(n21452), .Y(n10589) );
  sky130_fd_sc_hd__nand2_1 U26317 ( .A(n22330), .B(n21454), .Y(n22408) );
  sky130_fd_sc_hd__a21oi_1 U26318 ( .A1(n21456), .A2(n22408), .B1(n21455), .Y(
        n21460) );
  sky130_fd_sc_hd__o21ai_1 U26319 ( .A1(n22743), .A2(n21457), .B1(n24884), .Y(
        n21458) );
  sky130_fd_sc_hd__nor4_1 U26320 ( .A(n21461), .B(n21460), .C(n21459), .D(
        n21458), .Y(n21462) );
  sky130_fd_sc_hd__nand2_1 U26321 ( .A(j202_soc_core_j22_cpu_opst[0]), .B(
        n21465), .Y(n21466) );
  sky130_fd_sc_hd__nor2_1 U26322 ( .A(n22402), .B(n22401), .Y(n21468) );
  sky130_fd_sc_hd__a21oi_1 U26323 ( .A1(n24858), .A2(n21469), .B1(n21468), .Y(
        n21470) );
  sky130_fd_sc_hd__o211ai_1 U26324 ( .A1(n22416), .A2(n22417), .B1(n21644), 
        .C1(n21470), .Y(n10588) );
  sky130_fd_sc_hd__nand2b_1 U26325 ( .A_N(n21473), .B(n24858), .Y(n24843) );
  sky130_fd_sc_hd__nand2_1 U26326 ( .A(n21490), .B(n21583), .Y(n21559) );
  sky130_fd_sc_hd__a21oi_1 U26327 ( .A1(n24858), .A2(n24833), .B1(n21559), .Y(
        n21472) );
  sky130_fd_sc_hd__nand4_1 U26328 ( .A(n24843), .B(n21472), .C(n24874), .D(
        n21471), .Y(n10500) );
  sky130_fd_sc_hd__nor4_1 U26330 ( .A(n21589), .B(n21477), .C(n21476), .D(
        n21475), .Y(n21479) );
  sky130_fd_sc_hd__nor2_1 U26331 ( .A(n24863), .B(n21501), .Y(n21478) );
  sky130_fd_sc_hd__o21ai_1 U26332 ( .A1(n24882), .A2(n21479), .B1(n21478), .Y(
        n10600) );
  sky130_fd_sc_hd__nand2_1 U26333 ( .A(n21592), .B(n21599), .Y(n10604) );
  sky130_fd_sc_hd__nor4_1 U26335 ( .A(n21482), .B(n21589), .C(n21494), .D(
        n21481), .Y(n21484) );
  sky130_fd_sc_hd__nor2_1 U26336 ( .A(n21501), .B(n21483), .Y(n22340) );
  sky130_fd_sc_hd__o21ai_1 U26337 ( .A1(n21484), .A2(n24882), .B1(n22340), .Y(
        n10576) );
  sky130_fd_sc_hd__nor3_1 U26339 ( .A(n21573), .B(n21572), .C(n21486), .Y(
        n21641) );
  sky130_fd_sc_hd__nand2_1 U26340 ( .A(n21487), .B(n21641), .Y(n22395) );
  sky130_fd_sc_hd__nand2_1 U26341 ( .A(n21580), .B(n22395), .Y(n21488) );
  sky130_fd_sc_hd__nor4_1 U26342 ( .A(n21608), .B(n21489), .C(n21571), .D(
        n21488), .Y(n21491) );
  sky130_fd_sc_hd__o21ai_1 U26343 ( .A1(n24882), .A2(n21491), .B1(n21490), .Y(
        n10596) );
  sky130_fd_sc_hd__nor2_1 U26344 ( .A(n21492), .B(n24841), .Y(n24829) );
  sky130_fd_sc_hd__nand4b_1 U26345 ( .A_N(n21494), .B(n22332), .C(n21493), .D(
        n24829), .Y(n21495) );
  sky130_fd_sc_hd__nor4_1 U26346 ( .A(n21498), .B(n21497), .C(n21496), .D(
        n21495), .Y(n21503) );
  sky130_fd_sc_hd__a21oi_1 U26347 ( .A1(n22402), .A2(n21499), .B1(n22401), .Y(
        n21500) );
  sky130_fd_sc_hd__nor2_1 U26348 ( .A(n21501), .B(n21500), .Y(n21502) );
  sky130_fd_sc_hd__o21ai_1 U26349 ( .A1(n21607), .A2(n21503), .B1(n21502), .Y(
        n10580) );
  sky130_fd_sc_hd__nor2_1 U26350 ( .A(n21505), .B(n22409), .Y(n24853) );
  sky130_fd_sc_hd__nand4_1 U26351 ( .A(n21507), .B(n21537), .C(n21506), .D(
        n21631), .Y(n21508) );
  sky130_fd_sc_hd__nor2_1 U26352 ( .A(n21509), .B(n21508), .Y(n21587) );
  sky130_fd_sc_hd__nor2_1 U26353 ( .A(n21510), .B(n24848), .Y(n21585) );
  sky130_fd_sc_hd__nand4_1 U26354 ( .A(n21587), .B(n21585), .C(n21534), .D(
        n22413), .Y(n21511) );
  sky130_fd_sc_hd__nor4_1 U26355 ( .A(n21590), .B(n21513), .C(n21512), .D(
        n21511), .Y(n21514) );
  sky130_fd_sc_hd__o21ai_1 U26356 ( .A1(n24882), .A2(n21514), .B1(n21644), .Y(
        n10603) );
  sky130_fd_sc_hd__nand3_1 U26357 ( .A(n21516), .B(n24861), .C(n21515), .Y(
        n21517) );
  sky130_fd_sc_hd__or4_1 U26358 ( .A(n21554), .B(n21519), .C(n21518), .D(
        n21517), .X(n21541) );
  sky130_fd_sc_hd__nor3_1 U26359 ( .A(n24863), .B(n21559), .C(n21530), .Y(
        n21520) );
  sky130_fd_sc_hd__nand2_1 U26361 ( .A(n21523), .B(n21522), .Y(n21539) );
  sky130_fd_sc_hd__or3_1 U26362 ( .A(n21540), .B(n21539), .C(n21524), .X(
        n21525) );
  sky130_fd_sc_hd__o21ai_1 U26363 ( .A1(n21525), .A2(n21541), .B1(n24858), .Y(
        n21531) );
  sky130_fd_sc_hd__nor3b_1 U26364 ( .C_N(n22804), .A(n21527), .B(n21526), .Y(
        n21529) );
  sky130_fd_sc_hd__a21oi_1 U26365 ( .A1(n21529), .A2(n21528), .B1(n22401), .Y(
        n21552) );
  sky130_fd_sc_hd__nor2_1 U26366 ( .A(n22418), .B(n21644), .Y(n24877) );
  sky130_fd_sc_hd__nor3_1 U26367 ( .A(n21552), .B(n24877), .C(n21530), .Y(
        n21544) );
  sky130_fd_sc_hd__nand2_1 U26368 ( .A(n21531), .B(n21544), .Y(n10581) );
  sky130_fd_sc_hd__a21oi_1 U26369 ( .A1(n24869), .A2(n21533), .B1(n21532), .Y(
        n21535) );
  sky130_fd_sc_hd__nand3_1 U26370 ( .A(n21535), .B(n22741), .C(n21534), .Y(
        n22281) );
  sky130_fd_sc_hd__nand2_1 U26371 ( .A(n21537), .B(n21536), .Y(n21538) );
  sky130_fd_sc_hd__or4_1 U26372 ( .A(n21540), .B(n22281), .C(n21539), .D(
        n21538), .X(n21542) );
  sky130_fd_sc_hd__nor3_1 U26373 ( .A(n21543), .B(n21542), .C(n21541), .Y(
        n21545) );
  sky130_fd_sc_hd__o21ai_1 U26374 ( .A1(n24882), .A2(n21545), .B1(n21544), .Y(
        n10579) );
  sky130_fd_sc_hd__a21oi_1 U26375 ( .A1(n21548), .A2(n21547), .B1(n21546), .Y(
        n21550) );
  sky130_fd_sc_hd__a21oi_1 U26376 ( .A1(n21550), .A2(n21549), .B1(n24882), .Y(
        n21551) );
  sky130_fd_sc_hd__or3_1 U26377 ( .A(n21552), .B(n21551), .C(n23225), .X(
        n10485) );
  sky130_fd_sc_hd__nor2_1 U26378 ( .A(n21554), .B(n21553), .Y(n21557) );
  sky130_fd_sc_hd__nand3_1 U26379 ( .A(n21557), .B(n21556), .C(n21555), .Y(
        n21558) );
  sky130_fd_sc_hd__nand2_1 U26380 ( .A(n21558), .B(n24858), .Y(n21561) );
  sky130_fd_sc_hd__nand4_1 U26381 ( .A(n21561), .B(n21560), .C(n22339), .D(
        n24844), .Y(n10486) );
  sky130_fd_sc_hd__a21oi_1 U26382 ( .A1(n21564), .A2(n21563), .B1(n21562), .Y(
        n21579) );
  sky130_fd_sc_hd__nor4b_1 U26383 ( .D_N(n22413), .A(n21608), .B(n22732), .C(
        n21565), .Y(n21567) );
  sky130_fd_sc_hd__nand2_1 U26384 ( .A(n21567), .B(n21566), .Y(n22398) );
  sky130_fd_sc_hd__o22ai_1 U26385 ( .A1(n22342), .A2(n22412), .B1(n21569), 
        .B2(n21568), .Y(n21570) );
  sky130_fd_sc_hd__nor4_1 U26386 ( .A(n22746), .B(n22398), .C(n21571), .D(
        n21570), .Y(n21578) );
  sky130_fd_sc_hd__o22ai_1 U26387 ( .A1(n21575), .A2(n21574), .B1(n21573), 
        .B2(n21572), .Y(n21576) );
  sky130_fd_sc_hd__o21ai_1 U26388 ( .A1(n21634), .A2(n21576), .B1(n22735), .Y(
        n21577) );
  sky130_fd_sc_hd__nand4_1 U26389 ( .A(n21580), .B(n21579), .C(n21578), .D(
        n21577), .Y(n21581) );
  sky130_fd_sc_hd__a21oi_1 U26390 ( .A1(n21582), .A2(n21641), .B1(n21581), .Y(
        n21584) );
  sky130_fd_sc_hd__o21ai_1 U26391 ( .A1(n24882), .A2(n21584), .B1(n21583), .Y(
        n10591) );
  sky130_fd_sc_hd__nand2_1 U26393 ( .A(n21633), .B(n21585), .Y(n24859) );
  sky130_fd_sc_hd__a21oi_1 U26394 ( .A1(n21735), .A2(n21586), .B1(n24833), .Y(
        n24839) );
  sky130_fd_sc_hd__nand3_1 U26395 ( .A(n21587), .B(n24839), .C(n24860), .Y(
        n21588) );
  sky130_fd_sc_hd__nor4_1 U26396 ( .A(n21590), .B(n24859), .C(n21589), .D(
        n21588), .Y(n21591) );
  sky130_fd_sc_hd__o21ai_1 U26397 ( .A1(n24882), .A2(n21591), .B1(n21644), .Y(
        n10569) );
  sky130_fd_sc_hd__o21ai_1 U26398 ( .A1(n21592), .A2(n22309), .B1(n22401), .Y(
        n10571) );
  sky130_fd_sc_hd__a31oi_1 U26399 ( .A1(n21595), .A2(n24849), .A3(n21594), 
        .B1(n24882), .Y(j202_soc_core_j22_cpu_id_idec_N857) );
  sky130_fd_sc_hd__nand2_1 U26400 ( .A(n22734), .B(n21635), .Y(n21597) );
  sky130_fd_sc_hd__nor2_1 U26402 ( .A(n21598), .B(n22281), .Y(n22327) );
  sky130_fd_sc_hd__nor2_1 U26403 ( .A(n22333), .B(n22327), .Y(n21602) );
  sky130_fd_sc_hd__o21ai_0 U26404 ( .A1(n22332), .A2(n22330), .B1(n21599), .Y(
        n21601) );
  sky130_fd_sc_hd__nor4_1 U26405 ( .A(n21603), .B(n21602), .C(n21601), .D(
        n21600), .Y(n21606) );
  sky130_fd_sc_hd__nand2_1 U26406 ( .A(n21605), .B(n21604), .Y(n22796) );
  sky130_fd_sc_hd__o21ai_1 U26407 ( .A1(n21607), .A2(n21606), .B1(n22796), .Y(
        n10499) );
  sky130_fd_sc_hd__nand2_1 U26408 ( .A(n21990), .B(n25372), .Y(n21611) );
  sky130_fd_sc_hd__a31oi_1 U26409 ( .A1(n22733), .A2(n21609), .A3(n22734), 
        .B1(n21608), .Y(n21610) );
  sky130_fd_sc_hd__a21oi_1 U26410 ( .A1(n21611), .A2(n21610), .B1(n24882), .Y(
        j202_soc_core_j22_cpu_id_idec_N917) );
  sky130_fd_sc_hd__nand2_1 U26411 ( .A(n21613), .B(n22344), .Y(n21612) );
  sky130_fd_sc_hd__o21ai_0 U26412 ( .A1(n22723), .A2(n22344), .B1(n21612), .Y(
        j202_soc_core_j22_cpu_rf_N3270) );
  sky130_fd_sc_hd__nand2_1 U26413 ( .A(n21613), .B(n22345), .Y(n21615) );
  sky130_fd_sc_hd__a22oi_1 U26414 ( .A1(j202_soc_core_j22_cpu_pc[0]), .A2(
        n22367), .B1(n22725), .B2(n22369), .Y(n21614) );
  sky130_fd_sc_hd__nand2_1 U26415 ( .A(n21615), .B(n21614), .Y(
        j202_soc_core_j22_cpu_rf_N3345) );
  sky130_fd_sc_hd__o22ai_1 U26416 ( .A1(n21627), .A2(n22753), .B1(n22752), 
        .B2(n21626), .Y(n21628) );
  sky130_fd_sc_hd__a21oi_1 U26417 ( .A1(n22725), .A2(n22756), .B1(n21628), .Y(
        n21629) );
  sky130_fd_sc_hd__a31oi_1 U26419 ( .A1(n21633), .A2(n21632), .A3(n21631), 
        .B1(n24827), .Y(n21639) );
  sky130_fd_sc_hd__nand2_1 U26420 ( .A(n21635), .B(n21634), .Y(n21637) );
  sky130_fd_sc_hd__nand3_1 U26421 ( .A(n24849), .B(n21637), .C(n21636), .Y(
        n21638) );
  sky130_fd_sc_hd__a211oi_1 U26422 ( .A1(n21641), .A2(n21640), .B1(n21639), 
        .C1(n21638), .Y(n21642) );
  sky130_fd_sc_hd__o21ai_1 U26423 ( .A1(n24882), .A2(n21642), .B1(n22796), .Y(
        n10583) );
  sky130_fd_sc_hd__o21ai_1 U26424 ( .A1(n24882), .A2(n21645), .B1(n21644), .Y(
        n10602) );
  sky130_fd_sc_hd__nand2_1 U26425 ( .A(n22122), .B(n22344), .Y(n21646) );
  sky130_fd_sc_hd__o21ai_0 U26426 ( .A1(n22662), .A2(n22344), .B1(n21646), .Y(
        j202_soc_core_j22_cpu_rf_N3271) );
  sky130_fd_sc_hd__nand2_1 U26427 ( .A(n22122), .B(n22345), .Y(n21649) );
  sky130_fd_sc_hd__a22oi_1 U26428 ( .A1(n22367), .A2(n21647), .B1(n22757), 
        .B2(n22369), .Y(n21648) );
  sky130_fd_sc_hd__nand2_1 U26429 ( .A(n21649), .B(n21648), .Y(
        j202_soc_core_j22_cpu_rf_N3346) );
  sky130_fd_sc_hd__or3_1 U26430 ( .A(n21653), .B(n22125), .C(n21650), .X(
        n22920) );
  sky130_fd_sc_hd__nand4_1 U26431 ( .A(n21652), .B(n21651), .C(
        j202_soc_core_ahbcs_6__HREADY_), .D(n22920), .Y(n23248) );
  sky130_fd_sc_hd__nor3_1 U26432 ( .A(n21654), .B(n21653), .C(n21680), .Y(
        n21655) );
  sky130_fd_sc_hd__nand4_1 U26433 ( .A(j202_soc_core_ahbcs_6__HREADY_), .B(
        n21655), .C(n22125), .D(n23247), .Y(n22922) );
  sky130_fd_sc_hd__nand2_1 U26435 ( .A(n23239), .B(n21656), .Y(n21674) );
  sky130_fd_sc_hd__nand2_1 U26436 ( .A(n22153), .B(n21671), .Y(n21658) );
  sky130_fd_sc_hd__nor2_1 U26437 ( .A(n21658), .B(n21657), .Y(n21668) );
  sky130_fd_sc_hd__a21oi_1 U26439 ( .A1(n21668), .A2(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]), .B1(n21660), .Y(n21661) );
  sky130_fd_sc_hd__o21ai_1 U26440 ( .A1(n22125), .A2(n21674), .B1(n21661), .Y(
        j202_soc_core_j22_cpu_ml_N152) );
  sky130_fd_sc_hd__o21ai_1 U26441 ( .A1(n21680), .A2(n23248), .B1(n22922), .Y(
        j202_soc_core_j22_cpu_ml_N193) );
  sky130_fd_sc_hd__nand2_1 U26442 ( .A(n21668), .B(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[2]), .Y(n21662) );
  sky130_fd_sc_hd__o211ai_1 U26443 ( .A1(n21680), .A2(n21674), .B1(n21663), 
        .C1(n21662), .Y(j202_soc_core_j22_cpu_ml_N154) );
  sky130_fd_sc_hd__a21oi_1 U26445 ( .A1(n21668), .A2(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .B1(n21666), .Y(n21667) );
  sky130_fd_sc_hd__o21ai_1 U26446 ( .A1(n22923), .A2(n21674), .B1(n21667), .Y(
        j202_soc_core_j22_cpu_ml_N153) );
  sky130_fd_sc_hd__o22ai_1 U26447 ( .A1(n22128), .A2(n21670), .B1(n21669), 
        .B2(n21674), .Y(j202_soc_core_j22_cpu_ml_N155) );
  sky130_fd_sc_hd__a31oi_1 U26448 ( .A1(n21672), .A2(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[4]), .A3(n21671), .B1(n22187), 
        .Y(n21673) );
  sky130_fd_sc_hd__nor3_1 U26450 ( .A(j202_soc_core_j22_cpu_macop_MAC_[2]), 
        .B(n21676), .C(n22145), .Y(n22126) );
  sky130_fd_sc_hd__nand3_1 U26451 ( .A(n21680), .B(n22125), .C(n21679), .Y(
        n22150) );
  sky130_fd_sc_hd__nand2_1 U26452 ( .A(n22270), .B(n21681), .Y(n21682) );
  sky130_fd_sc_hd__a21oi_1 U26453 ( .A1(n21683), .A2(n22132), .B1(n22131), .Y(
        n21684) );
  sky130_fd_sc_hd__o21ai_1 U26454 ( .A1(n23303), .A2(n22135), .B1(n21684), .Y(
        j202_soc_core_j22_cpu_ml_N320) );
  sky130_fd_sc_hd__nand4_1 U26455 ( .A(n21695), .B(n21698), .C(n21697), .D(
        n21696), .Y(n21690) );
  sky130_fd_sc_hd__nand2_1 U26456 ( .A(n21731), .B(n21699), .Y(n21689) );
  sky130_fd_sc_hd__nand3_1 U26457 ( .A(n21700), .B(n21702), .C(n21701), .Y(
        n21686) );
  sky130_fd_sc_hd__nand2_1 U26458 ( .A(n21703), .B(n21704), .Y(n21685) );
  sky130_fd_sc_hd__nor2_1 U26459 ( .A(n21686), .B(n21685), .Y(n21687) );
  sky130_fd_sc_hd__nand3_1 U26460 ( .A(n21708), .B(n21709), .C(n21687), .Y(
        n21688) );
  sky130_fd_sc_hd__nor3_1 U26461 ( .A(n21690), .B(n21689), .C(n21688), .Y(
        n21691) );
  sky130_fd_sc_hd__nand4_1 U26462 ( .A(n21715), .B(n21717), .C(n21694), .D(
        n21691), .Y(n21693) );
  sky130_fd_sc_hd__nor2_1 U26463 ( .A(n21693), .B(n21719), .Y(n21722) );
  sky130_fd_sc_hd__nor4_1 U26464 ( .A(n21698), .B(n21697), .C(n21696), .D(
        n21695), .Y(n21713) );
  sky130_fd_sc_hd__nor2_1 U26465 ( .A(n21699), .B(n21731), .Y(n21712) );
  sky130_fd_sc_hd__nor3_1 U26466 ( .A(n21702), .B(n21701), .C(n21700), .Y(
        n21707) );
  sky130_fd_sc_hd__nand3_1 U26467 ( .A(n21707), .B(n21706), .C(n21705), .Y(
        n21710) );
  sky130_fd_sc_hd__nor3_1 U26468 ( .A(n21710), .B(n21709), .C(n21708), .Y(
        n21711) );
  sky130_fd_sc_hd__nand4_1 U26469 ( .A(n21714), .B(n21713), .C(n21712), .D(
        n21711), .Y(n21716) );
  sky130_fd_sc_hd__nor3_1 U26470 ( .A(n21717), .B(n21716), .C(n21715), .Y(
        n21718) );
  sky130_fd_sc_hd__nand2_1 U26471 ( .A(n21719), .B(n21718), .Y(n21720) );
  sky130_fd_sc_hd__nor2_1 U26472 ( .A(n21724), .B(n21723), .Y(n21725) );
  sky130_fd_sc_hd__nor2_1 U26473 ( .A(n22216), .B(n22198), .Y(n22195) );
  sky130_fd_sc_hd__a22oi_1 U26474 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[17]), .B1(n22219), .B2(n21726), .Y(
        n21727) );
  sky130_fd_sc_hd__nand2_1 U26475 ( .A(n22206), .B(n21727), .Y(
        j202_soc_core_j22_cpu_ml_machj[17]) );
  sky130_fd_sc_hd__a22oi_1 U26476 ( .A1(n22225), .A2(
        j202_soc_core_j22_cpu_ml_bufa[17]), .B1(n22224), .B2(n21730), .Y(
        n21732) );
  sky130_fd_sc_hd__nand2_1 U26477 ( .A(n21732), .B(n22245), .Y(
        j202_soc_core_j22_cpu_ml_maclj[17]) );
  sky130_fd_sc_hd__a222oi_1 U26478 ( .A1(n22280), .A2(n25386), .B1(n25382), 
        .B2(n22282), .C1(n25384), .C2(n22281), .Y(n21733) );
  sky130_fd_sc_hd__o21ai_1 U26479 ( .A1(n21733), .A2(n24882), .B1(n22283), .Y(
        n10494) );
  sky130_fd_sc_hd__a21oi_1 U26480 ( .A1(n21735), .A2(n21734), .B1(n24826), .Y(
        n22329) );
  sky130_fd_sc_hd__a222oi_1 U26481 ( .A1(n22281), .A2(n25382), .B1(n25386), 
        .B2(n22282), .C1(n25380), .C2(n22108), .Y(n21736) );
  sky130_fd_sc_hd__o21ai_1 U26482 ( .A1(n21736), .A2(n24882), .B1(n22283), .Y(
        n10495) );
  sky130_fd_sc_hd__o21ai_0 U26483 ( .A1(n21737), .A2(n22198), .B1(n22206), .Y(
        j202_soc_core_j22_cpu_ml_machj[20]) );
  sky130_fd_sc_hd__nand2_1 U26484 ( .A(n22132), .B(n22577), .Y(n21738) );
  sky130_fd_sc_hd__o211ai_1 U26485 ( .A1(n23312), .A2(n22135), .B1(n21738), 
        .C1(n22084), .Y(j202_soc_core_j22_cpu_ml_N324) );
  sky130_fd_sc_hd__o21ai_0 U26486 ( .A1(n21740), .A2(n22221), .B1(n22245), .Y(
        j202_soc_core_j22_cpu_ml_maclj[20]) );
  sky130_fd_sc_hd__nand2_1 U26487 ( .A(n22132), .B(n22575), .Y(n21741) );
  sky130_fd_sc_hd__o211ai_1 U26488 ( .A1(n23338), .A2(n22135), .B1(n21741), 
        .C1(n22084), .Y(j202_soc_core_j22_cpu_ml_N333) );
  sky130_fd_sc_hd__a21oi_1 U26489 ( .A1(j202_soc_core_j22_cpu_ml_bufa[29]), 
        .A2(n22204), .B1(n22195), .Y(n21743) );
  sky130_fd_sc_hd__a22oi_1 U26491 ( .A1(n22225), .A2(
        j202_soc_core_j22_cpu_ml_bufa[29]), .B1(n22224), .B2(n21745), .Y(
        n21746) );
  sky130_fd_sc_hd__nand2_1 U26492 ( .A(n21746), .B(n22245), .Y(
        j202_soc_core_j22_cpu_ml_maclj[29]) );
  sky130_fd_sc_hd__nand2_1 U26493 ( .A(n22132), .B(n22578), .Y(n21747) );
  sky130_fd_sc_hd__o211ai_1 U26494 ( .A1(n23315), .A2(n22135), .B1(n21747), 
        .C1(n22084), .Y(j202_soc_core_j22_cpu_ml_N325) );
  sky130_fd_sc_hd__a22oi_1 U26495 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[21]), .B1(n22219), .B2(n21748), .Y(
        n21749) );
  sky130_fd_sc_hd__nand2_1 U26496 ( .A(n22206), .B(n21749), .Y(
        j202_soc_core_j22_cpu_ml_machj[21]) );
  sky130_fd_sc_hd__o21ai_0 U26497 ( .A1(n21750), .A2(n22221), .B1(n22245), .Y(
        j202_soc_core_j22_cpu_ml_maclj[21]) );
  sky130_fd_sc_hd__nand2_1 U26498 ( .A(n21752), .B(n22344), .Y(n21751) );
  sky130_fd_sc_hd__o21ai_0 U26499 ( .A1(n22344), .A2(n23309), .B1(n21751), .Y(
        j202_soc_core_j22_cpu_rf_N3291) );
  sky130_fd_sc_hd__nand2_1 U26500 ( .A(n21752), .B(n22345), .Y(n21755) );
  sky130_fd_sc_hd__a22oi_1 U26501 ( .A1(n22369), .A2(n21753), .B1(n21758), 
        .B2(n22367), .Y(n21754) );
  sky130_fd_sc_hd__nand2_1 U26502 ( .A(n21755), .B(n21754), .Y(
        j202_soc_core_j22_cpu_rf_N3366) );
  sky130_fd_sc_hd__o22ai_1 U26503 ( .A1(n22642), .A2(n22753), .B1(n22374), 
        .B2(n23309), .Y(n21757) );
  sky130_fd_sc_hd__a21oi_1 U26504 ( .A1(n22378), .A2(n21758), .B1(n21757), .Y(
        n21759) );
  sky130_fd_sc_hd__o21ai_1 U26505 ( .A1(n22752), .A2(n21760), .B1(n21759), .Y(
        j202_soc_core_j22_cpu_rf_N317) );
  sky130_fd_sc_hd__nand2_1 U26506 ( .A(n21761), .B(n22344), .Y(n21762) );
  sky130_fd_sc_hd__o21ai_0 U26507 ( .A1(n22344), .A2(n23326), .B1(n21762), .Y(
        j202_soc_core_j22_cpu_rf_N3298) );
  sky130_fd_sc_hd__a22oi_1 U26508 ( .A1(n22369), .A2(n21079), .B1(n21767), 
        .B2(n22367), .Y(n21763) );
  sky130_fd_sc_hd__o21ai_0 U26509 ( .A1(n22372), .A2(n21764), .B1(n21763), .Y(
        j202_soc_core_j22_cpu_rf_N3373) );
  sky130_fd_sc_hd__o22ai_1 U26510 ( .A1(n22605), .A2(n22753), .B1(n22374), 
        .B2(n23326), .Y(n21766) );
  sky130_fd_sc_hd__a21oi_1 U26511 ( .A1(n21767), .A2(n22378), .B1(n21766), .Y(
        n21768) );
  sky130_fd_sc_hd__nand2_1 U26513 ( .A(n22132), .B(n22574), .Y(n21770) );
  sky130_fd_sc_hd__o211ai_1 U26514 ( .A1(n23326), .A2(n22135), .B1(n21770), 
        .C1(n22084), .Y(j202_soc_core_j22_cpu_ml_N329) );
  sky130_fd_sc_hd__a22oi_1 U26515 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[25]), .B1(n22219), .B2(n21771), .Y(
        n21772) );
  sky130_fd_sc_hd__nand2_1 U26516 ( .A(n22206), .B(n21772), .Y(
        j202_soc_core_j22_cpu_ml_machj[25]) );
  sky130_fd_sc_hd__o21ai_0 U26517 ( .A1(n21774), .A2(n22221), .B1(n22245), .Y(
        j202_soc_core_j22_cpu_ml_maclj[25]) );
  sky130_fd_sc_hd__a21oi_1 U26518 ( .A1(n21775), .A2(n22132), .B1(n22131), .Y(
        n21776) );
  sky130_fd_sc_hd__o21ai_1 U26519 ( .A1(n23306), .A2(n22135), .B1(n21776), .Y(
        j202_soc_core_j22_cpu_ml_N321) );
  sky130_fd_sc_hd__a22oi_1 U26520 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[18]), .B1(n22219), .B2(n21777), .Y(
        n21778) );
  sky130_fd_sc_hd__nand2_1 U26521 ( .A(n22206), .B(n21778), .Y(
        j202_soc_core_j22_cpu_ml_machj[18]) );
  sky130_fd_sc_hd__nand2_1 U26522 ( .A(n22225), .B(
        j202_soc_core_j22_cpu_ml_bufa[18]), .Y(n21779) );
  sky130_fd_sc_hd__o211ai_1 U26523 ( .A1(n21780), .A2(n22221), .B1(n21779), 
        .C1(n22245), .Y(j202_soc_core_j22_cpu_ml_maclj[18]) );
  sky130_fd_sc_hd__nand2_1 U26524 ( .A(n21782), .B(n22344), .Y(n21781) );
  sky130_fd_sc_hd__o21ai_0 U26525 ( .A1(n22344), .A2(n23306), .B1(n21781), .Y(
        j202_soc_core_j22_cpu_rf_N3290) );
  sky130_fd_sc_hd__nand2_1 U26526 ( .A(n21782), .B(n22345), .Y(n21785) );
  sky130_fd_sc_hd__a22oi_1 U26527 ( .A1(n22369), .A2(n21783), .B1(n21789), 
        .B2(n22367), .Y(n21784) );
  sky130_fd_sc_hd__nand2_1 U26528 ( .A(n21785), .B(n21784), .Y(
        j202_soc_core_j22_cpu_rf_N3365) );
  sky130_fd_sc_hd__o22ai_1 U26529 ( .A1(n21787), .A2(n22753), .B1(n22374), 
        .B2(n23306), .Y(n21788) );
  sky130_fd_sc_hd__a21oi_1 U26530 ( .A1(n22378), .A2(n21789), .B1(n21788), .Y(
        n21790) );
  sky130_fd_sc_hd__o21ai_1 U26531 ( .A1(n22752), .A2(n21791), .B1(n21790), .Y(
        j202_soc_core_j22_cpu_rf_N316) );
  sky130_fd_sc_hd__nand2_1 U26532 ( .A(n21803), .B(n22145), .Y(n21792) );
  sky130_fd_sc_hd__o21ai_1 U26533 ( .A1(n22557), .A2(n22145), .B1(n21792), .Y(
        j202_soc_core_j22_cpu_ml_N313) );
  sky130_fd_sc_hd__o21ai_0 U26534 ( .A1(n21794), .A2(n22213), .B1(n22219), .Y(
        j202_soc_core_j22_cpu_ml_machj[10]) );
  sky130_fd_sc_hd__nor2_1 U26535 ( .A(n21795), .B(n22221), .Y(n22243) );
  sky130_fd_sc_hd__nor2_1 U26536 ( .A(n21796), .B(n22221), .Y(n22241) );
  sky130_fd_sc_hd__a22oi_1 U26537 ( .A1(n22243), .A2(n21797), .B1(
        j202_soc_core_j22_cpu_ml_macl[10]), .B2(n22241), .Y(n21798) );
  sky130_fd_sc_hd__o211ai_1 U26538 ( .A1(n21799), .A2(n22246), .B1(n22245), 
        .C1(n21798), .Y(j202_soc_core_j22_cpu_ml_maclj[10]) );
  sky130_fd_sc_hd__nand2_1 U26539 ( .A(n25385), .B(n24858), .Y(n23222) );
  sky130_fd_sc_hd__o21a_1 U26540 ( .A1(n21800), .A2(n22308), .B1(n22283), .X(
        n22760) );
  sky130_fd_sc_hd__o21ai_1 U26541 ( .A1(n21801), .A2(n23222), .B1(n22760), .Y(
        n10490) );
  sky130_fd_sc_hd__nand2_1 U26542 ( .A(n21803), .B(n22366), .Y(n21802) );
  sky130_fd_sc_hd__o21ai_0 U26543 ( .A1(n22366), .A2(n21805), .B1(n21802), .Y(
        j202_soc_core_j22_cpu_rf_N3281) );
  sky130_fd_sc_hd__a22oi_1 U26544 ( .A1(n21806), .A2(n22367), .B1(n21803), 
        .B2(n22369), .Y(n21804) );
  sky130_fd_sc_hd__o21ai_0 U26545 ( .A1(n22372), .A2(n21805), .B1(n21804), .Y(
        j202_soc_core_j22_cpu_rf_N3356) );
  sky130_fd_sc_hd__o22ai_1 U26546 ( .A1(n21807), .A2(n22753), .B1(n22374), 
        .B2(n22168), .Y(n21808) );
  sky130_fd_sc_hd__a21oi_1 U26547 ( .A1(n21809), .A2(n22360), .B1(n21808), .Y(
        n21810) );
  sky130_fd_sc_hd__nand2_1 U26549 ( .A(n22322), .B(n22145), .Y(n21812) );
  sky130_fd_sc_hd__o21ai_0 U26551 ( .A1(n21814), .A2(n22213), .B1(n22219), .Y(
        j202_soc_core_j22_cpu_ml_machj[9]) );
  sky130_fd_sc_hd__a22oi_1 U26552 ( .A1(n22243), .A2(n21815), .B1(
        j202_soc_core_j22_cpu_ml_macl[9]), .B2(n22241), .Y(n21816) );
  sky130_fd_sc_hd__o211ai_1 U26553 ( .A1(n21817), .A2(n22246), .B1(n22245), 
        .C1(n21816), .Y(j202_soc_core_j22_cpu_ml_maclj[9]) );
  sky130_fd_sc_hd__nand2_1 U26554 ( .A(n21819), .B(n22344), .Y(n21818) );
  sky130_fd_sc_hd__o21ai_0 U26555 ( .A1(n22344), .A2(n23321), .B1(n21818), .Y(
        j202_soc_core_j22_cpu_rf_N3296) );
  sky130_fd_sc_hd__nand2_1 U26556 ( .A(n21819), .B(n22345), .Y(n21822) );
  sky130_fd_sc_hd__a22oi_1 U26557 ( .A1(n22369), .A2(n21820), .B1(n21825), 
        .B2(n22367), .Y(n21821) );
  sky130_fd_sc_hd__nand2_1 U26558 ( .A(n21822), .B(n21821), .Y(
        j202_soc_core_j22_cpu_rf_N3370) );
  sky130_fd_sc_hd__o22ai_1 U26559 ( .A1(n22613), .A2(n22753), .B1(n22374), 
        .B2(n23321), .Y(n21824) );
  sky130_fd_sc_hd__a21oi_1 U26560 ( .A1(n21825), .A2(n22378), .B1(n21824), .Y(
        n21826) );
  sky130_fd_sc_hd__a21oi_1 U26562 ( .A1(n21828), .A2(n22132), .B1(n22131), .Y(
        n21829) );
  sky130_fd_sc_hd__a22oi_1 U26564 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[23]), .B1(n22219), .B2(n21830), .Y(
        n21831) );
  sky130_fd_sc_hd__nand2_1 U26565 ( .A(n22206), .B(n21831), .Y(
        j202_soc_core_j22_cpu_ml_machj[23]) );
  sky130_fd_sc_hd__nand2_1 U26566 ( .A(n22225), .B(
        j202_soc_core_j22_cpu_ml_bufa[23]), .Y(n21832) );
  sky130_fd_sc_hd__o211ai_1 U26567 ( .A1(n21833), .A2(n22221), .B1(n21832), 
        .C1(n22245), .Y(j202_soc_core_j22_cpu_ml_maclj[23]) );
  sky130_fd_sc_hd__nand2_1 U26568 ( .A(n21834), .B(n22344), .Y(n21835) );
  sky130_fd_sc_hd__o21ai_0 U26569 ( .A1(n22344), .A2(n21937), .B1(n21835), .Y(
        j202_soc_core_j22_cpu_rf_N3297) );
  sky130_fd_sc_hd__a22oi_1 U26570 ( .A1(n22369), .A2(n21836), .B1(n21842), 
        .B2(n22367), .Y(n21837) );
  sky130_fd_sc_hd__o22ai_1 U26572 ( .A1(n21840), .A2(n22753), .B1(n22374), 
        .B2(n21937), .Y(n21841) );
  sky130_fd_sc_hd__a21oi_1 U26573 ( .A1(n21842), .A2(n22378), .B1(n21841), .Y(
        n21843) );
  sky130_fd_sc_hd__o22ai_1 U26575 ( .A1(n22611), .A2(n22753), .B1(n22374), 
        .B2(n22520), .Y(n21845) );
  sky130_fd_sc_hd__a21oi_1 U26576 ( .A1(n21846), .A2(n22360), .B1(n21845), .Y(
        n21847) );
  sky130_fd_sc_hd__nand2_1 U26578 ( .A(n21850), .B(n22344), .Y(n21849) );
  sky130_fd_sc_hd__o21ai_0 U26579 ( .A1(n22520), .A2(n22344), .B1(n21849), .Y(
        j202_soc_core_j22_cpu_rf_N3276) );
  sky130_fd_sc_hd__nand2_1 U26580 ( .A(n21850), .B(n22345), .Y(n21853) );
  sky130_fd_sc_hd__a22oi_1 U26581 ( .A1(n21851), .A2(n22367), .B1(n22045), 
        .B2(n22369), .Y(n21852) );
  sky130_fd_sc_hd__nand2_1 U26582 ( .A(n21853), .B(n21852), .Y(
        j202_soc_core_j22_cpu_rf_N3351) );
  sky130_fd_sc_hd__nand2_1 U26583 ( .A(n25390), .B(n21854), .Y(n21855) );
  sky130_fd_sc_hd__nand2_1 U26585 ( .A(n22729), .B(n22898), .Y(
        j202_soc_core_j22_cpu_rf_N3391) );
  sky130_fd_sc_hd__nand2_1 U26586 ( .A(n21858), .B(n22344), .Y(n21857) );
  sky130_fd_sc_hd__o21ai_0 U26587 ( .A1(n22158), .A2(n22344), .B1(n21857), .Y(
        j202_soc_core_j22_cpu_rf_N3286) );
  sky130_fd_sc_hd__nand2_1 U26588 ( .A(n21858), .B(n22345), .Y(n21860) );
  sky130_fd_sc_hd__a22oi_1 U26589 ( .A1(n22369), .A2(n22514), .B1(n21864), 
        .B2(n22367), .Y(n21859) );
  sky130_fd_sc_hd__nand2_1 U26590 ( .A(n21860), .B(n21859), .Y(
        j202_soc_core_j22_cpu_rf_N3360) );
  sky130_fd_sc_hd__o22ai_1 U26591 ( .A1(n21862), .A2(n22753), .B1(n22374), 
        .B2(n22158), .Y(n21863) );
  sky130_fd_sc_hd__a21oi_1 U26592 ( .A1(n22378), .A2(n21864), .B1(n21863), .Y(
        n21865) );
  sky130_fd_sc_hd__o21ai_1 U26593 ( .A1(n22752), .A2(n21866), .B1(n21865), .Y(
        j202_soc_core_j22_cpu_rf_N312) );
  sky130_fd_sc_hd__nand2_1 U26594 ( .A(n22132), .B(n21867), .Y(n21868) );
  sky130_fd_sc_hd__o211ai_1 U26595 ( .A1(n23318), .A2(n22135), .B1(n21868), 
        .C1(n22084), .Y(j202_soc_core_j22_cpu_ml_N326) );
  sky130_fd_sc_hd__a22oi_1 U26596 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[22]), .B1(n22219), .B2(n21869), .Y(
        n21870) );
  sky130_fd_sc_hd__nand2_1 U26597 ( .A(n22206), .B(n21870), .Y(
        j202_soc_core_j22_cpu_ml_machj[22]) );
  sky130_fd_sc_hd__nand2_1 U26598 ( .A(n22225), .B(
        j202_soc_core_j22_cpu_ml_bufa[22]), .Y(n21871) );
  sky130_fd_sc_hd__o211ai_1 U26599 ( .A1(n21872), .A2(n22221), .B1(n21871), 
        .C1(n22245), .Y(j202_soc_core_j22_cpu_ml_maclj[22]) );
  sky130_fd_sc_hd__nand2_1 U26600 ( .A(n21874), .B(n22344), .Y(n21873) );
  sky130_fd_sc_hd__o21ai_0 U26601 ( .A1(n23318), .A2(n22344), .B1(n21873), .Y(
        j202_soc_core_j22_cpu_rf_N3295) );
  sky130_fd_sc_hd__nand2_1 U26602 ( .A(n21874), .B(n22345), .Y(n21876) );
  sky130_fd_sc_hd__a22oi_1 U26603 ( .A1(n22369), .A2(n22513), .B1(n21880), 
        .B2(n22367), .Y(n21875) );
  sky130_fd_sc_hd__nand2_1 U26604 ( .A(n21876), .B(n21875), .Y(
        j202_soc_core_j22_cpu_rf_N3369) );
  sky130_fd_sc_hd__o22ai_1 U26605 ( .A1(n21878), .A2(n22753), .B1(n22374), 
        .B2(n23318), .Y(n21879) );
  sky130_fd_sc_hd__a21oi_1 U26606 ( .A1(n21880), .A2(n22378), .B1(n21879), .Y(
        n21881) );
  sky130_fd_sc_hd__o21ai_1 U26607 ( .A1(n22752), .A2(n21882), .B1(n21881), .Y(
        j202_soc_core_j22_cpu_rf_N320) );
  sky130_fd_sc_hd__nand2_1 U26608 ( .A(n22132), .B(n22579), .Y(n21883) );
  sky130_fd_sc_hd__o211ai_1 U26609 ( .A1(n23342), .A2(n22135), .B1(n21883), 
        .C1(n22084), .Y(j202_soc_core_j22_cpu_ml_N334) );
  sky130_fd_sc_hd__a21oi_1 U26610 ( .A1(j202_soc_core_j22_cpu_ml_bufa[30]), 
        .A2(n22204), .B1(n22195), .Y(n21885) );
  sky130_fd_sc_hd__o21ai_1 U26611 ( .A1(n22198), .A2(n21886), .B1(n21885), .Y(
        j202_soc_core_j22_cpu_ml_machj[30]) );
  sky130_fd_sc_hd__a22oi_1 U26612 ( .A1(n22225), .A2(
        j202_soc_core_j22_cpu_ml_bufa[30]), .B1(n22224), .B2(n21887), .Y(
        n21888) );
  sky130_fd_sc_hd__nand2_1 U26613 ( .A(n21888), .B(n22245), .Y(
        j202_soc_core_j22_cpu_ml_maclj[30]) );
  sky130_fd_sc_hd__nand2_1 U26614 ( .A(n21890), .B(n22366), .Y(n21889) );
  sky130_fd_sc_hd__o21ai_1 U26615 ( .A1(n22366), .A2(n11199), .B1(n21889), .Y(
        j202_soc_core_j22_cpu_rf_N3304) );
  sky130_fd_sc_hd__a22oi_1 U26616 ( .A1(n22369), .A2(n21890), .B1(n21894), 
        .B2(n22367), .Y(n21891) );
  sky130_fd_sc_hd__o21ai_1 U26617 ( .A1(n22372), .A2(n11199), .B1(n21891), .Y(
        j202_soc_core_j22_cpu_rf_N3378) );
  sky130_fd_sc_hd__o22ai_1 U26618 ( .A1(n22603), .A2(n22753), .B1(n22374), 
        .B2(n23342), .Y(n21893) );
  sky130_fd_sc_hd__a21oi_1 U26619 ( .A1(n21894), .A2(n22378), .B1(n21893), .Y(
        n21895) );
  sky130_fd_sc_hd__nand2_1 U26621 ( .A(n22514), .B(n22145), .Y(n21897) );
  sky130_fd_sc_hd__a22oi_1 U26623 ( .A1(n22243), .A2(n21898), .B1(
        j202_soc_core_j22_cpu_ml_macl[14]), .B2(n22241), .Y(n21899) );
  sky130_fd_sc_hd__o211ai_1 U26624 ( .A1(n21900), .A2(n22246), .B1(n22245), 
        .C1(n21899), .Y(j202_soc_core_j22_cpu_ml_maclj[14]) );
  sky130_fd_sc_hd__a22oi_1 U26625 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[14]), .B1(n22216), .B2(n21901), .Y(
        n21902) );
  sky130_fd_sc_hd__nand2_1 U26626 ( .A(n22219), .B(n21902), .Y(
        j202_soc_core_j22_cpu_ml_machj[14]) );
  sky130_fd_sc_hd__nor2_1 U26627 ( .A(j202_soc_core_ahb2aqu_00_aqu_st_0_), .B(
        j202_soc_core_rst), .Y(n21905) );
  sky130_fd_sc_hd__nand2_1 U26628 ( .A(n21904), .B(n21903), .Y(
        j202_soc_core_ahb2aqu_00_N93) );
  sky130_fd_sc_hd__nand2b_1 U26629 ( .A_N(n22099), .B(n21905), .Y(
        j202_soc_core_ahb2aqu_00_N95) );
  sky130_fd_sc_hd__nand2_1 U26630 ( .A(n22099), .B(n21906), .Y(n22830) );
  sky130_fd_sc_hd__o31a_1 U26631 ( .A1(n21908), .A2(n21907), .A3(n22403), .B1(
        n22830), .X(n22103) );
  sky130_fd_sc_hd__o21ai_0 U26633 ( .A1(n25379), .A2(n22403), .B1(n21909), .Y(
        n21910) );
  sky130_fd_sc_hd__nand2_1 U26634 ( .A(n21910), .B(n22816), .Y(n21912) );
  sky130_fd_sc_hd__nand2_1 U26635 ( .A(n10979), .B(n22827), .Y(n21911) );
  sky130_fd_sc_hd__nor4_1 U26636 ( .A(n25375), .B(n25374), .C(n25373), .D(
        n21913), .Y(n21914) );
  sky130_fd_sc_hd__nand2_1 U26637 ( .A(n25376), .B(n21914), .Y(n22025) );
  sky130_fd_sc_hd__nand3_1 U26638 ( .A(j202_soc_core_aquc_WE_), .B(
        j202_soc_core_aquc_SEL__3_), .C(j202_soc_core_aquc_CE__1_), .Y(n22815)
         );
  sky130_fd_sc_hd__nand2_1 U26639 ( .A(n22815), .B(j202_soc_core_uart_div0[6]), 
        .Y(n21916) );
  sky130_fd_sc_hd__o21ai_1 U26640 ( .A1(n22815), .A2(n24053), .B1(n21916), .Y(
        n43) );
  sky130_fd_sc_hd__nand2_1 U26641 ( .A(n21925), .B(n22145), .Y(n21917) );
  sky130_fd_sc_hd__o21ai_1 U26642 ( .A1(n22558), .A2(n22145), .B1(n21917), .Y(
        j202_soc_core_j22_cpu_ml_N311) );
  sky130_fd_sc_hd__o21ai_0 U26643 ( .A1(n21919), .A2(n22213), .B1(n22219), .Y(
        j202_soc_core_j22_cpu_ml_machj[8]) );
  sky130_fd_sc_hd__a22oi_1 U26644 ( .A1(n22243), .A2(n21920), .B1(
        j202_soc_core_j22_cpu_ml_macl[8]), .B2(n22241), .Y(n21921) );
  sky130_fd_sc_hd__o211ai_1 U26645 ( .A1(n21922), .A2(n22246), .B1(n22245), 
        .C1(n21921), .Y(j202_soc_core_j22_cpu_ml_maclj[8]) );
  sky130_fd_sc_hd__nand2_1 U26646 ( .A(n21924), .B(n22344), .Y(n21923) );
  sky130_fd_sc_hd__o21ai_0 U26647 ( .A1(n22344), .A2(n22173), .B1(n21923), .Y(
        j202_soc_core_j22_cpu_rf_N3279) );
  sky130_fd_sc_hd__nand2_1 U26648 ( .A(n21924), .B(n22345), .Y(n21928) );
  sky130_fd_sc_hd__a22oi_1 U26649 ( .A1(n21926), .A2(n22367), .B1(n21925), 
        .B2(n22369), .Y(n21927) );
  sky130_fd_sc_hd__nand2_1 U26650 ( .A(n21928), .B(n21927), .Y(
        j202_soc_core_j22_cpu_rf_N3354) );
  sky130_fd_sc_hd__o22ai_1 U26651 ( .A1(n21929), .A2(n22753), .B1(n22374), 
        .B2(n22173), .Y(n21930) );
  sky130_fd_sc_hd__a21oi_1 U26652 ( .A1(n21931), .A2(n22360), .B1(n21930), .Y(
        n21932) );
  sky130_fd_sc_hd__o21ai_1 U26653 ( .A1(n21933), .A2(n22759), .B1(n21932), .Y(
        j202_soc_core_j22_cpu_rf_N306) );
  sky130_fd_sc_hd__nand2_1 U26654 ( .A(n22729), .B(n21934), .Y(
        j202_soc_core_j22_cpu_rf_N2637) );
  sky130_fd_sc_hd__nand2_1 U26655 ( .A(n22132), .B(n21935), .Y(n21936) );
  sky130_fd_sc_hd__o211ai_1 U26656 ( .A1(n21937), .A2(n22135), .B1(n21936), 
        .C1(n22084), .Y(j202_soc_core_j22_cpu_ml_N328) );
  sky130_fd_sc_hd__a22oi_1 U26657 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[24]), .B1(n22219), .B2(n21938), .Y(
        n21939) );
  sky130_fd_sc_hd__nand2_1 U26658 ( .A(n22206), .B(n21939), .Y(
        j202_soc_core_j22_cpu_ml_machj[24]) );
  sky130_fd_sc_hd__o21ai_0 U26659 ( .A1(n21941), .A2(n22221), .B1(n22245), .Y(
        j202_soc_core_j22_cpu_ml_maclj[24]) );
  sky130_fd_sc_hd__a21oi_1 U26660 ( .A1(n22576), .A2(n22132), .B1(n22131), .Y(
        n21942) );
  sky130_fd_sc_hd__o21ai_1 U26661 ( .A1(n23332), .A2(n22135), .B1(n21942), .Y(
        j202_soc_core_j22_cpu_ml_N331) );
  sky130_fd_sc_hd__a22oi_1 U26662 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[27]), .B1(n22219), .B2(n21943), .Y(
        n21944) );
  sky130_fd_sc_hd__nand2_1 U26663 ( .A(n22206), .B(n21944), .Y(
        j202_soc_core_j22_cpu_ml_machj[27]) );
  sky130_fd_sc_hd__o21ai_0 U26664 ( .A1(n21946), .A2(n22221), .B1(n22245), .Y(
        j202_soc_core_j22_cpu_ml_maclj[27]) );
  sky130_fd_sc_hd__nand2_1 U26665 ( .A(n21947), .B(n22344), .Y(n21948) );
  sky130_fd_sc_hd__o21ai_0 U26666 ( .A1(n22344), .A2(n23332), .B1(n21948), .Y(
        j202_soc_core_j22_cpu_rf_N3300) );
  sky130_fd_sc_hd__a22oi_1 U26667 ( .A1(n22369), .A2(n21949), .B1(n21954), 
        .B2(n22367), .Y(n21950) );
  sky130_fd_sc_hd__o22ai_1 U26669 ( .A1(n22609), .A2(n22753), .B1(n22374), 
        .B2(n23332), .Y(n21953) );
  sky130_fd_sc_hd__a21oi_1 U26670 ( .A1(n21954), .A2(n22378), .B1(n21953), .Y(
        n21955) );
  sky130_fd_sc_hd__nand2_1 U26672 ( .A(n22515), .B(n22145), .Y(n21957) );
  sky130_fd_sc_hd__o21ai_1 U26673 ( .A1(n22564), .A2(n22145), .B1(n21957), .Y(
        j202_soc_core_j22_cpu_ml_N314) );
  sky130_fd_sc_hd__a22oi_1 U26674 ( .A1(n22243), .A2(n21958), .B1(
        j202_soc_core_j22_cpu_ml_macl[11]), .B2(n22241), .Y(n21959) );
  sky130_fd_sc_hd__o211ai_1 U26675 ( .A1(n21960), .A2(n22246), .B1(n22245), 
        .C1(n21959), .Y(j202_soc_core_j22_cpu_ml_maclj[11]) );
  sky130_fd_sc_hd__a22oi_1 U26676 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[11]), .B1(n22216), .B2(n21961), .Y(
        n21962) );
  sky130_fd_sc_hd__nand2_1 U26677 ( .A(n22219), .B(n21962), .Y(
        j202_soc_core_j22_cpu_ml_machj[11]) );
  sky130_fd_sc_hd__a21oi_1 U26678 ( .A1(n21963), .A2(n22132), .B1(n22131), .Y(
        n21964) );
  sky130_fd_sc_hd__a22oi_1 U26680 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[19]), .B1(n22219), .B2(n21965), .Y(
        n21966) );
  sky130_fd_sc_hd__nand2_1 U26681 ( .A(n22206), .B(n21966), .Y(
        j202_soc_core_j22_cpu_ml_machj[19]) );
  sky130_fd_sc_hd__nand2_1 U26682 ( .A(n22225), .B(
        j202_soc_core_j22_cpu_ml_bufa[19]), .Y(n21967) );
  sky130_fd_sc_hd__o211ai_1 U26683 ( .A1(n21968), .A2(n22221), .B1(n21967), 
        .C1(n22245), .Y(j202_soc_core_j22_cpu_ml_maclj[19]) );
  sky130_fd_sc_hd__nand2_1 U26684 ( .A(n21970), .B(n22344), .Y(n21969) );
  sky130_fd_sc_hd__o21ai_0 U26685 ( .A1(n22344), .A2(n23315), .B1(n21969), .Y(
        j202_soc_core_j22_cpu_rf_N3294) );
  sky130_fd_sc_hd__nand2_1 U26686 ( .A(n21970), .B(n22345), .Y(n21973) );
  sky130_fd_sc_hd__a22oi_1 U26687 ( .A1(n22369), .A2(n21971), .B1(n21976), 
        .B2(n22367), .Y(n21972) );
  sky130_fd_sc_hd__nand2_1 U26688 ( .A(n21973), .B(n21972), .Y(
        j202_soc_core_j22_cpu_rf_N3368) );
  sky130_fd_sc_hd__o22ai_1 U26689 ( .A1(n22599), .A2(n22753), .B1(n22374), 
        .B2(n23315), .Y(n21975) );
  sky130_fd_sc_hd__a21oi_1 U26690 ( .A1(n21976), .A2(n22378), .B1(n21975), .Y(
        n21977) );
  sky130_fd_sc_hd__o21ai_1 U26691 ( .A1(n22752), .A2(n21978), .B1(n21977), .Y(
        j202_soc_core_j22_cpu_rf_N319) );
  sky130_fd_sc_hd__nand2_1 U26692 ( .A(n21980), .B(n22344), .Y(n21979) );
  sky130_fd_sc_hd__o21ai_0 U26693 ( .A1(n22344), .A2(n23338), .B1(n21979), .Y(
        j202_soc_core_j22_cpu_rf_N3303) );
  sky130_fd_sc_hd__nand2_1 U26694 ( .A(n21980), .B(n22345), .Y(n21983) );
  sky130_fd_sc_hd__a22oi_1 U26695 ( .A1(n22369), .A2(n21981), .B1(n21987), 
        .B2(n22367), .Y(n21982) );
  sky130_fd_sc_hd__nand2_1 U26696 ( .A(n21983), .B(n21982), .Y(
        j202_soc_core_j22_cpu_rf_N3377) );
  sky130_fd_sc_hd__nand2_1 U26697 ( .A(n21984), .B(n22360), .Y(n21989) );
  sky130_fd_sc_hd__o22ai_1 U26698 ( .A1(n21985), .A2(n22753), .B1(n22374), 
        .B2(n23338), .Y(n21986) );
  sky130_fd_sc_hd__a21oi_1 U26699 ( .A1(n21987), .A2(n22378), .B1(n21986), .Y(
        n21988) );
  sky130_fd_sc_hd__nand2_1 U26700 ( .A(n21989), .B(n21988), .Y(
        j202_soc_core_j22_cpu_rf_N327) );
  sky130_fd_sc_hd__a222oi_1 U26701 ( .A1(n25380), .A2(n21990), .B1(n25381), 
        .B2(n22107), .C1(n22108), .C2(n25377), .Y(n21991) );
  sky130_fd_sc_hd__o21ai_1 U26702 ( .A1(n21991), .A2(n24882), .B1(n22283), .Y(
        n10497) );
  sky130_fd_sc_hd__o21ai_0 U26703 ( .A1(n21992), .A2(n22213), .B1(n22219), .Y(
        j202_soc_core_j22_cpu_ml_machj[4]) );
  sky130_fd_sc_hd__nand2_1 U26704 ( .A(n22484), .B(n22145), .Y(n21993) );
  sky130_fd_sc_hd__o21ai_1 U26705 ( .A1(n22647), .A2(n22145), .B1(n21993), .Y(
        j202_soc_core_j22_cpu_ml_N307) );
  sky130_fd_sc_hd__o21ai_0 U26706 ( .A1(n21995), .A2(n22221), .B1(n22245), .Y(
        j202_soc_core_j22_cpu_ml_maclj[4]) );
  sky130_fd_sc_hd__nand2_1 U26707 ( .A(n22057), .B(n21996), .Y(n21998) );
  sky130_fd_sc_hd__nand2_1 U26708 ( .A(n21998), .B(n21997), .Y(
        j202_soc_core_j22_cpu_rf_N2646) );
  sky130_fd_sc_hd__nand2_1 U26709 ( .A(n22013), .B(n22145), .Y(n21999) );
  sky130_fd_sc_hd__o21ai_1 U26710 ( .A1(n22488), .A2(n22145), .B1(n21999), .Y(
        j202_soc_core_j22_cpu_ml_N306) );
  sky130_fd_sc_hd__a22oi_1 U26711 ( .A1(n22243), .A2(n22000), .B1(
        j202_soc_core_j22_cpu_ml_macl[3]), .B2(n22241), .Y(n22001) );
  sky130_fd_sc_hd__o211ai_1 U26712 ( .A1(n22002), .A2(n22246), .B1(n22245), 
        .C1(n22001), .Y(j202_soc_core_j22_cpu_ml_maclj[3]) );
  sky130_fd_sc_hd__a22oi_1 U26713 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[3]), .B1(n22216), .B2(n22003), .Y(n22004) );
  sky130_fd_sc_hd__nand2_1 U26714 ( .A(n22219), .B(n22004), .Y(
        j202_soc_core_j22_cpu_ml_machj[3]) );
  sky130_fd_sc_hd__nand2_1 U26715 ( .A(n22006), .B(n22344), .Y(n22005) );
  sky130_fd_sc_hd__o21ai_1 U26716 ( .A1(n22519), .A2(n22344), .B1(n22005), .Y(
        j202_soc_core_j22_cpu_rf_N3273) );
  sky130_fd_sc_hd__nand2_1 U26717 ( .A(n22006), .B(n22345), .Y(n22008) );
  sky130_fd_sc_hd__a22oi_1 U26718 ( .A1(n22009), .A2(n22367), .B1(n22013), 
        .B2(n22369), .Y(n22007) );
  sky130_fd_sc_hd__nand2_1 U26719 ( .A(n22008), .B(n22007), .Y(
        j202_soc_core_j22_cpu_rf_N3348) );
  sky130_fd_sc_hd__o22ai_1 U26720 ( .A1(n22711), .A2(n22753), .B1(n22752), 
        .B2(n22011), .Y(n22012) );
  sky130_fd_sc_hd__a21oi_1 U26721 ( .A1(n22756), .A2(n22013), .B1(n22012), .Y(
        n22014) );
  sky130_fd_sc_hd__nand2_1 U26723 ( .A(n22017), .B(n22344), .Y(n22016) );
  sky130_fd_sc_hd__nand2_1 U26725 ( .A(n22017), .B(n22345), .Y(n22019) );
  sky130_fd_sc_hd__a22oi_1 U26726 ( .A1(n22369), .A2(n20409), .B1(n22022), 
        .B2(n22367), .Y(n22018) );
  sky130_fd_sc_hd__nand2_1 U26727 ( .A(n22019), .B(n22018), .Y(
        j202_soc_core_j22_cpu_rf_N3367) );
  sky130_fd_sc_hd__o22ai_1 U26728 ( .A1(n22640), .A2(n22753), .B1(n22374), 
        .B2(n23312), .Y(n22021) );
  sky130_fd_sc_hd__a21oi_1 U26729 ( .A1(n22022), .A2(n22378), .B1(n22021), .Y(
        n22023) );
  sky130_fd_sc_hd__o21ai_1 U26730 ( .A1(n22752), .A2(n22024), .B1(n22023), .Y(
        j202_soc_core_j22_cpu_rf_N318) );
  sky130_fd_sc_hd__nand2_1 U26731 ( .A(n22555), .B(n22145), .Y(n22026) );
  sky130_fd_sc_hd__o21ai_1 U26732 ( .A1(n22580), .A2(n22145), .B1(n22026), .Y(
        j202_soc_core_j22_cpu_ml_N308) );
  sky130_fd_sc_hd__o21ai_0 U26733 ( .A1(n22028), .A2(n22213), .B1(n22219), .Y(
        j202_soc_core_j22_cpu_ml_machj[5]) );
  sky130_fd_sc_hd__a22oi_1 U26734 ( .A1(n22243), .A2(n22029), .B1(
        j202_soc_core_j22_cpu_ml_macl[5]), .B2(n22241), .Y(n22030) );
  sky130_fd_sc_hd__o211ai_1 U26735 ( .A1(n22031), .A2(n22246), .B1(n22245), 
        .C1(n22030), .Y(j202_soc_core_j22_cpu_ml_maclj[5]) );
  sky130_fd_sc_hd__nand2_1 U26736 ( .A(n22033), .B(n22344), .Y(n22032) );
  sky130_fd_sc_hd__o21ai_0 U26737 ( .A1(n22492), .A2(n22344), .B1(n22032), .Y(
        j202_soc_core_j22_cpu_rf_N3275) );
  sky130_fd_sc_hd__nand2_1 U26738 ( .A(n22033), .B(n22345), .Y(n22036) );
  sky130_fd_sc_hd__a22oi_1 U26739 ( .A1(n22034), .A2(n22367), .B1(n22555), 
        .B2(n22369), .Y(n22035) );
  sky130_fd_sc_hd__nand2_1 U26740 ( .A(n22036), .B(n22035), .Y(
        j202_soc_core_j22_cpu_rf_N3350) );
  sky130_fd_sc_hd__o22ai_1 U26741 ( .A1(n22037), .A2(n22753), .B1(n22374), 
        .B2(n22492), .Y(n22038) );
  sky130_fd_sc_hd__a21oi_1 U26742 ( .A1(n22039), .A2(n22360), .B1(n22038), .Y(
        n22040) );
  sky130_fd_sc_hd__o21ai_1 U26743 ( .A1(n22041), .A2(n22759), .B1(n22040), .Y(
        j202_soc_core_j22_cpu_rf_N303) );
  sky130_fd_sc_hd__nand2_1 U26744 ( .A(n25390), .B(n22042), .Y(n22043) );
  sky130_fd_sc_hd__o21ai_1 U26745 ( .A1(n22044), .A2(n22785), .B1(n22043), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N4) );
  sky130_fd_sc_hd__nand2_1 U26746 ( .A(n22045), .B(n22145), .Y(n22046) );
  sky130_fd_sc_hd__o21ai_1 U26747 ( .A1(n22612), .A2(n22145), .B1(n22046), .Y(
        j202_soc_core_j22_cpu_ml_N309) );
  sky130_fd_sc_hd__a22oi_1 U26748 ( .A1(n22243), .A2(n22047), .B1(
        j202_soc_core_j22_cpu_ml_macl[6]), .B2(n22241), .Y(n22048) );
  sky130_fd_sc_hd__o211ai_1 U26749 ( .A1(n22049), .A2(n22246), .B1(n22245), 
        .C1(n22048), .Y(j202_soc_core_j22_cpu_ml_maclj[6]) );
  sky130_fd_sc_hd__a22oi_1 U26750 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[6]), .B1(n22216), .B2(n22050), .Y(n22051) );
  sky130_fd_sc_hd__nand2_1 U26751 ( .A(n22219), .B(n22051), .Y(
        j202_soc_core_j22_cpu_ml_machj[6]) );
  sky130_fd_sc_hd__o22ai_1 U26752 ( .A1(n22646), .A2(n22753), .B1(n22374), 
        .B2(n22536), .Y(n22052) );
  sky130_fd_sc_hd__a21oi_1 U26753 ( .A1(n22053), .A2(n22360), .B1(n22052), .Y(
        n22054) );
  sky130_fd_sc_hd__nand2_1 U26755 ( .A(n22057), .B(n22344), .Y(n22056) );
  sky130_fd_sc_hd__o21ai_0 U26756 ( .A1(n22536), .A2(n22344), .B1(n22056), .Y(
        j202_soc_core_j22_cpu_rf_N3274) );
  sky130_fd_sc_hd__nand2_1 U26757 ( .A(n22057), .B(n22345), .Y(n22060) );
  sky130_fd_sc_hd__a22oi_1 U26758 ( .A1(n22058), .A2(n22367), .B1(n22484), 
        .B2(n22369), .Y(n22059) );
  sky130_fd_sc_hd__nand2_1 U26759 ( .A(n22060), .B(n22059), .Y(
        j202_soc_core_j22_cpu_rf_N3349) );
  sky130_fd_sc_hd__nand2_1 U26760 ( .A(n25390), .B(n22061), .Y(n22062) );
  sky130_fd_sc_hd__o21ai_1 U26761 ( .A1(n22063), .A2(n22785), .B1(n22062), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N3) );
  sky130_fd_sc_hd__o22ai_1 U26762 ( .A1(n22064), .A2(n22753), .B1(n22374), 
        .B2(n22163), .Y(n22065) );
  sky130_fd_sc_hd__a21oi_1 U26763 ( .A1(n22066), .A2(n22360), .B1(n22065), .Y(
        n22067) );
  sky130_fd_sc_hd__nand2_1 U26765 ( .A(n22093), .B(n22366), .Y(n22069) );
  sky130_fd_sc_hd__o21ai_0 U26766 ( .A1(n22366), .A2(n22072), .B1(n22069), .Y(
        j202_soc_core_j22_cpu_rf_N3283) );
  sky130_fd_sc_hd__a22oi_1 U26767 ( .A1(n22070), .A2(n22367), .B1(n22093), 
        .B2(n22369), .Y(n22071) );
  sky130_fd_sc_hd__o21ai_0 U26768 ( .A1(n22372), .A2(n22072), .B1(n22071), .Y(
        j202_soc_core_j22_cpu_rf_N3358) );
  sky130_fd_sc_hd__nand2_1 U26769 ( .A(n22073), .B(n22360), .Y(n22077) );
  sky130_fd_sc_hd__o22ai_1 U26770 ( .A1(n22074), .A2(n22753), .B1(n22374), 
        .B2(n23335), .Y(n22075) );
  sky130_fd_sc_hd__a21oi_1 U26771 ( .A1(n22080), .A2(n22378), .B1(n22075), .Y(
        n22076) );
  sky130_fd_sc_hd__nand2_1 U26772 ( .A(n22077), .B(n22076), .Y(
        j202_soc_core_j22_cpu_rf_N326) );
  sky130_fd_sc_hd__nand2_1 U26773 ( .A(n22079), .B(n22344), .Y(n22078) );
  sky130_fd_sc_hd__o21ai_0 U26774 ( .A1(n22344), .A2(n23335), .B1(n22078), .Y(
        j202_soc_core_j22_cpu_rf_N3302) );
  sky130_fd_sc_hd__nand2_1 U26775 ( .A(n22079), .B(n22345), .Y(n22083) );
  sky130_fd_sc_hd__a22oi_1 U26776 ( .A1(n22369), .A2(n22081), .B1(n22080), 
        .B2(n22367), .Y(n22082) );
  sky130_fd_sc_hd__nand2_1 U26777 ( .A(n22083), .B(n22082), .Y(
        j202_soc_core_j22_cpu_rf_N3376) );
  sky130_fd_sc_hd__nand2_1 U26778 ( .A(n22132), .B(n22631), .Y(n22085) );
  sky130_fd_sc_hd__o211ai_1 U26779 ( .A1(n23335), .A2(n22135), .B1(n22085), 
        .C1(n22084), .Y(j202_soc_core_j22_cpu_ml_N332) );
  sky130_fd_sc_hd__a21oi_1 U26780 ( .A1(j202_soc_core_j22_cpu_ml_bufa[28]), 
        .A2(n22204), .B1(n22195), .Y(n22087) );
  sky130_fd_sc_hd__o21ai_1 U26781 ( .A1(n22088), .A2(n22198), .B1(n22087), .Y(
        j202_soc_core_j22_cpu_ml_machj[28]) );
  sky130_fd_sc_hd__a22oi_1 U26782 ( .A1(n22225), .A2(
        j202_soc_core_j22_cpu_ml_bufa[28]), .B1(n22224), .B2(n22089), .Y(
        n22090) );
  sky130_fd_sc_hd__nand2_1 U26783 ( .A(n22090), .B(n22245), .Y(
        j202_soc_core_j22_cpu_ml_maclj[28]) );
  sky130_fd_sc_hd__clkinv_1 U26784 ( .A(j202_soc_core_qspi_wb_wdat[28]), .Y(
        n22092) );
  sky130_fd_sc_hd__nand2_1 U26785 ( .A(n22815), .B(j202_soc_core_uart_div0[4]), 
        .Y(n22091) );
  sky130_fd_sc_hd__o21ai_1 U26786 ( .A1(n22815), .A2(n22092), .B1(n22091), .Y(
        n42) );
  sky130_fd_sc_hd__nand2_1 U26787 ( .A(n22093), .B(n22145), .Y(n22094) );
  sky130_fd_sc_hd__o21ai_1 U26788 ( .A1(n22560), .A2(n22145), .B1(n22094), .Y(
        j202_soc_core_j22_cpu_ml_N315) );
  sky130_fd_sc_hd__o21ai_0 U26789 ( .A1(n22095), .A2(n22213), .B1(n22219), .Y(
        j202_soc_core_j22_cpu_ml_machj[12]) );
  sky130_fd_sc_hd__a22oi_1 U26790 ( .A1(n22243), .A2(n22096), .B1(
        j202_soc_core_j22_cpu_ml_macl[12]), .B2(n22241), .Y(n22097) );
  sky130_fd_sc_hd__o211ai_1 U26791 ( .A1(n22098), .A2(n22246), .B1(n22245), 
        .C1(n22097), .Y(j202_soc_core_j22_cpu_ml_maclj[12]) );
  sky130_fd_sc_hd__o22a_1 U26792 ( .A1(n25379), .A2(n22100), .B1(n22829), .B2(
        n22099), .X(n22826) );
  sky130_fd_sc_hd__nand2_1 U26793 ( .A(n22826), .B(n22816), .Y(n22102) );
  sky130_fd_sc_hd__nand2_1 U26794 ( .A(n10976), .B(n22827), .Y(n22101) );
  sky130_fd_sc_hd__nand3_1 U26795 ( .A(n22103), .B(n22102), .C(n22101), .Y(
        j202_soc_core_ahb2aqu_00_N163) );
  sky130_fd_sc_hd__nand2_1 U26796 ( .A(n22813), .B(j202_soc_core_uart_div1[3]), 
        .Y(n22105) );
  sky130_fd_sc_hd__nand2_1 U26798 ( .A(n25193), .B(
        j202_soc_core_bldc_core_00_wdata[19]), .Y(n22106) );
  sky130_fd_sc_hd__o21ai_1 U26799 ( .A1(n25126), .A2(n25193), .B1(n22106), .Y(
        n27) );
  sky130_fd_sc_hd__a222oi_1 U26800 ( .A1(n25381), .A2(n22108), .B1(n25380), 
        .B2(n22107), .C1(n25386), .C2(n22281), .Y(n22109) );
  sky130_fd_sc_hd__o21ai_1 U26801 ( .A1(n22109), .A2(n24882), .B1(n22283), .Y(
        n10496) );
  sky130_fd_sc_hd__nand2_1 U26802 ( .A(n22111), .B(n22344), .Y(n22110) );
  sky130_fd_sc_hd__o21ai_0 U26803 ( .A1(n22344), .A2(n23303), .B1(n22110), .Y(
        j202_soc_core_j22_cpu_rf_N3289) );
  sky130_fd_sc_hd__nand2_1 U26804 ( .A(n22111), .B(n22345), .Y(n22114) );
  sky130_fd_sc_hd__a22oi_1 U26805 ( .A1(n22369), .A2(n22112), .B1(n22118), 
        .B2(n22367), .Y(n22113) );
  sky130_fd_sc_hd__nand2_1 U26806 ( .A(n22114), .B(n22113), .Y(
        j202_soc_core_j22_cpu_rf_N3364) );
  sky130_fd_sc_hd__o22ai_1 U26807 ( .A1(n22116), .A2(n22753), .B1(n22374), 
        .B2(n23303), .Y(n22117) );
  sky130_fd_sc_hd__a21oi_1 U26808 ( .A1(n22378), .A2(n22118), .B1(n22117), .Y(
        n22119) );
  sky130_fd_sc_hd__nand2_1 U26810 ( .A(n22813), .B(j202_soc_core_uart_div1[1]), 
        .Y(n22121) );
  sky130_fd_sc_hd__nand2_1 U26812 ( .A(n22122), .B(n22124), .Y(n22123) );
  sky130_fd_sc_hd__o21ai_0 U26813 ( .A1(n22662), .A2(n22124), .B1(n22123), .Y(
        j202_soc_core_j22_cpu_rf_N2628) );
  sky130_fd_sc_hd__o21ai_1 U26814 ( .A1(n22125), .A2(n23248), .B1(n22922), .Y(
        j202_soc_core_j22_cpu_ml_N191) );
  sky130_fd_sc_hd__a21oi_1 U26815 ( .A1(n22126), .A2(n22591), .B1(n22131), .Y(
        n22127) );
  sky130_fd_sc_hd__o31ai_1 U26816 ( .A1(n22128), .A2(n23348), .A3(n22135), 
        .B1(n22127), .Y(j202_soc_core_j22_cpu_ml_N336) );
  sky130_fd_sc_hd__a21oi_1 U26817 ( .A1(n22591), .A2(n22132), .B1(n22131), .Y(
        n22129) );
  sky130_fd_sc_hd__o21ai_1 U26818 ( .A1(n23348), .A2(n22135), .B1(n22129), .Y(
        j202_soc_core_j22_cpu_ml_N335) );
  sky130_fd_sc_hd__a21oi_1 U26819 ( .A1(n22573), .A2(n22132), .B1(n22131), .Y(
        n22130) );
  sky130_fd_sc_hd__o21ai_1 U26820 ( .A1(n23329), .A2(n22135), .B1(n22130), .Y(
        j202_soc_core_j22_cpu_ml_N330) );
  sky130_fd_sc_hd__a21oi_1 U26821 ( .A1(n22133), .A2(n22132), .B1(n22131), .Y(
        n22134) );
  sky130_fd_sc_hd__o21ai_1 U26822 ( .A1(n23300), .A2(n22135), .B1(n22134), .Y(
        j202_soc_core_j22_cpu_ml_N319) );
  sky130_fd_sc_hd__nand2_1 U26823 ( .A(n22136), .B(n22143), .Y(n22137) );
  sky130_fd_sc_hd__o21ai_1 U26824 ( .A1(n22143), .A2(n22274), .B1(n22137), .Y(
        j202_soc_core_j22_cpu_ml_N318) );
  sky130_fd_sc_hd__nand2_1 U26825 ( .A(n22554), .B(n22145), .Y(n22138) );
  sky130_fd_sc_hd__o21ai_1 U26826 ( .A1(n22561), .A2(n22145), .B1(n22138), .Y(
        j202_soc_core_j22_cpu_ml_N316) );
  sky130_fd_sc_hd__nand2_1 U26827 ( .A(n22495), .B(n22145), .Y(n22139) );
  sky130_fd_sc_hd__o21ai_1 U26828 ( .A1(n22645), .A2(n22145), .B1(n22139), .Y(
        j202_soc_core_j22_cpu_ml_N310) );
  sky130_fd_sc_hd__nand2_1 U26829 ( .A(n22547), .B(n22145), .Y(n22140) );
  sky130_fd_sc_hd__o21ai_1 U26830 ( .A1(n22487), .A2(n22145), .B1(n22140), .Y(
        j202_soc_core_j22_cpu_ml_N305) );
  sky130_fd_sc_hd__nand2_1 U26831 ( .A(n22141), .B(n22143), .Y(n22142) );
  sky130_fd_sc_hd__o21ai_1 U26832 ( .A1(n22143), .A2(n22662), .B1(n22142), .Y(
        j202_soc_core_j22_cpu_ml_N304) );
  sky130_fd_sc_hd__nand2_1 U26833 ( .A(n22725), .B(n22145), .Y(n22144) );
  sky130_fd_sc_hd__o21ai_1 U26834 ( .A1(n22146), .A2(n22145), .B1(n22144), .Y(
        j202_soc_core_j22_cpu_ml_N303) );
  sky130_fd_sc_hd__o21ai_0 U26835 ( .A1(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[1]), .A2(
        j202_soc_core_j22_cpu_ml_M_macop_MAC_[0]), .B1(n22147), .Y(n22148) );
  sky130_fd_sc_hd__nor3_1 U26836 ( .A(n22150), .B(n22275), .C(n22149), .Y(
        n22151) );
  sky130_fd_sc_hd__a31oi_1 U26837 ( .A1(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[1]), .A2(
        j202_soc_core_j22_cpu_ml_bufb[31]), .A3(n22187), .B1(n22151), .Y(
        n22152) );
  sky130_fd_sc_hd__nand2b_1 U26839 ( .A_N(n23345), .B(n22153), .Y(n22189) );
  sky130_fd_sc_hd__a22oi_1 U26840 ( .A1(j202_soc_core_j22_cpu_ml_bufb[31]), 
        .A2(n22187), .B1(n22186), .B2(n22154), .Y(n22155) );
  sky130_fd_sc_hd__o21ai_1 U26841 ( .A1(n22189), .A2(n22274), .B1(n22155), .Y(
        j202_soc_core_j22_cpu_ml_N427) );
  sky130_fd_sc_hd__a22oi_1 U26842 ( .A1(j202_soc_core_j22_cpu_ml_bufb[30]), 
        .A2(n22187), .B1(n22186), .B2(n22156), .Y(n22157) );
  sky130_fd_sc_hd__o21ai_1 U26843 ( .A1(n22189), .A2(n22158), .B1(n22157), .Y(
        j202_soc_core_j22_cpu_ml_N426) );
  sky130_fd_sc_hd__a22oi_1 U26844 ( .A1(j202_soc_core_j22_cpu_ml_bufb[29]), 
        .A2(n22187), .B1(n22186), .B2(n22159), .Y(n22160) );
  sky130_fd_sc_hd__a22oi_1 U26846 ( .A1(j202_soc_core_j22_cpu_ml_bufb[28]), 
        .A2(n22187), .B1(n22186), .B2(n22161), .Y(n22162) );
  sky130_fd_sc_hd__o21ai_1 U26847 ( .A1(n22189), .A2(n22163), .B1(n22162), .Y(
        j202_soc_core_j22_cpu_ml_N424) );
  sky130_fd_sc_hd__a22oi_1 U26848 ( .A1(j202_soc_core_j22_cpu_ml_bufb[27]), 
        .A2(n22187), .B1(n22186), .B2(n22164), .Y(n22165) );
  sky130_fd_sc_hd__o21ai_1 U26849 ( .A1(n22189), .A2(n22350), .B1(n22165), .Y(
        j202_soc_core_j22_cpu_ml_N423) );
  sky130_fd_sc_hd__a22oi_1 U26850 ( .A1(j202_soc_core_j22_cpu_ml_bufb[26]), 
        .A2(n22187), .B1(n22186), .B2(n22166), .Y(n22167) );
  sky130_fd_sc_hd__o21ai_1 U26851 ( .A1(n22189), .A2(n22168), .B1(n22167), .Y(
        j202_soc_core_j22_cpu_ml_N422) );
  sky130_fd_sc_hd__a22oi_1 U26852 ( .A1(j202_soc_core_j22_cpu_ml_bufb[25]), 
        .A2(n22187), .B1(n22186), .B2(n22169), .Y(n22170) );
  sky130_fd_sc_hd__a22oi_1 U26854 ( .A1(j202_soc_core_j22_cpu_ml_bufb[24]), 
        .A2(n22187), .B1(n22186), .B2(n22171), .Y(n22172) );
  sky130_fd_sc_hd__o21ai_1 U26855 ( .A1(n22189), .A2(n22173), .B1(n22172), .Y(
        j202_soc_core_j22_cpu_ml_N420) );
  sky130_fd_sc_hd__a22oi_1 U26856 ( .A1(j202_soc_core_j22_cpu_ml_bufb[23]), 
        .A2(n22187), .B1(n22186), .B2(n22704), .Y(n22174) );
  sky130_fd_sc_hd__o21ai_1 U26857 ( .A1(n22189), .A2(n22290), .B1(n22174), .Y(
        j202_soc_core_j22_cpu_ml_N419) );
  sky130_fd_sc_hd__a22oi_1 U26858 ( .A1(j202_soc_core_j22_cpu_ml_bufb[22]), 
        .A2(n22187), .B1(n22186), .B2(n22708), .Y(n22175) );
  sky130_fd_sc_hd__o21ai_1 U26859 ( .A1(n22189), .A2(n22520), .B1(n22175), .Y(
        j202_soc_core_j22_cpu_ml_N418) );
  sky130_fd_sc_hd__a22oi_1 U26860 ( .A1(j202_soc_core_j22_cpu_ml_bufb[21]), 
        .A2(n22187), .B1(n22186), .B2(n22176), .Y(n22177) );
  sky130_fd_sc_hd__o21ai_1 U26861 ( .A1(n22189), .A2(n22492), .B1(n22177), .Y(
        j202_soc_core_j22_cpu_ml_N417) );
  sky130_fd_sc_hd__a22oi_1 U26862 ( .A1(j202_soc_core_j22_cpu_ml_bufb[20]), 
        .A2(n22187), .B1(n22186), .B2(n22705), .Y(n22178) );
  sky130_fd_sc_hd__o21ai_1 U26863 ( .A1(n22189), .A2(n22536), .B1(n22178), .Y(
        j202_soc_core_j22_cpu_ml_N416) );
  sky130_fd_sc_hd__a22oi_1 U26864 ( .A1(j202_soc_core_j22_cpu_ml_bufb[19]), 
        .A2(n22187), .B1(n22186), .B2(n22179), .Y(n22180) );
  sky130_fd_sc_hd__o21ai_1 U26865 ( .A1(n22189), .A2(n22519), .B1(n22180), .Y(
        j202_soc_core_j22_cpu_ml_N415) );
  sky130_fd_sc_hd__a22oi_1 U26866 ( .A1(j202_soc_core_j22_cpu_ml_bufb[18]), 
        .A2(n22187), .B1(n22186), .B2(n22181), .Y(n22182) );
  sky130_fd_sc_hd__a22oi_1 U26868 ( .A1(j202_soc_core_j22_cpu_ml_bufb[17]), 
        .A2(n22187), .B1(n22186), .B2(n22183), .Y(n22184) );
  sky130_fd_sc_hd__o21ai_1 U26869 ( .A1(n22189), .A2(n22662), .B1(n22184), .Y(
        j202_soc_core_j22_cpu_ml_N413) );
  sky130_fd_sc_hd__a22oi_1 U26870 ( .A1(j202_soc_core_j22_cpu_ml_bufb[16]), 
        .A2(n22187), .B1(n22186), .B2(n22185), .Y(n22188) );
  sky130_fd_sc_hd__o21ai_1 U26871 ( .A1(n22189), .A2(n22723), .B1(n22188), .Y(
        j202_soc_core_j22_cpu_ml_N412) );
  sky130_fd_sc_hd__o22ai_1 U26872 ( .A1(n22246), .A2(n22191), .B1(n22190), 
        .B2(n22218), .Y(n22192) );
  sky130_fd_sc_hd__a211o_1 U26873 ( .A1(n22224), .A2(n22193), .B1(n22198), 
        .C1(n22192), .X(j202_soc_core_j22_cpu_ml_maclj[31]) );
  sky130_fd_sc_hd__a21oi_1 U26874 ( .A1(j202_soc_core_j22_cpu_ml_bufa[31]), 
        .A2(n22204), .B1(n22195), .Y(n22196) );
  sky130_fd_sc_hd__o21ai_1 U26875 ( .A1(n22198), .A2(n22197), .B1(n22196), .Y(
        j202_soc_core_j22_cpu_ml_machj[31]) );
  sky130_fd_sc_hd__a22oi_1 U26876 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[26]), .B1(n22219), .B2(n22199), .Y(
        n22200) );
  sky130_fd_sc_hd__nand2_1 U26877 ( .A(n22206), .B(n22200), .Y(
        j202_soc_core_j22_cpu_ml_machj[26]) );
  sky130_fd_sc_hd__a22oi_1 U26878 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[16]), .B1(n22219), .B2(n22201), .Y(
        n22202) );
  sky130_fd_sc_hd__nand2_1 U26879 ( .A(n22206), .B(n22202), .Y(
        j202_soc_core_j22_cpu_ml_machj[16]) );
  sky130_fd_sc_hd__a22oi_1 U26880 ( .A1(n22204), .A2(
        j202_soc_core_j22_cpu_ml_bufa[15]), .B1(n22219), .B2(n22203), .Y(
        n22205) );
  sky130_fd_sc_hd__nand2_1 U26881 ( .A(n22206), .B(n22205), .Y(
        j202_soc_core_j22_cpu_ml_machj[15]) );
  sky130_fd_sc_hd__o21ai_0 U26882 ( .A1(n22207), .A2(n22213), .B1(n22219), .Y(
        j202_soc_core_j22_cpu_ml_machj[13]) );
  sky130_fd_sc_hd__o21ai_0 U26883 ( .A1(n22209), .A2(n22213), .B1(n22219), .Y(
        j202_soc_core_j22_cpu_ml_machj[7]) );
  sky130_fd_sc_hd__o21ai_0 U26884 ( .A1(n22211), .A2(n22213), .B1(n22219), .Y(
        j202_soc_core_j22_cpu_ml_machj[2]) );
  sky130_fd_sc_hd__o21ai_0 U26885 ( .A1(n22214), .A2(n22213), .B1(n22219), .Y(
        j202_soc_core_j22_cpu_ml_machj[1]) );
  sky130_fd_sc_hd__nand2_1 U26886 ( .A(n22216), .B(n22215), .Y(n22217) );
  sky130_fd_sc_hd__nand3_1 U26887 ( .A(n22219), .B(n22218), .C(n22217), .Y(
        j202_soc_core_j22_cpu_ml_machj[0]) );
  sky130_fd_sc_hd__o21ai_0 U26888 ( .A1(n22222), .A2(n22221), .B1(n22245), .Y(
        j202_soc_core_j22_cpu_ml_maclj[26]) );
  sky130_fd_sc_hd__a22oi_1 U26889 ( .A1(n22225), .A2(
        j202_soc_core_j22_cpu_ml_bufa[16]), .B1(n22224), .B2(n22223), .Y(
        n22226) );
  sky130_fd_sc_hd__nand2_1 U26890 ( .A(n22226), .B(n22245), .Y(
        j202_soc_core_j22_cpu_ml_maclj[16]) );
  sky130_fd_sc_hd__a22oi_1 U26891 ( .A1(n22243), .A2(n22227), .B1(
        j202_soc_core_j22_cpu_ml_macl[15]), .B2(n22241), .Y(n22228) );
  sky130_fd_sc_hd__o211ai_1 U26892 ( .A1(n22229), .A2(n22246), .B1(n22245), 
        .C1(n22228), .Y(j202_soc_core_j22_cpu_ml_maclj[15]) );
  sky130_fd_sc_hd__a22oi_1 U26893 ( .A1(n22243), .A2(n22230), .B1(
        j202_soc_core_j22_cpu_ml_macl[13]), .B2(n22241), .Y(n22231) );
  sky130_fd_sc_hd__o211ai_1 U26894 ( .A1(n22232), .A2(n22246), .B1(n22245), 
        .C1(n22231), .Y(j202_soc_core_j22_cpu_ml_maclj[13]) );
  sky130_fd_sc_hd__a22oi_1 U26895 ( .A1(n22243), .A2(n22233), .B1(
        j202_soc_core_j22_cpu_ml_macl[7]), .B2(n22241), .Y(n22234) );
  sky130_fd_sc_hd__o211ai_1 U26896 ( .A1(n22235), .A2(n22246), .B1(n22245), 
        .C1(n22234), .Y(j202_soc_core_j22_cpu_ml_maclj[7]) );
  sky130_fd_sc_hd__a22oi_1 U26897 ( .A1(n22243), .A2(n22236), .B1(
        j202_soc_core_j22_cpu_ml_macl[2]), .B2(n22241), .Y(n22237) );
  sky130_fd_sc_hd__o211ai_1 U26898 ( .A1(n22238), .A2(n22246), .B1(n22245), 
        .C1(n22237), .Y(j202_soc_core_j22_cpu_ml_maclj[2]) );
  sky130_fd_sc_hd__a22oi_1 U26899 ( .A1(n22243), .A2(n22239), .B1(
        j202_soc_core_j22_cpu_ml_macl[1]), .B2(n22241), .Y(n22240) );
  sky130_fd_sc_hd__o211ai_1 U26900 ( .A1(n15666), .A2(n22246), .B1(n22245), 
        .C1(n22240), .Y(j202_soc_core_j22_cpu_ml_maclj[1]) );
  sky130_fd_sc_hd__a22oi_1 U26901 ( .A1(n22243), .A2(n22242), .B1(
        j202_soc_core_j22_cpu_ml_macl[0]), .B2(n22241), .Y(n22244) );
  sky130_fd_sc_hd__o211ai_1 U26902 ( .A1(n22247), .A2(n22246), .B1(n22245), 
        .C1(n22244), .Y(j202_soc_core_j22_cpu_ml_maclj[0]) );
  sky130_fd_sc_hd__nand2_1 U26903 ( .A(n22248), .B(n22344), .Y(n22249) );
  sky130_fd_sc_hd__o21ai_0 U26904 ( .A1(n22344), .A2(n23329), .B1(n22249), .Y(
        j202_soc_core_j22_cpu_rf_N3299) );
  sky130_fd_sc_hd__a22oi_1 U26905 ( .A1(n22512), .A2(n22369), .B1(n22254), 
        .B2(n22367), .Y(n22250) );
  sky130_fd_sc_hd__o21ai_1 U26906 ( .A1(n22372), .A2(n22251), .B1(n22250), .Y(
        j202_soc_core_j22_cpu_rf_N3374) );
  sky130_fd_sc_hd__o22ai_1 U26907 ( .A1(n22602), .A2(n22753), .B1(n22374), 
        .B2(n23329), .Y(n22253) );
  sky130_fd_sc_hd__a21oi_1 U26908 ( .A1(n22254), .A2(n22378), .B1(n22253), .Y(
        n22255) );
  sky130_fd_sc_hd__nand2_1 U26910 ( .A(n22258), .B(n22344), .Y(n22257) );
  sky130_fd_sc_hd__nand2_1 U26912 ( .A(n22258), .B(n22345), .Y(n22261) );
  sky130_fd_sc_hd__a22oi_1 U26913 ( .A1(n22259), .A2(n22367), .B1(n22547), 
        .B2(n22369), .Y(n22260) );
  sky130_fd_sc_hd__nand2_1 U26914 ( .A(n22261), .B(n22260), .Y(
        j202_soc_core_j22_cpu_rf_N3347) );
  sky130_fd_sc_hd__o22ai_1 U26915 ( .A1(n22264), .A2(n22753), .B1(n22752), 
        .B2(n22263), .Y(n22265) );
  sky130_fd_sc_hd__a21oi_1 U26916 ( .A1(n22756), .A2(n22547), .B1(n22265), .Y(
        n22266) );
  sky130_fd_sc_hd__o21ai_1 U26917 ( .A1(n22267), .A2(n22759), .B1(n22266), .Y(
        j202_soc_core_j22_cpu_rf_N300) );
  sky130_fd_sc_hd__nand2_1 U26918 ( .A(n22269), .B(n22344), .Y(n22268) );
  sky130_fd_sc_hd__o21ai_0 U26919 ( .A1(n22344), .A2(n22274), .B1(n22268), .Y(
        j202_soc_core_j22_cpu_rf_N3287) );
  sky130_fd_sc_hd__nand2_1 U26920 ( .A(n22269), .B(n22345), .Y(n22272) );
  sky130_fd_sc_hd__a22oi_1 U26921 ( .A1(n22369), .A2(n22270), .B1(n22277), 
        .B2(n22367), .Y(n22271) );
  sky130_fd_sc_hd__nand2_1 U26922 ( .A(n22272), .B(n22271), .Y(
        j202_soc_core_j22_cpu_rf_N3361) );
  sky130_fd_sc_hd__o22ai_1 U26923 ( .A1(n22275), .A2(n22753), .B1(n22374), 
        .B2(n22274), .Y(n22276) );
  sky130_fd_sc_hd__a21oi_1 U26924 ( .A1(n22378), .A2(n22277), .B1(n22276), .Y(
        n22278) );
  sky130_fd_sc_hd__o21ai_1 U26925 ( .A1(n22752), .A2(n22279), .B1(n22278), .Y(
        j202_soc_core_j22_cpu_rf_N313) );
  sky130_fd_sc_hd__a222oi_1 U26926 ( .A1(n25384), .A2(n22282), .B1(n22281), 
        .B2(n25383), .C1(n25382), .C2(n22280), .Y(n22284) );
  sky130_fd_sc_hd__o21ai_1 U26927 ( .A1(n22284), .A2(n24882), .B1(n22283), .Y(
        n10493) );
  sky130_fd_sc_hd__nand2_1 U26928 ( .A(n22286), .B(n22344), .Y(n22285) );
  sky130_fd_sc_hd__o21ai_0 U26929 ( .A1(n22290), .A2(n22344), .B1(n22285), .Y(
        j202_soc_core_j22_cpu_rf_N3278) );
  sky130_fd_sc_hd__nand2_1 U26930 ( .A(n22286), .B(n22345), .Y(n22288) );
  sky130_fd_sc_hd__a22oi_1 U26931 ( .A1(n22289), .A2(n22367), .B1(n22495), 
        .B2(n22369), .Y(n22287) );
  sky130_fd_sc_hd__nand2_1 U26932 ( .A(n22288), .B(n22287), .Y(
        j202_soc_core_j22_cpu_rf_N3352) );
  sky130_fd_sc_hd__o22ai_1 U26933 ( .A1(n22644), .A2(n22753), .B1(n22374), 
        .B2(n22290), .Y(n22291) );
  sky130_fd_sc_hd__a21oi_1 U26934 ( .A1(n22292), .A2(n22360), .B1(n22291), .Y(
        n22293) );
  sky130_fd_sc_hd__o21ai_1 U26935 ( .A1(n22294), .A2(n22759), .B1(n22293), .Y(
        j202_soc_core_j22_cpu_rf_N305) );
  sky130_fd_sc_hd__nand2_1 U26936 ( .A(n22554), .B(n22366), .Y(n22295) );
  sky130_fd_sc_hd__o21ai_0 U26937 ( .A1(n22366), .A2(n22297), .B1(n22295), .Y(
        j202_soc_core_j22_cpu_rf_N3284) );
  sky130_fd_sc_hd__a22oi_1 U26938 ( .A1(n22554), .A2(n22369), .B1(n22298), 
        .B2(n22367), .Y(n22296) );
  sky130_fd_sc_hd__o21ai_1 U26939 ( .A1(n22372), .A2(n22297), .B1(n22296), .Y(
        j202_soc_core_j22_cpu_rf_N3359) );
  sky130_fd_sc_hd__o22ai_1 U26940 ( .A1(n22300), .A2(n22753), .B1(n22374), 
        .B2(n22299), .Y(n22301) );
  sky130_fd_sc_hd__a21oi_1 U26941 ( .A1(n22302), .A2(n22360), .B1(n22301), .Y(
        n22303) );
  sky130_fd_sc_hd__o21ai_1 U26942 ( .A1(n22759), .A2(n22304), .B1(n22303), .Y(
        j202_soc_core_j22_cpu_rf_N311) );
  sky130_fd_sc_hd__nand2_1 U26943 ( .A(n22813), .B(j202_soc_core_uart_div1[7]), 
        .Y(n22305) );
  sky130_fd_sc_hd__o21ai_1 U26944 ( .A1(n24011), .A2(n22813), .B1(n22305), .Y(
        n111) );
  sky130_fd_sc_hd__nand2_1 U26945 ( .A(n22306), .B(n24858), .Y(n22761) );
  sky130_fd_sc_hd__o22a_1 U26946 ( .A1(n22309), .A2(n22761), .B1(n22308), .B2(
        n22307), .X(n22310) );
  sky130_fd_sc_hd__nand2_1 U26947 ( .A(n22760), .B(n22310), .Y(n10491) );
  sky130_fd_sc_hd__nand2_1 U26948 ( .A(n22322), .B(n22366), .Y(n22311) );
  sky130_fd_sc_hd__o21ai_0 U26949 ( .A1(n22366), .A2(n22319), .B1(n22311), .Y(
        j202_soc_core_j22_cpu_rf_N3280) );
  sky130_fd_sc_hd__a22oi_1 U26950 ( .A1(n22313), .A2(n22367), .B1(n22322), 
        .B2(n22369), .Y(n22312) );
  sky130_fd_sc_hd__o21ai_0 U26951 ( .A1(n22372), .A2(n22319), .B1(n22312), .Y(
        j202_soc_core_j22_cpu_rf_N3355) );
  sky130_fd_sc_hd__o22ai_1 U26952 ( .A1(n22314), .A2(n22753), .B1(n22374), 
        .B2(n20705), .Y(n22315) );
  sky130_fd_sc_hd__a21oi_1 U26953 ( .A1(n22316), .A2(n22360), .B1(n22315), .Y(
        n22317) );
  sky130_fd_sc_hd__o22ai_1 U26955 ( .A1(n22722), .A2(n20705), .B1(n22721), 
        .B2(n22319), .Y(n22320) );
  sky130_fd_sc_hd__nand2_1 U26956 ( .A(n22501), .B(n22715), .Y(n22325) );
  sky130_fd_sc_hd__nand2_1 U26957 ( .A(n22320), .B(n22325), .Y(n22324) );
  sky130_fd_sc_hd__nor3_1 U26958 ( .A(n22607), .B(n22596), .C(n24894), .Y(
        n22321) );
  sky130_fd_sc_hd__a21oi_1 U26959 ( .A1(n22322), .A2(n24894), .B1(n22321), .Y(
        n22323) );
  sky130_fd_sc_hd__nand2_1 U26960 ( .A(n22324), .B(n22323), .Y(
        j202_soc_core_j22_cpu_rf_N2640) );
  sky130_fd_sc_hd__nand2_1 U26962 ( .A(n22813), .B(j202_soc_core_uart_div1[2]), 
        .Y(n22326) );
  sky130_fd_sc_hd__o22ai_1 U26964 ( .A1(n22330), .A2(n22329), .B1(n22328), 
        .B2(n22327), .Y(n22335) );
  sky130_fd_sc_hd__o21ai_1 U26965 ( .A1(n22333), .A2(n22332), .B1(n22331), .Y(
        n22334) );
  sky130_fd_sc_hd__nor2_1 U26967 ( .A(n22336), .B(n22416), .Y(n24857) );
  sky130_fd_sc_hd__nand4_1 U26968 ( .A(n22340), .B(n22339), .C(n22338), .D(
        n22337), .Y(n10498) );
  sky130_fd_sc_hd__nand2_1 U26969 ( .A(n22815), .B(j202_soc_core_uart_div0[2]), 
        .Y(n22341) );
  sky130_fd_sc_hd__o21ai_1 U26970 ( .A1(n22815), .A2(n24026), .B1(n22341), .Y(
        n73) );
  sky130_fd_sc_hd__o21ai_1 U26971 ( .A1(n22342), .A2(n22761), .B1(n22760), .Y(
        n10489) );
  sky130_fd_sc_hd__nand2_1 U26972 ( .A(n22346), .B(n22344), .Y(n22343) );
  sky130_fd_sc_hd__o21ai_0 U26973 ( .A1(n22350), .A2(n22344), .B1(n22343), .Y(
        j202_soc_core_j22_cpu_rf_N3282) );
  sky130_fd_sc_hd__nand2_1 U26974 ( .A(n22346), .B(n22345), .Y(n22348) );
  sky130_fd_sc_hd__a22oi_1 U26975 ( .A1(n22349), .A2(n22367), .B1(n22515), 
        .B2(n22369), .Y(n22347) );
  sky130_fd_sc_hd__nand2_1 U26976 ( .A(n22348), .B(n22347), .Y(
        j202_soc_core_j22_cpu_rf_N3357) );
  sky130_fd_sc_hd__o22ai_1 U26977 ( .A1(n22351), .A2(n22753), .B1(n22374), 
        .B2(n22350), .Y(n22352) );
  sky130_fd_sc_hd__a21oi_1 U26978 ( .A1(n22353), .A2(n22360), .B1(n22352), .Y(
        n22354) );
  sky130_fd_sc_hd__o21ai_1 U26979 ( .A1(n22355), .A2(n22759), .B1(n22354), .Y(
        j202_soc_core_j22_cpu_rf_N309) );
  sky130_fd_sc_hd__nand2_1 U26980 ( .A(n22815), .B(j202_soc_core_uart_div0[3]), 
        .Y(n22356) );
  sky130_fd_sc_hd__o21ai_1 U26982 ( .A1(n24882), .A2(n22762), .B1(n22401), .Y(
        n10574) );
  sky130_fd_sc_hd__nand2_1 U26983 ( .A(n22358), .B(n22366), .Y(n22357) );
  sky130_fd_sc_hd__o21ai_1 U26984 ( .A1(n22366), .A2(n11201), .B1(n22357), .Y(
        j202_soc_core_j22_cpu_rf_N3305) );
  sky130_fd_sc_hd__a22oi_1 U26985 ( .A1(n22358), .A2(n22369), .B1(n22362), 
        .B2(n22367), .Y(n22359) );
  sky130_fd_sc_hd__o21ai_1 U26986 ( .A1(n22372), .A2(n11201), .B1(n22359), .Y(
        j202_soc_core_j22_cpu_rf_N3379) );
  sky130_fd_sc_hd__nand2_1 U26987 ( .A(n22426), .B(n22360), .Y(n22364) );
  sky130_fd_sc_hd__o22ai_1 U26988 ( .A1(n22607), .A2(n22753), .B1(n22374), 
        .B2(n23348), .Y(n22361) );
  sky130_fd_sc_hd__a21oi_1 U26989 ( .A1(n22362), .A2(n22378), .B1(n22361), .Y(
        n22363) );
  sky130_fd_sc_hd__nand2_1 U26990 ( .A(n22364), .B(n22363), .Y(
        j202_soc_core_j22_cpu_rf_N329) );
  sky130_fd_sc_hd__nand2_1 U26991 ( .A(n22368), .B(n22366), .Y(n22365) );
  sky130_fd_sc_hd__o21ai_0 U26992 ( .A1(n22366), .A2(n22371), .B1(n22365), .Y(
        j202_soc_core_j22_cpu_rf_N3288) );
  sky130_fd_sc_hd__a22oi_1 U26993 ( .A1(n22369), .A2(n22368), .B1(n22377), 
        .B2(n22367), .Y(n22370) );
  sky130_fd_sc_hd__o21ai_0 U26994 ( .A1(n22372), .A2(n22371), .B1(n22370), .Y(
        j202_soc_core_j22_cpu_rf_N3363) );
  sky130_fd_sc_hd__o22ai_1 U26995 ( .A1(n22375), .A2(n22753), .B1(n22374), 
        .B2(n23300), .Y(n22376) );
  sky130_fd_sc_hd__a21oi_1 U26996 ( .A1(n22378), .A2(n22377), .B1(n22376), .Y(
        n22379) );
  sky130_fd_sc_hd__o21ai_1 U26997 ( .A1(n22752), .A2(n22380), .B1(n22379), .Y(
        j202_soc_core_j22_cpu_rf_N314) );
  sky130_fd_sc_hd__o21a_1 U26998 ( .A1(j202_soc_core_rst), .A2(n22381), .B1(
        n10559), .X(n10538) );
  sky130_fd_sc_hd__nand2_1 U26999 ( .A(n23222), .B(n22401), .Y(n10572) );
  sky130_fd_sc_hd__clkinv_1 U27000 ( .A(j202_soc_core_qspi_wb_wdat[20]), .Y(
        n22383) );
  sky130_fd_sc_hd__nand2_1 U27001 ( .A(n22813), .B(j202_soc_core_uart_div1[4]), 
        .Y(n22382) );
  sky130_fd_sc_hd__o21ai_1 U27002 ( .A1(n22383), .A2(n22813), .B1(n22382), .Y(
        n109) );
  sky130_fd_sc_hd__a31oi_1 U27003 ( .A1(n22386), .A2(n22385), .A3(n22384), 
        .B1(n22742), .Y(n22394) );
  sky130_fd_sc_hd__a21oi_1 U27004 ( .A1(n22387), .A2(n22408), .B1(n22407), .Y(
        n22393) );
  sky130_fd_sc_hd__nand2_1 U27005 ( .A(n25385), .B(n25387), .Y(n24866) );
  sky130_fd_sc_hd__o22ai_1 U27007 ( .A1(n22390), .A2(n22409), .B1(n24866), 
        .B2(n22419), .Y(n22391) );
  sky130_fd_sc_hd__nor4_1 U27008 ( .A(n22394), .B(n22393), .C(n22392), .D(
        n22391), .Y(n22399) );
  sky130_fd_sc_hd__nor2_1 U27009 ( .A(n25386), .B(n22395), .Y(n22397) );
  sky130_fd_sc_hd__nor4b_1 U27010 ( .D_N(n22399), .A(n22398), .B(n22397), .C(
        n22396), .Y(n22400) );
  sky130_fd_sc_hd__o22ai_1 U27011 ( .A1(n22402), .A2(n22401), .B1(n24882), 
        .B2(n22400), .Y(n10592) );
  sky130_fd_sc_hd__nand3_1 U27012 ( .A(n11036), .B(
        j202_soc_core_ahbcs_6__HREADY_), .C(n22403), .Y(n22404) );
  sky130_fd_sc_hd__nand2_1 U27013 ( .A(n22404), .B(n25732), .Y(n10537) );
  sky130_fd_sc_hd__clkinv_1 U27014 ( .A(j202_soc_core_qspi_wb_wdat[24]), .Y(
        n22406) );
  sky130_fd_sc_hd__nand2_1 U27015 ( .A(n22815), .B(j202_soc_core_uart_div0[0]), 
        .Y(n22405) );
  sky130_fd_sc_hd__o21ai_1 U27016 ( .A1(n22815), .A2(n22406), .B1(n22405), .Y(
        n69) );
  sky130_fd_sc_hd__a21oi_1 U27017 ( .A1(n22409), .A2(n22408), .B1(n22407), .Y(
        n22410) );
  sky130_fd_sc_hd__nor2_1 U27018 ( .A(n22411), .B(n22410), .Y(n22414) );
  sky130_fd_sc_hd__nand4_1 U27019 ( .A(n22415), .B(n22414), .C(n22413), .D(
        n22412), .Y(n22422) );
  sky130_fd_sc_hd__nor3_1 U27020 ( .A(n22418), .B(n22417), .C(n22416), .Y(
        n22421) );
  sky130_fd_sc_hd__nor3_1 U27021 ( .A(n22419), .B(n23222), .C(n25387), .Y(
        n22420) );
  sky130_fd_sc_hd__a211o_1 U27022 ( .A1(n22422), .A2(n24858), .B1(n22421), 
        .C1(n22420), .X(n10595) );
  sky130_fd_sc_hd__xor2_1 U27023 ( .A(n22424), .B(n22423), .X(n22425) );
  sky130_fd_sc_hd__xnor2_1 U27024 ( .A(n22425), .B(n22511), .Y(n22506) );
  sky130_fd_sc_hd__xnor2_1 U27025 ( .A(n22506), .B(n22426), .Y(n22669) );
  sky130_fd_sc_hd__nand3_1 U27026 ( .A(n22669), .B(n22706), .C(n22687), .Y(
        n22504) );
  sky130_fd_sc_hd__xnor2_1 U27027 ( .A(j202_soc_core_j22_cpu_rfuo_sr__m_), .B(
        n22427), .Y(n22502) );
  sky130_fd_sc_hd__nand2_1 U27028 ( .A(n22428), .B(n22687), .Y(n22692) );
  sky130_fd_sc_hd__nor2_1 U27029 ( .A(n22697), .B(n22429), .Y(n22671) );
  sky130_fd_sc_hd__nand2_1 U27030 ( .A(n22430), .B(n22620), .Y(n22431) );
  sky130_fd_sc_hd__nand2_1 U27031 ( .A(n22432), .B(n22431), .Y(n22434) );
  sky130_fd_sc_hd__nor2_1 U27032 ( .A(n22434), .B(n22433), .Y(n22445) );
  sky130_fd_sc_hd__clkinv_1 U27033 ( .A(n22436), .Y(n22440) );
  sky130_fd_sc_hd__nand2_1 U27034 ( .A(n22437), .B(n22619), .Y(n22438) );
  sky130_fd_sc_hd__o211a_2 U27035 ( .A1(n22441), .A2(n22440), .B1(n22439), 
        .C1(n22438), .X(n22442) );
  sky130_fd_sc_hd__nand4_1 U27036 ( .A(n22445), .B(n22444), .C(n22443), .D(
        n22442), .Y(n22674) );
  sky130_fd_sc_hd__nand4_1 U27037 ( .A(n22449), .B(n22448), .C(n22447), .D(
        n22446), .Y(n22455) );
  sky130_fd_sc_hd__clkinv_1 U27038 ( .A(n22632), .Y(n22450) );
  sky130_fd_sc_hd__a2bb2oi_1 U27039 ( .B1(n22452), .B2(n22633), .A1_N(n22451), 
        .A2_N(n22450), .Y(n22454) );
  sky130_fd_sc_hd__nand4b_1 U27040 ( .A_N(n22455), .B(n22454), .C(n22595), .D(
        n22453), .Y(n22676) );
  sky130_fd_sc_hd__nand2_1 U27041 ( .A(n22457), .B(n22456), .Y(n22469) );
  sky130_fd_sc_hd__nand2_1 U27042 ( .A(n22458), .B(n22634), .Y(n22465) );
  sky130_fd_sc_hd__nand2_1 U27043 ( .A(n22459), .B(n22624), .Y(n22464) );
  sky130_fd_sc_hd__nand2_1 U27044 ( .A(n22460), .B(n22650), .Y(n22463) );
  sky130_fd_sc_hd__nand2_1 U27045 ( .A(n22461), .B(n22623), .Y(n22462) );
  sky130_fd_sc_hd__nand4_1 U27046 ( .A(n22465), .B(n22464), .C(n22463), .D(
        n22462), .Y(n22468) );
  sky130_fd_sc_hd__a22oi_1 U27047 ( .A1(n22625), .A2(n22471), .B1(n22626), 
        .B2(n22470), .Y(n22482) );
  sky130_fd_sc_hd__a22oi_1 U27048 ( .A1(n22473), .A2(n22621), .B1(n22472), 
        .B2(n22622), .Y(n22481) );
  sky130_fd_sc_hd__a2bb2oi_1 U27049 ( .B1(n22476), .B2(n22630), .A1_N(n22475), 
        .A2_N(n22474), .Y(n22480) );
  sky130_fd_sc_hd__a22oi_1 U27050 ( .A1(n22629), .A2(n22478), .B1(n22628), 
        .B2(n22477), .Y(n22479) );
  sky130_fd_sc_hd__nand4_1 U27051 ( .A(n22482), .B(n22481), .C(n22480), .D(
        n22479), .Y(n22673) );
  sky130_fd_sc_hd__nand4_1 U27052 ( .A(n22674), .B(n22676), .C(n22675), .D(
        n22673), .Y(n22498) );
  sky130_fd_sc_hd__a21oi_1 U27053 ( .A1(n22484), .A2(n22483), .B1(n22688), .Y(
        n22485) );
  sky130_fd_sc_hd__o21ai_1 U27054 ( .A1(n22487), .A2(n22486), .B1(n22485), .Y(
        n22490) );
  sky130_fd_sc_hd__o22ai_1 U27055 ( .A1(n22612), .A2(n22520), .B1(n22488), 
        .B2(n22519), .Y(n22489) );
  sky130_fd_sc_hd__a211oi_1 U27056 ( .A1(n22725), .A2(n22584), .B1(n22490), 
        .C1(n22489), .Y(n22491) );
  sky130_fd_sc_hd__a211oi_1 U27058 ( .A1(n22496), .A2(n22495), .B1(n22494), 
        .C1(n22493), .Y(n22497) );
  sky130_fd_sc_hd__a21oi_1 U27059 ( .A1(n22671), .A2(n22498), .B1(n22497), .Y(
        n22499) );
  sky130_fd_sc_hd__a21oi_1 U27061 ( .A1(n22502), .A2(n22501), .B1(n22500), .Y(
        n22503) );
  sky130_fd_sc_hd__nand2_1 U27062 ( .A(n22504), .B(n22503), .Y(n22505) );
  sky130_fd_sc_hd__nand3_1 U27063 ( .A(n22505), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[1]), .C(n22790), .Y(n22686) );
  sky130_fd_sc_hd__nand3_1 U27064 ( .A(n22511), .B(
        j202_soc_core_j22_cpu_exuop_EXU_[4]), .C(n22790), .Y(n22507) );
  sky130_fd_sc_hd__a21oi_1 U27066 ( .A1(n22511), .A2(n22510), .B1(n22707), .Y(
        n22665) );
  sky130_fd_sc_hd__nor4_1 U27067 ( .A(n22515), .B(n22514), .C(n22513), .D(
        n22512), .Y(n22663) );
  sky130_fd_sc_hd__nand4_1 U27069 ( .A(n22723), .B(n22520), .C(n22519), .D(
        n22518), .Y(n22553) );
  sky130_fd_sc_hd__nor4_1 U27070 ( .A(n22524), .B(n22523), .C(n22522), .D(
        n22521), .Y(n22550) );
  sky130_fd_sc_hd__a31oi_1 U27071 ( .A1(n22527), .A2(n22526), .A3(n22525), 
        .B1(n22551), .Y(n22529) );
  sky130_fd_sc_hd__nor4_1 U27072 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[0]), 
        .B(n22529), .C(n22688), .D(n22528), .Y(n22535) );
  sky130_fd_sc_hd__nand2_1 U27073 ( .A(n22531), .B(n22530), .Y(n22532) );
  sky130_fd_sc_hd__nand4_1 U27074 ( .A(n22535), .B(n22534), .C(n22533), .D(
        n22532), .Y(n22546) );
  sky130_fd_sc_hd__nand2_1 U27075 ( .A(n22537), .B(n22536), .Y(n22545) );
  sky130_fd_sc_hd__nor4_1 U27076 ( .A(n22541), .B(n22540), .C(n22539), .D(
        n25388), .Y(n22543) );
  sky130_fd_sc_hd__a21oi_1 U27077 ( .A1(n22543), .A2(n22542), .B1(n22551), .Y(
        n22544) );
  sky130_fd_sc_hd__nor4_1 U27078 ( .A(n22547), .B(n22546), .C(n22545), .D(
        n22544), .Y(n22548) );
  sky130_fd_sc_hd__o211ai_1 U27079 ( .A1(n22551), .A2(n22550), .B1(n22549), 
        .C1(n22548), .Y(n22552) );
  sky130_fd_sc_hd__nor4_1 U27080 ( .A(n22555), .B(n22554), .C(n22553), .D(
        n22552), .Y(n22661) );
  sky130_fd_sc_hd__nand4_1 U27081 ( .A(n22558), .B(n22557), .C(
        j202_soc_core_j22_cpu_exuop_EXU_[0]), .D(n22556), .Y(n22572) );
  sky130_fd_sc_hd__nand4_1 U27082 ( .A(n22562), .B(n22561), .C(n22560), .D(
        n22559), .Y(n22571) );
  sky130_fd_sc_hd__nand4_1 U27083 ( .A(n22566), .B(n22565), .C(n22564), .D(
        n22563), .Y(n22570) );
  sky130_fd_sc_hd__nand4_1 U27084 ( .A(n22568), .B(n22614), .C(n22643), .D(
        n22567), .Y(n22569) );
  sky130_fd_sc_hd__nor4_1 U27085 ( .A(n22572), .B(n22571), .C(n22570), .D(
        n22569), .Y(n22588) );
  sky130_fd_sc_hd__nor4_1 U27086 ( .A(n22576), .B(n22575), .C(n22574), .D(
        n22573), .Y(n22587) );
  sky130_fd_sc_hd__nor4_1 U27087 ( .A(n22631), .B(n22579), .C(n22578), .D(
        n22577), .Y(n22586) );
  sky130_fd_sc_hd__nand4_1 U27088 ( .A(n22647), .B(n22580), .C(n22612), .D(
        n22645), .Y(n22582) );
  sky130_fd_sc_hd__nor4_1 U27089 ( .A(n22584), .B(n22583), .C(n22582), .D(
        n22581), .Y(n22585) );
  sky130_fd_sc_hd__nand4_1 U27090 ( .A(n22588), .B(n22587), .C(n22586), .D(
        n22585), .Y(n22598) );
  sky130_fd_sc_hd__nor2_1 U27091 ( .A(j202_soc_core_j22_cpu_exuop_EXU_[1]), 
        .B(n22589), .Y(n22696) );
  sky130_fd_sc_hd__a21oi_1 U27092 ( .A1(n22592), .A2(n22591), .B1(n22590), .Y(
        n22593) );
  sky130_fd_sc_hd__o22ai_1 U27093 ( .A1(n22596), .A2(n22595), .B1(n22594), 
        .B2(n22593), .Y(n22597) );
  sky130_fd_sc_hd__a31oi_1 U27094 ( .A1(n22598), .A2(n22608), .A3(n22696), 
        .B1(n22597), .Y(n22659) );
  sky130_fd_sc_hd__o22ai_1 U27095 ( .A1(n22602), .A2(n22601), .B1(n22600), 
        .B2(n22599), .Y(n22618) );
  sky130_fd_sc_hd__o22ai_1 U27096 ( .A1(n22606), .A2(n22605), .B1(n22604), 
        .B2(n22603), .Y(n22617) );
  sky130_fd_sc_hd__o22ai_1 U27097 ( .A1(n22610), .A2(n22609), .B1(n22608), 
        .B2(n22607), .Y(n22616) );
  sky130_fd_sc_hd__o22ai_1 U27098 ( .A1(n22614), .A2(n22613), .B1(n22612), 
        .B2(n22611), .Y(n22615) );
  sky130_fd_sc_hd__nor4_1 U27099 ( .A(n22618), .B(n22617), .C(n22616), .D(
        n22615), .Y(n22657) );
  sky130_fd_sc_hd__nand4_1 U27100 ( .A(n22622), .B(n22621), .C(n22620), .D(
        n22619), .Y(n22639) );
  sky130_fd_sc_hd__nand4_1 U27101 ( .A(n22626), .B(n22625), .C(n22624), .D(
        n22623), .Y(n22638) );
  sky130_fd_sc_hd__nand4_1 U27102 ( .A(n22630), .B(n22629), .C(n22628), .D(
        n22627), .Y(n22637) );
  sky130_fd_sc_hd__a211oi_1 U27103 ( .A1(n23333), .A2(n22631), .B1(n22688), 
        .C1(n22695), .Y(n22635) );
  sky130_fd_sc_hd__nand4_1 U27104 ( .A(n22635), .B(n22634), .C(n22633), .D(
        n22632), .Y(n22636) );
  sky130_fd_sc_hd__nor4_1 U27105 ( .A(n22639), .B(n22638), .C(n22637), .D(
        n22636), .Y(n22656) );
  sky130_fd_sc_hd__o22ai_1 U27106 ( .A1(n22643), .A2(n22642), .B1(n22641), 
        .B2(n22640), .Y(n22654) );
  sky130_fd_sc_hd__o22ai_1 U27107 ( .A1(n22647), .A2(n22646), .B1(n22645), 
        .B2(n22644), .Y(n22653) );
  sky130_fd_sc_hd__nand4_1 U27108 ( .A(n22651), .B(n22650), .C(n22649), .D(
        n22648), .Y(n22652) );
  sky130_fd_sc_hd__nor3_1 U27109 ( .A(n22654), .B(n22653), .C(n22652), .Y(
        n22655) );
  sky130_fd_sc_hd__nand3_1 U27110 ( .A(n22657), .B(n22656), .C(n22655), .Y(
        n22658) );
  sky130_fd_sc_hd__nand2_1 U27111 ( .A(n22659), .B(n22658), .Y(n22660) );
  sky130_fd_sc_hd__a31oi_1 U27112 ( .A1(n22663), .A2(n22662), .A3(n22661), 
        .B1(n22660), .Y(n22664) );
  sky130_fd_sc_hd__o21ai_1 U27113 ( .A1(n22694), .A2(n22665), .B1(n22664), .Y(
        n22666) );
  sky130_fd_sc_hd__a21oi_1 U27114 ( .A1(n22667), .A2(n22697), .B1(n22666), .Y(
        n22685) );
  sky130_fd_sc_hd__nand2_1 U27115 ( .A(n22669), .B(n22668), .Y(n22682) );
  sky130_fd_sc_hd__nor2_1 U27116 ( .A(n22670), .B(n22694), .Y(n22672) );
  sky130_fd_sc_hd__nor2_1 U27117 ( .A(n22672), .B(n22671), .Y(n22716) );
  sky130_fd_sc_hd__nor2_1 U27118 ( .A(n22716), .B(n22673), .Y(n22680) );
  sky130_fd_sc_hd__clkinv_1 U27119 ( .A(n22674), .Y(n22679) );
  sky130_fd_sc_hd__clkinv_1 U27120 ( .A(n22675), .Y(n22678) );
  sky130_fd_sc_hd__clkinv_1 U27121 ( .A(n22676), .Y(n22677) );
  sky130_fd_sc_hd__nand4_1 U27122 ( .A(n22680), .B(n22679), .C(n22678), .D(
        n22677), .Y(n22681) );
  sky130_fd_sc_hd__nand2_1 U27123 ( .A(n22682), .B(n22681), .Y(n22683) );
  sky130_fd_sc_hd__nand2_1 U27124 ( .A(n22683), .B(n22689), .Y(n22684) );
  sky130_fd_sc_hd__nand3_1 U27125 ( .A(n22686), .B(n22685), .C(n22684), .Y(
        n22719) );
  sky130_fd_sc_hd__o22ai_1 U27126 ( .A1(n22691), .A2(n22690), .B1(n22689), 
        .B2(n22688), .Y(n22703) );
  sky130_fd_sc_hd__o22ai_1 U27127 ( .A1(n22695), .A2(n22694), .B1(n22693), 
        .B2(n22692), .Y(n22702) );
  sky130_fd_sc_hd__a21oi_1 U27128 ( .A1(j202_soc_core_j22_cpu_exuop_EXU_[4]), 
        .A2(n22697), .B1(n22696), .Y(n22699) );
  sky130_fd_sc_hd__nor3_1 U27130 ( .A(n22703), .B(n22702), .C(n22701), .Y(
        n22714) );
  sky130_fd_sc_hd__nor2_1 U27131 ( .A(n22705), .B(n22704), .Y(n22712) );
  sky130_fd_sc_hd__nand2_1 U27132 ( .A(n22707), .B(n22706), .Y(n22709) );
  sky130_fd_sc_hd__nor2_1 U27133 ( .A(n22709), .B(n22708), .Y(n22710) );
  sky130_fd_sc_hd__nand4_1 U27134 ( .A(n22712), .B(n22754), .C(n22711), .D(
        n22710), .Y(n22713) );
  sky130_fd_sc_hd__o211ai_1 U27135 ( .A1(n22716), .A2(n22715), .B1(n22714), 
        .C1(n22713), .Y(n22717) );
  sky130_fd_sc_hd__nand2_1 U27136 ( .A(n23239), .B(n22717), .Y(n22728) );
  sky130_fd_sc_hd__nand2_1 U27137 ( .A(n22719), .B(n22718), .Y(n22727) );
  sky130_fd_sc_hd__o22ai_1 U27138 ( .A1(n22723), .A2(n22722), .B1(n22721), 
        .B2(n22720), .Y(n22724) );
  sky130_fd_sc_hd__a22oi_1 U27139 ( .A1(n24894), .A2(n22725), .B1(n22724), 
        .B2(n22728), .Y(n22726) );
  sky130_fd_sc_hd__nand2_1 U27140 ( .A(n22727), .B(n22726), .Y(
        j202_soc_core_j22_cpu_rf_N2626) );
  sky130_fd_sc_hd__nand2_1 U27141 ( .A(n22729), .B(n22728), .Y(
        j202_soc_core_j22_cpu_rf_N2625) );
  sky130_fd_sc_hd__clkinv_1 U27142 ( .A(j202_soc_core_qspi_wb_wdat[16]), .Y(
        n22731) );
  sky130_fd_sc_hd__nand2_1 U27143 ( .A(n22813), .B(j202_soc_core_uart_div1[0]), 
        .Y(n22730) );
  sky130_fd_sc_hd__a31oi_1 U27145 ( .A1(n22735), .A2(n22734), .A3(n22733), 
        .B1(n22732), .Y(n22737) );
  sky130_fd_sc_hd__o211ai_1 U27146 ( .A1(n22739), .A2(n22738), .B1(n22737), 
        .C1(n22736), .Y(n22747) );
  sky130_fd_sc_hd__o211ai_1 U27147 ( .A1(n22743), .A2(n22742), .B1(n22741), 
        .C1(n22740), .Y(n22745) );
  sky130_fd_sc_hd__nor4_1 U27148 ( .A(n22747), .B(n22746), .C(n22745), .D(
        n22744), .Y(n22749) );
  sky130_fd_sc_hd__o22ai_1 U27150 ( .A1(n22754), .A2(n22753), .B1(n22752), 
        .B2(n22751), .Y(n22755) );
  sky130_fd_sc_hd__a21oi_1 U27151 ( .A1(n22757), .A2(n22756), .B1(n22755), .Y(
        n22758) );
  sky130_fd_sc_hd__o21ai_1 U27152 ( .A1(j202_soc_core_j22_cpu_pc[1]), .A2(
        n22759), .B1(n22758), .Y(j202_soc_core_j22_cpu_rf_N299) );
  sky130_fd_sc_hd__nor3_1 U27154 ( .A(j202_soc_core_ahb2apb_00_state[2]), .B(
        n22763), .C(n22824), .Y(j202_soc_core_ahb2apb_00_N89) );
  sky130_fd_sc_hd__nor4_1 U27155 ( .A(j202_soc_core_ahb2apb_00_state[2]), .B(
        j202_soc_core_rst), .C(n22764), .D(n22767), .Y(
        j202_soc_core_ahb2apb_00_N91) );
  sky130_fd_sc_hd__nand2b_1 U27156 ( .A_N(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[1]), .B(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[0]), .Y(n22765) );
  sky130_fd_sc_hd__nand3_1 U27157 ( .A(n22766), .B(n22765), .C(n22768), .Y(
        n22769) );
  sky130_fd_sc_hd__nand3_1 U27158 ( .A(n22768), .B(
        j202_soc_core_ahb2apb_00_state[0]), .C(n22767), .Y(n24783) );
  sky130_fd_sc_hd__a21oi_1 U27159 ( .A1(n22769), .A2(n24783), .B1(
        j202_soc_core_rst), .Y(j202_soc_core_ahb2apb_00_N90) );
  sky130_fd_sc_hd__nor2_1 U27160 ( .A(j202_soc_core_wbqspiflash_00_spif_cmd), 
        .B(j202_soc_core_wbqspiflash_00_spif_ctrl), .Y(n25043) );
  sky130_fd_sc_hd__nor2_1 U27161 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(n23529), .Y(n23514) );
  sky130_fd_sc_hd__nand3_1 U27162 ( .A(n23514), .B(n22770), .C(n23513), .Y(
        n23561) );
  sky130_fd_sc_hd__o22ai_1 U27163 ( .A1(n23760), .A2(
        j202_soc_core_wbqspiflash_00_spif_cmd), .B1(
        j202_soc_core_wbqspiflash_00_spif_ctrl), .B2(
        j202_soc_core_wbqspiflash_00_write_protect), .Y(n22773) );
  sky130_fd_sc_hd__nor2_1 U27164 ( .A(n23412), .B(n22843), .Y(n25042) );
  sky130_fd_sc_hd__nor2_1 U27165 ( .A(n25046), .B(n24995), .Y(n23480) );
  sky130_fd_sc_hd__nor2_1 U27166 ( .A(n23513), .B(n24899), .Y(n25116) );
  sky130_fd_sc_hd__nand2_1 U27167 ( .A(n25027), .B(n25116), .Y(n23417) );
  sky130_fd_sc_hd__clkinv_1 U27168 ( .A(n25086), .Y(n23251) );
  sky130_fd_sc_hd__clkinv_1 U27169 ( .A(n25100), .Y(n23370) );
  sky130_fd_sc_hd__o22ai_1 U27170 ( .A1(j202_soc_core_wbqspiflash_00_spi_busy), 
        .A2(n23251), .B1(n25099), .B2(n23370), .Y(n23520) );
  sky130_fd_sc_hd__a211oi_1 U27171 ( .A1(n23480), .A2(n22838), .B1(n23520), 
        .C1(n22771), .Y(n22772) );
  sky130_fd_sc_hd__o31ai_1 U27172 ( .A1(n25043), .A2(n23561), .A3(n22773), 
        .B1(n22772), .Y(n22780) );
  sky130_fd_sc_hd__clkinv_1 U27173 ( .A(n23428), .Y(n22774) );
  sky130_fd_sc_hd__nand2_1 U27174 ( .A(n22774), .B(n23494), .Y(n22776) );
  sky130_fd_sc_hd__a31oi_1 U27175 ( .A1(n22776), .A2(
        j202_soc_core_qspi_wb_addr[24]), .A3(n23289), .B1(n22775), .Y(n22777)
         );
  sky130_fd_sc_hd__nand2_1 U27176 ( .A(n23404), .B(n23364), .Y(n25035) );
  sky130_fd_sc_hd__o22ai_1 U27177 ( .A1(n22777), .A2(n23523), .B1(n23758), 
        .B2(n25035), .Y(n22778) );
  sky130_fd_sc_hd__a211oi_1 U27178 ( .A1(j202_soc_core_wbqspiflash_00_spif_req), .A2(n22780), .B1(n22779), .C1(n22778), .Y(n22782) );
  sky130_fd_sc_hd__nand2_1 U27179 ( .A(n23364), .B(n23403), .Y(n25036) );
  sky130_fd_sc_hd__clkinv_1 U27180 ( .A(n25036), .Y(n22781) );
  sky130_fd_sc_hd__nand2_1 U27181 ( .A(n25389), .B(n22781), .Y(n23474) );
  sky130_fd_sc_hd__o21ai_1 U27182 ( .A1(j202_soc_core_rst), .A2(n22782), .B1(
        n23474), .Y(j202_soc_core_wbqspiflash_00_N730) );
  sky130_fd_sc_hd__nand2_1 U27183 ( .A(n25390), .B(n22783), .Y(n22784) );
  sky130_fd_sc_hd__o21ai_0 U27184 ( .A1(n22786), .A2(n22785), .B1(n22784), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N6) );
  sky130_fd_sc_hd__a21oi_1 U27185 ( .A1(n24879), .A2(n22788), .B1(n22787), .Y(
        n22795) );
  sky130_fd_sc_hd__a21oi_1 U27186 ( .A1(n22791), .A2(n22790), .B1(n22789), .Y(
        n22794) );
  sky130_fd_sc_hd__nand3_1 U27187 ( .A(n23239), .B(n22794), .C(n22793), .Y(
        n23224) );
  sky130_fd_sc_hd__o21ai_1 U27188 ( .A1(n23232), .A2(n22795), .B1(n23224), .Y(
        n10567) );
  sky130_fd_sc_hd__o21ai_0 U27189 ( .A1(n22797), .A2(n24882), .B1(n22796), .Y(
        n10587) );
  sky130_fd_sc_hd__nand4b_1 U27190 ( .A_N(n22801), .B(n22800), .C(n22799), .D(
        n22798), .Y(n22806) );
  sky130_fd_sc_hd__a21oi_1 U27191 ( .A1(n22804), .A2(n22803), .B1(n22802), .Y(
        n22805) );
  sky130_fd_sc_hd__nand2_1 U27193 ( .A(n22808), .B(n22807), .Y(n10605) );
  sky130_fd_sc_hd__nand2_1 U27194 ( .A(n22815), .B(j202_soc_core_uart_div0[5]), 
        .Y(n22809) );
  sky130_fd_sc_hd__o21ai_1 U27195 ( .A1(n22815), .A2(n24046), .B1(n22809), .Y(
        n72) );
  sky130_fd_sc_hd__nand2_1 U27196 ( .A(n22815), .B(j202_soc_core_uart_div0[1]), 
        .Y(n22810) );
  sky130_fd_sc_hd__o21ai_1 U27197 ( .A1(n22815), .A2(n24019), .B1(n22810), .Y(
        n135) );
  sky130_fd_sc_hd__nand2_1 U27198 ( .A(n22813), .B(j202_soc_core_uart_div1[5]), 
        .Y(n22811) );
  sky130_fd_sc_hd__o21ai_1 U27199 ( .A1(n23997), .A2(n22813), .B1(n22811), .Y(
        n110) );
  sky130_fd_sc_hd__nand2_1 U27200 ( .A(n22813), .B(j202_soc_core_uart_div1[6]), 
        .Y(n22812) );
  sky130_fd_sc_hd__o21ai_1 U27201 ( .A1(n24000), .A2(n22813), .B1(n22812), .Y(
        n74) );
  sky130_fd_sc_hd__nand2_1 U27202 ( .A(n22815), .B(j202_soc_core_uart_div0[7]), 
        .Y(n22814) );
  sky130_fd_sc_hd__nor2_1 U27204 ( .A(n22816), .B(n22824), .Y(
        j202_soc_core_ahb2apb_00_N24) );
  sky130_fd_sc_hd__nor2_1 U27205 ( .A(n22818), .B(n22824), .Y(
        j202_soc_core_ahb2apb_00_N29) );
  sky130_fd_sc_hd__nor2_1 U27206 ( .A(n22819), .B(n22824), .Y(
        j202_soc_core_ahb2apb_00_N30) );
  sky130_fd_sc_hd__nor2_1 U27207 ( .A(n22821), .B(n22824), .Y(
        j202_soc_core_ahb2apb_00_N55) );
  sky130_fd_sc_hd__nor2_1 U27208 ( .A(n22823), .B(n22824), .Y(
        j202_soc_core_ahb2apb_00_N26) );
  sky130_fd_sc_hd__nor2_1 U27209 ( .A(n22825), .B(n22824), .Y(
        j202_soc_core_ahb2apb_00_N25) );
  sky130_fd_sc_hd__nand2_1 U27210 ( .A(n22826), .B(n25391), .Y(n22832) );
  sky130_fd_sc_hd__a22oi_1 U27211 ( .A1(n22829), .A2(n22828), .B1(n10994), 
        .B2(n22827), .Y(n22831) );
  sky130_fd_sc_hd__nand3_1 U27212 ( .A(n22832), .B(n22831), .C(n22830), .Y(
        j202_soc_core_ahb2aqu_00_N161) );
  sky130_fd_sc_hd__nor3_1 U27213 ( .A(j202_soc_core_wbqspiflash_00_state[3]), 
        .B(j202_soc_core_wbqspiflash_00_state[0]), .C(n23513), .Y(n23490) );
  sky130_fd_sc_hd__nor2_1 U27214 ( .A(j202_soc_core_wbqspiflash_00_spif_cmd), 
        .B(n25015), .Y(n25051) );
  sky130_fd_sc_hd__nand2_1 U27215 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .B(n25051), .Y(n25032)
         );
  sky130_fd_sc_hd__nor2_1 U27216 ( .A(n24901), .B(n25032), .Y(n25094) );
  sky130_fd_sc_hd__nor2_1 U27217 ( .A(n24998), .B(n25094), .Y(n23456) );
  sky130_fd_sc_hd__nand2_1 U27218 ( .A(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled), .B(n25043), .Y(n23413) );
  sky130_fd_sc_hd__and3_1 U27219 ( .A(n23456), .B(n24995), .C(n23413), .X(
        n23441) );
  sky130_fd_sc_hd__nand2_1 U27220 ( .A(n23395), .B(n23541), .Y(n23445) );
  sky130_fd_sc_hd__nor2_1 U27221 ( .A(n23513), .B(n23445), .Y(n25025) );
  sky130_fd_sc_hd__clkinv_1 U27222 ( .A(n25025), .Y(n23466) );
  sky130_fd_sc_hd__a21oi_1 U27224 ( .A1(n23525), .A2(n23422), .B1(n23295), .Y(
        n22836) );
  sky130_fd_sc_hd__nand2_1 U27225 ( .A(n23382), .B(n23495), .Y(n23465) );
  sky130_fd_sc_hd__nor2_1 U27226 ( .A(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled), .B(n23465), .Y(n23408) );
  sky130_fd_sc_hd__clkinv_1 U27227 ( .A(n22833), .Y(n25048) );
  sky130_fd_sc_hd__nor2_1 U27228 ( .A(n22834), .B(n25048), .Y(n25024) );
  sky130_fd_sc_hd__o21ai_1 U27229 ( .A1(n23408), .A2(n23461), .B1(n23364), .Y(
        n22835) );
  sky130_fd_sc_hd__nand2b_1 U27230 ( .A_N(n23478), .B(n25102), .Y(n25072) );
  sky130_fd_sc_hd__nand4_1 U27231 ( .A(n22836), .B(n25107), .C(n22835), .D(
        n25072), .Y(n22837) );
  sky130_fd_sc_hd__a31oi_1 U27232 ( .A1(n23490), .A2(n22838), .A3(n23441), 
        .B1(n22837), .Y(n22842) );
  sky130_fd_sc_hd__nand2_1 U27233 ( .A(n25051), .B(n22839), .Y(n25013) );
  sky130_fd_sc_hd__nor3_1 U27234 ( .A(n23760), .B(n23445), .C(n25013), .Y(
        n23470) );
  sky130_fd_sc_hd__nor2_1 U27235 ( .A(n22847), .B(n22852), .Y(n23376) );
  sky130_fd_sc_hd__clkinv_1 U27236 ( .A(n23376), .Y(n23467) );
  sky130_fd_sc_hd__nand2_1 U27237 ( .A(n25011), .B(n23467), .Y(n22840) );
  sky130_fd_sc_hd__a21oi_1 U27238 ( .A1(n23470), .A2(n22847), .B1(n22840), .Y(
        n22841) );
  sky130_fd_sc_hd__nand2_1 U27239 ( .A(n23364), .B(n23463), .Y(n25004) );
  sky130_fd_sc_hd__a31oi_1 U27240 ( .A1(n22842), .A2(n22841), .A3(n25004), 
        .B1(j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N736) );
  sky130_fd_sc_hd__a21oi_1 U27241 ( .A1(n25116), .A2(n25070), .B1(n23395), .Y(
        n23355) );
  sky130_fd_sc_hd__nand2_1 U27242 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(n23526), .Y(n22846) );
  sky130_fd_sc_hd__a21oi_1 U27243 ( .A1(n25005), .A2(n22844), .B1(n22843), .Y(
        n22845) );
  sky130_fd_sc_hd__a31oi_1 U27244 ( .A1(n23355), .A2(n22847), .A3(n22846), 
        .B1(n22845), .Y(n22849) );
  sky130_fd_sc_hd__nand3_1 U27245 ( .A(n25116), .B(n23535), .C(n25070), .Y(
        n23577) );
  sky130_fd_sc_hd__nand2_1 U27246 ( .A(n23577), .B(n23467), .Y(n25104) );
  sky130_fd_sc_hd__clkinv_1 U27247 ( .A(n25104), .Y(n22848) );
  sky130_fd_sc_hd__nand4_1 U27248 ( .A(n22850), .B(n22849), .C(n25731), .D(
        n22848), .Y(j202_soc_core_wbqspiflash_00_N735) );
  sky130_fd_sc_hd__clkinv_1 U27249 ( .A(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled), .Y(n25061) );
  sky130_fd_sc_hd__nor2_1 U27250 ( .A(j202_soc_core_wbqspiflash_00_state[4]), 
        .B(n25011), .Y(n25077) );
  sky130_fd_sc_hd__nor2_1 U27251 ( .A(n24898), .B(n25077), .Y(n25112) );
  sky130_fd_sc_hd__nand4_1 U27253 ( .A(n25112), .B(n22852), .C(n23468), .D(
        n22851), .Y(n22853) );
  sky130_fd_sc_hd__a31oi_1 U27254 ( .A1(n25043), .A2(n22854), .A3(n25061), 
        .B1(n22853), .Y(n22855) );
  sky130_fd_sc_hd__nor2_1 U27255 ( .A(j202_soc_core_rst), .B(n22855), .Y(
        j202_soc_core_wbqspiflash_00_N737) );
  sky130_fd_sc_hd__nand2_1 U27256 ( .A(n22856), .B(
        j202_soc_core_wbqspiflash_00_spi_busy), .Y(n23354) );
  sky130_fd_sc_hd__a21oi_1 U27257 ( .A1(n23514), .A2(n23354), .B1(n25104), .Y(
        n22857) );
  sky130_fd_sc_hd__nand2_1 U27258 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(j202_soc_core_wbqspiflash_00_state[4]), .Y(n23505) );
  sky130_fd_sc_hd__nor2_1 U27259 ( .A(n23435), .B(n23505), .Y(n23420) );
  sky130_fd_sc_hd__nand2_1 U27260 ( .A(j202_soc_core_wbqspiflash_00_state[2]), 
        .B(n23420), .Y(n25073) );
  sky130_fd_sc_hd__nand4_1 U27261 ( .A(n22857), .B(n23528), .C(n25046), .D(
        n25073), .Y(n23351) );
  sky130_fd_sc_hd__o21a_1 U27262 ( .A1(n22858), .A2(n23351), .B1(n25734), .X(
        j202_soc_core_wbqspiflash_00_N746) );
  sky130_fd_sc_hd__nor2_1 U27263 ( .A(n23697), .B(n23597), .Y(n22859) );
  sky130_fd_sc_hd__nand2_1 U27264 ( .A(n23593), .B(n23740), .Y(n23753) );
  sky130_fd_sc_hd__nor2_1 U27265 ( .A(j202_soc_core_wbqspiflash_00_spi_hold), 
        .B(n23753), .Y(n23596) );
  sky130_fd_sc_hd__or4_1 U27266 ( .A(n23690), .B(n22860), .C(n22859), .D(
        n23596), .X(j202_soc_core_wbqspiflash_00_lldriver_N308) );
  sky130_fd_sc_hd__nand2_1 U27267 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B(n23734), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N423) );
  sky130_fd_sc_hd__a211o_1 U27268 ( .A1(U7_RSOP_1488_C3_DATA3_2), .A2(n23747), 
        .B1(n22880), .C1(n25392), .X(
        j202_soc_core_wbqspiflash_00_lldriver_N427) );
  sky130_fd_sc_hd__nand2_1 U27269 ( .A(n23590), .B(n23690), .Y(n23609) );
  sky130_fd_sc_hd__nand4_1 U27270 ( .A(n23609), .B(n23731), .C(n22862), .D(
        n23608), .Y(j202_soc_core_wbqspiflash_00_lldriver_N424) );
  sky130_fd_sc_hd__o21ai_1 U27271 ( .A1(j202_soc_core_wbqspiflash_00_spi_spd), 
        .A2(n22862), .B1(n22861), .Y(n23742) );
  sky130_fd_sc_hd__xnor2_1 U27272 ( .A(n22864), .B(n22866), .Y(n22865) );
  sky130_fd_sc_hd__or2_0 U27273 ( .A(n23742), .B(n22865), .X(
        j202_soc_core_wbqspiflash_00_lldriver_N426) );
  sky130_fd_sc_hd__o211ai_1 U27274 ( .A1(n22868), .A2(n22867), .B1(n23694), 
        .C1(n22866), .Y(j202_soc_core_wbqspiflash_00_lldriver_N425) );
  sky130_fd_sc_hd__nor2_1 U27275 ( .A(j202_soc_core_wbqspiflash_00_spi_len[0]), 
        .B(j202_soc_core_wbqspiflash_00_lldriver_N311), .Y(n22873) );
  sky130_fd_sc_hd__clkinv_1 U27276 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[3]), .Y(n22869) );
  sky130_fd_sc_hd__o22ai_1 U27277 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_len[0]), .A2(n23699), .B1(n23612), 
        .B2(n22869), .Y(n22870) );
  sky130_fd_sc_hd__nor2_1 U27278 ( .A(n22870), .B(DP_OP_1501J1_126_8405_n3), 
        .Y(n22874) );
  sky130_fd_sc_hd__a21oi_1 U27279 ( .A1(DP_OP_1501J1_126_8405_n3), .A2(n22870), 
        .B1(n22874), .Y(n22871) );
  sky130_fd_sc_hd__a21oi_1 U27280 ( .A1(n23612), .A2(n23699), .B1(n22871), .Y(
        n22872) );
  sky130_fd_sc_hd__a211o_1 U27281 ( .A1(n22880), .A2(
        j202_soc_core_wbqspiflash_00_spi_len[0]), .B1(n22873), .C1(n22872), 
        .X(j202_soc_core_wbqspiflash_00_lldriver_N428) );
  sky130_fd_sc_hd__xor2_1 U27282 ( .A(j202_soc_core_wbqspiflash_00_spi_len[0]), 
        .B(j202_soc_core_wbqspiflash_00_spi_len[1]), .X(n22879) );
  sky130_fd_sc_hd__a22oi_1 U27283 ( .A1(n25392), .A2(n22879), .B1(n23747), 
        .B2(j202_soc_core_wbqspiflash_00_lldriver_spi_len[4]), .Y(n22875) );
  sky130_fd_sc_hd__nand2_1 U27284 ( .A(n22874), .B(n22875), .Y(n22883) );
  sky130_fd_sc_hd__a21oi_1 U27285 ( .A1(n22883), .A2(n22875), .B1(n22886), .Y(
        n22876) );
  sky130_fd_sc_hd__a22oi_1 U27287 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_len[1]), .A2(n22880), .B1(n23690), 
        .B2(n22879), .Y(n22881) );
  sky130_fd_sc_hd__nand2_1 U27288 ( .A(n22882), .B(n22881), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N429) );
  sky130_fd_sc_hd__nand2_1 U27289 ( .A(j202_soc_core_wbqspiflash_00_spi_len[1]), .B(j202_soc_core_wbqspiflash_00_spi_len[0]), .Y(n22887) );
  sky130_fd_sc_hd__clkinv_1 U27290 ( .A(n22887), .Y(n23533) );
  sky130_fd_sc_hd__a22oi_1 U27291 ( .A1(n25392), .A2(n23533), .B1(n23747), 
        .B2(j202_soc_core_wbqspiflash_00_lldriver_spi_len[5]), .Y(n22884) );
  sky130_fd_sc_hd__xnor2_1 U27292 ( .A(n22884), .B(n22883), .Y(n22885) );
  sky130_fd_sc_hd__o22ai_1 U27293 ( .A1(n22887), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B1(n22886), .B2(n22885), 
        .Y(j202_soc_core_wbqspiflash_00_lldriver_N430) );
  sky130_fd_sc_hd__nand2_1 U27294 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[0]), 
        .B(j202_soc_core_ahb2apb_02_hsize_buf[1]), .Y(
        j202_soc_core_ahb2apb_02_N123) );
  sky130_fd_sc_hd__clkinv_1 U27295 ( .A(j202_soc_core_gpio_core_00_reg_addr[1]), .Y(n22891) );
  sky130_fd_sc_hd__clkinv_1 U27296 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[0]), 
        .Y(n22889) );
  sky130_fd_sc_hd__nand2_1 U27297 ( .A(n22891), .B(n22889), .Y(n22894) );
  sky130_fd_sc_hd__nor2_1 U27298 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[1]), 
        .B(n22889), .Y(n22892) );
  sky130_fd_sc_hd__clkinv_1 U27299 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[1]), 
        .Y(n22888) );
  sky130_fd_sc_hd__nor2_1 U27300 ( .A(j202_soc_core_ahb2apb_02_hsize_buf[0]), 
        .B(n22888), .Y(n22890) );
  sky130_fd_sc_hd__a21oi_1 U27301 ( .A1(j202_soc_core_gpio_core_00_reg_addr[1]), .A2(n22892), .B1(n22890), .Y(n22893) );
  sky130_fd_sc_hd__o21ai_0 U27302 ( .A1(j202_soc_core_gpio_core_00_reg_addr[0]), .A2(n22894), .B1(n22893), .Y(n10904) );
  sky130_fd_sc_hd__nand2_1 U27303 ( .A(j202_soc_core_gpio_core_00_reg_addr[1]), 
        .B(n22889), .Y(n22897) );
  sky130_fd_sc_hd__a21oi_1 U27304 ( .A1(n22892), .A2(n22891), .B1(n22890), .Y(
        n22895) );
  sky130_fd_sc_hd__o21ai_0 U27305 ( .A1(j202_soc_core_gpio_core_00_reg_addr[0]), .A2(n22897), .B1(n22895), .Y(n10902) );
  sky130_fd_sc_hd__clkinv_1 U27306 ( .A(j202_soc_core_gpio_core_00_reg_addr[0]), .Y(n22896) );
  sky130_fd_sc_hd__o21ai_0 U27307 ( .A1(n22894), .A2(n22896), .B1(n22893), .Y(
        n10903) );
  sky130_fd_sc_hd__o21ai_0 U27308 ( .A1(n22897), .A2(n22896), .B1(n22895), .Y(
        n10901) );
  sky130_fd_sc_hd__a22o_1 U27309 ( .A1(n25393), .A2(j202_soc_core_intr_vec__6_), .B1(n22898), .B2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[6]), .X(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N9) );
  sky130_fd_sc_hd__clkinv_1 U27310 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[1]), .Y(n24244) );
  sky130_fd_sc_hd__o22ai_1 U27311 ( .A1(n22906), .A2(n24244), .B1(n22899), 
        .B2(n22904), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N4) );
  sky130_fd_sc_hd__clkinv_1 U27312 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[4]), .Y(n24189) );
  sky130_fd_sc_hd__o22ai_1 U27313 ( .A1(n22906), .A2(n24189), .B1(n22900), 
        .B2(n22904), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N7) );
  sky130_fd_sc_hd__clkinv_1 U27314 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .Y(n22902) );
  sky130_fd_sc_hd__o22ai_1 U27315 ( .A1(n22906), .A2(n22902), .B1(n22901), 
        .B2(n22904), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N3) );
  sky130_fd_sc_hd__clkinv_1 U27316 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]), .Y(n24238) );
  sky130_fd_sc_hd__o22ai_1 U27317 ( .A1(n22906), .A2(n24238), .B1(n22903), 
        .B2(n22904), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N5) );
  sky130_fd_sc_hd__clkinv_1 U27318 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[3]), .Y(n24237) );
  sky130_fd_sc_hd__o22ai_1 U27319 ( .A1(n22906), .A2(n24237), .B1(n22905), 
        .B2(n22904), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_bs_intr_vec_1_N6) );
  sky130_fd_sc_hd__nand2_1 U27320 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[0]), 
        .B(j202_soc_core_ahb2apb_01_hsize_buf[1]), .Y(
        j202_soc_core_ahb2apb_01_N123) );
  sky130_fd_sc_hd__clkinv_1 U27321 ( .A(j202_soc_core_intc_core_00_bs_addr[0]), 
        .Y(n22915) );
  sky130_fd_sc_hd__clkinv_1 U27322 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[0]), 
        .Y(n22909) );
  sky130_fd_sc_hd__nor2_1 U27323 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[1]), 
        .B(n22909), .Y(n22912) );
  sky130_fd_sc_hd__clkinv_1 U27324 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[1]), 
        .Y(n22907) );
  sky130_fd_sc_hd__nor2_1 U27325 ( .A(j202_soc_core_ahb2apb_01_hsize_buf[0]), 
        .B(n22907), .Y(n22910) );
  sky130_fd_sc_hd__a21oi_1 U27326 ( .A1(j202_soc_core_intc_core_00_bs_addr[1]), 
        .A2(n22912), .B1(n22910), .Y(n22908) );
  sky130_fd_sc_hd__o31ai_1 U27327 ( .A1(j202_soc_core_intc_core_00_bs_addr[1]), 
        .A2(j202_soc_core_ahb2apb_01_hsize_buf[0]), .A3(n22915), .B1(n22908), 
        .Y(n10744) );
  sky130_fd_sc_hd__o21ai_0 U27328 ( .A1(j202_soc_core_ahb2apb_01_hsize_buf[0]), 
        .A2(n24446), .B1(n22908), .Y(n10745) );
  sky130_fd_sc_hd__nand2_1 U27329 ( .A(j202_soc_core_intc_core_00_bs_addr[1]), 
        .B(n22909), .Y(n22914) );
  sky130_fd_sc_hd__clkinv_1 U27330 ( .A(j202_soc_core_intc_core_00_bs_addr[1]), 
        .Y(n22911) );
  sky130_fd_sc_hd__a21oi_1 U27331 ( .A1(n22912), .A2(n22911), .B1(n22910), .Y(
        n22913) );
  sky130_fd_sc_hd__o21ai_0 U27332 ( .A1(j202_soc_core_intc_core_00_bs_addr[0]), 
        .A2(n22914), .B1(n22913), .Y(n10743) );
  sky130_fd_sc_hd__o21ai_0 U27333 ( .A1(n22915), .A2(n22914), .B1(n22913), .Y(
        n10742) );
  sky130_fd_sc_hd__nand2_1 U27334 ( .A(n23254), .B(j202_soc_core_uart_din_i[1]), .Y(n22916) );
  sky130_fd_sc_hd__clkinv_1 U27336 ( .A(n23417), .Y(n25106) );
  sky130_fd_sc_hd__nand2_1 U27337 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(n25106), .Y(n23583) );
  sky130_fd_sc_hd__o21ai_1 U27338 ( .A1(n23756), .A2(n23494), .B1(n23583), .Y(
        j202_soc_core_wbqspiflash_00_N663) );
  sky130_fd_sc_hd__nand2_1 U27339 ( .A(n23254), .B(j202_soc_core_uart_din_i[2]), .Y(n22917) );
  sky130_fd_sc_hd__clkinv_1 U27341 ( .A(j202_soc_core_qspi_wb_wdat[0]), .Y(
        n22919) );
  sky130_fd_sc_hd__nand2_1 U27342 ( .A(n23254), .B(j202_soc_core_uart_din_i[0]), .Y(n22918) );
  sky130_fd_sc_hd__clkinv_1 U27344 ( .A(n22920), .Y(n22921) );
  sky130_fd_sc_hd__nand2_1 U27345 ( .A(j202_soc_core_ahbcs_6__HREADY_), .B(
        n22921), .Y(n23246) );
  sky130_fd_sc_hd__o211ai_1 U27346 ( .A1(n22923), .A2(n23248), .B1(n22922), 
        .C1(n23246), .Y(j202_soc_core_j22_cpu_ml_N192) );
  sky130_fd_sc_hd__nand2_1 U27347 ( .A(n23254), .B(j202_soc_core_uart_din_i[3]), .Y(n22924) );
  sky130_fd_sc_hd__clkinv_1 U27349 ( .A(j202_soc_core_qspi_wb_wdat[4]), .Y(
        n22926) );
  sky130_fd_sc_hd__nand2_1 U27350 ( .A(n23254), .B(j202_soc_core_uart_din_i[4]), .Y(n22925) );
  sky130_fd_sc_hd__o21ai_1 U27351 ( .A1(n22926), .A2(n23254), .B1(n22925), .Y(
        n91) );
  sky130_fd_sc_hd__nand2_1 U27352 ( .A(n23254), .B(j202_soc_core_uart_din_i[5]), .Y(n22927) );
  sky130_fd_sc_hd__o21ai_1 U27353 ( .A1(n23897), .A2(n23254), .B1(n22927), .Y(
        n90) );
  sky130_fd_sc_hd__nand2_1 U27354 ( .A(n23254), .B(j202_soc_core_uart_din_i[6]), .Y(n22928) );
  sky130_fd_sc_hd__o21ai_1 U27355 ( .A1(n23903), .A2(n23254), .B1(n22928), .Y(
        n89) );
  sky130_fd_sc_hd__nand2_1 U27356 ( .A(n23254), .B(j202_soc_core_uart_din_i[7]), .Y(n22929) );
  sky130_fd_sc_hd__clkinv_1 U27358 ( .A(j202_soc_core_pwrite[0]), .Y(n22930)
         );
  sky130_fd_sc_hd__nor2_1 U27359 ( .A(n22930), .B(n24783), .Y(
        j202_soc_core_cmt_core_00_cmt_apb_00_reg_wen) );
  sky130_fd_sc_hd__clkinv_1 U27360 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]), .Y(n22954) );
  sky130_fd_sc_hd__clkinv_1 U27361 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[4]), .Y(n22957) );
  sky130_fd_sc_hd__clkinv_1 U27362 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[2]), .Y(n25138) );
  sky130_fd_sc_hd__nand2_1 U27363 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .Y(n22961) );
  sky130_fd_sc_hd__nor2_1 U27364 ( .A(n25138), .B(n22961), .Y(n22960) );
  sky130_fd_sc_hd__nand2_1 U27365 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[3]), .B(n22960), .Y(
        n22958) );
  sky130_fd_sc_hd__nor2_1 U27366 ( .A(n22957), .B(n22958), .Y(n22944) );
  sky130_fd_sc_hd__clkinv_1 U27367 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[6]), .Y(n25178) );
  sky130_fd_sc_hd__o22ai_1 U27368 ( .A1(n25172), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .B1(n25178), .B2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .Y(n22931) );
  sky130_fd_sc_hd__a221oi_1 U27369 ( .A1(n25172), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .B1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .B2(n25178), .C1(
        n22931), .Y(n22943) );
  sky130_fd_sc_hd__clkinv_1 U27370 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[3]), .Y(n25140) );
  sky130_fd_sc_hd__o22ai_1 U27371 ( .A1(n25156), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .B1(n25140), .B2(
        j202_soc_core_bldc_core_00_pwm_period[3]), .Y(n22932) );
  sky130_fd_sc_hd__a221oi_1 U27372 ( .A1(n25156), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .B1(
        j202_soc_core_bldc_core_00_pwm_period[3]), .B2(n25140), .C1(n22932), 
        .Y(n22942) );
  sky130_fd_sc_hd__clkinv_1 U27373 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .Y(n25129) );
  sky130_fd_sc_hd__o22ai_1 U27374 ( .A1(n25180), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]), .B1(n25129), .B2(
        j202_soc_core_bldc_core_00_pwm_period[10]), .Y(n22933) );
  sky130_fd_sc_hd__a221oi_1 U27375 ( .A1(n25180), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]), .B1(
        j202_soc_core_bldc_core_00_pwm_period[10]), .B2(n25129), .C1(n22933), 
        .Y(n22941) );
  sky130_fd_sc_hd__o22ai_1 U27376 ( .A1(
        j202_soc_core_bldc_core_00_pwm_period[4]), .A2(n22957), .B1(n25174), 
        .B2(j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[4]), .Y(n22939) );
  sky130_fd_sc_hd__o2bb2ai_1 U27377 ( .B1(
        j202_soc_core_bldc_core_00_pwm_period[2]), .B2(n25138), .A1_N(
        j202_soc_core_bldc_core_00_pwm_period[2]), .A2_N(n25138), .Y(n22938)
         );
  sky130_fd_sc_hd__clkinv_1 U27378 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[11]), .Y(n25125) );
  sky130_fd_sc_hd__o22ai_1 U27379 ( .A1(
        j202_soc_core_bldc_core_00_pwm_period[11]), .A2(n25125), .B1(n25184), 
        .B2(j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[11]), .Y(n22937) );
  sky130_fd_sc_hd__clkinv_1 U27380 ( .A(
        j202_soc_core_bldc_core_00_pwm_period[5]), .Y(n25176) );
  sky130_fd_sc_hd__o22ai_1 U27381 ( .A1(n25182), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .B1(n25153), .B2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]), .Y(n22934) );
  sky130_fd_sc_hd__a221oi_1 U27382 ( .A1(n25182), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .B1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]), .B2(n25153), .C1(
        n22934), .Y(n22935) );
  sky130_fd_sc_hd__o221ai_1 U27383 ( .A1(
        j202_soc_core_bldc_core_00_pwm_period[5]), .A2(n22954), .B1(n25176), 
        .B2(j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]), .C1(n22935), 
        .Y(n22936) );
  sky130_fd_sc_hd__nor4_1 U27384 ( .A(n22939), .B(n22938), .C(n22937), .D(
        n22936), .Y(n22940) );
  sky130_fd_sc_hd__nand4_1 U27385 ( .A(n22943), .B(n22942), .C(n22941), .D(
        n22940), .Y(n25149) );
  sky130_fd_sc_hd__nand2_1 U27386 ( .A(n22944), .B(n25149), .Y(n22955) );
  sky130_fd_sc_hd__nor2_1 U27387 ( .A(n22954), .B(n22955), .Y(n22951) );
  sky130_fd_sc_hd__nand2_1 U27388 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .B(n22951), .Y(
        n22953) );
  sky130_fd_sc_hd__nand2_1 U27389 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]), .B(n25149), .Y(
        n22950) );
  sky130_fd_sc_hd__nor2_1 U27390 ( .A(n22953), .B(n22950), .Y(n22949) );
  sky130_fd_sc_hd__nand2_1 U27391 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .B(n22949), .Y(
        n22948) );
  sky130_fd_sc_hd__nand2_1 U27392 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]), .B(n25149), .Y(
        n22946) );
  sky130_fd_sc_hd__nor2_1 U27393 ( .A(n22948), .B(n22946), .Y(n22964) );
  sky130_fd_sc_hd__a21oi_1 U27394 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .A2(n25149), .B1(
        n22964), .Y(n22945) );
  sky130_fd_sc_hd__a21oi_1 U27395 ( .A1(n22964), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .B1(n22945), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[10]) );
  sky130_fd_sc_hd__a21oi_1 U27396 ( .A1(n22948), .A2(n22946), .B1(n22964), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[9]) );
  sky130_fd_sc_hd__a21oi_1 U27397 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .A2(n25149), .B1(
        n22949), .Y(n22947) );
  sky130_fd_sc_hd__nor2b_1 U27398 ( .B_N(n22948), .A(n22947), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[8]) );
  sky130_fd_sc_hd__a21oi_1 U27399 ( .A1(n22953), .A2(n22950), .B1(n22949), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[7]) );
  sky130_fd_sc_hd__a21oi_1 U27400 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .A2(n25149), .B1(
        n22951), .Y(n22952) );
  sky130_fd_sc_hd__nor2b_1 U27401 ( .B_N(n22953), .A(n22952), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[6]) );
  sky130_fd_sc_hd__o22ai_1 U27403 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]), .A2(n22955), .B1(
        n22954), .B2(n22956), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[5]) );
  sky130_fd_sc_hd__a21oi_1 U27404 ( .A1(n22957), .A2(n22958), .B1(n22956), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[4]) );
  sky130_fd_sc_hd__o21ai_1 U27405 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[3]), .A2(n22960), .B1(
        n22958), .Y(n22959) );
  sky130_fd_sc_hd__nor2_1 U27406 ( .A(n22963), .B(n22959), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[3]) );
  sky130_fd_sc_hd__a211oi_1 U27407 ( .A1(n25138), .A2(n22961), .B1(n22960), 
        .C1(n22963), .Y(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[2])
         );
  sky130_fd_sc_hd__o21ai_1 U27408 ( .A1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .B1(n22961), .Y(
        n22962) );
  sky130_fd_sc_hd__nor2_1 U27409 ( .A(n22963), .B(n22962), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[1]) );
  sky130_fd_sc_hd__nand2_1 U27410 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .B(n25149), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[0]) );
  sky130_fd_sc_hd__nand2_1 U27411 ( .A(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .B(n22964), .Y(
        n22966) );
  sky130_fd_sc_hd__nand2_1 U27412 ( .A(n25149), .B(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[11]), .Y(n22965) );
  sky130_fd_sc_hd__xor2_1 U27413 ( .A(n22966), .B(n22965), .X(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_clkcnt[11]) );
  sky130_fd_sc_hd__or3_1 U27414 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[0]), .C(n24784), .X(io_oeb[11]) );
  sky130_fd_sc_hd__nor2_1 U27415 ( .A(j202_soc_core_pwrite[0]), .B(n24783), 
        .Y(n22973) );
  sky130_fd_sc_hd__nand3_1 U27416 ( .A(n22968), .B(n22973), .C(n22967), .Y(
        n22976) );
  sky130_fd_sc_hd__nor2_1 U27417 ( .A(n22976), .B(n22971), .Y(n23002) );
  sky130_fd_sc_hd__or3_1 U27418 ( .A(j202_soc_core_cmt_core_00_reg_addr[3]), 
        .B(j202_soc_core_cmt_core_00_reg_addr[2]), .C(n22972), .X(n23102) );
  sky130_fd_sc_hd__clkinv_1 U27419 ( .A(n22973), .Y(n22969) );
  sky130_fd_sc_hd__nor2_1 U27420 ( .A(n23102), .B(n22969), .Y(n23020) );
  sky130_fd_sc_hd__a22oi_1 U27421 ( .A1(j202_soc_core_cmt_core_00_cks0[0]), 
        .A2(n23002), .B1(n23020), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[0]), .Y(
        n22980) );
  sky130_fd_sc_hd__nand2_1 U27422 ( .A(j202_soc_core_cmt_core_00_reg_addr[3]), 
        .B(j202_soc_core_cmt_core_00_reg_addr[2]), .Y(n22970) );
  sky130_fd_sc_hd__nor2_1 U27423 ( .A(n22970), .B(n22976), .Y(n23022) );
  sky130_fd_sc_hd__a22oi_1 U27424 ( .A1(j202_soc_core_cmt_core_00_const1[0]), 
        .A2(n23021), .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[0]), .Y(
        n22979) );
  sky130_fd_sc_hd__nor3_1 U27425 ( .A(j202_soc_core_cmt_core_00_reg_addr[3]), 
        .B(j202_soc_core_cmt_core_00_reg_addr[2]), .C(n22976), .Y(n22981) );
  sky130_fd_sc_hd__nor2_1 U27426 ( .A(n22972), .B(n22971), .Y(n22974) );
  sky130_fd_sc_hd__nor2_1 U27427 ( .A(n22976), .B(n22975), .Y(n23001) );
  sky130_fd_sc_hd__a22o_1 U27428 ( .A1(j202_soc_core_cmt_core_00_const0[0]), 
        .A2(n23023), .B1(j202_soc_core_cmt_core_00_cks1[0]), .B2(n23001), .X(
        n22977) );
  sky130_fd_sc_hd__a21oi_1 U27429 ( .A1(j202_soc_core_cmt_core_00_str0), .A2(
        n22981), .B1(n22977), .Y(n22978) );
  sky130_fd_sc_hd__nand3_1 U27430 ( .A(n22980), .B(n22979), .C(n22978), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[0]) );
  sky130_fd_sc_hd__a22oi_1 U27431 ( .A1(j202_soc_core_cmt_core_00_const0[1]), 
        .A2(n23023), .B1(n23020), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[1]), .Y(
        n22985) );
  sky130_fd_sc_hd__a22oi_1 U27432 ( .A1(j202_soc_core_cmt_core_00_cks1[1]), 
        .A2(n23001), .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[1]), .Y(
        n22984) );
  sky130_fd_sc_hd__a22oi_1 U27433 ( .A1(j202_soc_core_cmt_core_00_cks0[1]), 
        .A2(n23002), .B1(j202_soc_core_cmt_core_00_str1), .B2(n22981), .Y(
        n22983) );
  sky130_fd_sc_hd__nand2_1 U27434 ( .A(j202_soc_core_cmt_core_00_const1[1]), 
        .B(n23021), .Y(n22982) );
  sky130_fd_sc_hd__nand4_1 U27435 ( .A(n22985), .B(n22984), .C(n22983), .D(
        n22982), .Y(j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[1]) );
  sky130_fd_sc_hd__a22oi_1 U27436 ( .A1(j202_soc_core_cmt_core_00_const1[2]), 
        .A2(n23021), .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[2]), .Y(
        n22988) );
  sky130_fd_sc_hd__a22oi_1 U27437 ( .A1(n23002), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[2]), .B1(n23001), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[2]), .Y(n22987) );
  sky130_fd_sc_hd__a22oi_1 U27438 ( .A1(j202_soc_core_cmt_core_00_const0[2]), 
        .A2(n23023), .B1(n23020), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[2]), .Y(
        n22986) );
  sky130_fd_sc_hd__nand3_1 U27439 ( .A(n22988), .B(n22987), .C(n22986), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[2]) );
  sky130_fd_sc_hd__a22oi_1 U27440 ( .A1(j202_soc_core_cmt_core_00_const1[3]), 
        .A2(n23021), .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[3]), .Y(
        n22991) );
  sky130_fd_sc_hd__a22oi_1 U27441 ( .A1(j202_soc_core_cmt_core_00_const0[3]), 
        .A2(n23023), .B1(n23002), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[3]), .Y(n22990) );
  sky130_fd_sc_hd__a22oi_1 U27442 ( .A1(n23020), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[3]), 
        .B1(n23001), .B2(j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[3]), .Y(
        n22989) );
  sky130_fd_sc_hd__nand3_1 U27443 ( .A(n22991), .B(n22990), .C(n22989), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[3]) );
  sky130_fd_sc_hd__a22oi_1 U27444 ( .A1(n23020), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[4]), 
        .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[4]), .Y(
        n22994) );
  sky130_fd_sc_hd__a22oi_1 U27445 ( .A1(j202_soc_core_cmt_core_00_const0[4]), 
        .A2(n23023), .B1(n23001), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[4]), .Y(n22993) );
  sky130_fd_sc_hd__a22oi_1 U27446 ( .A1(j202_soc_core_cmt_core_00_const1[4]), 
        .A2(n23021), .B1(n23002), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[4]), .Y(n22992) );
  sky130_fd_sc_hd__nand3_1 U27447 ( .A(n22994), .B(n22993), .C(n22992), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[4]) );
  sky130_fd_sc_hd__a22oi_1 U27448 ( .A1(n23020), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[5]), 
        .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[5]), .Y(
        n22997) );
  sky130_fd_sc_hd__a22oi_1 U27449 ( .A1(j202_soc_core_cmt_core_00_const0[5]), 
        .A2(n23023), .B1(j202_soc_core_cmt_core_00_const1[5]), .B2(n23021), 
        .Y(n22996) );
  sky130_fd_sc_hd__a22oi_1 U27450 ( .A1(n23002), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[5]), .B1(n23001), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[5]), .Y(n22995) );
  sky130_fd_sc_hd__nand3_1 U27451 ( .A(n22997), .B(n22996), .C(n22995), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[5]) );
  sky130_fd_sc_hd__a22oi_1 U27452 ( .A1(n23002), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[6]), .B1(n23020), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[6]), .Y(
        n23000) );
  sky130_fd_sc_hd__a22oi_1 U27453 ( .A1(j202_soc_core_cmt_core_00_const0[6]), 
        .A2(n23023), .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[6]), .Y(
        n22999) );
  sky130_fd_sc_hd__a22oi_1 U27454 ( .A1(j202_soc_core_cmt_core_00_const1[6]), 
        .A2(n23021), .B1(n23001), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[6]), .Y(n22998) );
  sky130_fd_sc_hd__nand3_1 U27455 ( .A(n23000), .B(n22999), .C(n22998), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[6]) );
  sky130_fd_sc_hd__a22oi_1 U27456 ( .A1(j202_soc_core_cmt_core_00_const1[7]), 
        .A2(n23021), .B1(n23001), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_0_), .Y(
        n23005) );
  sky130_fd_sc_hd__a22oi_1 U27457 ( .A1(n23002), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_0_), .B1(
        n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[7]), .Y(
        n23004) );
  sky130_fd_sc_hd__a22oi_1 U27458 ( .A1(j202_soc_core_cmt_core_00_const0[7]), 
        .A2(n23023), .B1(n23020), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[7]), .Y(
        n23003) );
  sky130_fd_sc_hd__nand3_1 U27459 ( .A(n23005), .B(n23004), .C(n23003), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[7]) );
  sky130_fd_sc_hd__a22oi_1 U27460 ( .A1(j202_soc_core_cmt_core_00_const0[8]), 
        .A2(n23023), .B1(n23020), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[8]), .Y(
        n23007) );
  sky130_fd_sc_hd__a22oi_1 U27461 ( .A1(j202_soc_core_cmt_core_00_const1[8]), 
        .A2(n23021), .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[8]), .Y(
        n23006) );
  sky130_fd_sc_hd__nand2_1 U27462 ( .A(n23007), .B(n23006), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[8]) );
  sky130_fd_sc_hd__a22oi_1 U27463 ( .A1(n23020), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[9]), 
        .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[9]), .Y(
        n23009) );
  sky130_fd_sc_hd__a22oi_1 U27464 ( .A1(j202_soc_core_cmt_core_00_const0[9]), 
        .A2(n23023), .B1(j202_soc_core_cmt_core_00_const1[9]), .B2(n23021), 
        .Y(n23008) );
  sky130_fd_sc_hd__nand2_1 U27465 ( .A(n23009), .B(n23008), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[9]) );
  sky130_fd_sc_hd__a22oi_1 U27466 ( .A1(j202_soc_core_cmt_core_00_const1[10]), 
        .A2(n23021), .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[10]), 
        .Y(n23011) );
  sky130_fd_sc_hd__a22oi_1 U27467 ( .A1(j202_soc_core_cmt_core_00_const0[10]), 
        .A2(n23023), .B1(n23020), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[10]), 
        .Y(n23010) );
  sky130_fd_sc_hd__nand2_1 U27468 ( .A(n23011), .B(n23010), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[10]) );
  sky130_fd_sc_hd__a22oi_1 U27469 ( .A1(j202_soc_core_cmt_core_00_const1[11]), 
        .A2(n23021), .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[11]), 
        .Y(n23013) );
  sky130_fd_sc_hd__a22oi_1 U27470 ( .A1(j202_soc_core_cmt_core_00_const0[11]), 
        .A2(n23023), .B1(n23020), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[11]), 
        .Y(n23012) );
  sky130_fd_sc_hd__nand2_1 U27471 ( .A(n23013), .B(n23012), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[11]) );
  sky130_fd_sc_hd__a22oi_1 U27472 ( .A1(n23020), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[12]), 
        .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[12]), 
        .Y(n23015) );
  sky130_fd_sc_hd__a22oi_1 U27473 ( .A1(j202_soc_core_cmt_core_00_const0[12]), 
        .A2(n23023), .B1(j202_soc_core_cmt_core_00_const1[12]), .B2(n23021), 
        .Y(n23014) );
  sky130_fd_sc_hd__nand2_1 U27474 ( .A(n23015), .B(n23014), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[12]) );
  sky130_fd_sc_hd__a22oi_1 U27475 ( .A1(j202_soc_core_cmt_core_00_const1[13]), 
        .A2(n23021), .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[13]), 
        .Y(n23017) );
  sky130_fd_sc_hd__a22oi_1 U27476 ( .A1(j202_soc_core_cmt_core_00_const0[13]), 
        .A2(n23023), .B1(n23020), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[13]), 
        .Y(n23016) );
  sky130_fd_sc_hd__nand2_1 U27477 ( .A(n23017), .B(n23016), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[13]) );
  sky130_fd_sc_hd__a22oi_1 U27478 ( .A1(n23020), .A2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[14]), 
        .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[14]), 
        .Y(n23019) );
  sky130_fd_sc_hd__a22oi_1 U27479 ( .A1(j202_soc_core_cmt_core_00_const0[14]), 
        .A2(n23023), .B1(j202_soc_core_cmt_core_00_const1[14]), .B2(n23021), 
        .Y(n23018) );
  sky130_fd_sc_hd__nand2_1 U27480 ( .A(n23019), .B(n23018), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[14]) );
  sky130_fd_sc_hd__a22oi_1 U27481 ( .A1(j202_soc_core_cmt_core_00_const1[15]), 
        .A2(n23021), .B1(n23020), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt1_reg_latch_status[15]), 
        .Y(n23025) );
  sky130_fd_sc_hd__a22oi_1 U27482 ( .A1(j202_soc_core_cmt_core_00_const0[15]), 
        .A2(n23023), .B1(n23022), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcnt0_reg_latch_status[15]), 
        .Y(n23024) );
  sky130_fd_sc_hd__nand2_1 U27483 ( .A(n23025), .B(n23024), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_nxt_rdata[15]) );
  sky130_fd_sc_hd__nand2_1 U27484 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[0]), .B(
        j202_soc_core_cmt_core_00_str0), .Y(n23027) );
  sky130_fd_sc_hd__o21ai_1 U27485 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[0]), .A2(
        j202_soc_core_cmt_core_00_str0), .B1(n23027), .Y(n23026) );
  sky130_fd_sc_hd__clkinv_1 U27486 ( .A(n23076), .Y(n23050) );
  sky130_fd_sc_hd__nand2_1 U27487 ( .A(n23026), .B(n23050), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[0]) );
  sky130_fd_sc_hd__clkinv_1 U27488 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[1]), .Y(n23028) );
  sky130_fd_sc_hd__nor2_1 U27489 ( .A(n23028), .B(n23027), .Y(n23029) );
  sky130_fd_sc_hd__a211oi_1 U27490 ( .A1(n23028), .A2(n23027), .B1(n23029), 
        .C1(n23076), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[1])
         );
  sky130_fd_sc_hd__nand2_1 U27491 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[2]), .B(n23029), .Y(
        n23031) );
  sky130_fd_sc_hd__o21ai_1 U27492 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[2]), .A2(n23029), .B1(
        n23031), .Y(n23030) );
  sky130_fd_sc_hd__nor2_1 U27493 ( .A(n23076), .B(n23030), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[2]) );
  sky130_fd_sc_hd__clkinv_1 U27494 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[3]), .Y(n23032) );
  sky130_fd_sc_hd__nor2_1 U27495 ( .A(n23032), .B(n23031), .Y(n23033) );
  sky130_fd_sc_hd__a211oi_1 U27496 ( .A1(n23032), .A2(n23031), .B1(n23033), 
        .C1(n23076), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[3])
         );
  sky130_fd_sc_hd__nand2_1 U27497 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[4]), .B(n23033), .Y(
        n23035) );
  sky130_fd_sc_hd__nor2_1 U27499 ( .A(n23076), .B(n23034), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[4]) );
  sky130_fd_sc_hd__nor2_1 U27500 ( .A(n23036), .B(n23035), .Y(n23037) );
  sky130_fd_sc_hd__a211oi_1 U27501 ( .A1(n23036), .A2(n23035), .B1(n23037), 
        .C1(n23076), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[5])
         );
  sky130_fd_sc_hd__nand2_1 U27502 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[6]), .B(n23037), .Y(
        n23039) );
  sky130_fd_sc_hd__o21ai_1 U27503 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[6]), .A2(n23037), .B1(
        n23039), .Y(n23038) );
  sky130_fd_sc_hd__nor2_1 U27504 ( .A(n23076), .B(n23038), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[6]) );
  sky130_fd_sc_hd__nor2_1 U27505 ( .A(n23040), .B(n23039), .Y(n23041) );
  sky130_fd_sc_hd__a211oi_1 U27506 ( .A1(n23040), .A2(n23039), .B1(n23041), 
        .C1(n23076), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[7])
         );
  sky130_fd_sc_hd__nand2_1 U27507 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[8]), .B(n23041), .Y(
        n23044) );
  sky130_fd_sc_hd__o21ai_1 U27508 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[8]), .A2(n23041), .B1(
        n23044), .Y(n23042) );
  sky130_fd_sc_hd__nor2_1 U27509 ( .A(n23076), .B(n23042), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[8]) );
  sky130_fd_sc_hd__o21ai_1 U27510 ( .A1(n23045), .A2(n23044), .B1(n23050), .Y(
        n23043) );
  sky130_fd_sc_hd__a21oi_1 U27511 ( .A1(n23045), .A2(n23044), .B1(n23043), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt0[9]) );
  sky130_fd_sc_hd__clkinv_1 U27512 ( .A(n23046), .Y(n23070) );
  sky130_fd_sc_hd__clkinv_1 U27513 ( .A(j202_soc_core_cmt_core_00_cnt0[0]), 
        .Y(n23048) );
  sky130_fd_sc_hd__clkinv_1 U27514 ( .A(n23086), .Y(n23088) );
  sky130_fd_sc_hd__o221ai_1 U27516 ( .A1(j202_soc_core_cmt_core_00_cnt0[0]), 
        .A2(n23070), .B1(n23048), .B2(n23076), .C1(n23047), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[0]) );
  sky130_fd_sc_hd__nor2_1 U27517 ( .A(n23050), .B(n23049), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt0_to1) );
  sky130_fd_sc_hd__a22oi_1 U27519 ( .A1(n23074), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[1]), .B1(
        j202_soc_core_cmt_core_00_cnt0[1]), .B2(n23050), .Y(n23051) );
  sky130_fd_sc_hd__a211oi_1 U27521 ( .A1(n23057), .A2(n23054), .B1(n23053), 
        .C1(n23070), .Y(n23055) );
  sky130_fd_sc_hd__a21oi_1 U27522 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[2]), .A2(n23074), .B1(n23055), 
        .Y(n23056) );
  sky130_fd_sc_hd__o21ai_1 U27523 ( .A1(n23057), .A2(n23076), .B1(n23056), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[2]) );
  sky130_fd_sc_hd__a21oi_1 U27524 ( .A1(j202_soc_core_cmt_core_00_cnt0[4]), 
        .A2(n23086), .B1(n23058), .Y(n23059) );
  sky130_fd_sc_hd__o22ai_1 U27525 ( .A1(n23060), .A2(n23059), .B1(n23101), 
        .B2(n25207), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[4])
         );
  sky130_fd_sc_hd__nand2_1 U27526 ( .A(j202_soc_core_cmt_core_00_cnt0[5]), .B(
        n23060), .Y(n23062) );
  sky130_fd_sc_hd__clkinv_1 U27527 ( .A(n23062), .Y(n23064) );
  sky130_fd_sc_hd__a21oi_1 U27528 ( .A1(j202_soc_core_cmt_core_00_cnt0[5]), 
        .A2(n23086), .B1(n23060), .Y(n23061) );
  sky130_fd_sc_hd__o22ai_1 U27529 ( .A1(n23064), .A2(n23061), .B1(n23101), 
        .B2(n25210), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[5])
         );
  sky130_fd_sc_hd__clkinv_1 U27530 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[6]), .Y(n25215) );
  sky130_fd_sc_hd__nor2_1 U27531 ( .A(n23063), .B(n23062), .Y(n23068) );
  sky130_fd_sc_hd__nor2_1 U27532 ( .A(n23088), .B(n23068), .Y(n23066) );
  sky130_fd_sc_hd__o22ai_1 U27535 ( .A1(j202_soc_core_cmt_core_00_cnt0[7]), 
        .A2(n23068), .B1(n23067), .B2(n23066), .Y(n23069) );
  sky130_fd_sc_hd__o21ai_1 U27536 ( .A1(n23101), .A2(n25217), .B1(n23069), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[7]) );
  sky130_fd_sc_hd__a211oi_1 U27537 ( .A1(n23077), .A2(n23072), .B1(n23071), 
        .C1(n23070), .Y(n23073) );
  sky130_fd_sc_hd__a21oi_1 U27538 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[8]), .A2(n23074), .B1(n23073), 
        .Y(n23075) );
  sky130_fd_sc_hd__o21ai_1 U27539 ( .A1(n23077), .A2(n23076), .B1(n23075), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[8]) );
  sky130_fd_sc_hd__a21o_1 U27540 ( .A1(n23079), .A2(n23078), .B1(n23088), .X(
        n23080) );
  sky130_fd_sc_hd__o22ai_1 U27541 ( .A1(n23081), .A2(n23080), .B1(n23101), 
        .B2(n25150), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[9])
         );
  sky130_fd_sc_hd__a21oi_1 U27542 ( .A1(j202_soc_core_cmt_core_00_cnt0[10]), 
        .A2(n23086), .B1(n23081), .Y(n23082) );
  sky130_fd_sc_hd__o22ai_1 U27543 ( .A1(n23083), .A2(n23082), .B1(n23101), 
        .B2(n25225), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[10])
         );
  sky130_fd_sc_hd__nor2b_1 U27544 ( .B_N(n23085), .A(n23084), .Y(n23089) );
  sky130_fd_sc_hd__a21oi_1 U27545 ( .A1(j202_soc_core_cmt_core_00_cnt0[12]), 
        .A2(n23086), .B1(n23085), .Y(n23087) );
  sky130_fd_sc_hd__o22ai_1 U27546 ( .A1(n23089), .A2(n23087), .B1(n23101), 
        .B2(n23200), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[12])
         );
  sky130_fd_sc_hd__nand2_1 U27547 ( .A(j202_soc_core_cmt_core_00_cnt0[13]), 
        .B(n23089), .Y(n23096) );
  sky130_fd_sc_hd__clkinv_1 U27548 ( .A(n23096), .Y(n23092) );
  sky130_fd_sc_hd__nor2_1 U27549 ( .A(n23092), .B(n23088), .Y(n23098) );
  sky130_fd_sc_hd__o21ai_1 U27551 ( .A1(n23091), .A2(n23101), .B1(n23090), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[13]) );
  sky130_fd_sc_hd__o22ai_1 U27552 ( .A1(j202_soc_core_cmt_core_00_cnt0[14]), 
        .A2(n23092), .B1(n23095), .B2(n23098), .Y(n23093) );
  sky130_fd_sc_hd__o21ai_1 U27553 ( .A1(n23101), .A2(n23094), .B1(n23093), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[14]) );
  sky130_fd_sc_hd__nor2_1 U27554 ( .A(n23096), .B(n23095), .Y(n23099) );
  sky130_fd_sc_hd__a21oi_1 U27555 ( .A1(j202_soc_core_cmt_core_00_cnt0[14]), 
        .A2(j202_soc_core_cmt_core_00_cnt0[15]), .B1(n23096), .Y(n23097) );
  sky130_fd_sc_hd__o22ai_1 U27556 ( .A1(n23099), .A2(
        j202_soc_core_cmt_core_00_cnt0[15]), .B1(n23098), .B2(n23097), .Y(
        n23100) );
  sky130_fd_sc_hd__nand2_1 U27558 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[0]), .B(
        j202_soc_core_cmt_core_00_str1), .Y(n23112) );
  sky130_fd_sc_hd__nor2_1 U27560 ( .A(n23103), .B(n23102), .Y(n23209) );
  sky130_fd_sc_hd__clkinv_1 U27561 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[7]), .Y(n23125) );
  sky130_fd_sc_hd__clkinv_1 U27562 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[3]), .Y(n23117) );
  sky130_fd_sc_hd__o32ai_1 U27563 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[3]), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[5]), .A3(
        j202_soc_core_cmt_core_00_cks1[1]), .B1(n23125), .B2(n23117), .Y(
        n23110) );
  sky130_fd_sc_hd__nor4_1 U27564 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[8]), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[2]), .C(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[0]), .D(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[1]), .Y(n23108) );
  sky130_fd_sc_hd__clkinv_1 U27565 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[9]), .Y(n23130) );
  sky130_fd_sc_hd__clkinv_1 U27566 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[5]), .Y(n23121) );
  sky130_fd_sc_hd__a21oi_1 U27567 ( .A1(n23121), .A2(n23130), .B1(
        j202_soc_core_cmt_core_00_cks1[0]), .Y(n23104) );
  sky130_fd_sc_hd__a31oi_1 U27568 ( .A1(j202_soc_core_cmt_core_00_cks1[1]), 
        .A2(n23130), .A3(n23125), .B1(n23104), .Y(n23107) );
  sky130_fd_sc_hd__nor2_1 U27569 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[4]), .B(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[6]), .Y(n23106) );
  sky130_fd_sc_hd__nand4_1 U27571 ( .A(n23108), .B(n23107), .C(n23106), .D(
        n23105), .Y(n23109) );
  sky130_fd_sc_hd__a211oi_1 U27572 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[5]), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[9]), .B1(n23110), .C1(
        n23109), .Y(n23152) );
  sky130_fd_sc_hd__nor2_1 U27573 ( .A(n23209), .B(n23152), .Y(n23198) );
  sky130_fd_sc_hd__nand2_1 U27574 ( .A(n23111), .B(n23198), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[0]) );
  sky130_fd_sc_hd__clkinv_1 U27575 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[1]), .Y(n23113) );
  sky130_fd_sc_hd__nor2_1 U27576 ( .A(n23113), .B(n23112), .Y(n23114) );
  sky130_fd_sc_hd__a211oi_1 U27577 ( .A1(n23113), .A2(n23112), .B1(n23114), 
        .C1(n23196), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[1])
         );
  sky130_fd_sc_hd__nand2_1 U27578 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[2]), .B(n23114), .Y(
        n23116) );
  sky130_fd_sc_hd__o21ai_1 U27579 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[2]), .A2(n23114), .B1(
        n23116), .Y(n23115) );
  sky130_fd_sc_hd__nor2_1 U27580 ( .A(n23196), .B(n23115), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[2]) );
  sky130_fd_sc_hd__nor2_1 U27581 ( .A(n23117), .B(n23116), .Y(n23118) );
  sky130_fd_sc_hd__a211oi_1 U27582 ( .A1(n23117), .A2(n23116), .B1(n23118), 
        .C1(n23196), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[3])
         );
  sky130_fd_sc_hd__nand2_1 U27583 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[4]), .B(n23118), .Y(
        n23120) );
  sky130_fd_sc_hd__o21ai_1 U27584 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[4]), .A2(n23118), .B1(
        n23120), .Y(n23119) );
  sky130_fd_sc_hd__nor2_1 U27585 ( .A(n23196), .B(n23119), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[4]) );
  sky130_fd_sc_hd__nor2_1 U27586 ( .A(n23121), .B(n23120), .Y(n23122) );
  sky130_fd_sc_hd__a211oi_1 U27587 ( .A1(n23121), .A2(n23120), .B1(n23122), 
        .C1(n23196), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[5])
         );
  sky130_fd_sc_hd__nand2_1 U27588 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[6]), .B(n23122), .Y(
        n23124) );
  sky130_fd_sc_hd__o21ai_1 U27589 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[6]), .A2(n23122), .B1(
        n23124), .Y(n23123) );
  sky130_fd_sc_hd__nor2_1 U27590 ( .A(n23196), .B(n23123), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[6]) );
  sky130_fd_sc_hd__nor2_1 U27591 ( .A(n23125), .B(n23124), .Y(n23126) );
  sky130_fd_sc_hd__a211oi_1 U27592 ( .A1(n23125), .A2(n23124), .B1(n23126), 
        .C1(n23196), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[7])
         );
  sky130_fd_sc_hd__nand2_1 U27593 ( .A(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[8]), .B(n23126), .Y(
        n23129) );
  sky130_fd_sc_hd__o21ai_1 U27594 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[8]), .A2(n23126), .B1(
        n23129), .Y(n23127) );
  sky130_fd_sc_hd__nor2_1 U27595 ( .A(n23196), .B(n23127), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[8]) );
  sky130_fd_sc_hd__o21ai_1 U27596 ( .A1(n23130), .A2(n23129), .B1(n23198), .Y(
        n23128) );
  sky130_fd_sc_hd__a21oi_1 U27597 ( .A1(n23130), .A2(n23129), .B1(n23128), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_clkcnt1[9]) );
  sky130_fd_sc_hd__clkinv_1 U27598 ( .A(j202_soc_core_cmt_core_00_const1[8]), 
        .Y(n25224) );
  sky130_fd_sc_hd__clkinv_1 U27599 ( .A(j202_soc_core_cmt_core_00_const1[1]), 
        .Y(n25155) );
  sky130_fd_sc_hd__o22ai_1 U27600 ( .A1(n25224), .A2(
        j202_soc_core_cmt_core_00_cnt1[8]), .B1(n25155), .B2(
        j202_soc_core_cmt_core_00_cnt1[1]), .Y(n23131) );
  sky130_fd_sc_hd__a221oi_1 U27601 ( .A1(n25224), .A2(
        j202_soc_core_cmt_core_00_cnt1[8]), .B1(
        j202_soc_core_cmt_core_00_cnt1[1]), .B2(n25155), .C1(n23131), .Y(
        n23139) );
  sky130_fd_sc_hd__clkinv_1 U27602 ( .A(j202_soc_core_cmt_core_00_const1[6]), 
        .Y(n25216) );
  sky130_fd_sc_hd__clkinv_1 U27603 ( .A(j202_soc_core_cmt_core_00_const1[0]), 
        .Y(n25199) );
  sky130_fd_sc_hd__o22ai_1 U27604 ( .A1(n25216), .A2(
        j202_soc_core_cmt_core_00_cnt1[6]), .B1(n25199), .B2(
        j202_soc_core_cmt_core_00_cnt1[0]), .Y(n23132) );
  sky130_fd_sc_hd__a221oi_1 U27605 ( .A1(n25216), .A2(
        j202_soc_core_cmt_core_00_cnt1[6]), .B1(
        j202_soc_core_cmt_core_00_cnt1[0]), .B2(n25199), .C1(n23132), .Y(
        n23138) );
  sky130_fd_sc_hd__clkinv_1 U27606 ( .A(j202_soc_core_cmt_core_00_const1[7]), 
        .Y(n25218) );
  sky130_fd_sc_hd__clkinv_1 U27607 ( .A(j202_soc_core_cmt_core_00_const1[9]), 
        .Y(n25151) );
  sky130_fd_sc_hd__o22ai_1 U27608 ( .A1(n25218), .A2(
        j202_soc_core_cmt_core_00_cnt1[7]), .B1(n25151), .B2(
        j202_soc_core_cmt_core_00_cnt1[9]), .Y(n23133) );
  sky130_fd_sc_hd__a221oi_1 U27609 ( .A1(n25218), .A2(
        j202_soc_core_cmt_core_00_cnt1[7]), .B1(
        j202_soc_core_cmt_core_00_cnt1[9]), .B2(n25151), .C1(n23133), .Y(
        n23137) );
  sky130_fd_sc_hd__clkinv_1 U27610 ( .A(j202_soc_core_cmt_core_00_cnt1[14]), 
        .Y(n23211) );
  sky130_fd_sc_hd__clkinv_1 U27611 ( .A(j202_soc_core_cmt_core_00_cnt1[4]), 
        .Y(n23135) );
  sky130_fd_sc_hd__o22ai_1 U27612 ( .A1(n23211), .A2(
        j202_soc_core_cmt_core_00_const1[14]), .B1(n23135), .B2(
        j202_soc_core_cmt_core_00_const1[4]), .Y(n23134) );
  sky130_fd_sc_hd__a221oi_1 U27613 ( .A1(n23211), .A2(
        j202_soc_core_cmt_core_00_const1[14]), .B1(
        j202_soc_core_cmt_core_00_const1[4]), .B2(n23135), .C1(n23134), .Y(
        n23136) );
  sky130_fd_sc_hd__nand4_1 U27614 ( .A(n23139), .B(n23138), .C(n23137), .D(
        n23136), .Y(n23151) );
  sky130_fd_sc_hd__clkinv_1 U27615 ( .A(j202_soc_core_cmt_core_00_const1[2]), 
        .Y(n25196) );
  sky130_fd_sc_hd__clkinv_1 U27616 ( .A(j202_soc_core_cmt_core_00_const1[3]), 
        .Y(n25221) );
  sky130_fd_sc_hd__o22ai_1 U27617 ( .A1(n25196), .A2(
        j202_soc_core_cmt_core_00_cnt1[2]), .B1(n25221), .B2(
        j202_soc_core_cmt_core_00_cnt1[3]), .Y(n23140) );
  sky130_fd_sc_hd__a221oi_1 U27618 ( .A1(n25196), .A2(
        j202_soc_core_cmt_core_00_cnt1[2]), .B1(
        j202_soc_core_cmt_core_00_cnt1[3]), .B2(n25221), .C1(n23140), .Y(
        n23149) );
  sky130_fd_sc_hd__clkinv_1 U27619 ( .A(j202_soc_core_cmt_core_00_cnt1[12]), 
        .Y(n23142) );
  sky130_fd_sc_hd__clkinv_1 U27620 ( .A(j202_soc_core_cmt_core_00_cnt1[11]), 
        .Y(n23197) );
  sky130_fd_sc_hd__o22ai_1 U27621 ( .A1(n23142), .A2(
        j202_soc_core_cmt_core_00_const1[12]), .B1(n23197), .B2(
        j202_soc_core_cmt_core_00_const1[11]), .Y(n23141) );
  sky130_fd_sc_hd__a221oi_1 U27622 ( .A1(n23142), .A2(
        j202_soc_core_cmt_core_00_const1[12]), .B1(
        j202_soc_core_cmt_core_00_const1[11]), .B2(n23197), .C1(n23141), .Y(
        n23148) );
  sky130_fd_sc_hd__clkinv_1 U27623 ( .A(j202_soc_core_cmt_core_00_cnt1[15]), 
        .Y(n23144) );
  sky130_fd_sc_hd__clkinv_1 U27624 ( .A(j202_soc_core_cmt_core_00_const1[5]), 
        .Y(n25211) );
  sky130_fd_sc_hd__o22ai_1 U27625 ( .A1(n23144), .A2(
        j202_soc_core_cmt_core_00_const1[15]), .B1(n25211), .B2(
        j202_soc_core_cmt_core_00_cnt1[5]), .Y(n23143) );
  sky130_fd_sc_hd__a221oi_1 U27626 ( .A1(n23144), .A2(
        j202_soc_core_cmt_core_00_const1[15]), .B1(
        j202_soc_core_cmt_core_00_cnt1[5]), .B2(n25211), .C1(n23143), .Y(
        n23147) );
  sky130_fd_sc_hd__clkinv_1 U27627 ( .A(j202_soc_core_cmt_core_00_cnt1[13]), 
        .Y(n23205) );
  sky130_fd_sc_hd__clkinv_1 U27628 ( .A(j202_soc_core_cmt_core_00_const1[10]), 
        .Y(n25226) );
  sky130_fd_sc_hd__o22ai_1 U27629 ( .A1(n23205), .A2(
        j202_soc_core_cmt_core_00_const1[13]), .B1(n25226), .B2(
        j202_soc_core_cmt_core_00_cnt1[10]), .Y(n23145) );
  sky130_fd_sc_hd__a221oi_1 U27630 ( .A1(n23205), .A2(
        j202_soc_core_cmt_core_00_const1[13]), .B1(
        j202_soc_core_cmt_core_00_cnt1[10]), .B2(n25226), .C1(n23145), .Y(
        n23146) );
  sky130_fd_sc_hd__nand4_1 U27631 ( .A(n23149), .B(n23148), .C(n23147), .D(
        n23146), .Y(n23150) );
  sky130_fd_sc_hd__nor2_1 U27632 ( .A(n23151), .B(n23150), .Y(n23157) );
  sky130_fd_sc_hd__clkinv_1 U27633 ( .A(n23157), .Y(n23155) );
  sky130_fd_sc_hd__nand2_1 U27634 ( .A(n23152), .B(n23217), .Y(n23156) );
  sky130_fd_sc_hd__a21oi_1 U27635 ( .A1(n23155), .A2(
        j202_soc_core_cmt_core_00_cnt1[0]), .B1(n23156), .Y(n23153) );
  sky130_fd_sc_hd__a21oi_1 U27636 ( .A1(j202_soc_core_cmt_core_00_cnt1[0]), 
        .A2(n23198), .B1(n23153), .Y(n23154) );
  sky130_fd_sc_hd__nor2_1 U27638 ( .A(n23198), .B(n23155), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_set_cmpcnt1_to1) );
  sky130_fd_sc_hd__nor2_1 U27639 ( .A(n23157), .B(n23156), .Y(n23202) );
  sky130_fd_sc_hd__nand2_1 U27640 ( .A(j202_soc_core_cmt_core_00_cnt1[0]), .B(
        j202_soc_core_cmt_core_00_cnt1[1]), .Y(n23158) );
  sky130_fd_sc_hd__a22oi_1 U27642 ( .A1(j202_soc_core_cmt_core_00_cnt1[1]), 
        .A2(n23198), .B1(n23209), .B2(j202_soc_core_cmt_core_00_wdata_cnt0[1]), 
        .Y(n23159) );
  sky130_fd_sc_hd__nand3_1 U27644 ( .A(j202_soc_core_cmt_core_00_cnt1[2]), .B(
        j202_soc_core_cmt_core_00_cnt1[0]), .C(
        j202_soc_core_cmt_core_00_cnt1[1]), .Y(n23165) );
  sky130_fd_sc_hd__a21oi_1 U27645 ( .A1(n23202), .A2(n23165), .B1(n23198), .Y(
        n23164) );
  sky130_fd_sc_hd__a31oi_1 U27646 ( .A1(j202_soc_core_cmt_core_00_cnt1[0]), 
        .A2(j202_soc_core_cmt_core_00_cnt1[1]), .A3(n23202), .B1(
        j202_soc_core_cmt_core_00_cnt1[2]), .Y(n23161) );
  sky130_fd_sc_hd__o22ai_1 U27647 ( .A1(n23164), .A2(n23161), .B1(n23217), 
        .B2(n25195), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[2])
         );
  sky130_fd_sc_hd__clkinv_1 U27648 ( .A(j202_soc_core_cmt_core_00_cnt1[3]), 
        .Y(n23166) );
  sky130_fd_sc_hd__nor3_1 U27649 ( .A(j202_soc_core_cmt_core_00_cnt1[3]), .B(
        n23192), .C(n23165), .Y(n23162) );
  sky130_fd_sc_hd__a21oi_1 U27650 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[3]), .A2(n23209), .B1(n23162), 
        .Y(n23163) );
  sky130_fd_sc_hd__o21ai_1 U27651 ( .A1(n23164), .A2(n23166), .B1(n23163), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[3]) );
  sky130_fd_sc_hd__nor2_1 U27652 ( .A(n23166), .B(n23165), .Y(n23167) );
  sky130_fd_sc_hd__nand2_1 U27653 ( .A(j202_soc_core_cmt_core_00_cnt1[4]), .B(
        n23167), .Y(n23170) );
  sky130_fd_sc_hd__o21ai_1 U27654 ( .A1(j202_soc_core_cmt_core_00_cnt1[4]), 
        .A2(n23167), .B1(n23170), .Y(n23169) );
  sky130_fd_sc_hd__a22oi_1 U27655 ( .A1(j202_soc_core_cmt_core_00_cnt1[4]), 
        .A2(n23198), .B1(n23209), .B2(j202_soc_core_cmt_core_00_wdata_cnt0[4]), 
        .Y(n23168) );
  sky130_fd_sc_hd__o21ai_1 U27656 ( .A1(n23192), .A2(n23169), .B1(n23168), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[4]) );
  sky130_fd_sc_hd__clkinv_1 U27657 ( .A(j202_soc_core_cmt_core_00_cnt1[5]), 
        .Y(n23173) );
  sky130_fd_sc_hd__nor2_1 U27658 ( .A(n23173), .B(n23170), .Y(n23174) );
  sky130_fd_sc_hd__a211oi_1 U27659 ( .A1(n23173), .A2(n23170), .B1(n23174), 
        .C1(n23192), .Y(n23171) );
  sky130_fd_sc_hd__a21oi_1 U27660 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[5]), .A2(n23209), .B1(n23171), 
        .Y(n23172) );
  sky130_fd_sc_hd__o21ai_1 U27661 ( .A1(n23173), .A2(n23196), .B1(n23172), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[5]) );
  sky130_fd_sc_hd__nand2_1 U27662 ( .A(j202_soc_core_cmt_core_00_cnt1[6]), .B(
        n23174), .Y(n23179) );
  sky130_fd_sc_hd__o21ai_1 U27663 ( .A1(j202_soc_core_cmt_core_00_cnt1[6]), 
        .A2(n23174), .B1(n23179), .Y(n23176) );
  sky130_fd_sc_hd__a22oi_1 U27664 ( .A1(j202_soc_core_cmt_core_00_cnt1[6]), 
        .A2(n23198), .B1(n23209), .B2(j202_soc_core_cmt_core_00_wdata_cnt0[6]), 
        .Y(n23175) );
  sky130_fd_sc_hd__nor2_1 U27666 ( .A(n23192), .B(n23179), .Y(n23177) );
  sky130_fd_sc_hd__clkinv_1 U27667 ( .A(j202_soc_core_cmt_core_00_cnt1[7]), 
        .Y(n23180) );
  sky130_fd_sc_hd__nor2_1 U27668 ( .A(n23180), .B(n23179), .Y(n23184) );
  sky130_fd_sc_hd__o21ai_1 U27669 ( .A1(n23184), .A2(n23192), .B1(n23196), .Y(
        n23181) );
  sky130_fd_sc_hd__o21ai_1 U27671 ( .A1(n25217), .A2(n23217), .B1(n23178), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[7]) );
  sky130_fd_sc_hd__clkinv_1 U27672 ( .A(
        j202_soc_core_cmt_core_00_wdata_cnt0[8]), .Y(n25223) );
  sky130_fd_sc_hd__nor3_1 U27673 ( .A(n23180), .B(n23192), .C(n23179), .Y(
        n23185) );
  sky130_fd_sc_hd__clkinv_1 U27674 ( .A(j202_soc_core_cmt_core_00_cnt1[8]), 
        .Y(n23182) );
  sky130_fd_sc_hd__o22ai_1 U27675 ( .A1(j202_soc_core_cmt_core_00_cnt1[8]), 
        .A2(n23185), .B1(n23182), .B2(n23181), .Y(n23183) );
  sky130_fd_sc_hd__o21ai_1 U27676 ( .A1(n23217), .A2(n25223), .B1(n23183), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[8]) );
  sky130_fd_sc_hd__nand3_1 U27677 ( .A(j202_soc_core_cmt_core_00_cnt1[8]), .B(
        j202_soc_core_cmt_core_00_cnt1[9]), .C(n23184), .Y(n23191) );
  sky130_fd_sc_hd__a21oi_1 U27678 ( .A1(n23202), .A2(n23191), .B1(n23198), .Y(
        n23190) );
  sky130_fd_sc_hd__a21oi_1 U27679 ( .A1(j202_soc_core_cmt_core_00_cnt1[8]), 
        .A2(n23185), .B1(j202_soc_core_cmt_core_00_cnt1[9]), .Y(n23186) );
  sky130_fd_sc_hd__o22ai_1 U27680 ( .A1(n23190), .A2(n23186), .B1(n23217), 
        .B2(n25150), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[9])
         );
  sky130_fd_sc_hd__clkinv_1 U27681 ( .A(j202_soc_core_cmt_core_00_cnt1[10]), 
        .Y(n23189) );
  sky130_fd_sc_hd__nor3_1 U27682 ( .A(j202_soc_core_cmt_core_00_cnt1[10]), .B(
        n23192), .C(n23191), .Y(n23187) );
  sky130_fd_sc_hd__a21oi_1 U27683 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[10]), .A2(n23209), .B1(n23187), 
        .Y(n23188) );
  sky130_fd_sc_hd__o21ai_1 U27684 ( .A1(n23190), .A2(n23189), .B1(n23188), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[10]) );
  sky130_fd_sc_hd__nand2b_1 U27685 ( .A_N(n23191), .B(
        j202_soc_core_cmt_core_00_cnt1[10]), .Y(n23193) );
  sky130_fd_sc_hd__nor2_1 U27686 ( .A(n23197), .B(n23193), .Y(n23199) );
  sky130_fd_sc_hd__a211oi_1 U27687 ( .A1(n23197), .A2(n23193), .B1(n23199), 
        .C1(n23192), .Y(n23194) );
  sky130_fd_sc_hd__a21oi_1 U27688 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[11]), .A2(n23209), .B1(n23194), 
        .Y(n23195) );
  sky130_fd_sc_hd__nand2_1 U27690 ( .A(j202_soc_core_cmt_core_00_cnt1[12]), 
        .B(n23199), .Y(n23203) );
  sky130_fd_sc_hd__a21oi_1 U27691 ( .A1(n23202), .A2(n23203), .B1(n23198), .Y(
        n23208) );
  sky130_fd_sc_hd__nor2_1 U27692 ( .A(j202_soc_core_cmt_core_00_cnt1[12]), .B(
        n23206), .Y(n23201) );
  sky130_fd_sc_hd__o22ai_1 U27693 ( .A1(n23208), .A2(n23201), .B1(n23217), 
        .B2(n23200), .Y(j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[12])
         );
  sky130_fd_sc_hd__nand2_1 U27694 ( .A(n23202), .B(n23205), .Y(n23207) );
  sky130_fd_sc_hd__a2bb2oi_1 U27695 ( .B1(
        j202_soc_core_cmt_core_00_wdata_cnt0[13]), .B2(n23209), .A1_N(n23207), 
        .A2_N(n23203), .Y(n23204) );
  sky130_fd_sc_hd__nand3_1 U27697 ( .A(j202_soc_core_cmt_core_00_cnt1[12]), 
        .B(j202_soc_core_cmt_core_00_cnt1[13]), .C(n23206), .Y(n23212) );
  sky130_fd_sc_hd__nand2_1 U27698 ( .A(n23208), .B(n23207), .Y(n23214) );
  sky130_fd_sc_hd__a22oi_1 U27699 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[14]), .A2(n23209), .B1(
        j202_soc_core_cmt_core_00_cnt1[14]), .B2(n23214), .Y(n23210) );
  sky130_fd_sc_hd__o21ai_1 U27700 ( .A1(j202_soc_core_cmt_core_00_cnt1[14]), 
        .A2(n23212), .B1(n23210), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[14]) );
  sky130_fd_sc_hd__nor2_1 U27701 ( .A(n23212), .B(n23211), .Y(n23215) );
  sky130_fd_sc_hd__a21oi_1 U27702 ( .A1(j202_soc_core_cmt_core_00_cnt1[14]), 
        .A2(j202_soc_core_cmt_core_00_cnt1[15]), .B1(n23212), .Y(n23213) );
  sky130_fd_sc_hd__o22ai_1 U27703 ( .A1(n23215), .A2(
        j202_soc_core_cmt_core_00_cnt1[15]), .B1(n23214), .B2(n23213), .Y(
        n23216) );
  sky130_fd_sc_hd__nor2b_1 U27705 ( .B_N(j202_soc_core_uart_TOP_rx_sio_ce_r1), 
        .A(j202_soc_core_uart_TOP_rx_sio_ce_r2), .Y(
        j202_soc_core_uart_TOP_N118) );
  sky130_fd_sc_hd__nor2_1 U27706 ( .A(j202_soc_core_uart_TOP_shift_en), .B(
        j202_soc_core_uart_TOP_txf_empty_r), .Y(j202_soc_core_uart_TOP_N137)
         );
  sky130_fd_sc_hd__nand3_1 U27707 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[1]), 
        .B(n23219), .C(n23816), .Y(j202_soc_core_uart_TOP_N128) );
  sky130_fd_sc_hd__clkinv_1 U27708 ( .A(j202_soc_core_uart_TOP_tx_bit_cnt[2]), 
        .Y(n23824) );
  sky130_fd_sc_hd__nand4b_1 U27709 ( .A_N(j202_soc_core_uart_TOP_tx_bit_cnt[1]), .B(j202_soc_core_uart_TOP_tx_bit_cnt[0]), .C(
        j202_soc_core_uart_TOP_tx_bit_cnt[3]), .D(n23824), .Y(
        j202_soc_core_uart_TOP_N123) );
  sky130_fd_sc_hd__nor2b_1 U27710 ( .B_N(n25399), .A(
        j202_soc_core_uart_BRG_sio_ce_r), .Y(j202_soc_core_uart_BRG_N59) );
  sky130_fd_sc_hd__nor2_1 U27711 ( .A(n24882), .B(n23220), .Y(
        j202_soc_core_j22_cpu_id_idec_N900) );
  sky130_fd_sc_hd__nor2_1 U27713 ( .A(n23232), .B(n23227), .Y(n24880) );
  sky130_fd_sc_hd__o21ai_1 U27714 ( .A1(n23226), .A2(n23225), .B1(n24880), .Y(
        n23233) );
  sky130_fd_sc_hd__nor2_1 U27715 ( .A(n25734), .B(n23227), .Y(n23231) );
  sky130_fd_sc_hd__nand2_1 U27716 ( .A(n23228), .B(j202_soc_core_intr_vec__1_), 
        .Y(n23230) );
  sky130_fd_sc_hd__a21oi_1 U27717 ( .A1(n23232), .A2(n23230), .B1(n23229), .Y(
        n24864) );
  sky130_fd_sc_hd__nand2_1 U27719 ( .A(n23233), .B(n24889), .Y(
        j202_soc_core_j22_cpu_id_idec_N894) );
  sky130_fd_sc_hd__o31ai_1 U27720 ( .A1(n23239), .A2(n23237), .A3(n23236), 
        .B1(n23235), .Y(n24892) );
  sky130_fd_sc_hd__nor2_1 U27721 ( .A(n23238), .B(n24892), .Y(
        j202_soc_core_j22_cpu_id_idec_N960) );
  sky130_fd_sc_hd__and3_1 U27722 ( .A(n23239), .B(
        j202_soc_core_j22_cpu_id_idec_N960), .C(
        j202_soc_core_j22_cpu_regop_Wm__0_), .X(
        j202_soc_core_j22_cpu_id_idec_N956) );
  sky130_fd_sc_hd__and3_1 U27723 ( .A(n23239), .B(
        j202_soc_core_j22_cpu_id_idec_N960), .C(
        j202_soc_core_j22_cpu_regop_Wm__1_), .X(
        j202_soc_core_j22_cpu_id_idec_N957) );
  sky130_fd_sc_hd__and3_1 U27724 ( .A(n23239), .B(
        j202_soc_core_j22_cpu_id_idec_N960), .C(
        j202_soc_core_j22_cpu_regop_Wm__2_), .X(
        j202_soc_core_j22_cpu_id_idec_N958) );
  sky130_fd_sc_hd__and3_1 U27725 ( .A(n23239), .B(
        j202_soc_core_j22_cpu_id_idec_N960), .C(
        j202_soc_core_j22_cpu_regop_Wm__3_), .X(
        j202_soc_core_j22_cpu_id_idec_N959) );
  sky130_fd_sc_hd__nand2_1 U27727 ( .A(n25543), .B(n23241), .Y(n23244) );
  sky130_fd_sc_hd__nor2_1 U27728 ( .A(n23242), .B(n23244), .Y(
        j202_soc_core_j22_cpu_ma_N54) );
  sky130_fd_sc_hd__nor2_1 U27729 ( .A(n23243), .B(n23244), .Y(
        j202_soc_core_j22_cpu_ma_N55) );
  sky130_fd_sc_hd__nor2_1 U27730 ( .A(n23245), .B(n23244), .Y(
        j202_soc_core_j22_cpu_ma_N56) );
  sky130_fd_sc_hd__o21ai_1 U27731 ( .A1(n23248), .A2(n23247), .B1(n23246), .Y(
        j202_soc_core_j22_cpu_ml_N195) );
  sky130_fd_sc_hd__nor3_1 U27732 ( .A(n24894), .B(n23250), .C(n23249), .Y(
        j202_soc_core_j22_cpu_N8) );
  sky130_fd_sc_hd__clkinv_1 U27733 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[0]), .Y(n24938) );
  sky130_fd_sc_hd__nor2_1 U27734 ( .A(n23251), .B(n24938), .Y(
        j202_soc_core_wbqspiflash_00_N628) );
  sky130_fd_sc_hd__clkinv_1 U27735 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[1]), .Y(n23793) );
  sky130_fd_sc_hd__nor2_1 U27736 ( .A(n23251), .B(n23793), .Y(
        j202_soc_core_wbqspiflash_00_N629) );
  sky130_fd_sc_hd__nand2b_1 U27738 ( .A_N(j202_soc_core_cmt_core_00_cmf0), .B(
        n23252), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_nxt_latch_status_0_) );
  sky130_fd_sc_hd__nand2b_1 U27740 ( .A_N(j202_soc_core_cmt_core_00_cmf1), .B(
        n23253), .Y(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_nxt_latch_status_0_) );
  sky130_fd_sc_hd__xnor2_1 U27741 ( .A(j202_soc_core_uart_TOP_rxd_s), .B(
        j202_soc_core_uart_TOP_rxd_r), .Y(n23814) );
  sky130_fd_sc_hd__nor2_1 U27742 ( .A(j202_soc_core_rst), .B(n23814), .Y(
        j202_soc_core_uart_TOP_N102) );
  sky130_fd_sc_hd__clkinv_1 U27743 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[0]), 
        .Y(n23811) );
  sky130_fd_sc_hd__nor2_1 U27744 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[0]), 
        .B(n23811), .Y(n23257) );
  sky130_fd_sc_hd__o211ai_1 U27745 ( .A1(n23257), .A2(n23256), .B1(n25201), 
        .C1(n23255), .Y(n23258) );
  sky130_fd_sc_hd__nand3_1 U27746 ( .A(n25734), .B(n25122), .C(n23258), .Y(
        j202_soc_core_uart_TOP_tx_fifo_N41) );
  sky130_fd_sc_hd__nor2_1 U27747 ( .A(j202_soc_core_rst), .B(n23258), .Y(
        j202_soc_core_uart_TOP_tx_fifo_N42) );
  sky130_fd_sc_hd__clkinv_1 U27748 ( .A(n25394), .Y(n23259) );
  sky130_fd_sc_hd__nand2_1 U27749 ( .A(j202_soc_core_uart_RDRXD1), .B(n23259), 
        .Y(n25205) );
  sky130_fd_sc_hd__o22ai_1 U27750 ( .A1(j202_soc_core_uart_TOP_rx_fifo_rp[0]), 
        .A2(n23261), .B1(n25206), .B2(j202_soc_core_uart_TOP_rx_fifo_wp[0]), 
        .Y(n23260) );
  sky130_fd_sc_hd__o211ai_1 U27751 ( .A1(j202_soc_core_uart_TOP_rx_fifo_wp[0]), 
        .A2(n23261), .B1(n25235), .C1(n23260), .Y(n23262) );
  sky130_fd_sc_hd__nand3_1 U27752 ( .A(n25734), .B(n25205), .C(n23262), .Y(
        j202_soc_core_uart_TOP_rx_fifo_N41) );
  sky130_fd_sc_hd__nor2_1 U27753 ( .A(j202_soc_core_rst), .B(n23262), .Y(
        j202_soc_core_uart_TOP_rx_fifo_N42) );
  sky130_fd_sc_hd__nor2_1 U27754 ( .A(j202_soc_core_rst), .B(
        j202_soc_core_uart_BRG_ps_clr), .Y(n24824) );
  sky130_fd_sc_hd__clkinv_1 U27755 ( .A(n24824), .Y(n23271) );
  sky130_fd_sc_hd__nor2_1 U27756 ( .A(j202_soc_core_uart_BRG_ps[0]), .B(n23271), .Y(j202_soc_core_uart_BRG_N12) );
  sky130_fd_sc_hd__nand2_1 U27757 ( .A(j202_soc_core_uart_BRG_ps[0]), .B(
        j202_soc_core_uart_BRG_ps[1]), .Y(n23264) );
  sky130_fd_sc_hd__o21ai_1 U27758 ( .A1(j202_soc_core_uart_BRG_ps[0]), .A2(
        j202_soc_core_uart_BRG_ps[1]), .B1(n23264), .Y(n23263) );
  sky130_fd_sc_hd__nor2_1 U27759 ( .A(n23271), .B(n23263), .Y(
        j202_soc_core_uart_BRG_N13) );
  sky130_fd_sc_hd__clkinv_1 U27760 ( .A(j202_soc_core_uart_BRG_ps[2]), .Y(
        n24816) );
  sky130_fd_sc_hd__nor2_1 U27761 ( .A(n24816), .B(n23264), .Y(n23265) );
  sky130_fd_sc_hd__a211oi_1 U27762 ( .A1(n24816), .A2(n23264), .B1(n23265), 
        .C1(n23271), .Y(j202_soc_core_uart_BRG_N14) );
  sky130_fd_sc_hd__nand2_1 U27763 ( .A(j202_soc_core_uart_BRG_ps[3]), .B(
        n23265), .Y(n23267) );
  sky130_fd_sc_hd__o21ai_1 U27764 ( .A1(j202_soc_core_uart_BRG_ps[3]), .A2(
        n23265), .B1(n23267), .Y(n23266) );
  sky130_fd_sc_hd__nor2_1 U27765 ( .A(n23271), .B(n23266), .Y(
        j202_soc_core_uart_BRG_N15) );
  sky130_fd_sc_hd__clkinv_1 U27766 ( .A(j202_soc_core_uart_BRG_ps[4]), .Y(
        n23268) );
  sky130_fd_sc_hd__nor2_1 U27767 ( .A(n23268), .B(n23267), .Y(n23269) );
  sky130_fd_sc_hd__a211oi_1 U27768 ( .A1(n23268), .A2(n23267), .B1(n23269), 
        .C1(n23271), .Y(j202_soc_core_uart_BRG_N16) );
  sky130_fd_sc_hd__nand2_1 U27769 ( .A(j202_soc_core_uart_BRG_ps[5]), .B(
        n23269), .Y(n23272) );
  sky130_fd_sc_hd__o21ai_1 U27770 ( .A1(j202_soc_core_uart_BRG_ps[5]), .A2(
        n23269), .B1(n23272), .Y(n23270) );
  sky130_fd_sc_hd__nor2_1 U27771 ( .A(n23271), .B(n23270), .Y(
        j202_soc_core_uart_BRG_N17) );
  sky130_fd_sc_hd__clkinv_1 U27772 ( .A(j202_soc_core_uart_BRG_ps[6]), .Y(
        n24820) );
  sky130_fd_sc_hd__nor2_1 U27773 ( .A(n24820), .B(n23272), .Y(n23274) );
  sky130_fd_sc_hd__a211oi_1 U27774 ( .A1(n24820), .A2(n23272), .B1(n23274), 
        .C1(n23271), .Y(j202_soc_core_uart_BRG_N18) );
  sky130_fd_sc_hd__a21oi_1 U27776 ( .A1(j202_soc_core_uart_BRG_ps[7]), .A2(
        n23274), .B1(n23273), .Y(j202_soc_core_uart_BRG_N19) );
  sky130_fd_sc_hd__nand3_1 U27777 ( .A(n25734), .B(n24823), .C(
        j202_soc_core_uart_BRG_ps_clr), .Y(n23284) );
  sky130_fd_sc_hd__nor2_1 U27778 ( .A(j202_soc_core_uart_BRG_br_cnt[0]), .B(
        n23284), .Y(j202_soc_core_uart_BRG_N35) );
  sky130_fd_sc_hd__nand2_1 U27779 ( .A(j202_soc_core_uart_BRG_br_cnt[1]), .B(
        j202_soc_core_uart_BRG_br_cnt[0]), .Y(n23276) );
  sky130_fd_sc_hd__o21ai_1 U27780 ( .A1(j202_soc_core_uart_BRG_br_cnt[1]), 
        .A2(j202_soc_core_uart_BRG_br_cnt[0]), .B1(n23276), .Y(n23275) );
  sky130_fd_sc_hd__nor2_1 U27781 ( .A(n23284), .B(n23275), .Y(
        j202_soc_core_uart_BRG_N36) );
  sky130_fd_sc_hd__clkinv_1 U27782 ( .A(j202_soc_core_uart_BRG_br_cnt[2]), .Y(
        n24798) );
  sky130_fd_sc_hd__nor2_1 U27783 ( .A(n24798), .B(n23276), .Y(n23277) );
  sky130_fd_sc_hd__a211oi_1 U27784 ( .A1(n24798), .A2(n23276), .B1(n23277), 
        .C1(n23284), .Y(j202_soc_core_uart_BRG_N37) );
  sky130_fd_sc_hd__nand2_1 U27785 ( .A(j202_soc_core_uart_BRG_br_cnt[3]), .B(
        n23277), .Y(n23279) );
  sky130_fd_sc_hd__o21ai_1 U27786 ( .A1(j202_soc_core_uart_BRG_br_cnt[3]), 
        .A2(n23277), .B1(n23279), .Y(n23278) );
  sky130_fd_sc_hd__nor2_1 U27787 ( .A(n23284), .B(n23278), .Y(
        j202_soc_core_uart_BRG_N38) );
  sky130_fd_sc_hd__clkinv_1 U27788 ( .A(j202_soc_core_uart_BRG_br_cnt[4]), .Y(
        n23280) );
  sky130_fd_sc_hd__nor2_1 U27789 ( .A(n23280), .B(n23279), .Y(n23281) );
  sky130_fd_sc_hd__a211oi_1 U27790 ( .A1(n23280), .A2(n23279), .B1(n23281), 
        .C1(n23284), .Y(j202_soc_core_uart_BRG_N39) );
  sky130_fd_sc_hd__nand2_1 U27791 ( .A(j202_soc_core_uart_BRG_br_cnt[5]), .B(
        n23281), .Y(n23283) );
  sky130_fd_sc_hd__nor2_1 U27793 ( .A(n23284), .B(n23282), .Y(
        j202_soc_core_uart_BRG_N40) );
  sky130_fd_sc_hd__clkinv_1 U27794 ( .A(j202_soc_core_uart_BRG_br_cnt[6]), .Y(
        n24802) );
  sky130_fd_sc_hd__nor2_1 U27795 ( .A(n24802), .B(n23283), .Y(n23286) );
  sky130_fd_sc_hd__a211oi_1 U27796 ( .A1(n24802), .A2(n23283), .B1(n23286), 
        .C1(n23284), .Y(j202_soc_core_uart_BRG_N41) );
  sky130_fd_sc_hd__o21bai_1 U27797 ( .A1(j202_soc_core_uart_BRG_br_cnt[7]), 
        .A2(n23286), .B1_N(n23284), .Y(n23285) );
  sky130_fd_sc_hd__a21oi_1 U27798 ( .A1(j202_soc_core_uart_BRG_br_cnt[7]), 
        .A2(n23286), .B1(n23285), .Y(j202_soc_core_uart_BRG_N42) );
  sky130_fd_sc_hd__nand2_1 U27799 ( .A(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_), .B(
        j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_1), .Y(n23288)
         );
  sky130_fd_sc_hd__clkinv_1 U27800 ( .A(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_wen), .Y(
        n25162) );
  sky130_fd_sc_hd__a2bb2oi_1 U27801 ( .B1(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_latch_status_0_), .B2(n25162), .A1_N(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_0_), .A2_N(
        n23809), .Y(n23287) );
  sky130_fd_sc_hd__o21ai_1 U27802 ( .A1(
        j202_soc_core_bldc_core_00_bldc_hall_00_latch_data_en_2), .A2(n23288), 
        .B1(n23287), .Y(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_00_nxt_latch_status_0_) );
  sky130_fd_sc_hd__a21oi_1 U27803 ( .A1(n23291), .A2(n23290), .B1(n25111), .Y(
        n23547) );
  sky130_fd_sc_hd__clkinv_1 U27804 ( .A(n23583), .Y(n23548) );
  sky130_fd_sc_hd__nor2_1 U27805 ( .A(n25111), .B(n23292), .Y(n23540) );
  sky130_fd_sc_hd__a21oi_1 U27806 ( .A1(n23292), .A2(n23396), .B1(n23540), .Y(
        n23293) );
  sky130_fd_sc_hd__clkinv_1 U27807 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[0]), .Y(n23792) );
  sky130_fd_sc_hd__nand4_1 U27808 ( .A(n23788), .B(
        j202_soc_core_wbqspiflash_00_spi_valid), .C(n23789), .D(n23792), .Y(
        n23582) );
  sky130_fd_sc_hd__nand2_1 U27810 ( .A(n23478), .B(n23466), .Y(n23436) );
  sky130_fd_sc_hd__nand2b_1 U27811 ( .A_N(n23349), .B(n23436), .Y(n23373) );
  sky130_fd_sc_hd__o22ai_1 U27812 ( .A1(n23293), .A2(n25107), .B1(n23505), 
        .B2(n23373), .Y(n23294) );
  sky130_fd_sc_hd__a211o_1 U27813 ( .A1(n23547), .A2(n23548), .B1(n23295), 
        .C1(n23294), .X(j202_soc_core_wbqspiflash_00_N590) );
  sky130_fd_sc_hd__nand2_1 U27814 ( .A(j202_soc_core_wbqspiflash_00_spi_busy), 
        .B(n24898), .Y(n23539) );
  sky130_fd_sc_hd__a22oi_1 U27815 ( .A1(n25070), .A2(n25068), .B1(n23528), 
        .B2(n23539), .Y(j202_soc_core_wbqspiflash_00_N592) );
  sky130_fd_sc_hd__a21oi_1 U27816 ( .A1(n25011), .A2(n23467), .B1(
        j202_soc_core_wbqspiflash_00_state[4]), .Y(n23371) );
  sky130_fd_sc_hd__nand3b_1 U27817 ( .A_N(n23371), .B(n25107), .C(n23577), .Y(
        j202_soc_core_wbqspiflash_00_N594) );
  sky130_fd_sc_hd__o21ai_1 U27818 ( .A1(n23343), .A2(n23298), .B1(n23339), .Y(
        n23299) );
  sky130_fd_sc_hd__o21ai_0 U27819 ( .A1(n23300), .A2(n23347), .B1(n23299), .Y(
        j202_soc_core_j22_cpu_ml_N354) );
  sky130_fd_sc_hd__o21ai_0 U27821 ( .A1(n23303), .A2(n23347), .B1(n23302), .Y(
        j202_soc_core_j22_cpu_ml_N355) );
  sky130_fd_sc_hd__o21ai_0 U27823 ( .A1(n23306), .A2(n23347), .B1(n23305), .Y(
        j202_soc_core_j22_cpu_ml_N356) );
  sky130_fd_sc_hd__o21ai_1 U27824 ( .A1(n23343), .A2(n23307), .B1(n23339), .Y(
        n23308) );
  sky130_fd_sc_hd__o21ai_0 U27825 ( .A1(n23309), .A2(n23347), .B1(n23308), .Y(
        j202_soc_core_j22_cpu_ml_N357) );
  sky130_fd_sc_hd__o21ai_1 U27826 ( .A1(n23343), .A2(n23310), .B1(n23339), .Y(
        n23311) );
  sky130_fd_sc_hd__o21ai_0 U27827 ( .A1(n23312), .A2(n23347), .B1(n23311), .Y(
        j202_soc_core_j22_cpu_ml_N359) );
  sky130_fd_sc_hd__o21ai_1 U27828 ( .A1(n23343), .A2(n23313), .B1(n23339), .Y(
        n23314) );
  sky130_fd_sc_hd__o21ai_0 U27829 ( .A1(n23315), .A2(n23347), .B1(n23314), .Y(
        j202_soc_core_j22_cpu_ml_N360) );
  sky130_fd_sc_hd__a21oi_1 U27830 ( .A1(n23345), .A2(n23316), .B1(n23343), .Y(
        n23317) );
  sky130_fd_sc_hd__o21ai_0 U27831 ( .A1(n23318), .A2(n23347), .B1(n23317), .Y(
        j202_soc_core_j22_cpu_ml_N361) );
  sky130_fd_sc_hd__o21ai_0 U27833 ( .A1(n23321), .A2(n23347), .B1(n23320), .Y(
        j202_soc_core_j22_cpu_ml_N362) );
  sky130_fd_sc_hd__o21ai_1 U27834 ( .A1(n23343), .A2(n23322), .B1(n23339), .Y(
        n23323) );
  sky130_fd_sc_hd__o21ai_0 U27835 ( .A1(n21937), .A2(n23347), .B1(n23323), .Y(
        j202_soc_core_j22_cpu_ml_N363) );
  sky130_fd_sc_hd__o21ai_1 U27836 ( .A1(n23343), .A2(n23324), .B1(n23339), .Y(
        n23325) );
  sky130_fd_sc_hd__o21ai_0 U27837 ( .A1(n23326), .A2(n23347), .B1(n23325), .Y(
        j202_soc_core_j22_cpu_ml_N364) );
  sky130_fd_sc_hd__o21ai_1 U27838 ( .A1(n23343), .A2(n23327), .B1(n23339), .Y(
        n23328) );
  sky130_fd_sc_hd__o21ai_0 U27839 ( .A1(n23329), .A2(n23347), .B1(n23328), .Y(
        j202_soc_core_j22_cpu_ml_N365) );
  sky130_fd_sc_hd__o21ai_0 U27841 ( .A1(n23332), .A2(n23347), .B1(n23331), .Y(
        j202_soc_core_j22_cpu_ml_N366) );
  sky130_fd_sc_hd__o21ai_1 U27842 ( .A1(n23343), .A2(n23333), .B1(n23339), .Y(
        n23334) );
  sky130_fd_sc_hd__o21ai_0 U27843 ( .A1(n23335), .A2(n23347), .B1(n23334), .Y(
        j202_soc_core_j22_cpu_ml_N367) );
  sky130_fd_sc_hd__o21ai_0 U27845 ( .A1(n23338), .A2(n23347), .B1(n23337), .Y(
        j202_soc_core_j22_cpu_ml_N368) );
  sky130_fd_sc_hd__o21ai_1 U27846 ( .A1(n23343), .A2(n23340), .B1(n23339), .Y(
        n23341) );
  sky130_fd_sc_hd__o21ai_0 U27847 ( .A1(n23342), .A2(n23347), .B1(n23341), .Y(
        j202_soc_core_j22_cpu_ml_N369) );
  sky130_fd_sc_hd__a21oi_1 U27848 ( .A1(n23345), .A2(n23344), .B1(n23343), .Y(
        n23346) );
  sky130_fd_sc_hd__o21ai_1 U27849 ( .A1(n23348), .A2(n23347), .B1(n23346), .Y(
        j202_soc_core_j22_cpu_ml_N370) );
  sky130_fd_sc_hd__nand2_1 U27850 ( .A(n23384), .B(
        j202_soc_core_wbqspiflash_00_state[4]), .Y(n25101) );
  sky130_fd_sc_hd__nor2_1 U27851 ( .A(n23398), .B(n25101), .Y(n24954) );
  sky130_fd_sc_hd__a21oi_1 U27852 ( .A1(n24954), .A2(n25100), .B1(n23349), .Y(
        n23522) );
  sky130_fd_sc_hd__nand2_1 U27853 ( .A(j202_soc_core_wbqspiflash_00_spi_valid), 
        .B(n25731), .Y(n23362) );
  sky130_fd_sc_hd__o22ai_1 U27854 ( .A1(j202_soc_core_rst), .A2(n23522), .B1(
        n23362), .B2(n25108), .Y(j202_soc_core_wbqspiflash_00_N749) );
  sky130_fd_sc_hd__o211ai_1 U27855 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_valid), .A2(
        j202_soc_core_wbqspiflash_00_state[4]), .B1(
        j202_soc_core_wbqspiflash_00_state[2]), .C1(n23450), .Y(n23350) );
  sky130_fd_sc_hd__a21oi_1 U27856 ( .A1(n23522), .A2(n23350), .B1(
        j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N750) );
  sky130_fd_sc_hd__nand2_1 U27857 ( .A(n23536), .B(n23788), .Y(n25002) );
  sky130_fd_sc_hd__clkinv_1 U27858 ( .A(n25002), .Y(n23393) );
  sky130_fd_sc_hd__nor2_1 U27859 ( .A(j202_soc_core_rst), .B(n23393), .Y(
        j202_soc_core_wbqspiflash_00_N748) );
  sky130_fd_sc_hd__a21oi_1 U27860 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), 
        .A2(n25000), .B1(n23351), .Y(n23353) );
  sky130_fd_sc_hd__nand2_1 U27861 ( .A(n23384), .B(n25005), .Y(n23352) );
  sky130_fd_sc_hd__a21oi_1 U27862 ( .A1(n23353), .A2(n23352), .B1(
        j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N747) );
  sky130_fd_sc_hd__nor2_1 U27863 ( .A(j202_soc_core_rst), .B(
        j202_soc_core_wbqspiflash_00_state[1]), .Y(n23394) );
  sky130_fd_sc_hd__a21oi_1 U27865 ( .A1(n25027), .A2(n23356), .B1(n23355), .Y(
        n23357) );
  sky130_fd_sc_hd__o22ai_1 U27866 ( .A1(n23536), .A2(n23358), .B1(
        j202_soc_core_rst), .B2(n23357), .Y(j202_soc_core_wbqspiflash_00_N745)
         );
  sky130_fd_sc_hd__nor3_1 U27867 ( .A(j202_soc_core_rst), .B(n23359), .C(
        n23756), .Y(j202_soc_core_wbqspiflash_00_N744) );
  sky130_fd_sc_hd__nand2_1 U27868 ( .A(n25734), .B(n23360), .Y(
        j202_soc_core_wbqspiflash_00_N743) );
  sky130_fd_sc_hd__nand2_1 U27869 ( .A(n25732), .B(n23361), .Y(
        j202_soc_core_wbqspiflash_00_N742) );
  sky130_fd_sc_hd__nor2_1 U27870 ( .A(n23577), .B(n23362), .Y(
        j202_soc_core_wbqspiflash_00_N741) );
  sky130_fd_sc_hd__a21oi_1 U27871 ( .A1(
        j202_soc_core_wbqspiflash_00_write_in_progress), .A2(n23792), .B1(
        n23363), .Y(n23365) );
  sky130_fd_sc_hd__nor2_1 U27872 ( .A(j202_soc_core_rst), .B(n23364), .Y(
        n23560) );
  sky130_fd_sc_hd__nand2_1 U27874 ( .A(j202_soc_core_wbqspiflash_00_spi_out[1]), .B(n23754), .Y(n23367) );
  sky130_fd_sc_hd__nor2_1 U27875 ( .A(n23412), .B(n23366), .Y(n24991) );
  sky130_fd_sc_hd__nand2_1 U27876 ( .A(n24991), .B(
        j202_soc_core_wbqspiflash_00_spif_data[1]), .Y(n24917) );
  sky130_fd_sc_hd__a21oi_1 U27877 ( .A1(n23367), .A2(n24917), .B1(
        j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N739) );
  sky130_fd_sc_hd__nand2_1 U27878 ( .A(n25100), .B(n24991), .Y(n23369) );
  sky130_fd_sc_hd__nand3_1 U27879 ( .A(n25734), .B(n23369), .C(n23368), .Y(
        j202_soc_core_wbqspiflash_00_N738) );
  sky130_fd_sc_hd__a211oi_1 U27880 ( .A1(j202_soc_core_qspi_wb_cyc), .A2(
        j202_soc_core_ahb2wbqspi_00_stb_o), .B1(n23495), .C1(n23577), .Y(
        n23390) );
  sky130_fd_sc_hd__clkinv_1 U27881 ( .A(n24991), .Y(n25010) );
  sky130_fd_sc_hd__a21oi_1 U27882 ( .A1(n24960), .A2(n25010), .B1(n23370), .Y(
        n23580) );
  sky130_fd_sc_hd__a21oi_1 U27883 ( .A1(n23372), .A2(n25070), .B1(n23371), .Y(
        n23374) );
  sky130_fd_sc_hd__nand4_1 U27884 ( .A(n23375), .B(n23374), .C(n25073), .D(
        n23373), .Y(n23389) );
  sky130_fd_sc_hd__clkinv_1 U27885 ( .A(n23445), .Y(n23378) );
  sky130_fd_sc_hd__a21oi_1 U27886 ( .A1(n23378), .A2(n23377), .B1(n23376), .Y(
        n23387) );
  sky130_fd_sc_hd__a21oi_1 U27887 ( .A1(n23381), .A2(n23380), .B1(n23379), .Y(
        n23386) );
  sky130_fd_sc_hd__nand4_1 U27888 ( .A(n23384), .B(n25005), .C(n23383), .D(
        n23382), .Y(n23385) );
  sky130_fd_sc_hd__o22ai_1 U27889 ( .A1(n23387), .A2(n23515), .B1(n23386), 
        .B2(n23385), .Y(n23388) );
  sky130_fd_sc_hd__nor4_1 U27890 ( .A(n23390), .B(n23580), .C(n23389), .D(
        n23388), .Y(n23391) );
  sky130_fd_sc_hd__a21oi_1 U27891 ( .A1(n23392), .A2(n23391), .B1(
        j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N734) );
  sky130_fd_sc_hd__nand3_1 U27892 ( .A(n23393), .B(n25734), .C(n23785), .Y(
        j202_soc_core_wbqspiflash_00_N733) );
  sky130_fd_sc_hd__o211ai_1 U27893 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), .A2(n23395), .B1(n25116), .C1(n23394), .Y(j202_soc_core_wbqspiflash_00_N729)
         );
  sky130_fd_sc_hd__nor2_1 U27894 ( .A(n23396), .B(n25109), .Y(n23449) );
  sky130_fd_sc_hd__nor2_1 U27895 ( .A(n23540), .B(
        j202_soc_core_wbqspiflash_00_spi_spd), .Y(n23397) );
  sky130_fd_sc_hd__o21ai_1 U27896 ( .A1(n23449), .A2(n23397), .B1(n23455), .Y(
        n23424) );
  sky130_fd_sc_hd__nor2_1 U27897 ( .A(j202_soc_core_wbqspiflash_00_state[1]), 
        .B(n23398), .Y(n23421) );
  sky130_fd_sc_hd__nor2_1 U27898 ( .A(n23451), .B(
        j202_soc_core_wbqspiflash_00_state[0]), .Y(n23493) );
  sky130_fd_sc_hd__clkinv_1 U27899 ( .A(n23493), .Y(n23400) );
  sky130_fd_sc_hd__clkinv_1 U27900 ( .A(n23468), .Y(n24911) );
  sky130_fd_sc_hd__a31oi_1 U27901 ( .A1(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled), .A2(n25027), .A3(
        n23789), .B1(n24911), .Y(n23399) );
  sky130_fd_sc_hd__o211ai_1 U27903 ( .A1(n23402), .A2(n23562), .B1(n25032), 
        .C1(n23401), .Y(n23415) );
  sky130_fd_sc_hd__nand2_1 U27904 ( .A(n23409), .B(
        j202_soc_core_qspi_wb_addr[2]), .Y(n25066) );
  sky130_fd_sc_hd__clkinv_1 U27905 ( .A(n23403), .Y(n23405) );
  sky130_fd_sc_hd__nand3_1 U27906 ( .A(n23404), .B(n23495), .C(n23758), .Y(
        n23430) );
  sky130_fd_sc_hd__a21oi_1 U27908 ( .A1(n23425), .A2(n25066), .B1(n23406), .Y(
        n23411) );
  sky130_fd_sc_hd__clkinv_1 U27909 ( .A(n23407), .Y(n23429) );
  sky130_fd_sc_hd__a31oi_1 U27910 ( .A1(n23429), .A2(n23495), .A3(n23409), 
        .B1(n23408), .Y(n23410) );
  sky130_fd_sc_hd__nand2_1 U27911 ( .A(n23411), .B(n23410), .Y(n23414) );
  sky130_fd_sc_hd__nor2_1 U27912 ( .A(j202_soc_core_wbqspiflash_00_state[0]), 
        .B(n23412), .Y(n24996) );
  sky130_fd_sc_hd__a222oi_1 U27913 ( .A1(n23415), .A2(n23479), .B1(n23414), 
        .B2(n23493), .C1(n23413), .C2(n24996), .Y(n23416) );
  sky130_fd_sc_hd__o22ai_1 U27914 ( .A1(n23547), .A2(n23417), .B1(
        j202_soc_core_wbqspiflash_00_state[3]), .B2(n23416), .Y(n23418) );
  sky130_fd_sc_hd__nor4_1 U27915 ( .A(n23421), .B(n23420), .C(n23419), .D(
        n23418), .Y(n23423) );
  sky130_fd_sc_hd__nor2_1 U27916 ( .A(n25070), .B(n23422), .Y(n25063) );
  sky130_fd_sc_hd__nand2_1 U27917 ( .A(n23762), .B(n25063), .Y(n25055) );
  sky130_fd_sc_hd__a31oi_1 U27918 ( .A1(n23424), .A2(n23423), .A3(n25055), 
        .B1(j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N724) );
  sky130_fd_sc_hd__clkinv_1 U27919 ( .A(n23425), .Y(n23426) );
  sky130_fd_sc_hd__o22ai_1 U27920 ( .A1(n23465), .A2(n25061), .B1(n25053), 
        .B2(n23426), .Y(n23427) );
  sky130_fd_sc_hd__a21oi_1 U27921 ( .A1(n23429), .A2(n23428), .B1(n23427), .Y(
        n23432) );
  sky130_fd_sc_hd__a31oi_1 U27922 ( .A1(n23432), .A2(n23431), .A3(n23430), 
        .B1(n23464), .Y(n23444) );
  sky130_fd_sc_hd__nor2_1 U27923 ( .A(n23542), .B(n23433), .Y(n23512) );
  sky130_fd_sc_hd__nor2_1 U27924 ( .A(
        j202_soc_core_wbqspiflash_00_last_status[6]), .B(
        j202_soc_core_wbqspiflash_00_last_status[5]), .Y(n23434) );
  sky130_fd_sc_hd__nor3_1 U27925 ( .A(n23434), .B(
        j202_soc_core_wbqspiflash_00_spif_data[6]), .C(
        j202_soc_core_wbqspiflash_00_spif_data[5]), .Y(n23504) );
  sky130_fd_sc_hd__nor3_1 U27926 ( .A(n25005), .B(n23504), .C(n23435), .Y(
        n23439) );
  sky130_fd_sc_hd__clkinv_1 U27927 ( .A(n23541), .Y(n23527) );
  sky130_fd_sc_hd__a21oi_1 U27928 ( .A1(n25064), .A2(n25063), .B1(n23436), .Y(
        n23437) );
  sky130_fd_sc_hd__o22ai_1 U27929 ( .A1(n23788), .A2(n23527), .B1(n23526), 
        .B2(n23437), .Y(n23438) );
  sky130_fd_sc_hd__nor4_1 U27930 ( .A(n25106), .B(n23512), .C(n23439), .D(
        n23438), .Y(n23440) );
  sky130_fd_sc_hd__o21ai_1 U27931 ( .A1(n23442), .A2(n23441), .B1(n23440), .Y(
        n23443) );
  sky130_fd_sc_hd__nor2_1 U27932 ( .A(n23444), .B(n23443), .Y(n23454) );
  sky130_fd_sc_hd__a31oi_1 U27934 ( .A1(
        j202_soc_core_wbqspiflash_00_write_in_progress), .A2(n24998), .A3(
        n23758), .B1(n23445), .Y(n23446) );
  sky130_fd_sc_hd__o21ai_1 U27935 ( .A1(n23448), .A2(n23447), .B1(n23446), .Y(
        n23453) );
  sky130_fd_sc_hd__nor2_1 U27936 ( .A(n23449), .B(n23540), .Y(n23458) );
  sky130_fd_sc_hd__o21ai_1 U27937 ( .A1(n23458), .A2(n23451), .B1(n23450), .Y(
        n23452) );
  sky130_fd_sc_hd__a31oi_1 U27938 ( .A1(n23454), .A2(n23453), .A3(n23452), 
        .B1(j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N725) );
  sky130_fd_sc_hd__nor2b_1 U27939 ( .B_N(n23455), .A(
        j202_soc_core_wbqspiflash_00_spi_spd), .Y(n23459) );
  sky130_fd_sc_hd__a22oi_1 U27940 ( .A1(n23459), .A2(n23458), .B1(n23457), 
        .B2(n23456), .Y(n23473) );
  sky130_fd_sc_hd__o22ai_1 U27941 ( .A1(n23541), .A2(n25101), .B1(n23526), 
        .B2(n23476), .Y(n23460) );
  sky130_fd_sc_hd__a221oi_1 U27942 ( .A1(n23463), .A2(n23462), .B1(n23461), 
        .B2(n23462), .C1(n23460), .Y(n23472) );
  sky130_fd_sc_hd__nor2_1 U27943 ( .A(n23465), .B(n23464), .Y(n24910) );
  sky130_fd_sc_hd__nand4_1 U27944 ( .A(n23468), .B(n23467), .C(n23466), .D(
        n25072), .Y(n23469) );
  sky130_fd_sc_hd__nor3_1 U27945 ( .A(n23470), .B(n24910), .C(n23469), .Y(
        n23471) );
  sky130_fd_sc_hd__a31oi_1 U27946 ( .A1(n23473), .A2(n23472), .A3(n23471), 
        .B1(j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N726) );
  sky130_fd_sc_hd__clkinv_1 U27947 ( .A(n23474), .Y(n23475) );
  sky130_fd_sc_hd__nand2_1 U27948 ( .A(n23475), .B(n25053), .Y(n23489) );
  sky130_fd_sc_hd__nor3_1 U27949 ( .A(n23547), .B(n23476), .C(n24899), .Y(
        n23487) );
  sky130_fd_sc_hd__o22ai_1 U27950 ( .A1(j202_soc_core_wbqspiflash_00_state[4]), 
        .A2(n23478), .B1(n23477), .B2(n23523), .Y(n23486) );
  sky130_fd_sc_hd__nand2_1 U27951 ( .A(n23479), .B(n23788), .Y(n23559) );
  sky130_fd_sc_hd__clkinv_1 U27952 ( .A(n23559), .Y(n25093) );
  sky130_fd_sc_hd__a21oi_1 U27953 ( .A1(n23498), .A2(n25093), .B1(n23480), .Y(
        n23484) );
  sky130_fd_sc_hd__nand3_1 U27955 ( .A(n23484), .B(n23483), .C(n23482), .Y(
        n23485) );
  sky130_fd_sc_hd__nor4_1 U27956 ( .A(n23487), .B(n25085), .C(n23486), .D(
        n23485), .Y(n23488) );
  sky130_fd_sc_hd__o22ai_1 U27957 ( .A1(
        j202_soc_core_wbqspiflash_00_write_in_progress), .A2(n23489), .B1(
        j202_soc_core_rst), .B2(n23488), .Y(j202_soc_core_wbqspiflash_00_N727)
         );
  sky130_fd_sc_hd__o21ai_1 U27958 ( .A1(j202_soc_core_wbqspiflash_00_state[2]), 
        .A2(n24998), .B1(n23490), .Y(n23492) );
  sky130_fd_sc_hd__clkinv_1 U27959 ( .A(n25044), .Y(n24974) );
  sky130_fd_sc_hd__nand4_1 U27960 ( .A(n25004), .B(n23492), .C(n23491), .D(
        n24974), .Y(n23503) );
  sky130_fd_sc_hd__nand2_1 U27961 ( .A(n23493), .B(
        j202_soc_core_ahb2wbqspi_00_stb_o), .Y(n25023) );
  sky130_fd_sc_hd__clkinv_1 U27962 ( .A(n25023), .Y(n23497) );
  sky130_fd_sc_hd__a21oi_1 U27964 ( .A1(n23497), .A2(n23496), .B1(n23789), .Y(
        n23501) );
  sky130_fd_sc_hd__a21oi_1 U27965 ( .A1(n24998), .A2(n23758), .B1(n23498), .Y(
        n23499) );
  sky130_fd_sc_hd__nand2_1 U27966 ( .A(j202_soc_core_wbqspiflash_00_state[2]), 
        .B(n23514), .Y(n25029) );
  sky130_fd_sc_hd__o22ai_1 U27967 ( .A1(n23501), .A2(n23500), .B1(n23499), 
        .B2(n25029), .Y(n23502) );
  sky130_fd_sc_hd__a211oi_1 U27968 ( .A1(n24954), .A2(n23504), .B1(n23503), 
        .C1(n23502), .Y(n23508) );
  sky130_fd_sc_hd__or3_1 U27969 ( .A(j202_soc_core_wbqspiflash_00_state[3]), 
        .B(n23506), .C(n23505), .X(n23507) );
  sky130_fd_sc_hd__a21oi_1 U27970 ( .A1(n23508), .A2(n23507), .B1(
        j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N728) );
  sky130_fd_sc_hd__a21o_1 U27971 ( .A1(j202_soc_core_wbqspiflash_00_spi_valid), 
        .A2(n23510), .B1(n23509), .X(n25098) );
  sky130_fd_sc_hd__a21oi_1 U27972 ( .A1(n25046), .A2(n25098), .B1(n23511), .Y(
        n23557) );
  sky130_fd_sc_hd__a21oi_1 U27973 ( .A1(n23789), .A2(
        j202_soc_core_wbqspiflash_00_state[1]), .B1(n23512), .Y(n23517) );
  sky130_fd_sc_hd__nand2_1 U27974 ( .A(n23514), .B(n23513), .Y(n23516) );
  sky130_fd_sc_hd__a21oi_1 U27975 ( .A1(n23517), .A2(n23516), .B1(n23515), .Y(
        n23556) );
  sky130_fd_sc_hd__a21oi_1 U27976 ( .A1(
        j202_soc_core_wbqspiflash_00_write_in_progress), .A2(n23519), .B1(
        n23518), .Y(n23524) );
  sky130_fd_sc_hd__a31oi_1 U27977 ( .A1(j202_soc_core_wbqspiflash_00_spi_valid), .A2(n23533), .A3(n25077), .B1(n23520), .Y(n23521) );
  sky130_fd_sc_hd__o211ai_1 U27978 ( .A1(n23524), .A2(n23523), .B1(n23522), 
        .C1(n23521), .Y(n23555) );
  sky130_fd_sc_hd__a21oi_1 U27979 ( .A1(n23787), .A2(n25100), .B1(n23525), .Y(
        n23553) );
  sky130_fd_sc_hd__clkinv_1 U27980 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[31]), .Y(n23733) );
  sky130_fd_sc_hd__nor3_1 U27981 ( .A(j202_soc_core_wbqspiflash_00_spi_in[28]), 
        .B(j202_soc_core_wbqspiflash_00_spi_in[30]), .C(n23733), .Y(n23532) );
  sky130_fd_sc_hd__a31oi_1 U27982 ( .A1(n23526), .A2(
        j202_soc_core_wbqspiflash_00_state[0]), .A3(n23534), .B1(n25001), .Y(
        n23530) );
  sky130_fd_sc_hd__nor2_1 U27983 ( .A(n23528), .B(n23527), .Y(n25080) );
  sky130_fd_sc_hd__clkinv_1 U27984 ( .A(n25080), .Y(n25090) );
  sky130_fd_sc_hd__o22ai_1 U27985 ( .A1(n23530), .A2(n23529), .B1(n23735), 
        .B2(n25090), .Y(n23531) );
  sky130_fd_sc_hd__a31oi_1 U27986 ( .A1(n25085), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[29]), .A3(n23532), .B1(n23531), 
        .Y(n23538) );
  sky130_fd_sc_hd__nand4_1 U27987 ( .A(n23536), .B(n23535), .C(n23534), .D(
        n23533), .Y(n23537) );
  sky130_fd_sc_hd__a21oi_1 U27988 ( .A1(n23538), .A2(n23537), .B1(
        j202_soc_core_wbqspiflash_00_spi_busy), .Y(n23546) );
  sky130_fd_sc_hd__o21ai_1 U27990 ( .A1(n23542), .A2(n23541), .B1(n25100), .Y(
        n23543) );
  sky130_fd_sc_hd__o22ai_1 U27991 ( .A1(n25101), .A2(n23543), .B1(n25073), 
        .B2(n23593), .Y(n23544) );
  sky130_fd_sc_hd__nor3_1 U27992 ( .A(n23546), .B(n23545), .C(n23544), .Y(
        n23552) );
  sky130_fd_sc_hd__nand4_1 U27994 ( .A(n23553), .B(n23552), .C(n25731), .D(
        n23551), .Y(n23554) );
  sky130_fd_sc_hd__nor4_1 U27995 ( .A(n23557), .B(n23556), .C(n23555), .D(
        n23554), .Y(n23558) );
  sky130_fd_sc_hd__o22ai_1 U27997 ( .A1(n25395), .A2(n23560), .B1(
        j202_soc_core_wbqspiflash_00_spif_data[28]), .B2(n23559), .Y(
        j202_soc_core_wbqspiflash_00_N722) );
  sky130_fd_sc_hd__o31a_1 U27998 ( .A1(n23757), .A2(n23562), .A3(n23561), .B1(
        n25734), .X(n23563) );
  sky130_fd_sc_hd__o22ai_1 U28000 ( .A1(n25052), .A2(
        j202_soc_core_wbqspiflash_00_erased_sector[4]), .B1(n25089), .B2(
        j202_soc_core_wbqspiflash_00_erased_sector[7]), .Y(n23565) );
  sky130_fd_sc_hd__a221o_1 U28001 ( .A1(n25052), .A2(
        j202_soc_core_wbqspiflash_00_erased_sector[4]), .B1(
        j202_soc_core_wbqspiflash_00_erased_sector[7]), .B2(n25089), .C1(
        n23565), .X(n23576) );
  sky130_fd_sc_hd__o22ai_1 U28002 ( .A1(n23567), .A2(
        j202_soc_core_wbqspiflash_00_erased_sector[3]), .B1(n25069), .B2(
        j202_soc_core_wbqspiflash_00_erased_sector[5]), .Y(n23566) );
  sky130_fd_sc_hd__a221oi_1 U28003 ( .A1(n23567), .A2(
        j202_soc_core_wbqspiflash_00_erased_sector[3]), .B1(
        j202_soc_core_wbqspiflash_00_erased_sector[5]), .B2(n25069), .C1(
        n23566), .Y(n23574) );
  sky130_fd_sc_hd__o22ai_1 U28004 ( .A1(n25019), .A2(
        j202_soc_core_wbqspiflash_00_erased_sector[1]), .B1(n23569), .B2(
        j202_soc_core_wbqspiflash_00_erased_sector[2]), .Y(n23568) );
  sky130_fd_sc_hd__a221oi_1 U28005 ( .A1(n25019), .A2(
        j202_soc_core_wbqspiflash_00_erased_sector[1]), .B1(
        j202_soc_core_wbqspiflash_00_erased_sector[2]), .B2(n23569), .C1(
        n23568), .Y(n23573) );
  sky130_fd_sc_hd__o22ai_1 U28006 ( .A1(n24944), .A2(
        j202_soc_core_wbqspiflash_00_erased_sector[0]), .B1(n23571), .B2(
        j202_soc_core_wbqspiflash_00_erased_sector[6]), .Y(n23570) );
  sky130_fd_sc_hd__a221oi_1 U28007 ( .A1(n24944), .A2(
        j202_soc_core_wbqspiflash_00_erased_sector[0]), .B1(
        j202_soc_core_wbqspiflash_00_erased_sector[6]), .B2(n23571), .C1(
        n23570), .Y(n23572) );
  sky130_fd_sc_hd__nand4_1 U28008 ( .A(n24898), .B(n23574), .C(n23573), .D(
        n23572), .Y(n23575) );
  sky130_fd_sc_hd__clkinv_1 U28010 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[14]), .Y(n24942) );
  sky130_fd_sc_hd__nor2_1 U28011 ( .A(j202_soc_core_rst), .B(n24942), .Y(
        j202_soc_core_wbqspiflash_00_N711) );
  sky130_fd_sc_hd__clkinv_1 U28012 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[18]), .Y(n24966) );
  sky130_fd_sc_hd__nor2_1 U28013 ( .A(j202_soc_core_rst), .B(n24966), .Y(
        j202_soc_core_wbqspiflash_00_N715) );
  sky130_fd_sc_hd__clkinv_1 U28014 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[19]), .Y(n24973) );
  sky130_fd_sc_hd__nor2_1 U28015 ( .A(j202_soc_core_rst), .B(n24973), .Y(
        j202_soc_core_wbqspiflash_00_N716) );
  sky130_fd_sc_hd__nand2_1 U28016 ( .A(n25108), .B(n23577), .Y(n23581) );
  sky130_fd_sc_hd__a22oi_1 U28017 ( .A1(j202_soc_core_wbqspiflash_00_state[4]), 
        .A2(n23578), .B1(j202_soc_core_wbqspiflash_00_spi_out[0]), .B2(n23581), 
        .Y(n23579) );
  sky130_fd_sc_hd__a21oi_1 U28018 ( .A1(n23579), .A2(n23583), .B1(
        j202_soc_core_rst), .Y(j202_soc_core_wbqspiflash_00_N709) );
  sky130_fd_sc_hd__a21oi_1 U28019 ( .A1(j202_soc_core_wbqspiflash_00_spi_valid), .A2(n23581), .B1(n23580), .Y(n23584) );
  sky130_fd_sc_hd__nand4_1 U28020 ( .A(n23585), .B(n23584), .C(n23583), .D(
        n23582), .Y(j202_soc_core_wbqspiflash_00_N708) );
  sky130_fd_sc_hd__nand2_1 U28021 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .B(
        j202_soc_core_wbqspiflash_00_alt_ctrl), .Y(n23586) );
  sky130_fd_sc_hd__o21ai_0 U28022 ( .A1(n23587), .A2(
        j202_soc_core_wbqspiflash_00_spif_override), .B1(n23586), .Y(io_out[9]) );
  sky130_fd_sc_hd__nand2_1 U28023 ( .A(n23738), .B(n23588), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N356) );
  sky130_fd_sc_hd__nand3_1 U28025 ( .A(n23599), .B(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .C(n23591), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N354) );
  sky130_fd_sc_hd__a31oi_1 U28026 ( .A1(j202_soc_core_wbqspiflash_00_spi_wr), 
        .A2(n23592), .A3(j202_soc_core_wbqspiflash_00_lldriver_state[0]), .B1(
        n23750), .Y(n23595) );
  sky130_fd_sc_hd__or4_1 U28028 ( .A(n23596), .B(n23595), .C(n23594), .D(
        n25396), .X(j202_soc_core_wbqspiflash_00_lldriver_N321) );
  sky130_fd_sc_hd__nand2b_1 U28030 ( .A_N(n23741), .B(n23598), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N315) );
  sky130_fd_sc_hd__nand2b_1 U28031 ( .A_N(
        j202_soc_core_wbqspiflash_00_lldriver_N423), .B(n23599), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N313) );
  sky130_fd_sc_hd__nor4_1 U28032 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[3]), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[1]), .C(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[4]), .D(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[5]), .Y(n23607) );
  sky130_fd_sc_hd__nand2_1 U28033 ( .A(n23601), .B(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[2]), .Y(n23605) );
  sky130_fd_sc_hd__nand2_1 U28034 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[0]), .B(n23603), .Y(
        n23604) );
  sky130_fd_sc_hd__o22ai_1 U28035 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[0]), .A2(n23605), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_spi_len[2]), .B2(n23604), .Y(
        n23606) );
  sky130_fd_sc_hd__a21oi_1 U28036 ( .A1(n23607), .A2(n23606), .B1(n25529), .Y(
        n23611) );
  sky130_fd_sc_hd__nand4_1 U28037 ( .A(n23611), .B(n23610), .C(n23609), .D(
        n23608), .Y(j202_soc_core_wbqspiflash_00_lldriver_N307) );
  sky130_fd_sc_hd__nor2_1 U28038 ( .A(n23612), .B(
        j202_soc_core_wbqspiflash_00_lldriver_r_spd), .Y(n23743) );
  sky130_fd_sc_hd__a222oi_1 U28039 ( .A1(n23742), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[0]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[0]), .B2(n23743), .C1(
        n23690), .C2(j202_soc_core_wbqspiflash_00_spi_in[1]), .Y(n23613) );
  sky130_fd_sc_hd__a222oi_1 U28040 ( .A1(n23742), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[1]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[1]), .B2(n23743), .C1(
        n23690), .C2(j202_soc_core_wbqspiflash_00_spi_in[2]), .Y(n23614) );
  sky130_fd_sc_hd__clkinv_1 U28041 ( .A(j202_soc_core_wbqspiflash_00_spi_in[3]), .Y(n23624) );
  sky130_fd_sc_hd__a22oi_1 U28042 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[2]), .A2(n23743), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[2]), .B2(n23742), .Y(n23615) );
  sky130_fd_sc_hd__a22oi_1 U28044 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[3]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[0]), .B2(n23732), .Y(
        n23617) );
  sky130_fd_sc_hd__a22oi_1 U28045 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[4]), .B1(n23689), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[0]), .Y(n23616) );
  sky130_fd_sc_hd__o211ai_1 U28046 ( .A1(n23694), .A2(n23624), .B1(n23617), 
        .C1(n23616), .Y(j202_soc_core_wbqspiflash_00_lldriver_N395) );
  sky130_fd_sc_hd__clkinv_1 U28047 ( .A(j202_soc_core_wbqspiflash_00_spi_in[4]), .Y(n23627) );
  sky130_fd_sc_hd__a22oi_1 U28048 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[4]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[1]), .B2(n23732), .Y(
        n23619) );
  sky130_fd_sc_hd__a22oi_1 U28049 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[5]), .B1(n23689), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[1]), .Y(n23618) );
  sky130_fd_sc_hd__o211ai_1 U28050 ( .A1(n23694), .A2(n23627), .B1(n23619), 
        .C1(n23618), .Y(j202_soc_core_wbqspiflash_00_lldriver_N396) );
  sky130_fd_sc_hd__clkinv_1 U28051 ( .A(j202_soc_core_wbqspiflash_00_spi_in[5]), .Y(n23630) );
  sky130_fd_sc_hd__a22oi_1 U28052 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[5]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[2]), .B2(n23732), .Y(
        n23621) );
  sky130_fd_sc_hd__a22oi_1 U28053 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[6]), .B1(n23689), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[2]), .Y(n23620) );
  sky130_fd_sc_hd__o211ai_1 U28054 ( .A1(n23694), .A2(n23630), .B1(n23621), 
        .C1(n23620), .Y(j202_soc_core_wbqspiflash_00_lldriver_N397) );
  sky130_fd_sc_hd__a22oi_1 U28055 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[6]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[3]), .B2(n23732), .Y(
        n23623) );
  sky130_fd_sc_hd__a22oi_1 U28056 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[7]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[6]), .B2(n23742), .Y(n23622) );
  sky130_fd_sc_hd__o211ai_1 U28057 ( .A1(n23624), .A2(n23738), .B1(n23623), 
        .C1(n23622), .Y(j202_soc_core_wbqspiflash_00_lldriver_N398) );
  sky130_fd_sc_hd__a22oi_1 U28058 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[7]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[4]), .B2(n23732), .Y(
        n23626) );
  sky130_fd_sc_hd__a22oi_1 U28059 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[8]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[7]), .B2(n23742), .Y(n23625) );
  sky130_fd_sc_hd__o211ai_1 U28060 ( .A1(n23627), .A2(n23738), .B1(n23626), 
        .C1(n23625), .Y(j202_soc_core_wbqspiflash_00_lldriver_N399) );
  sky130_fd_sc_hd__a22oi_1 U28061 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[8]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[5]), .B2(n23732), .Y(
        n23629) );
  sky130_fd_sc_hd__a22oi_1 U28062 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[9]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[8]), .B2(n23742), .Y(n23628) );
  sky130_fd_sc_hd__o211ai_1 U28063 ( .A1(n23738), .A2(n23630), .B1(n23629), 
        .C1(n23628), .Y(j202_soc_core_wbqspiflash_00_lldriver_N400) );
  sky130_fd_sc_hd__a22oi_1 U28064 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[9]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[6]), .B2(n23732), .Y(
        n23633) );
  sky130_fd_sc_hd__a22oi_1 U28065 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[10]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[9]), .B2(n23742), .Y(n23632) );
  sky130_fd_sc_hd__nand2_1 U28066 ( .A(n23689), .B(
        j202_soc_core_wbqspiflash_00_spi_in[6]), .Y(n23631) );
  sky130_fd_sc_hd__nand3_1 U28067 ( .A(n23633), .B(n23632), .C(n23631), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N401) );
  sky130_fd_sc_hd__a22oi_1 U28068 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[10]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[7]), .B2(n23732), .Y(
        n23636) );
  sky130_fd_sc_hd__a22oi_1 U28069 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[11]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[10]), .B2(n23742), .Y(n23635) );
  sky130_fd_sc_hd__nand2_1 U28070 ( .A(n23689), .B(
        j202_soc_core_wbqspiflash_00_spi_in[7]), .Y(n23634) );
  sky130_fd_sc_hd__nand3_1 U28071 ( .A(n23636), .B(n23635), .C(n23634), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N402) );
  sky130_fd_sc_hd__a22oi_1 U28072 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[11]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[8]), .B2(n23732), .Y(
        n23639) );
  sky130_fd_sc_hd__a22oi_1 U28073 ( .A1(j202_soc_core_wbqspiflash_00_spi_in[8]), .A2(n23689), .B1(j202_soc_core_wbqspiflash_00_spi_in[11]), .B2(n23742), .Y(
        n23638) );
  sky130_fd_sc_hd__nand2_1 U28074 ( .A(n23690), .B(
        j202_soc_core_wbqspiflash_00_spi_in[12]), .Y(n23637) );
  sky130_fd_sc_hd__nand3_1 U28075 ( .A(n23639), .B(n23638), .C(n23637), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N403) );
  sky130_fd_sc_hd__a22oi_1 U28076 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[12]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[9]), .B2(n23732), .Y(
        n23642) );
  sky130_fd_sc_hd__a22oi_1 U28077 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[13]), .B1(n23689), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[9]), .Y(n23641) );
  sky130_fd_sc_hd__nand2_1 U28078 ( .A(j202_soc_core_wbqspiflash_00_spi_in[12]), .B(n23742), .Y(n23640) );
  sky130_fd_sc_hd__nand3_1 U28079 ( .A(n23642), .B(n23641), .C(n23640), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N404) );
  sky130_fd_sc_hd__a22oi_1 U28080 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[13]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[10]), .B2(n23732), .Y(
        n23645) );
  sky130_fd_sc_hd__a22oi_1 U28081 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_in[10]), .A2(n23689), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[13]), .B2(n23742), .Y(n23644) );
  sky130_fd_sc_hd__nand2_1 U28082 ( .A(n23690), .B(
        j202_soc_core_wbqspiflash_00_spi_in[14]), .Y(n23643) );
  sky130_fd_sc_hd__nand3_1 U28083 ( .A(n23645), .B(n23644), .C(n23643), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N405) );
  sky130_fd_sc_hd__a22oi_1 U28084 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[14]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[11]), .B2(n23732), .Y(
        n23648) );
  sky130_fd_sc_hd__a22oi_1 U28085 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[15]), .B1(n23689), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[11]), .Y(n23647) );
  sky130_fd_sc_hd__nand2_1 U28086 ( .A(j202_soc_core_wbqspiflash_00_spi_in[14]), .B(n23742), .Y(n23646) );
  sky130_fd_sc_hd__nand3_1 U28087 ( .A(n23648), .B(n23647), .C(n23646), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N406) );
  sky130_fd_sc_hd__a22oi_1 U28088 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[15]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[12]), .B2(n23732), .Y(
        n23651) );
  sky130_fd_sc_hd__a22oi_1 U28089 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[16]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[15]), .B2(n23742), .Y(n23650) );
  sky130_fd_sc_hd__nand2_1 U28090 ( .A(n23689), .B(
        j202_soc_core_wbqspiflash_00_spi_in[12]), .Y(n23649) );
  sky130_fd_sc_hd__nand3_1 U28091 ( .A(n23651), .B(n23650), .C(n23649), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N407) );
  sky130_fd_sc_hd__a22oi_1 U28092 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[16]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[13]), .B2(n23732), .Y(
        n23654) );
  sky130_fd_sc_hd__a22oi_1 U28093 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[17]), .B1(n23689), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[13]), .Y(n23653) );
  sky130_fd_sc_hd__nand2_1 U28094 ( .A(j202_soc_core_wbqspiflash_00_spi_in[16]), .B(n23742), .Y(n23652) );
  sky130_fd_sc_hd__nand3_1 U28095 ( .A(n23654), .B(n23653), .C(n23652), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N408) );
  sky130_fd_sc_hd__a22oi_1 U28096 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[17]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[14]), .B2(n23732), .Y(
        n23657) );
  sky130_fd_sc_hd__a22oi_1 U28097 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_in[14]), .A2(n23689), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[17]), .B2(n23742), .Y(n23656) );
  sky130_fd_sc_hd__nand2_1 U28098 ( .A(n23690), .B(
        j202_soc_core_wbqspiflash_00_spi_in[18]), .Y(n23655) );
  sky130_fd_sc_hd__nand3_1 U28099 ( .A(n23657), .B(n23656), .C(n23655), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N409) );
  sky130_fd_sc_hd__a22oi_1 U28100 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[18]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[15]), .B2(n23732), .Y(
        n23660) );
  sky130_fd_sc_hd__a22oi_1 U28101 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[19]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[18]), .B2(n23742), .Y(n23659) );
  sky130_fd_sc_hd__nand2_1 U28102 ( .A(n23689), .B(
        j202_soc_core_wbqspiflash_00_spi_in[15]), .Y(n23658) );
  sky130_fd_sc_hd__nand3_1 U28103 ( .A(n23660), .B(n23659), .C(n23658), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N410) );
  sky130_fd_sc_hd__a22oi_1 U28104 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[19]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[16]), .B2(n23732), .Y(
        n23663) );
  sky130_fd_sc_hd__a22oi_1 U28105 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_in[16]), .A2(n23689), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[19]), .B2(n23742), .Y(n23662) );
  sky130_fd_sc_hd__nand2_1 U28106 ( .A(n23690), .B(
        j202_soc_core_wbqspiflash_00_spi_in[20]), .Y(n23661) );
  sky130_fd_sc_hd__nand3_1 U28107 ( .A(n23663), .B(n23662), .C(n23661), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N411) );
  sky130_fd_sc_hd__a22oi_1 U28108 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[20]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[17]), .B2(n23732), .Y(
        n23666) );
  sky130_fd_sc_hd__a22oi_1 U28109 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[21]), .B1(n23689), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[17]), .Y(n23665) );
  sky130_fd_sc_hd__nand2_1 U28110 ( .A(j202_soc_core_wbqspiflash_00_spi_in[20]), .B(n23742), .Y(n23664) );
  sky130_fd_sc_hd__nand3_1 U28111 ( .A(n23666), .B(n23665), .C(n23664), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N412) );
  sky130_fd_sc_hd__a22oi_1 U28112 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[21]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[18]), .B2(n23732), .Y(
        n23669) );
  sky130_fd_sc_hd__a22oi_1 U28113 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[22]), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[21]), .B2(n23742), .Y(n23668) );
  sky130_fd_sc_hd__nand2_1 U28114 ( .A(n23689), .B(
        j202_soc_core_wbqspiflash_00_spi_in[18]), .Y(n23667) );
  sky130_fd_sc_hd__nand3_1 U28115 ( .A(n23669), .B(n23668), .C(n23667), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N413) );
  sky130_fd_sc_hd__a22oi_1 U28116 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[22]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[19]), .B2(n23732), .Y(
        n23672) );
  sky130_fd_sc_hd__a22oi_1 U28117 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_in[19]), .A2(n23689), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[22]), .B2(n23742), .Y(n23671) );
  sky130_fd_sc_hd__nand2_1 U28118 ( .A(n23690), .B(
        j202_soc_core_wbqspiflash_00_spi_in[23]), .Y(n23670) );
  sky130_fd_sc_hd__nand3_1 U28119 ( .A(n23672), .B(n23671), .C(n23670), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N414) );
  sky130_fd_sc_hd__a22oi_1 U28120 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[23]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[20]), .B2(n23732), .Y(
        n23675) );
  sky130_fd_sc_hd__a22oi_1 U28121 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_in[20]), .A2(n23689), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[23]), .B2(n23742), .Y(n23674) );
  sky130_fd_sc_hd__nand2_1 U28122 ( .A(n23690), .B(
        j202_soc_core_wbqspiflash_00_spi_in[24]), .Y(n23673) );
  sky130_fd_sc_hd__nand3_1 U28123 ( .A(n23675), .B(n23674), .C(n23673), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N415) );
  sky130_fd_sc_hd__a22oi_1 U28124 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[24]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[21]), .B2(n23732), .Y(
        n23678) );
  sky130_fd_sc_hd__a22oi_1 U28125 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[25]), .B1(n23689), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[21]), .Y(n23677) );
  sky130_fd_sc_hd__nand2_1 U28126 ( .A(j202_soc_core_wbqspiflash_00_spi_in[24]), .B(n23742), .Y(n23676) );
  sky130_fd_sc_hd__nand3_1 U28127 ( .A(n23678), .B(n23677), .C(n23676), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N416) );
  sky130_fd_sc_hd__a22oi_1 U28128 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[25]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[22]), .B2(n23732), .Y(
        n23681) );
  sky130_fd_sc_hd__a22oi_1 U28129 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[26]), .B1(n23689), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[22]), .Y(n23680) );
  sky130_fd_sc_hd__nand2_1 U28130 ( .A(j202_soc_core_wbqspiflash_00_spi_in[25]), .B(n23742), .Y(n23679) );
  sky130_fd_sc_hd__nand3_1 U28131 ( .A(n23681), .B(n23680), .C(n23679), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N417) );
  sky130_fd_sc_hd__a22oi_1 U28132 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[26]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[23]), .B2(n23732), .Y(
        n23684) );
  sky130_fd_sc_hd__a22oi_1 U28133 ( .A1(n23690), .A2(
        j202_soc_core_wbqspiflash_00_spi_in[27]), .B1(n23689), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[23]), .Y(n23683) );
  sky130_fd_sc_hd__nand2_1 U28134 ( .A(j202_soc_core_wbqspiflash_00_spi_in[26]), .B(n23742), .Y(n23682) );
  sky130_fd_sc_hd__nand3_1 U28135 ( .A(n23684), .B(n23683), .C(n23682), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N418) );
  sky130_fd_sc_hd__clkinv_1 U28136 ( .A(
        j202_soc_core_wbqspiflash_00_spi_in[28]), .Y(n23739) );
  sky130_fd_sc_hd__a22oi_1 U28137 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[27]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[24]), .B2(n23732), .Y(
        n23686) );
  sky130_fd_sc_hd__a22oi_1 U28138 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_in[24]), .A2(n23689), .B1(
        j202_soc_core_wbqspiflash_00_spi_in[27]), .B2(n23742), .Y(n23685) );
  sky130_fd_sc_hd__o211ai_1 U28139 ( .A1(n23739), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B1(n23686), .C1(n23685), 
        .Y(j202_soc_core_wbqspiflash_00_lldriver_N419) );
  sky130_fd_sc_hd__a22oi_1 U28140 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[28]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[25]), .B2(n23732), .Y(
        n23688) );
  sky130_fd_sc_hd__a22oi_1 U28141 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_in[29]), .A2(n23690), .B1(n23689), 
        .B2(j202_soc_core_wbqspiflash_00_spi_in[25]), .Y(n23687) );
  sky130_fd_sc_hd__o211ai_1 U28142 ( .A1(n23694), .A2(n23739), .B1(n23688), 
        .C1(n23687), .Y(j202_soc_core_wbqspiflash_00_lldriver_N420) );
  sky130_fd_sc_hd__a22oi_1 U28143 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[29]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[26]), .B2(n23732), .Y(
        n23692) );
  sky130_fd_sc_hd__a22oi_1 U28144 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_in[30]), .A2(n23690), .B1(n23689), 
        .B2(j202_soc_core_wbqspiflash_00_spi_in[26]), .Y(n23691) );
  sky130_fd_sc_hd__o211ai_1 U28145 ( .A1(n23694), .A2(n23693), .B1(n23692), 
        .C1(n23691), .Y(j202_soc_core_wbqspiflash_00_lldriver_N421) );
  sky130_fd_sc_hd__a22oi_1 U28146 ( .A1(n23743), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[30]), .B1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[27]), .B2(n23732), .Y(
        n23696) );
  sky130_fd_sc_hd__o221ai_1 U28147 ( .A1(j202_soc_core_wbqspiflash_00_spi_spd), 
        .A2(j202_soc_core_wbqspiflash_00_spi_in[30]), .B1(n23735), .B2(
        j202_soc_core_wbqspiflash_00_spi_in[27]), .C1(n23740), .Y(n23695) );
  sky130_fd_sc_hd__o211ai_1 U28148 ( .A1(n23733), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B1(n23696), .C1(n23695), 
        .Y(j202_soc_core_wbqspiflash_00_lldriver_N422) );
  sky130_fd_sc_hd__o22ai_1 U28149 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(io_in[11]), .B1(
        n24784), .B2(io_in[10]), .Y(n23700) );
  sky130_fd_sc_hd__nor2_1 U28150 ( .A(n23700), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N358) );
  sky130_fd_sc_hd__o22ai_1 U28151 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[0]), .B1(n24784), .B2(
        io_in[11]), .Y(n23701) );
  sky130_fd_sc_hd__nor2_1 U28152 ( .A(n23701), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N359) );
  sky130_fd_sc_hd__o22ai_1 U28153 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[1]), .B1(n24784), .B2(
        io_in[12]), .Y(n23702) );
  sky130_fd_sc_hd__nor2_1 U28154 ( .A(n23702), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N360) );
  sky130_fd_sc_hd__o22ai_1 U28155 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[2]), .B1(n24784), .B2(
        io_in[13]), .Y(n23703) );
  sky130_fd_sc_hd__nor2_1 U28156 ( .A(n23703), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N361) );
  sky130_fd_sc_hd__o22ai_1 U28157 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[3]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[0]), .Y(n23704) );
  sky130_fd_sc_hd__nor2_1 U28158 ( .A(n23704), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N362) );
  sky130_fd_sc_hd__o22ai_1 U28159 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[4]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[1]), .Y(n23705) );
  sky130_fd_sc_hd__nor2_1 U28160 ( .A(n23705), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N363) );
  sky130_fd_sc_hd__o22ai_1 U28161 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[5]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[2]), .Y(n23706) );
  sky130_fd_sc_hd__nor2_1 U28162 ( .A(n23706), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N364) );
  sky130_fd_sc_hd__o22ai_1 U28163 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[6]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[3]), .Y(n23707) );
  sky130_fd_sc_hd__nor2_1 U28164 ( .A(n23707), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N365) );
  sky130_fd_sc_hd__o22ai_1 U28165 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[7]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[4]), .Y(n23708) );
  sky130_fd_sc_hd__nor2_1 U28166 ( .A(n23708), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N366) );
  sky130_fd_sc_hd__o22ai_1 U28167 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[8]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[5]), .Y(n23709) );
  sky130_fd_sc_hd__nor2_1 U28168 ( .A(n23709), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N367) );
  sky130_fd_sc_hd__o22ai_1 U28169 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[9]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[6]), .Y(n23710) );
  sky130_fd_sc_hd__nor2_1 U28170 ( .A(n23710), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N368) );
  sky130_fd_sc_hd__o22ai_1 U28171 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[10]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[7]), .Y(n23711) );
  sky130_fd_sc_hd__nor2_1 U28172 ( .A(n23711), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N369) );
  sky130_fd_sc_hd__o22ai_1 U28173 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[11]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[8]), .Y(n23712) );
  sky130_fd_sc_hd__nor2_1 U28174 ( .A(n23712), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N370) );
  sky130_fd_sc_hd__o22ai_1 U28175 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[12]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[9]), .Y(n23713) );
  sky130_fd_sc_hd__nor3_1 U28176 ( .A(n23731), .B(n23697), .C(n23713), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N371) );
  sky130_fd_sc_hd__o22ai_1 U28177 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[13]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[10]), .Y(n23714) );
  sky130_fd_sc_hd__nor3_1 U28178 ( .A(n23731), .B(n23697), .C(n23714), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N372) );
  sky130_fd_sc_hd__o22ai_1 U28179 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[14]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[11]), .Y(n23715) );
  sky130_fd_sc_hd__nor2_1 U28180 ( .A(n23715), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N373) );
  sky130_fd_sc_hd__o22ai_1 U28181 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[15]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[12]), .Y(n23716) );
  sky130_fd_sc_hd__nor2_1 U28182 ( .A(n23716), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N374) );
  sky130_fd_sc_hd__o22ai_1 U28183 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[16]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[13]), .Y(n23717) );
  sky130_fd_sc_hd__nor2_1 U28184 ( .A(n23717), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N375) );
  sky130_fd_sc_hd__o22ai_1 U28185 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[17]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[14]), .Y(n23718) );
  sky130_fd_sc_hd__nor2_1 U28186 ( .A(n23718), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N376) );
  sky130_fd_sc_hd__o22ai_1 U28187 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[18]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[15]), .Y(n23719) );
  sky130_fd_sc_hd__nor2_1 U28188 ( .A(n23719), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N377) );
  sky130_fd_sc_hd__o22ai_1 U28189 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[19]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[16]), .Y(n23720) );
  sky130_fd_sc_hd__nor2_1 U28190 ( .A(n23720), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N378) );
  sky130_fd_sc_hd__o22ai_1 U28191 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[20]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[17]), .Y(n23721) );
  sky130_fd_sc_hd__nor3_1 U28192 ( .A(n23731), .B(n23697), .C(n23721), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N379) );
  sky130_fd_sc_hd__o22ai_1 U28193 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[21]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[18]), .Y(n23722) );
  sky130_fd_sc_hd__nor3_1 U28194 ( .A(n23731), .B(n23697), .C(n23722), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N380) );
  sky130_fd_sc_hd__o22ai_1 U28195 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[22]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[19]), .Y(n23723) );
  sky130_fd_sc_hd__nor2_1 U28196 ( .A(n23723), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N381) );
  sky130_fd_sc_hd__o22ai_1 U28197 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[23]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[20]), .Y(n23724) );
  sky130_fd_sc_hd__nor2_1 U28198 ( .A(n23724), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N382) );
  sky130_fd_sc_hd__o22ai_1 U28199 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[24]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[21]), .Y(n23725) );
  sky130_fd_sc_hd__nor2_1 U28200 ( .A(n23725), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N383) );
  sky130_fd_sc_hd__o22ai_1 U28201 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[25]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[22]), .Y(n23726) );
  sky130_fd_sc_hd__nor2_1 U28202 ( .A(n23726), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N384) );
  sky130_fd_sc_hd__o22ai_1 U28203 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[26]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[23]), .Y(n23727) );
  sky130_fd_sc_hd__nor2_1 U28204 ( .A(n23727), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N385) );
  sky130_fd_sc_hd__o22ai_1 U28205 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[27]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[24]), .Y(n23728) );
  sky130_fd_sc_hd__nor2_1 U28206 ( .A(n23728), .B(n23699), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N386) );
  sky130_fd_sc_hd__o22ai_1 U28207 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[28]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[25]), .Y(n23729) );
  sky130_fd_sc_hd__nor3_1 U28208 ( .A(n23731), .B(n23697), .C(n23729), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N387) );
  sky130_fd_sc_hd__o22ai_1 U28209 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[29]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[26]), .Y(n23730) );
  sky130_fd_sc_hd__nor3_1 U28210 ( .A(n23731), .B(n23697), .C(n23730), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N388) );
  sky130_fd_sc_hd__o22ai_1 U28211 ( .A1(
        j202_soc_core_wbqspiflash_00_w_qspi_mod[1]), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[30]), .B1(n24784), .B2(
        j202_soc_core_wbqspiflash_00_lldriver_r_input[27]), .Y(n23698) );
  sky130_fd_sc_hd__nor2_1 U28212 ( .A(n23699), .B(n23698), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N389) );
  sky130_fd_sc_hd__nor2_1 U28213 ( .A(n23700), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N323) );
  sky130_fd_sc_hd__nor2_1 U28214 ( .A(n23701), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N324) );
  sky130_fd_sc_hd__nor2_1 U28215 ( .A(n23702), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N325) );
  sky130_fd_sc_hd__nor2_1 U28216 ( .A(n23703), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N326) );
  sky130_fd_sc_hd__nor2_1 U28217 ( .A(n23704), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N327) );
  sky130_fd_sc_hd__nor2_1 U28218 ( .A(n23705), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N328) );
  sky130_fd_sc_hd__nor2_1 U28219 ( .A(n23706), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N329) );
  sky130_fd_sc_hd__nor2_1 U28220 ( .A(n23707), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N330) );
  sky130_fd_sc_hd__nor2_1 U28221 ( .A(n23708), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N331) );
  sky130_fd_sc_hd__nor2_1 U28222 ( .A(n23709), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N332) );
  sky130_fd_sc_hd__nor2_1 U28223 ( .A(n23710), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N333) );
  sky130_fd_sc_hd__nor2_1 U28224 ( .A(n23711), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N334) );
  sky130_fd_sc_hd__nor2_1 U28225 ( .A(n23712), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N335) );
  sky130_fd_sc_hd__nor2_1 U28226 ( .A(n23731), .B(n23713), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N336) );
  sky130_fd_sc_hd__nor2_1 U28227 ( .A(n23731), .B(n23714), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N337) );
  sky130_fd_sc_hd__nor2_1 U28228 ( .A(n23715), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N338) );
  sky130_fd_sc_hd__nor2_1 U28229 ( .A(n23716), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N339) );
  sky130_fd_sc_hd__nor2_1 U28230 ( .A(n23717), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N340) );
  sky130_fd_sc_hd__nor2_1 U28231 ( .A(n23718), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N341) );
  sky130_fd_sc_hd__nor2_1 U28232 ( .A(n23719), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N342) );
  sky130_fd_sc_hd__nor2_1 U28233 ( .A(n23720), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N343) );
  sky130_fd_sc_hd__nor2_1 U28234 ( .A(n23731), .B(n23721), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N344) );
  sky130_fd_sc_hd__nor2_1 U28235 ( .A(n23731), .B(n23722), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N345) );
  sky130_fd_sc_hd__nor2_1 U28236 ( .A(n23723), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N346) );
  sky130_fd_sc_hd__nor2_1 U28237 ( .A(n23724), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N347) );
  sky130_fd_sc_hd__nor2_1 U28238 ( .A(n23725), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N348) );
  sky130_fd_sc_hd__nor2_1 U28239 ( .A(n23726), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N349) );
  sky130_fd_sc_hd__nor2_1 U28240 ( .A(n23727), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N350) );
  sky130_fd_sc_hd__nor2_1 U28241 ( .A(n23728), .B(n23731), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N351) );
  sky130_fd_sc_hd__nor2_1 U28242 ( .A(n23731), .B(n23729), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N352) );
  sky130_fd_sc_hd__nor2_1 U28243 ( .A(n23731), .B(n23730), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N353) );
  sky130_fd_sc_hd__a21oi_1 U28244 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[28]), .A2(n23732), .B1(
        n23741), .Y(n23737) );
  sky130_fd_sc_hd__nor2_1 U28245 ( .A(n23734), .B(n23733), .Y(n23746) );
  sky130_fd_sc_hd__a22oi_1 U28246 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[31]), .A2(n23743), .B1(
        n23746), .B2(n23735), .Y(n23736) );
  sky130_fd_sc_hd__o211ai_1 U28247 ( .A1(n23739), .A2(n23738), .B1(n23737), 
        .C1(n23736), .Y(j202_soc_core_wbqspiflash_00_lldriver_N316) );
  sky130_fd_sc_hd__nand2_1 U28248 ( .A(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[30]), .B(n23747), .Y(
        n23745) );
  sky130_fd_sc_hd__nand2_1 U28249 ( .A(j202_soc_core_wbqspiflash_00_spi_in[30]), .B(n23740), .Y(n23744) );
  sky130_fd_sc_hd__nor3_1 U28250 ( .A(n23743), .B(n23742), .C(n23741), .Y(
        n23749) );
  sky130_fd_sc_hd__nand3_1 U28251 ( .A(n23745), .B(n23744), .C(n23749), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N318) );
  sky130_fd_sc_hd__a21oi_1 U28252 ( .A1(n23747), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_r_word[31]), .B1(n23746), .Y(
        n23748) );
  sky130_fd_sc_hd__nand2_1 U28253 ( .A(n23749), .B(n23748), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N319) );
  sky130_fd_sc_hd__nand4_1 U28254 ( .A(n23751), .B(n23753), .C(n23750), .D(
        n23752), .Y(j202_soc_core_wbqspiflash_00_lldriver_N312) );
  sky130_fd_sc_hd__nand2_1 U28255 ( .A(n23753), .B(n23752), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N310) );
  sky130_fd_sc_hd__a211oi_1 U28256 ( .A1(n23787), .A2(n23757), .B1(n23754), 
        .C1(n23761), .Y(n23755) );
  sky130_fd_sc_hd__nor2_1 U28257 ( .A(n23755), .B(n23792), .Y(
        j202_soc_core_wbqspiflash_00_N667) );
  sky130_fd_sc_hd__clkinv_1 U28258 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[1]), .Y(n23794) );
  sky130_fd_sc_hd__nor2_1 U28259 ( .A(n23755), .B(n23794), .Y(
        j202_soc_core_wbqspiflash_00_N668) );
  sky130_fd_sc_hd__clkinv_1 U28260 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[2]), .Y(n23796) );
  sky130_fd_sc_hd__nor2_1 U28261 ( .A(n23755), .B(n23796), .Y(
        j202_soc_core_wbqspiflash_00_N669) );
  sky130_fd_sc_hd__clkinv_1 U28262 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[3]), .Y(n23797) );
  sky130_fd_sc_hd__nor2_1 U28263 ( .A(n23755), .B(n23797), .Y(
        j202_soc_core_wbqspiflash_00_N670) );
  sky130_fd_sc_hd__clkinv_1 U28264 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[4]), .Y(n23798) );
  sky130_fd_sc_hd__nor2_1 U28265 ( .A(n23755), .B(n23798), .Y(
        j202_soc_core_wbqspiflash_00_N671) );
  sky130_fd_sc_hd__clkinv_1 U28266 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[5]), .Y(n23790) );
  sky130_fd_sc_hd__nor2_1 U28267 ( .A(n23755), .B(n23790), .Y(
        j202_soc_core_wbqspiflash_00_N672) );
  sky130_fd_sc_hd__clkinv_1 U28268 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[6]), .Y(n23791) );
  sky130_fd_sc_hd__nor2_1 U28269 ( .A(n23755), .B(n23791), .Y(
        j202_soc_core_wbqspiflash_00_N673) );
  sky130_fd_sc_hd__clkinv_1 U28270 ( .A(
        j202_soc_core_wbqspiflash_00_spi_out[7]), .Y(n23799) );
  sky130_fd_sc_hd__nor2_1 U28271 ( .A(n23755), .B(n23799), .Y(
        j202_soc_core_wbqspiflash_00_N674) );
  sky130_fd_sc_hd__a22o_1 U28273 ( .A1(
        j202_soc_core_wbqspiflash_00_erased_sector[0]), .A2(n23759), .B1(
        j202_soc_core_wbqspiflash_00_spi_out[14]), .B2(n23761), .X(
        j202_soc_core_wbqspiflash_00_N681) );
  sky130_fd_sc_hd__a22o_1 U28274 ( .A1(
        j202_soc_core_wbqspiflash_00_erased_sector[1]), .A2(n23759), .B1(
        j202_soc_core_wbqspiflash_00_spi_out[15]), .B2(n23761), .X(
        j202_soc_core_wbqspiflash_00_N682) );
  sky130_fd_sc_hd__a22o_1 U28275 ( .A1(
        j202_soc_core_wbqspiflash_00_erased_sector[2]), .A2(n23759), .B1(
        j202_soc_core_wbqspiflash_00_spi_out[16]), .B2(n23761), .X(
        j202_soc_core_wbqspiflash_00_N683) );
  sky130_fd_sc_hd__a22o_1 U28276 ( .A1(
        j202_soc_core_wbqspiflash_00_erased_sector[3]), .A2(n23759), .B1(
        j202_soc_core_wbqspiflash_00_spi_out[17]), .B2(n23761), .X(
        j202_soc_core_wbqspiflash_00_N684) );
  sky130_fd_sc_hd__a22o_1 U28277 ( .A1(
        j202_soc_core_wbqspiflash_00_erased_sector[4]), .A2(n23759), .B1(
        j202_soc_core_wbqspiflash_00_spi_out[18]), .B2(n23761), .X(
        j202_soc_core_wbqspiflash_00_N685) );
  sky130_fd_sc_hd__a22o_1 U28278 ( .A1(
        j202_soc_core_wbqspiflash_00_erased_sector[5]), .A2(n23759), .B1(
        j202_soc_core_wbqspiflash_00_spi_out[19]), .B2(n23761), .X(
        j202_soc_core_wbqspiflash_00_N686) );
  sky130_fd_sc_hd__a22o_1 U28279 ( .A1(
        j202_soc_core_wbqspiflash_00_erased_sector[6]), .A2(n23759), .B1(
        j202_soc_core_wbqspiflash_00_spi_out[20]), .B2(n23761), .X(
        j202_soc_core_wbqspiflash_00_N687) );
  sky130_fd_sc_hd__a22o_1 U28280 ( .A1(
        j202_soc_core_wbqspiflash_00_erased_sector[7]), .A2(n23759), .B1(
        j202_soc_core_wbqspiflash_00_spi_out[21]), .B2(n23761), .X(
        j202_soc_core_wbqspiflash_00_N688) );
  sky130_fd_sc_hd__a22o_1 U28281 ( .A1(
        j202_soc_core_wbqspiflash_00_quad_mode_enabled), .A2(n23759), .B1(
        j202_soc_core_wbqspiflash_00_spi_out[27]), .B2(n23761), .X(
        j202_soc_core_wbqspiflash_00_N694) );
  sky130_fd_sc_hd__a22o_1 U28282 ( .A1(
        j202_soc_core_wbqspiflash_00_spi_out[28]), .A2(n23761), .B1(n23758), 
        .B2(n23759), .X(j202_soc_core_wbqspiflash_00_N695) );
  sky130_fd_sc_hd__a22o_1 U28283 ( .A1(j202_soc_core_wbqspiflash_00_spi_busy), 
        .A2(n23759), .B1(j202_soc_core_wbqspiflash_00_spi_out[29]), .B2(n23761), .X(j202_soc_core_wbqspiflash_00_N696) );
  sky130_fd_sc_hd__a22o_1 U28284 ( .A1(
        j202_soc_core_wbqspiflash_00_dirty_sector), .A2(n23759), .B1(
        j202_soc_core_wbqspiflash_00_spi_out[30]), .B2(n23761), .X(
        j202_soc_core_wbqspiflash_00_N697) );
  sky130_fd_sc_hd__nand2_1 U28285 ( .A(n23760), .B(n23787), .Y(n23764) );
  sky130_fd_sc_hd__a22oi_1 U28286 ( .A1(
        j202_soc_core_wbqspiflash_00_write_in_progress), .A2(n23762), .B1(
        j202_soc_core_wbqspiflash_00_spi_out[31]), .B2(n23761), .Y(n23763) );
  sky130_fd_sc_hd__nor2_1 U28288 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[0]), .B(n25002), .Y(
        j202_soc_core_wbqspiflash_00_N614) );
  sky130_fd_sc_hd__nor2_1 U28289 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[0]), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[1]), .Y(n23765) );
  sky130_fd_sc_hd__a21oi_1 U28290 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[0]), .A2(
        j202_soc_core_wbqspiflash_00_reset_counter[1]), .B1(n23765), .Y(n23766) );
  sky130_fd_sc_hd__nor2_1 U28291 ( .A(n25002), .B(n23766), .Y(
        j202_soc_core_wbqspiflash_00_N615) );
  sky130_fd_sc_hd__clkinv_1 U28292 ( .A(n23767), .Y(n23769) );
  sky130_fd_sc_hd__o21ai_1 U28293 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[0]), .A2(
        j202_soc_core_wbqspiflash_00_reset_counter[1]), .B1(
        j202_soc_core_wbqspiflash_00_reset_counter[2]), .Y(n23768) );
  sky130_fd_sc_hd__a31oi_1 U28294 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), 
        .A2(n23769), .A3(n23768), .B1(n23784), .Y(
        j202_soc_core_wbqspiflash_00_N616) );
  sky130_fd_sc_hd__a21oi_1 U28295 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[3]), .A2(n23769), .B1(
        n25070), .Y(n23770) );
  sky130_fd_sc_hd__a21oi_1 U28296 ( .A1(n23770), .A2(n23771), .B1(n23784), .Y(
        j202_soc_core_wbqspiflash_00_N617) );
  sky130_fd_sc_hd__a21oi_1 U28297 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[4]), .A2(n23771), .B1(
        n23773), .Y(n23772) );
  sky130_fd_sc_hd__a21oi_1 U28298 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), 
        .A2(n23772), .B1(n23784), .Y(j202_soc_core_wbqspiflash_00_N618) );
  sky130_fd_sc_hd__clkinv_1 U28299 ( .A(n23773), .Y(n23774) );
  sky130_fd_sc_hd__a21oi_1 U28300 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[5]), .A2(n23774), .B1(
        n25070), .Y(n23775) );
  sky130_fd_sc_hd__a21oi_1 U28301 ( .A1(n23775), .A2(n23776), .B1(n23784), .Y(
        j202_soc_core_wbqspiflash_00_N619) );
  sky130_fd_sc_hd__a21oi_1 U28302 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[6]), .A2(n23776), .B1(
        n23778), .Y(n23777) );
  sky130_fd_sc_hd__a21oi_1 U28303 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), 
        .A2(n23777), .B1(n23784), .Y(j202_soc_core_wbqspiflash_00_N620) );
  sky130_fd_sc_hd__clkinv_1 U28304 ( .A(n23778), .Y(n23779) );
  sky130_fd_sc_hd__a21oi_1 U28305 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[7]), .A2(n23779), .B1(
        n25070), .Y(n23780) );
  sky130_fd_sc_hd__a21oi_1 U28306 ( .A1(n23780), .A2(n23781), .B1(n23784), .Y(
        j202_soc_core_wbqspiflash_00_N621) );
  sky130_fd_sc_hd__a21oi_1 U28307 ( .A1(
        j202_soc_core_wbqspiflash_00_reset_counter[8]), .A2(n23781), .B1(
        n23783), .Y(n23782) );
  sky130_fd_sc_hd__a21oi_1 U28308 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), 
        .A2(n23782), .B1(n23784), .Y(j202_soc_core_wbqspiflash_00_N622) );
  sky130_fd_sc_hd__o21a_1 U28309 ( .A1(n23801), .A2(n23783), .B1(
        j202_soc_core_wbqspiflash_00_state[0]), .X(n23786) );
  sky130_fd_sc_hd__a21oi_1 U28310 ( .A1(n23786), .A2(n23785), .B1(n23784), .Y(
        j202_soc_core_wbqspiflash_00_N623) );
  sky130_fd_sc_hd__a21oi_1 U28311 ( .A1(n23789), .A2(n23788), .B1(n23787), .Y(
        n23800) );
  sky130_fd_sc_hd__nand2_1 U28312 ( .A(n24954), .B(
        j202_soc_core_wbqspiflash_00_spif_data[5]), .Y(n24977) );
  sky130_fd_sc_hd__o21ai_1 U28313 ( .A1(n23800), .A2(n23790), .B1(n24977), .Y(
        j202_soc_core_wbqspiflash_00_N611) );
  sky130_fd_sc_hd__nand2_1 U28314 ( .A(n24954), .B(
        j202_soc_core_wbqspiflash_00_spif_data[6]), .Y(n24982) );
  sky130_fd_sc_hd__o21ai_1 U28315 ( .A1(n23800), .A2(n23791), .B1(n24982), .Y(
        j202_soc_core_wbqspiflash_00_N612) );
  sky130_fd_sc_hd__o22ai_1 U28316 ( .A1(n23800), .A2(n23792), .B1(n24960), 
        .B2(n24938), .Y(j202_soc_core_wbqspiflash_00_N605) );
  sky130_fd_sc_hd__o22ai_1 U28317 ( .A1(n23800), .A2(n23794), .B1(n24960), 
        .B2(n23793), .Y(j202_soc_core_wbqspiflash_00_N606) );
  sky130_fd_sc_hd__clkinv_1 U28318 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[2]), .Y(n23795) );
  sky130_fd_sc_hd__o22ai_1 U28319 ( .A1(n23800), .A2(n23796), .B1(n24960), 
        .B2(n23795), .Y(j202_soc_core_wbqspiflash_00_N607) );
  sky130_fd_sc_hd__clkinv_1 U28320 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[3]), .Y(n24959) );
  sky130_fd_sc_hd__o22ai_1 U28321 ( .A1(n23800), .A2(n23797), .B1(n24960), 
        .B2(n24959), .Y(j202_soc_core_wbqspiflash_00_N608) );
  sky130_fd_sc_hd__nand2_1 U28322 ( .A(n24954), .B(
        j202_soc_core_wbqspiflash_00_spif_data[4]), .Y(n24969) );
  sky130_fd_sc_hd__o21ai_1 U28323 ( .A1(n23800), .A2(n23798), .B1(n24969), .Y(
        j202_soc_core_wbqspiflash_00_N609) );
  sky130_fd_sc_hd__nand2_1 U28324 ( .A(n24954), .B(
        j202_soc_core_wbqspiflash_00_spif_data[7]), .Y(n24993) );
  sky130_fd_sc_hd__o21ai_1 U28325 ( .A1(n23800), .A2(n23799), .B1(n24993), .Y(
        j202_soc_core_wbqspiflash_00_N613) );
  sky130_fd_sc_hd__or3_1 U28326 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[8]), .B(
        j202_soc_core_wbqspiflash_00_reset_counter[0]), .C(n23801), .X(
        j202_soc_core_wbqspiflash_00_N86) );
  sky130_fd_sc_hd__nor2_1 U28327 ( .A(
        j202_soc_core_wbqspiflash_00_reset_counter[8]), .B(n23801), .Y(n23803)
         );
  sky130_fd_sc_hd__nand2_1 U28328 ( .A(n23803), .B(n23802), .Y(
        j202_soc_core_wbqspiflash_00_N85) );
  sky130_fd_sc_hd__clkinv_1 U28329 ( .A(j202_soc_core_bldc_core_00_comm[0]), 
        .Y(n25169) );
  sky130_fd_sc_hd__o22ai_1 U28330 ( .A1(j202_soc_core_bldc_core_00_comm[1]), 
        .A2(j202_soc_core_bldc_core_00_comm[0]), .B1(n25161), .B2(n25169), .Y(
        n23808) );
  sky130_fd_sc_hd__nor2_1 U28331 ( .A(n23808), .B(n23805), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posc) );
  sky130_fd_sc_hd__nand2_1 U28332 ( .A(j202_soc_core_bldc_core_00_comm[1]), 
        .B(n25169), .Y(n23806) );
  sky130_fd_sc_hd__nand2_1 U28333 ( .A(j202_soc_core_bldc_core_00_comm[0]), 
        .B(n25161), .Y(n23804) );
  sky130_fd_sc_hd__o22ai_1 U28334 ( .A1(n23806), .A2(n23805), .B1(n23804), 
        .B2(n23807), .Y(j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_negb)
         );
  sky130_fd_sc_hd__o21a_1 U28335 ( .A1(n25398), .A2(n25397), .B1(n23808), .X(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posb) );
  sky130_fd_sc_hd__nor2_1 U28336 ( .A(n23808), .B(n23807), .Y(
        j202_soc_core_bldc_core_00_bldc_pwm_00_nxt_pwm_posa) );
  sky130_fd_sc_hd__nor2_1 U28337 ( .A(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bisr_wen), .B(
        n23809), .Y(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_nxt_bldc_int) );
  sky130_fd_sc_hd__nand2_1 U28338 ( .A(n25400), .B(n25732), .Y(n23810) );
  sky130_fd_sc_hd__a211oi_1 U28339 ( .A1(j202_soc_core_uart_BRG_cnt[0]), .A2(
        j202_soc_core_uart_BRG_cnt[1]), .B1(n25399), .C1(n23810), .Y(
        j202_soc_core_uart_BRG_N57) );
  sky130_fd_sc_hd__nor2_1 U28340 ( .A(j202_soc_core_uart_BRG_cnt[0]), .B(
        n23810), .Y(j202_soc_core_uart_BRG_N56) );
  sky130_fd_sc_hd__nand2b_1 U28341 ( .A_N(n25400), .B(n25734), .Y(
        j202_soc_core_uart_BRG_N55) );
  sky130_fd_sc_hd__nand2_1 U28342 ( .A(n25235), .B(n25234), .Y(n25233) );
  sky130_fd_sc_hd__nor2_1 U28343 ( .A(n25232), .B(n25233), .Y(
        j202_soc_core_uart_TOP_rx_fifo_N30) );
  sky130_fd_sc_hd__nor2_1 U28344 ( .A(j202_soc_core_uart_TOP_rx_fifo_wp[1]), 
        .B(n25231), .Y(j202_soc_core_uart_TOP_rx_fifo_N31) );
  sky130_fd_sc_hd__nor2_1 U28345 ( .A(j202_soc_core_uart_TOP_rx_fifo_wp[1]), 
        .B(n25233), .Y(j202_soc_core_uart_TOP_rx_fifo_N32) );
  sky130_fd_sc_hd__nor2_1 U28346 ( .A(n23812), .B(n25200), .Y(
        j202_soc_core_uart_TOP_tx_fifo_N29) );
  sky130_fd_sc_hd__nand2_1 U28347 ( .A(n25201), .B(n23811), .Y(n23813) );
  sky130_fd_sc_hd__nor2_1 U28348 ( .A(n23812), .B(n23813), .Y(
        j202_soc_core_uart_TOP_tx_fifo_N30) );
  sky130_fd_sc_hd__nor2_1 U28349 ( .A(j202_soc_core_uart_TOP_tx_fifo_wp[1]), 
        .B(n23813), .Y(j202_soc_core_uart_TOP_tx_fifo_N32) );
  sky130_fd_sc_hd__nand3b_1 U28350 ( .A_N(j202_soc_core_uart_sio_ce_x4), .B(
        n23814), .C(n25732), .Y(j202_soc_core_uart_TOP_N101) );
  sky130_fd_sc_hd__nor3_1 U28351 ( .A(j202_soc_core_rst), .B(
        j202_soc_core_uart_TOP_rx_bit_cnt[0]), .C(n23821), .Y(
        j202_soc_core_uart_TOP_N86) );
  sky130_fd_sc_hd__a21oi_1 U28352 ( .A1(j202_soc_core_uart_TOP_rx_bit_cnt[1]), 
        .A2(n23816), .B1(n23815), .Y(n23817) );
  sky130_fd_sc_hd__o21ai_1 U28353 ( .A1(n23817), .A2(n23821), .B1(n25734), .Y(
        j202_soc_core_uart_TOP_N87) );
  sky130_fd_sc_hd__and3_1 U28354 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[2]), 
        .B(j202_soc_core_uart_TOP_rx_bit_cnt[1]), .C(
        j202_soc_core_uart_TOP_rx_bit_cnt[0]), .X(n23819) );
  sky130_fd_sc_hd__a21oi_1 U28355 ( .A1(j202_soc_core_uart_TOP_rx_bit_cnt[1]), 
        .A2(j202_soc_core_uart_TOP_rx_bit_cnt[0]), .B1(
        j202_soc_core_uart_TOP_rx_bit_cnt[2]), .Y(n23818) );
  sky130_fd_sc_hd__nor4_1 U28356 ( .A(j202_soc_core_rst), .B(n23819), .C(
        n23818), .D(n23821), .Y(j202_soc_core_uart_TOP_N88) );
  sky130_fd_sc_hd__xnor2_1 U28357 ( .A(j202_soc_core_uart_TOP_rx_bit_cnt[3]), 
        .B(n23819), .Y(n23820) );
  sky130_fd_sc_hd__nand2b_1 U28359 ( .A_N(j202_soc_core_uart_TOP_rxd_s), .B(
        j202_soc_core_uart_TOP_rxd_r), .Y(n23822) );
  sky130_fd_sc_hd__o211ai_1 U28360 ( .A1(j202_soc_core_uart_TOP_rx_go), .A2(
        n23822), .B1(n25731), .C1(n23821), .Y(j202_soc_core_uart_TOP_N85) );
  sky130_fd_sc_hd__nand2b_1 U28361 ( .A_N(j202_soc_core_uart_TOP_load), .B(
        n25401), .Y(n23828) );
  sky130_fd_sc_hd__nand2_1 U28363 ( .A(j202_soc_core_uart_TOP_tx_bit_cnt[0]), 
        .B(j202_soc_core_uart_TOP_tx_bit_cnt[1]), .Y(n23825) );
  sky130_fd_sc_hd__nor2_1 U28365 ( .A(n23828), .B(n23823), .Y(
        j202_soc_core_uart_TOP_N59) );
  sky130_fd_sc_hd__and3_1 U28366 ( .A(j202_soc_core_uart_TOP_tx_bit_cnt[0]), 
        .B(j202_soc_core_uart_TOP_tx_bit_cnt[1]), .C(
        j202_soc_core_uart_TOP_tx_bit_cnt[2]), .X(n23826) );
  sky130_fd_sc_hd__a211oi_1 U28367 ( .A1(n23825), .A2(n23824), .B1(n23826), 
        .C1(n23828), .Y(j202_soc_core_uart_TOP_N60) );
  sky130_fd_sc_hd__xnor2_1 U28368 ( .A(j202_soc_core_uart_TOP_tx_bit_cnt[3]), 
        .B(n23826), .Y(n23827) );
  sky130_fd_sc_hd__clkinv_1 U28370 ( .A(j202_soc_core_uart_TOP_N24), .Y(n23858) );
  sky130_fd_sc_hd__nand2_1 U28371 ( .A(n23858), .B(n25731), .Y(
        j202_soc_core_uart_TOP_N57) );
  sky130_fd_sc_hd__nor2_1 U28372 ( .A(j202_soc_core_uart_TOP_shift_en), .B(
        j202_soc_core_uart_TOP_shift_en_r), .Y(n23829) );
  sky130_fd_sc_hd__nor2_1 U28373 ( .A(j202_soc_core_uart_TOP_hold_reg[0]), .B(
        n23829), .Y(n23830) );
  sky130_fd_sc_hd__clkinv_1 U28374 ( .A(j202_soc_core_uart_sio_ce), .Y(n24821)
         );
  sky130_fd_sc_hd__nor2_1 U28376 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[0]), 
        .B(j202_soc_core_uart_TOP_tx_fifo_rp[1]), .Y(n23857) );
  sky130_fd_sc_hd__nor2_1 U28377 ( .A(n25123), .B(n23831), .Y(n23855) );
  sky130_fd_sc_hd__a22oi_1 U28378 ( .A1(n23857), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[24]), .B1(n23855), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[0]), .Y(n23833) );
  sky130_fd_sc_hd__nor2_1 U28379 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[0]), 
        .B(n23831), .Y(n23856) );
  sky130_fd_sc_hd__nor2_1 U28380 ( .A(j202_soc_core_uart_TOP_tx_fifo_rp[1]), 
        .B(n25123), .Y(n23854) );
  sky130_fd_sc_hd__a22oi_1 U28381 ( .A1(n23856), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[8]), .B1(n23854), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[16]), .Y(n23832) );
  sky130_fd_sc_hd__a21oi_1 U28382 ( .A1(n23833), .A2(n23832), .B1(n25122), .Y(
        n23834) );
  sky130_fd_sc_hd__a21o_1 U28383 ( .A1(j202_soc_core_uart_TOP_hold_reg[2]), 
        .A2(n23853), .B1(n23834), .X(j202_soc_core_uart_TOP_N26) );
  sky130_fd_sc_hd__a22oi_1 U28384 ( .A1(n23854), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[17]), .B1(n23855), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[1]), .Y(n23836) );
  sky130_fd_sc_hd__a22oi_1 U28385 ( .A1(n23856), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[9]), .B1(n23857), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[25]), .Y(n23835) );
  sky130_fd_sc_hd__a21oi_1 U28386 ( .A1(n23836), .A2(n23835), .B1(n25122), .Y(
        n23837) );
  sky130_fd_sc_hd__a21o_1 U28387 ( .A1(j202_soc_core_uart_TOP_hold_reg[3]), 
        .A2(n23853), .B1(n23837), .X(j202_soc_core_uart_TOP_N27) );
  sky130_fd_sc_hd__a22oi_1 U28388 ( .A1(n23854), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[18]), .B1(n23855), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[2]), .Y(n23839) );
  sky130_fd_sc_hd__a22oi_1 U28389 ( .A1(n23856), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[10]), .B1(n23857), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[26]), .Y(n23838) );
  sky130_fd_sc_hd__a21oi_1 U28390 ( .A1(n23839), .A2(n23838), .B1(n25122), .Y(
        n23840) );
  sky130_fd_sc_hd__a21o_1 U28391 ( .A1(j202_soc_core_uart_TOP_hold_reg[4]), 
        .A2(n23853), .B1(n23840), .X(j202_soc_core_uart_TOP_N28) );
  sky130_fd_sc_hd__a22oi_1 U28392 ( .A1(n23856), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[11]), .B1(n23854), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[19]), .Y(n23842) );
  sky130_fd_sc_hd__a22oi_1 U28393 ( .A1(n23857), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[27]), .B1(n23855), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[3]), .Y(n23841) );
  sky130_fd_sc_hd__a21oi_1 U28394 ( .A1(n23842), .A2(n23841), .B1(n25122), .Y(
        n23843) );
  sky130_fd_sc_hd__a21o_1 U28395 ( .A1(j202_soc_core_uart_TOP_hold_reg[5]), 
        .A2(n23853), .B1(n23843), .X(j202_soc_core_uart_TOP_N29) );
  sky130_fd_sc_hd__a22oi_1 U28396 ( .A1(n23854), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[20]), .B1(n23855), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[4]), .Y(n23845) );
  sky130_fd_sc_hd__a22oi_1 U28397 ( .A1(n23856), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[12]), .B1(n23857), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[28]), .Y(n23844) );
  sky130_fd_sc_hd__a21oi_1 U28398 ( .A1(n23845), .A2(n23844), .B1(n25122), .Y(
        n23846) );
  sky130_fd_sc_hd__a21o_1 U28399 ( .A1(j202_soc_core_uart_TOP_hold_reg[6]), 
        .A2(n23853), .B1(n23846), .X(j202_soc_core_uart_TOP_N30) );
  sky130_fd_sc_hd__a22oi_1 U28400 ( .A1(n23856), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[13]), .B1(n23857), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[29]), .Y(n23848) );
  sky130_fd_sc_hd__a22oi_1 U28401 ( .A1(n23854), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[21]), .B1(n23855), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[5]), .Y(n23847) );
  sky130_fd_sc_hd__a21oi_1 U28402 ( .A1(n23848), .A2(n23847), .B1(n25122), .Y(
        n23849) );
  sky130_fd_sc_hd__a21o_1 U28403 ( .A1(j202_soc_core_uart_TOP_hold_reg[7]), 
        .A2(n23853), .B1(n23849), .X(j202_soc_core_uart_TOP_N31) );
  sky130_fd_sc_hd__a22oi_1 U28404 ( .A1(n23857), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[30]), .B1(n23855), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[6]), .Y(n23851) );
  sky130_fd_sc_hd__a22oi_1 U28405 ( .A1(n23856), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[14]), .B1(n23854), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[22]), .Y(n23850) );
  sky130_fd_sc_hd__a21oi_1 U28406 ( .A1(n23851), .A2(n23850), .B1(n25122), .Y(
        n23852) );
  sky130_fd_sc_hd__a21o_1 U28407 ( .A1(j202_soc_core_uart_TOP_hold_reg[8]), 
        .A2(n23853), .B1(n23852), .X(j202_soc_core_uart_TOP_N32) );
  sky130_fd_sc_hd__a21oi_1 U28408 ( .A1(n23854), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[23]), .B1(n25122), .Y(n23861) );
  sky130_fd_sc_hd__a22oi_1 U28409 ( .A1(n23856), .A2(
        j202_soc_core_uart_TOP_tx_fifo_mem[15]), .B1(n23855), .B2(
        j202_soc_core_uart_TOP_tx_fifo_mem[7]), .Y(n23860) );
  sky130_fd_sc_hd__nand2_1 U28410 ( .A(n23857), .B(
        j202_soc_core_uart_TOP_tx_fifo_mem[31]), .Y(n23859) );
  sky130_fd_sc_hd__a31oi_1 U28411 ( .A1(n23861), .A2(n23860), .A3(n23859), 
        .B1(n23858), .Y(j202_soc_core_uart_TOP_N33) );
  sky130_fd_sc_hd__nand2_1 U28412 ( .A(n23862), .B(j202_soc_core_uart_sio_ce), 
        .Y(n23863) );
  sky130_fd_sc_hd__o21ai_1 U28413 ( .A1(j202_soc_core_uart_TOP_tx_fifo_gb), 
        .A2(n23863), .B1(n25734), .Y(j202_soc_core_uart_TOP_N16) );
  sky130_fd_sc_hd__clkinv_1 U28414 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[2]), .Y(n23881) );
  sky130_fd_sc_hd__nor2_1 U28415 ( .A(j202_soc_core_rst), .B(n23881), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N5) );
  sky130_fd_sc_hd__clkinv_1 U28416 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[20]), .Y(n23988) );
  sky130_fd_sc_hd__nor2_1 U28417 ( .A(j202_soc_core_rst), .B(n23988), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N23) );
  sky130_fd_sc_hd__clkinv_1 U28418 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[28]), .Y(n24040) );
  sky130_fd_sc_hd__nor2_1 U28419 ( .A(j202_soc_core_rst), .B(n24040), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_3_N31) );
  sky130_fd_sc_hd__a21oi_1 U28420 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[0]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[0]), .B1(
        gpio_en_o[0]), .Y(n23864) );
  sky130_fd_sc_hd__nand3_1 U28421 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[0]), .B(n23864), .C(n25734), .Y(n23871) );
  sky130_fd_sc_hd__clkinv_1 U28422 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[0]), .Y(n23865) );
  sky130_fd_sc_hd__o22ai_1 U28423 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[0]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[0]), .B1(n23865), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[0]), .Y(n23870)
         );
  sky130_fd_sc_hd__nand2_1 U28424 ( .A(n24071), .B(n23866), .Y(n24075) );
  sky130_fd_sc_hd__nor2_1 U28425 ( .A(n23867), .B(n24075), .Y(n23872) );
  sky130_fd_sc_hd__nor2_1 U28426 ( .A(j202_soc_core_rst), .B(n23872), .Y(
        n24042) );
  sky130_fd_sc_hd__o21ai_1 U28428 ( .A1(n23871), .A2(n23870), .B1(n23869), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N40) );
  sky130_fd_sc_hd__clkinv_1 U28430 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[1]), .Y(n23874) );
  sky130_fd_sc_hd__o22ai_1 U28431 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[1]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]), .B1(n23874), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[1]), .Y(n23875)
         );
  sky130_fd_sc_hd__a21oi_1 U28432 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[1]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]), .B1(n23875), 
        .Y(n23876) );
  sky130_fd_sc_hd__nand3_1 U28433 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[1]), .B(n23876), .C(
        io_oeb[1]), .Y(n23877) );
  sky130_fd_sc_hd__a21oi_1 U28434 ( .A1(n23878), .A2(n23877), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N41) );
  sky130_fd_sc_hd__nand4_1 U28436 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[2]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[2]), .C(n25731), .D(
        n23881), .Y(n23880) );
  sky130_fd_sc_hd__o41ai_1 U28437 ( .A1(j202_soc_core_rst), .A2(n23881), .A3(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[2]), .A4(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[2]), .B1(n23880), .Y(
        n23882) );
  sky130_fd_sc_hd__nand3_1 U28438 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[2]), .B(n23882), .C(
        io_oeb[2]), .Y(n23883) );
  sky130_fd_sc_hd__o21ai_1 U28439 ( .A1(j202_soc_core_rst), .A2(n23884), .B1(
        n23883), .Y(j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N42) );
  sky130_fd_sc_hd__clkinv_1 U28441 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[3]), .Y(n23886) );
  sky130_fd_sc_hd__o22ai_1 U28442 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[3]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]), .B1(n23886), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[3]), .Y(n23887)
         );
  sky130_fd_sc_hd__a21oi_1 U28443 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[3]), .B1(n23887), 
        .Y(n23888) );
  sky130_fd_sc_hd__nand3_1 U28444 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[3]), .B(n23888), .C(
        io_oeb[3]), .Y(n23889) );
  sky130_fd_sc_hd__a21oi_1 U28445 ( .A1(n23890), .A2(n23889), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N43) );
  sky130_fd_sc_hd__o211ai_1 U28446 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[4]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[4]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[4]), .C1(n25734), .Y(
        n23896) );
  sky130_fd_sc_hd__clkinv_1 U28447 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[4]), .Y(n23892) );
  sky130_fd_sc_hd__a21oi_1 U28448 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[4]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[4]), .B1(
        gpio_en_o[4]), .Y(n23891) );
  sky130_fd_sc_hd__o21ai_1 U28449 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[4]), .A2(n23892), 
        .B1(n23891), .Y(n23895) );
  sky130_fd_sc_hd__o21ai_1 U28450 ( .A1(n23893), .A2(n24042), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[4]), .Y(n23894) );
  sky130_fd_sc_hd__o21ai_1 U28451 ( .A1(n23896), .A2(n23895), .B1(n23894), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N44) );
  sky130_fd_sc_hd__clkinv_1 U28453 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[5]), .Y(n23898) );
  sky130_fd_sc_hd__o22ai_1 U28454 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[5]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]), .B1(n23898), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[5]), .Y(n23899)
         );
  sky130_fd_sc_hd__a21oi_1 U28455 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[5]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]), .B1(n23899), 
        .Y(n23900) );
  sky130_fd_sc_hd__nand3_1 U28456 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[5]), .B(n23900), .C(
        io_oeb[7]), .Y(n23901) );
  sky130_fd_sc_hd__a21oi_1 U28457 ( .A1(n23902), .A2(n23901), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N45) );
  sky130_fd_sc_hd__o21ai_1 U28458 ( .A1(n23903), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[6]), .Y(n23908) );
  sky130_fd_sc_hd__clkinv_1 U28459 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[6]), .Y(n23904) );
  sky130_fd_sc_hd__o22ai_1 U28460 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[6]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]), .B1(n23904), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[6]), .Y(n23905)
         );
  sky130_fd_sc_hd__a21oi_1 U28461 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[6]), .B1(n23905), 
        .Y(n23906) );
  sky130_fd_sc_hd__nand3_1 U28462 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[6]), .B(n23906), .C(
        io_oeb[26]), .Y(n23907) );
  sky130_fd_sc_hd__a21oi_1 U28463 ( .A1(n23908), .A2(n23907), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N46) );
  sky130_fd_sc_hd__o21ai_1 U28464 ( .A1(n23909), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[7]), .Y(n23914) );
  sky130_fd_sc_hd__clkinv_1 U28465 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[7]), .Y(n23910) );
  sky130_fd_sc_hd__o22ai_1 U28466 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[7]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]), .B1(n23910), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[7]), .Y(n23911)
         );
  sky130_fd_sc_hd__a21oi_1 U28467 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[7]), .B1(n23911), 
        .Y(n23912) );
  sky130_fd_sc_hd__nand3_1 U28468 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[7]), .B(n23912), .C(
        io_oeb[27]), .Y(n23913) );
  sky130_fd_sc_hd__a21oi_1 U28469 ( .A1(n23914), .A2(n23913), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N47) );
  sky130_fd_sc_hd__clkinv_1 U28470 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[8]), .Y(n23915) );
  sky130_fd_sc_hd__o21ai_0 U28471 ( .A1(n23915), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[8]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[8]), .Y(n23916) );
  sky130_fd_sc_hd__a21oi_1 U28472 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[8]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]), .B1(n23916), 
        .Y(n23917) );
  sky130_fd_sc_hd__o21ai_1 U28474 ( .A1(n23918), .A2(n24042), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[8]), .Y(n23919) );
  sky130_fd_sc_hd__o31ai_1 U28475 ( .A1(j202_soc_core_rst), .A2(gpio_en_o[8]), 
        .A3(n23920), .B1(n23919), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N48) );
  sky130_fd_sc_hd__clkinv_1 U28476 ( .A(j202_soc_core_qspi_wb_wdat[9]), .Y(
        n23921) );
  sky130_fd_sc_hd__o21ai_1 U28477 ( .A1(n23921), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[9]), .Y(n23926) );
  sky130_fd_sc_hd__clkinv_1 U28478 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[9]), .Y(n23922) );
  sky130_fd_sc_hd__o22ai_1 U28479 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[9]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[9]), .B1(n23922), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[9]), .Y(n23923)
         );
  sky130_fd_sc_hd__a21oi_1 U28480 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[9]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[9]), .B1(n23923), 
        .Y(n23924) );
  sky130_fd_sc_hd__nand3_1 U28481 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[9]), .B(n23924), .C(
        io_oeb[29]), .Y(n23925) );
  sky130_fd_sc_hd__a21oi_1 U28482 ( .A1(n23926), .A2(n23925), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N49) );
  sky130_fd_sc_hd__clkinv_1 U28483 ( .A(j202_soc_core_qspi_wb_wdat[10]), .Y(
        n23927) );
  sky130_fd_sc_hd__o21ai_1 U28484 ( .A1(n23927), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[10]), .Y(n23932) );
  sky130_fd_sc_hd__clkinv_1 U28485 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[10]), .Y(n23928) );
  sky130_fd_sc_hd__o22ai_1 U28486 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[10]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[10]), .B1(n23928), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[10]), .Y(n23929)
         );
  sky130_fd_sc_hd__a21oi_1 U28487 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[10]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[10]), .B1(n23929), 
        .Y(n23930) );
  sky130_fd_sc_hd__nand3_1 U28488 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[10]), .B(n23930), .C(
        io_oeb[30]), .Y(n23931) );
  sky130_fd_sc_hd__a21oi_1 U28489 ( .A1(n23932), .A2(n23931), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N50) );
  sky130_fd_sc_hd__clkinv_1 U28490 ( .A(j202_soc_core_qspi_wb_wdat[11]), .Y(
        n23933) );
  sky130_fd_sc_hd__o21ai_1 U28491 ( .A1(n23933), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[11]), .Y(n23938) );
  sky130_fd_sc_hd__clkinv_1 U28492 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[11]), .Y(n23934) );
  sky130_fd_sc_hd__o22ai_1 U28493 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[11]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[11]), .B1(n23934), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[11]), .Y(n23935)
         );
  sky130_fd_sc_hd__a21oi_1 U28494 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[11]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[11]), .B1(n23935), 
        .Y(n23936) );
  sky130_fd_sc_hd__nand3_1 U28495 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[11]), .B(n23936), .C(
        io_oeb[31]), .Y(n23937) );
  sky130_fd_sc_hd__a21oi_1 U28496 ( .A1(n23938), .A2(n23937), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N51) );
  sky130_fd_sc_hd__a21oi_1 U28497 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[12]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[12]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[12]), .Y(n23943) );
  sky130_fd_sc_hd__nand4_1 U28499 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[12]), .B(n25734), .C(
        io_oeb[32]), .D(n23939), .Y(n23942) );
  sky130_fd_sc_hd__o21ai_1 U28500 ( .A1(n23940), .A2(n24042), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[12]), .Y(n23941) );
  sky130_fd_sc_hd__clkinv_1 U28502 ( .A(j202_soc_core_qspi_wb_wdat[13]), .Y(
        n23944) );
  sky130_fd_sc_hd__o21ai_1 U28503 ( .A1(n23944), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[13]), .Y(n23949) );
  sky130_fd_sc_hd__clkinv_1 U28504 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[13]), .Y(n23945) );
  sky130_fd_sc_hd__o22ai_1 U28505 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[13]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13]), .B1(n23945), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[13]), .Y(n23946)
         );
  sky130_fd_sc_hd__a21oi_1 U28506 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[13]), .B1(n23946), 
        .Y(n23947) );
  sky130_fd_sc_hd__nand3_1 U28507 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[13]), .B(n23947), .C(
        io_oeb[33]), .Y(n23948) );
  sky130_fd_sc_hd__a21oi_1 U28508 ( .A1(n23949), .A2(n23948), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N53) );
  sky130_fd_sc_hd__clkinv_1 U28509 ( .A(j202_soc_core_qspi_wb_wdat[14]), .Y(
        n23950) );
  sky130_fd_sc_hd__clkinv_1 U28511 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[14]), .Y(n23951) );
  sky130_fd_sc_hd__o22ai_1 U28512 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[14]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14]), .B1(n23951), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[14]), .Y(n23952)
         );
  sky130_fd_sc_hd__a21oi_1 U28513 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[14]), .B1(n23952), 
        .Y(n23953) );
  sky130_fd_sc_hd__nand3_1 U28514 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[14]), .B(n23953), .C(
        io_oeb[34]), .Y(n23954) );
  sky130_fd_sc_hd__a21oi_1 U28515 ( .A1(n23955), .A2(n23954), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N54) );
  sky130_fd_sc_hd__clkinv_1 U28516 ( .A(j202_soc_core_qspi_wb_wdat[15]), .Y(
        n23956) );
  sky130_fd_sc_hd__o21ai_1 U28517 ( .A1(n23956), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[15]), .Y(n23961) );
  sky130_fd_sc_hd__clkinv_1 U28518 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[15]), .Y(n23957) );
  sky130_fd_sc_hd__o22ai_1 U28519 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[15]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15]), .B1(n23957), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[15]), .Y(n23958)
         );
  sky130_fd_sc_hd__a21oi_1 U28520 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[15]), .B1(n23958), 
        .Y(n23959) );
  sky130_fd_sc_hd__nand3_1 U28521 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[15]), .B(n23959), .C(
        io_oeb[35]), .Y(n23960) );
  sky130_fd_sc_hd__a21oi_1 U28522 ( .A1(n23961), .A2(n23960), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N55) );
  sky130_fd_sc_hd__clkinv_1 U28523 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[16]), .Y(n23962) );
  sky130_fd_sc_hd__o21ai_0 U28524 ( .A1(n23962), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[16]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[16]), .Y(n23963) );
  sky130_fd_sc_hd__a21oi_1 U28525 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[16]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16]), .B1(n23963), 
        .Y(n23964) );
  sky130_fd_sc_hd__o21ai_1 U28526 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[16]), .B1(n23964), .Y(
        n23967) );
  sky130_fd_sc_hd__o21ai_1 U28527 ( .A1(n23965), .A2(n24042), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[16]), .Y(n23966) );
  sky130_fd_sc_hd__o31ai_1 U28528 ( .A1(j202_soc_core_rst), .A2(gpio_en_o[16]), 
        .A3(n23967), .B1(n23966), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N56) );
  sky130_fd_sc_hd__clkinv_1 U28530 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[17]), .Y(n23969) );
  sky130_fd_sc_hd__o22ai_1 U28531 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[17]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[17]), .B1(n23969), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[17]), .Y(n23970)
         );
  sky130_fd_sc_hd__a21oi_1 U28532 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[17]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[17]), .B1(n23970), 
        .Y(n23971) );
  sky130_fd_sc_hd__nand3_1 U28533 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[17]), .B(n23971), .C(
        io_oeb[37]), .Y(n23972) );
  sky130_fd_sc_hd__a21oi_1 U28534 ( .A1(n23973), .A2(n23972), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N57) );
  sky130_fd_sc_hd__o21ai_1 U28535 ( .A1(n23974), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[18]), .Y(n23980) );
  sky130_fd_sc_hd__clkinv_1 U28536 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[18]), .Y(n23977) );
  sky130_fd_sc_hd__a21oi_1 U28537 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[18]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[18]), .B1(gpio_en_o[18]), 
        .Y(n23975) );
  sky130_fd_sc_hd__nand2_1 U28538 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[18]), .B(n23975), .Y(
        n23976) );
  sky130_fd_sc_hd__a21oi_1 U28539 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[18]), .A2(n23977), 
        .B1(n23976), .Y(n23978) );
  sky130_fd_sc_hd__a21oi_1 U28541 ( .A1(n23980), .A2(n23979), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N58) );
  sky130_fd_sc_hd__o21ai_1 U28542 ( .A1(n23981), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[19]), .Y(n23987) );
  sky130_fd_sc_hd__clkinv_1 U28543 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[19]), .Y(n23982) );
  sky130_fd_sc_hd__a21oi_1 U28544 ( .A1(n23982), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[19]), .B1(
        gpio_en_o[19]), .Y(n23983) );
  sky130_fd_sc_hd__nand2_1 U28545 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[19]), .B(n23983), .Y(
        n23984) );
  sky130_fd_sc_hd__a21oi_1 U28546 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[19]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[19]), .B1(n23984), .Y(
        n23985) );
  sky130_fd_sc_hd__a21oi_1 U28548 ( .A1(n23987), .A2(n23986), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N59) );
  sky130_fd_sc_hd__nor2_1 U28549 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[20]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[20]), .Y(n23993) );
  sky130_fd_sc_hd__o2bb2ai_1 U28550 ( .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[20]), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[20]), .A1_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[20]), .A2_N(n23988), .Y(
        n23989) );
  sky130_fd_sc_hd__nand3_1 U28551 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[20]), .B(n23989), .C(
        n25732), .Y(n23992) );
  sky130_fd_sc_hd__o21ai_1 U28552 ( .A1(n23990), .A2(n24042), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[20]), .Y(n23991) );
  sky130_fd_sc_hd__o31ai_1 U28553 ( .A1(gpio_en_o[20]), .A2(n23993), .A3(
        n23992), .B1(n23991), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N60) );
  sky130_fd_sc_hd__clkinv_1 U28554 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[21]), .Y(n23994) );
  sky130_fd_sc_hd__o22ai_1 U28555 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[21]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[21]), .B1(n23994), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_dtr[21]), .Y(n23995) );
  sky130_fd_sc_hd__a211oi_1 U28556 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[21]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[21]), .B1(gpio_en_o[21]), 
        .C1(n23995), .Y(n23996) );
  sky130_fd_sc_hd__nand2_1 U28557 ( .A(n23996), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[21]), .Y(n23999) );
  sky130_fd_sc_hd__o21ai_1 U28558 ( .A1(n23997), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[21]), .Y(n23998) );
  sky130_fd_sc_hd__a21oi_1 U28559 ( .A1(n23999), .A2(n23998), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N61) );
  sky130_fd_sc_hd__o21ai_1 U28560 ( .A1(n24000), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[22]), .Y(n24006) );
  sky130_fd_sc_hd__clkinv_1 U28561 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[22]), .Y(n24003) );
  sky130_fd_sc_hd__a21oi_1 U28562 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[22]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[22]), .B1(gpio_en_o[22]), 
        .Y(n24001) );
  sky130_fd_sc_hd__nand2_1 U28563 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[22]), .B(n24001), .Y(
        n24002) );
  sky130_fd_sc_hd__a21oi_1 U28564 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[22]), .A2(n24003), 
        .B1(n24002), .Y(n24004) );
  sky130_fd_sc_hd__a21oi_1 U28566 ( .A1(n24006), .A2(n24005), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N62) );
  sky130_fd_sc_hd__clkinv_1 U28567 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[23]), .Y(n24007) );
  sky130_fd_sc_hd__a21oi_1 U28568 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[23]), .A2(n24007), 
        .B1(gpio_en_o[23]), .Y(n24008) );
  sky130_fd_sc_hd__a21oi_1 U28570 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[23]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[23]), .B1(n24009), .Y(
        n24010) );
  sky130_fd_sc_hd__nand2_1 U28571 ( .A(n24010), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[23]), .Y(n24013) );
  sky130_fd_sc_hd__o21ai_1 U28572 ( .A1(n24011), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[23]), .Y(n24012) );
  sky130_fd_sc_hd__a21oi_1 U28573 ( .A1(n24013), .A2(n24012), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N63) );
  sky130_fd_sc_hd__o211ai_1 U28574 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[24]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[24]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[24]), .C1(n25734), .Y(
        n24018) );
  sky130_fd_sc_hd__clkinv_1 U28575 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[24]), .Y(n24014) );
  sky130_fd_sc_hd__a221o_1 U28576 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[24]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[24]), .B1(n24014), 
        .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[24]), .C1(
        gpio_en_o[24]), .X(n24017) );
  sky130_fd_sc_hd__o21ai_1 U28577 ( .A1(n24015), .A2(n24042), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[24]), .Y(n24016) );
  sky130_fd_sc_hd__o21ai_1 U28579 ( .A1(n24019), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[25]), .Y(n24025) );
  sky130_fd_sc_hd__clkinv_1 U28580 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[25]), .Y(n24020) );
  sky130_fd_sc_hd__a21oi_1 U28581 ( .A1(n24020), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[25]), .B1(
        gpio_en_o[25]), .Y(n24021) );
  sky130_fd_sc_hd__nand2_1 U28582 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[25]), .B(n24021), .Y(
        n24022) );
  sky130_fd_sc_hd__a21oi_1 U28583 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[25]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[25]), .B1(n24022), .Y(
        n24023) );
  sky130_fd_sc_hd__a21oi_1 U28585 ( .A1(n24025), .A2(n24024), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N65) );
  sky130_fd_sc_hd__o21ai_1 U28586 ( .A1(n24026), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[26]), .Y(n24032) );
  sky130_fd_sc_hd__clkinv_1 U28587 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[26]), .Y(n24029) );
  sky130_fd_sc_hd__a21oi_1 U28588 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[26]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[26]), .B1(gpio_en_o[26]), 
        .Y(n24027) );
  sky130_fd_sc_hd__nand2_1 U28589 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[26]), .B(n24027), .Y(
        n24028) );
  sky130_fd_sc_hd__a21oi_1 U28590 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[26]), .A2(n24029), 
        .B1(n24028), .Y(n24030) );
  sky130_fd_sc_hd__a21oi_1 U28592 ( .A1(n24032), .A2(n24031), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N66) );
  sky130_fd_sc_hd__clkinv_1 U28593 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[27]), .Y(n24033) );
  sky130_fd_sc_hd__a21oi_1 U28594 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[27]), .A2(n24033), 
        .B1(gpio_en_o[27]), .Y(n24034) );
  sky130_fd_sc_hd__a21oi_1 U28596 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[27]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[27]), .B1(n24035), 
        .Y(n24036) );
  sky130_fd_sc_hd__nand2_1 U28597 ( .A(n24036), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[27]), .Y(n24039) );
  sky130_fd_sc_hd__a21oi_1 U28599 ( .A1(n24039), .A2(n24038), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N67) );
  sky130_fd_sc_hd__o2bb2ai_1 U28600 ( .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[28]), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[28]), .A1_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[28]), .A2_N(n24040), .Y(
        n24041) );
  sky130_fd_sc_hd__o211ai_1 U28601 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[28]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[28]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[28]), .C1(n24041), .Y(
        n24045) );
  sky130_fd_sc_hd__o21ai_1 U28602 ( .A1(n24043), .A2(n24042), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[28]), .Y(n24044) );
  sky130_fd_sc_hd__o31ai_1 U28603 ( .A1(j202_soc_core_rst), .A2(gpio_en_o[28]), 
        .A3(n24045), .B1(n24044), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N68) );
  sky130_fd_sc_hd__o21ai_1 U28604 ( .A1(n24046), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[29]), .Y(n24052) );
  sky130_fd_sc_hd__clkinv_1 U28605 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[29]), .Y(n24047) );
  sky130_fd_sc_hd__a21oi_1 U28606 ( .A1(n24047), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[29]), .B1(
        gpio_en_o[29]), .Y(n24048) );
  sky130_fd_sc_hd__nand2_1 U28607 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[29]), .B(n24048), .Y(
        n24049) );
  sky130_fd_sc_hd__a21oi_1 U28608 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[29]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[29]), .B1(n24049), .Y(
        n24050) );
  sky130_fd_sc_hd__o21ai_1 U28609 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[29]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[29]), .B1(n24050), 
        .Y(n24051) );
  sky130_fd_sc_hd__a21oi_1 U28610 ( .A1(n24052), .A2(n24051), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N69) );
  sky130_fd_sc_hd__o21ai_1 U28611 ( .A1(n24053), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[30]), .Y(n24059) );
  sky130_fd_sc_hd__clkinv_1 U28612 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[30]), .Y(n24054) );
  sky130_fd_sc_hd__a21oi_1 U28613 ( .A1(n24054), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[30]), .B1(
        gpio_en_o[30]), .Y(n24055) );
  sky130_fd_sc_hd__nand2_1 U28614 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[30]), .B(n24055), .Y(
        n24056) );
  sky130_fd_sc_hd__a21oi_1 U28615 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[30]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[30]), .B1(n24056), .Y(
        n24057) );
  sky130_fd_sc_hd__a21oi_1 U28617 ( .A1(n24059), .A2(n24058), .B1(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N70) );
  sky130_fd_sc_hd__a21oi_1 U28618 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[31]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[31]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[31]), .Y(n24065) );
  sky130_fd_sc_hd__nand4b_1 U28620 ( .A_N(gpio_en_o[31]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[31]), .C(n25732), .D(
        n24060), .Y(n24064) );
  sky130_fd_sc_hd__o21ai_1 U28621 ( .A1(n24062), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[31]), .Y(n24063) );
  sky130_fd_sc_hd__o22ai_1 U28622 ( .A1(n24065), .A2(n24064), .B1(
        j202_soc_core_rst), .B2(n24063), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N71) );
  sky130_fd_sc_hd__nor2b_1 U28623 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[0]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N3) );
  sky130_fd_sc_hd__nor2b_1 U28624 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[1]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N4) );
  sky130_fd_sc_hd__nor2b_1 U28625 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[2]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N5) );
  sky130_fd_sc_hd__nor2b_1 U28626 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[3]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N6) );
  sky130_fd_sc_hd__nor2b_1 U28627 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[4]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N7) );
  sky130_fd_sc_hd__nor2b_1 U28628 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[5]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N8) );
  sky130_fd_sc_hd__nor2b_1 U28629 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[6]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N9) );
  sky130_fd_sc_hd__nor2b_1 U28630 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[7]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N10) );
  sky130_fd_sc_hd__nor2b_1 U28631 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[8]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N11) );
  sky130_fd_sc_hd__nor2b_1 U28632 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[9]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N12) );
  sky130_fd_sc_hd__nor2b_1 U28633 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[10]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N13) );
  sky130_fd_sc_hd__nor2b_1 U28634 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[11]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N14) );
  sky130_fd_sc_hd__nor2b_1 U28635 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[12]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N15) );
  sky130_fd_sc_hd__nor2b_1 U28636 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[13]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N16) );
  sky130_fd_sc_hd__nor2b_1 U28637 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[14]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N17) );
  sky130_fd_sc_hd__nor2b_1 U28638 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[15]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N18) );
  sky130_fd_sc_hd__nor2b_1 U28639 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[16]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N19) );
  sky130_fd_sc_hd__nor2b_1 U28640 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[17]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N20) );
  sky130_fd_sc_hd__nor2b_1 U28641 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[18]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N21) );
  sky130_fd_sc_hd__nor2b_1 U28642 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[19]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N22) );
  sky130_fd_sc_hd__nor2b_1 U28643 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[20]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N23) );
  sky130_fd_sc_hd__nor2b_1 U28644 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[21]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N24) );
  sky130_fd_sc_hd__nor2b_1 U28645 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[25]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N28) );
  sky130_fd_sc_hd__nor2b_1 U28646 ( .B_N(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_1[29]), .A(
        j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_2_N32) );
  sky130_fd_sc_hd__nor2b_1 U28647 ( .B_N(io_in[0]), .A(j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N3) );
  sky130_fd_sc_hd__nor2b_1 U28648 ( .B_N(io_in[1]), .A(j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N4) );
  sky130_fd_sc_hd__nor2b_1 U28649 ( .B_N(io_in[2]), .A(j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N5) );
  sky130_fd_sc_hd__nor2b_1 U28650 ( .B_N(io_in[3]), .A(j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N6) );
  sky130_fd_sc_hd__nor2b_1 U28651 ( .B_N(io_in[4]), .A(j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N7) );
  sky130_fd_sc_hd__nor2b_1 U28652 ( .B_N(io_in[7]), .A(j202_soc_core_rst), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N8) );
  sky130_fd_sc_hd__nor2b_1 U28653 ( .B_N(io_in[26]), .A(j202_soc_core_rst), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N9) );
  sky130_fd_sc_hd__nor2b_1 U28654 ( .B_N(io_in[27]), .A(j202_soc_core_rst), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N10) );
  sky130_fd_sc_hd__nor2b_1 U28655 ( .B_N(io_in[28]), .A(j202_soc_core_rst), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N11) );
  sky130_fd_sc_hd__nor2b_1 U28656 ( .B_N(io_in[29]), .A(j202_soc_core_rst), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N12) );
  sky130_fd_sc_hd__nor2b_1 U28657 ( .B_N(io_in[30]), .A(j202_soc_core_rst), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N13) );
  sky130_fd_sc_hd__nor2b_1 U28658 ( .B_N(io_in[31]), .A(j202_soc_core_rst), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N14) );
  sky130_fd_sc_hd__nor2b_1 U28659 ( .B_N(io_in[32]), .A(j202_soc_core_rst), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N15) );
  sky130_fd_sc_hd__nor2b_1 U28660 ( .B_N(io_in[33]), .A(j202_soc_core_rst), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N16) );
  sky130_fd_sc_hd__nor2b_1 U28661 ( .B_N(io_in[34]), .A(j202_soc_core_rst), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N17) );
  sky130_fd_sc_hd__nor2b_1 U28662 ( .B_N(io_in[35]), .A(j202_soc_core_rst), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N18) );
  sky130_fd_sc_hd__nor2b_1 U28663 ( .B_N(io_in[36]), .A(j202_soc_core_rst), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N19) );
  sky130_fd_sc_hd__nor2b_1 U28664 ( .B_N(io_in[37]), .A(j202_soc_core_rst), 
        .Y(j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N20) );
  sky130_fd_sc_hd__nor3b_1 U28665 ( .C_N(la_data_in[18]), .A(j202_soc_core_rst), .B(la_oenb[18]), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N21) );
  sky130_fd_sc_hd__nor3b_1 U28666 ( .C_N(la_data_in[19]), .A(j202_soc_core_rst), .B(la_oenb[19]), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N22) );
  sky130_fd_sc_hd__nor3b_1 U28667 ( .C_N(la_data_in[20]), .A(j202_soc_core_rst), .B(la_oenb[20]), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N23) );
  sky130_fd_sc_hd__nor3b_1 U28668 ( .C_N(la_data_in[21]), .A(j202_soc_core_rst), .B(la_oenb[21]), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N24) );
  sky130_fd_sc_hd__nor3b_1 U28669 ( .C_N(la_data_in[22]), .A(j202_soc_core_rst), .B(la_oenb[22]), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N25) );
  sky130_fd_sc_hd__nor3b_1 U28670 ( .C_N(la_data_in[23]), .A(j202_soc_core_rst), .B(la_oenb[23]), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N26) );
  sky130_fd_sc_hd__nor3b_1 U28671 ( .C_N(la_data_in[24]), .A(j202_soc_core_rst), .B(la_oenb[24]), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N27) );
  sky130_fd_sc_hd__nor3b_1 U28672 ( .C_N(la_data_in[25]), .A(j202_soc_core_rst), .B(la_oenb[25]), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N28) );
  sky130_fd_sc_hd__nor3b_1 U28673 ( .C_N(la_data_in[26]), .A(j202_soc_core_rst), .B(la_oenb[26]), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N29) );
  sky130_fd_sc_hd__nor3b_1 U28674 ( .C_N(la_data_in[27]), .A(j202_soc_core_rst), .B(la_oenb[27]), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N30) );
  sky130_fd_sc_hd__nor3b_1 U28675 ( .C_N(la_data_in[28]), .A(j202_soc_core_rst), .B(la_oenb[28]), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N31) );
  sky130_fd_sc_hd__nor3b_1 U28676 ( .C_N(la_data_in[29]), .A(j202_soc_core_rst), .B(la_oenb[29]), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N32) );
  sky130_fd_sc_hd__nor3b_1 U28677 ( .C_N(la_data_in[30]), .A(j202_soc_core_rst), .B(la_oenb[30]), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N33) );
  sky130_fd_sc_hd__nor3b_1 U28678 ( .C_N(la_data_in[31]), .A(j202_soc_core_rst), .B(la_oenb[31]), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_dff_gpio_in_1_N34) );
  sky130_fd_sc_hd__nand2_1 U28679 ( .A(n24067), .B(n25731), .Y(n24068) );
  sky130_fd_sc_hd__nor2_1 U28680 ( .A(n24069), .B(n24068), .Y(n24074) );
  sky130_fd_sc_hd__nand2_1 U28681 ( .A(n24074), .B(n24070), .Y(n24072) );
  sky130_fd_sc_hd__nor2b_1 U28682 ( .B_N(n24071), .A(n24072), .Y(n24173) );
  sky130_fd_sc_hd__nor2_1 U28683 ( .A(n24073), .B(n24072), .Y(n24174) );
  sky130_fd_sc_hd__a22oi_1 U28684 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[0]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[0]), .Y(n24082) );
  sky130_fd_sc_hd__nor2_1 U28685 ( .A(n24075), .B(n24079), .Y(n24177) );
  sky130_fd_sc_hd__nor2_1 U28686 ( .A(n24079), .B(n24076), .Y(n24175) );
  sky130_fd_sc_hd__a22oi_1 U28687 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[0]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[0]), .B2(n24175), .Y(
        n24081) );
  sky130_fd_sc_hd__nor2_1 U28688 ( .A(n24077), .B(n24079), .Y(n24176) );
  sky130_fd_sc_hd__nor2_1 U28689 ( .A(n24079), .B(n24078), .Y(n24178) );
  sky130_fd_sc_hd__a22oi_1 U28690 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[0]), .A2(n24176), .B1(
        gpio_en_o[0]), .B2(n24178), .Y(n24080) );
  sky130_fd_sc_hd__nand3_1 U28691 ( .A(n24082), .B(n24081), .C(n24080), .Y(
        j202_soc_core_ahb2apb_02_N128) );
  sky130_fd_sc_hd__a22oi_1 U28692 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[1]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[1]), .Y(n24085) );
  sky130_fd_sc_hd__a22oi_1 U28693 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[1]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[1]), .B2(n24176), .Y(
        n24084) );
  sky130_fd_sc_hd__a22oi_1 U28694 ( .A1(gpio_en_o[1]), .A2(n24178), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[1]), .B2(n24175), .Y(
        n24083) );
  sky130_fd_sc_hd__nand3_1 U28695 ( .A(n24085), .B(n24084), .C(n24083), .Y(
        j202_soc_core_ahb2apb_02_N129) );
  sky130_fd_sc_hd__a22oi_1 U28696 ( .A1(n24174), .A2(la_data_out[2]), .B1(
        n24173), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[2]), 
        .Y(n24088) );
  sky130_fd_sc_hd__a22oi_1 U28697 ( .A1(n24176), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[2]), .B1(n24178), .B2(
        gpio_en_o[2]), .Y(n24087) );
  sky130_fd_sc_hd__a22oi_1 U28698 ( .A1(n24175), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[2]), .B1(n24177), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[2]), .Y(n24086) );
  sky130_fd_sc_hd__nand3_1 U28699 ( .A(n24088), .B(n24087), .C(n24086), .Y(
        j202_soc_core_ahb2apb_02_N130) );
  sky130_fd_sc_hd__a22oi_1 U28700 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[3]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[3]), .Y(n24091) );
  sky130_fd_sc_hd__a22oi_1 U28701 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[3]), .A2(n24176), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[3]), .B2(n24175), .Y(
        n24090) );
  sky130_fd_sc_hd__a22oi_1 U28702 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[3]), .A2(n24177), .B1(
        gpio_en_o[3]), .B2(n24178), .Y(n24089) );
  sky130_fd_sc_hd__nand3_1 U28703 ( .A(n24091), .B(n24090), .C(n24089), .Y(
        j202_soc_core_ahb2apb_02_N131) );
  sky130_fd_sc_hd__a22oi_1 U28704 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[4]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[4]), .Y(n24094) );
  sky130_fd_sc_hd__a22oi_1 U28705 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[4]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[4]), .B2(n24175), .Y(
        n24093) );
  sky130_fd_sc_hd__a22oi_1 U28706 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[4]), .A2(n24176), .B1(
        gpio_en_o[4]), .B2(n24178), .Y(n24092) );
  sky130_fd_sc_hd__nand3_1 U28707 ( .A(n24094), .B(n24093), .C(n24092), .Y(
        j202_soc_core_ahb2apb_02_N132) );
  sky130_fd_sc_hd__a22oi_1 U28708 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[5]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[5]), .Y(n24097) );
  sky130_fd_sc_hd__a22oi_1 U28709 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[5]), .A2(n24175), .B1(
        gpio_en_o[5]), .B2(n24178), .Y(n24096) );
  sky130_fd_sc_hd__a22oi_1 U28710 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[5]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[5]), .B2(n24176), .Y(
        n24095) );
  sky130_fd_sc_hd__nand3_1 U28711 ( .A(n24097), .B(n24096), .C(n24095), .Y(
        j202_soc_core_ahb2apb_02_N133) );
  sky130_fd_sc_hd__a22oi_1 U28712 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[6]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[6]), .Y(n24100) );
  sky130_fd_sc_hd__a22oi_1 U28713 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[6]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[6]), .B2(n24176), .Y(
        n24099) );
  sky130_fd_sc_hd__a22oi_1 U28714 ( .A1(gpio_en_o[6]), .A2(n24178), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[6]), .B2(n24175), .Y(
        n24098) );
  sky130_fd_sc_hd__nand3_1 U28715 ( .A(n24100), .B(n24099), .C(n24098), .Y(
        j202_soc_core_ahb2apb_02_N134) );
  sky130_fd_sc_hd__a22oi_1 U28716 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[7]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[7]), .Y(n24103) );
  sky130_fd_sc_hd__a22oi_1 U28717 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[7]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[7]), .B2(n24176), .Y(
        n24102) );
  sky130_fd_sc_hd__a22oi_1 U28718 ( .A1(gpio_en_o[7]), .A2(n24178), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[7]), .B2(n24175), .Y(
        n24101) );
  sky130_fd_sc_hd__nand3_1 U28719 ( .A(n24103), .B(n24102), .C(n24101), .Y(
        j202_soc_core_ahb2apb_02_N135) );
  sky130_fd_sc_hd__a22oi_1 U28720 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[8]), .Y(n24106) );
  sky130_fd_sc_hd__a22oi_1 U28721 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[8]), .A2(n24176), .B1(
        gpio_en_o[8]), .B2(n24178), .Y(n24105) );
  sky130_fd_sc_hd__a22oi_1 U28722 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[8]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[8]), .B2(n24175), .Y(
        n24104) );
  sky130_fd_sc_hd__nand3_1 U28723 ( .A(n24106), .B(n24105), .C(n24104), .Y(
        j202_soc_core_ahb2apb_02_N136) );
  sky130_fd_sc_hd__a22oi_1 U28724 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[9]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[9]), .Y(n24109) );
  sky130_fd_sc_hd__a22oi_1 U28725 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[9]), .A2(n24176), .B1(
        gpio_en_o[9]), .B2(n24178), .Y(n24108) );
  sky130_fd_sc_hd__a22oi_1 U28726 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[9]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[9]), .B2(n24175), .Y(
        n24107) );
  sky130_fd_sc_hd__nand3_1 U28727 ( .A(n24109), .B(n24108), .C(n24107), .Y(
        j202_soc_core_ahb2apb_02_N137) );
  sky130_fd_sc_hd__a22oi_1 U28728 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[10]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[10]), .Y(n24112) );
  sky130_fd_sc_hd__a22oi_1 U28729 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[10]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[10]), .B2(n24176), .Y(
        n24111) );
  sky130_fd_sc_hd__a22oi_1 U28730 ( .A1(gpio_en_o[10]), .A2(n24178), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[10]), .B2(n24175), .Y(
        n24110) );
  sky130_fd_sc_hd__nand3_1 U28731 ( .A(n24112), .B(n24111), .C(n24110), .Y(
        j202_soc_core_ahb2apb_02_N138) );
  sky130_fd_sc_hd__a22oi_1 U28732 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[11]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[11]), .Y(n24115) );
  sky130_fd_sc_hd__a22oi_1 U28733 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[11]), .A2(n24176), .B1(
        gpio_en_o[11]), .B2(n24178), .Y(n24114) );
  sky130_fd_sc_hd__a22oi_1 U28734 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[11]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[11]), .B2(n24175), .Y(
        n24113) );
  sky130_fd_sc_hd__nand3_1 U28735 ( .A(n24115), .B(n24114), .C(n24113), .Y(
        j202_soc_core_ahb2apb_02_N139) );
  sky130_fd_sc_hd__a22oi_1 U28736 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[12]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[12]), .Y(n24118) );
  sky130_fd_sc_hd__a22oi_1 U28737 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[12]), .A2(n24176), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[12]), .B2(n24175), .Y(
        n24117) );
  sky130_fd_sc_hd__a22oi_1 U28738 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[12]), .A2(n24177), .B1(
        gpio_en_o[12]), .B2(n24178), .Y(n24116) );
  sky130_fd_sc_hd__nand3_1 U28739 ( .A(n24118), .B(n24117), .C(n24116), .Y(
        j202_soc_core_ahb2apb_02_N140) );
  sky130_fd_sc_hd__a22oi_1 U28740 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[13]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[13]), .Y(n24121) );
  sky130_fd_sc_hd__a22oi_1 U28741 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[13]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[13]), .B2(n24175), .Y(
        n24120) );
  sky130_fd_sc_hd__a22oi_1 U28742 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[13]), .A2(n24176), .B1(
        gpio_en_o[13]), .B2(n24178), .Y(n24119) );
  sky130_fd_sc_hd__nand3_1 U28743 ( .A(n24121), .B(n24120), .C(n24119), .Y(
        j202_soc_core_ahb2apb_02_N141) );
  sky130_fd_sc_hd__a22oi_1 U28744 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[14]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[14]), .Y(n24124) );
  sky130_fd_sc_hd__a22oi_1 U28745 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[14]), .A2(n24176), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[14]), .B2(n24175), .Y(
        n24123) );
  sky130_fd_sc_hd__a22oi_1 U28746 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[14]), .A2(n24177), .B1(
        gpio_en_o[14]), .B2(n24178), .Y(n24122) );
  sky130_fd_sc_hd__nand3_1 U28747 ( .A(n24124), .B(n24123), .C(n24122), .Y(
        j202_soc_core_ahb2apb_02_N142) );
  sky130_fd_sc_hd__a22oi_1 U28748 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[15]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[15]), .Y(n24127) );
  sky130_fd_sc_hd__a22oi_1 U28749 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[15]), .A2(n24177), .B1(
        gpio_en_o[15]), .B2(n24178), .Y(n24126) );
  sky130_fd_sc_hd__a22oi_1 U28750 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[15]), .A2(n24176), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[15]), .B2(n24175), .Y(
        n24125) );
  sky130_fd_sc_hd__nand3_1 U28751 ( .A(n24127), .B(n24126), .C(n24125), .Y(
        j202_soc_core_ahb2apb_02_N143) );
  sky130_fd_sc_hd__a22oi_1 U28752 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[16]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[16]), .Y(n24130) );
  sky130_fd_sc_hd__a22oi_1 U28753 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[16]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[16]), .B2(n24176), .Y(
        n24129) );
  sky130_fd_sc_hd__a22oi_1 U28754 ( .A1(gpio_en_o[16]), .A2(n24178), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[16]), .B2(n24175), .Y(
        n24128) );
  sky130_fd_sc_hd__nand3_1 U28755 ( .A(n24130), .B(n24129), .C(n24128), .Y(
        j202_soc_core_ahb2apb_02_N144) );
  sky130_fd_sc_hd__a22oi_1 U28756 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[17]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[17]), .Y(n24133) );
  sky130_fd_sc_hd__a22oi_1 U28757 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[17]), .A2(n24176), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[17]), .B2(n24175), .Y(
        n24132) );
  sky130_fd_sc_hd__a22oi_1 U28758 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[17]), .A2(n24177), .B1(
        gpio_en_o[17]), .B2(n24178), .Y(n24131) );
  sky130_fd_sc_hd__nand3_1 U28759 ( .A(n24133), .B(n24132), .C(n24131), .Y(
        j202_soc_core_ahb2apb_02_N145) );
  sky130_fd_sc_hd__a22oi_1 U28760 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[18]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[18]), .Y(n24136) );
  sky130_fd_sc_hd__a22oi_1 U28761 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[18]), .A2(n24176), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[18]), .B2(n24175), .Y(
        n24135) );
  sky130_fd_sc_hd__a22oi_1 U28762 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[18]), .A2(n24177), .B1(
        gpio_en_o[18]), .B2(n24178), .Y(n24134) );
  sky130_fd_sc_hd__nand3_1 U28763 ( .A(n24136), .B(n24135), .C(n24134), .Y(
        j202_soc_core_ahb2apb_02_N146) );
  sky130_fd_sc_hd__a22oi_1 U28764 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[19]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[19]), .Y(n24139) );
  sky130_fd_sc_hd__a22oi_1 U28765 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[19]), .A2(n24176), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[19]), .B2(n24175), .Y(
        n24138) );
  sky130_fd_sc_hd__a22oi_1 U28766 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[19]), .A2(n24177), .B1(
        gpio_en_o[19]), .B2(n24178), .Y(n24137) );
  sky130_fd_sc_hd__nand3_1 U28767 ( .A(n24139), .B(n24138), .C(n24137), .Y(
        j202_soc_core_ahb2apb_02_N147) );
  sky130_fd_sc_hd__a22oi_1 U28768 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[20]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[20]), .Y(n24142) );
  sky130_fd_sc_hd__a22oi_1 U28769 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[20]), .A2(n24175), .B1(
        gpio_en_o[20]), .B2(n24178), .Y(n24141) );
  sky130_fd_sc_hd__a22oi_1 U28770 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[20]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[20]), .B2(n24176), .Y(
        n24140) );
  sky130_fd_sc_hd__nand3_1 U28771 ( .A(n24142), .B(n24141), .C(n24140), .Y(
        j202_soc_core_ahb2apb_02_N148) );
  sky130_fd_sc_hd__a22oi_1 U28772 ( .A1(n24174), .A2(la_data_out[21]), .B1(
        n24173), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[21]), 
        .Y(n24145) );
  sky130_fd_sc_hd__a22oi_1 U28773 ( .A1(n24176), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[21]), .B1(n24177), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[21]), .Y(n24144) );
  sky130_fd_sc_hd__a22oi_1 U28774 ( .A1(n24178), .A2(gpio_en_o[21]), .B1(
        n24175), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_ier[21]), .Y(
        n24143) );
  sky130_fd_sc_hd__nand3_1 U28775 ( .A(n24145), .B(n24144), .C(n24143), .Y(
        j202_soc_core_ahb2apb_02_N149) );
  sky130_fd_sc_hd__a22oi_1 U28776 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[22]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[22]), .Y(n24148) );
  sky130_fd_sc_hd__a22oi_1 U28777 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[22]), .A2(n24176), .B1(
        gpio_en_o[22]), .B2(n24178), .Y(n24147) );
  sky130_fd_sc_hd__a22oi_1 U28778 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[22]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[22]), .B2(n24175), .Y(
        n24146) );
  sky130_fd_sc_hd__nand3_1 U28779 ( .A(n24148), .B(n24147), .C(n24146), .Y(
        j202_soc_core_ahb2apb_02_N150) );
  sky130_fd_sc_hd__a22oi_1 U28780 ( .A1(n24174), .A2(la_data_out[23]), .B1(
        n24173), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[23]), 
        .Y(n24151) );
  sky130_fd_sc_hd__a22oi_1 U28781 ( .A1(n24176), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[23]), .B1(n24175), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[23]), .Y(n24150) );
  sky130_fd_sc_hd__a22oi_1 U28782 ( .A1(n24178), .A2(gpio_en_o[23]), .B1(
        n24177), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_isr[23]), .Y(
        n24149) );
  sky130_fd_sc_hd__nand3_1 U28783 ( .A(n24151), .B(n24150), .C(n24149), .Y(
        j202_soc_core_ahb2apb_02_N151) );
  sky130_fd_sc_hd__a22oi_1 U28784 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[24]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[24]), .Y(n24154) );
  sky130_fd_sc_hd__a22oi_1 U28785 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[24]), .A2(n24176), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[24]), .B2(n24175), .Y(
        n24153) );
  sky130_fd_sc_hd__a22oi_1 U28786 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[24]), .A2(n24177), .B1(
        gpio_en_o[24]), .B2(n24178), .Y(n24152) );
  sky130_fd_sc_hd__nand3_1 U28787 ( .A(n24154), .B(n24153), .C(n24152), .Y(
        j202_soc_core_ahb2apb_02_N152) );
  sky130_fd_sc_hd__a22oi_1 U28788 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[25]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[25]), .Y(n24157) );
  sky130_fd_sc_hd__a22oi_1 U28789 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[25]), .A2(n24176), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[25]), .B2(n24175), .Y(
        n24156) );
  sky130_fd_sc_hd__a22oi_1 U28790 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[25]), .A2(n24177), .B1(
        gpio_en_o[25]), .B2(n24178), .Y(n24155) );
  sky130_fd_sc_hd__nand3_1 U28791 ( .A(n24157), .B(n24156), .C(n24155), .Y(
        j202_soc_core_ahb2apb_02_N153) );
  sky130_fd_sc_hd__a22oi_1 U28792 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[26]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[26]), .Y(n24160) );
  sky130_fd_sc_hd__a22oi_1 U28793 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[26]), .A2(n24175), .B1(
        gpio_en_o[26]), .B2(n24178), .Y(n24159) );
  sky130_fd_sc_hd__a22oi_1 U28794 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[26]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[26]), .B2(n24176), .Y(
        n24158) );
  sky130_fd_sc_hd__nand3_1 U28795 ( .A(n24160), .B(n24159), .C(n24158), .Y(
        j202_soc_core_ahb2apb_02_N154) );
  sky130_fd_sc_hd__a22oi_1 U28796 ( .A1(n24174), .A2(la_data_out[27]), .B1(
        n24173), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[27]), 
        .Y(n24163) );
  sky130_fd_sc_hd__a22oi_1 U28797 ( .A1(n24175), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[27]), .B1(n24177), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[27]), .Y(n24162) );
  sky130_fd_sc_hd__a22oi_1 U28798 ( .A1(n24176), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[27]), .B1(n24178), .B2(
        gpio_en_o[27]), .Y(n24161) );
  sky130_fd_sc_hd__nand3_1 U28799 ( .A(n24163), .B(n24162), .C(n24161), .Y(
        j202_soc_core_ahb2apb_02_N155) );
  sky130_fd_sc_hd__a22oi_1 U28800 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[28]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[28]), .Y(n24166) );
  sky130_fd_sc_hd__a22oi_1 U28801 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[28]), .A2(n24176), .B1(
        gpio_en_o[28]), .B2(n24178), .Y(n24165) );
  sky130_fd_sc_hd__a22oi_1 U28802 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[28]), .A2(n24177), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[28]), .B2(n24175), .Y(
        n24164) );
  sky130_fd_sc_hd__nand3_1 U28803 ( .A(n24166), .B(n24165), .C(n24164), .Y(
        j202_soc_core_ahb2apb_02_N156) );
  sky130_fd_sc_hd__a22oi_1 U28804 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[29]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[29]), .Y(n24169) );
  sky130_fd_sc_hd__a22oi_1 U28805 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[29]), .A2(n24176), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[29]), .B2(n24175), .Y(
        n24168) );
  sky130_fd_sc_hd__a22oi_1 U28806 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[29]), .A2(n24177), .B1(
        gpio_en_o[29]), .B2(n24178), .Y(n24167) );
  sky130_fd_sc_hd__nand3_1 U28807 ( .A(n24169), .B(n24168), .C(n24167), .Y(
        j202_soc_core_ahb2apb_02_N157) );
  sky130_fd_sc_hd__a22oi_1 U28808 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[30]), .A2(n24173), 
        .B1(n24174), .B2(la_data_out[30]), .Y(n24172) );
  sky130_fd_sc_hd__a22oi_1 U28809 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[30]), .A2(n24176), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[30]), .B2(n24175), .Y(
        n24171) );
  sky130_fd_sc_hd__a22oi_1 U28810 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[30]), .A2(n24177), .B1(
        gpio_en_o[30]), .B2(n24178), .Y(n24170) );
  sky130_fd_sc_hd__nand3_1 U28811 ( .A(n24172), .B(n24171), .C(n24170), .Y(
        j202_soc_core_ahb2apb_02_N158) );
  sky130_fd_sc_hd__a22oi_1 U28812 ( .A1(n24174), .A2(la_data_out[31]), .B1(
        n24173), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[31]), 
        .Y(n24181) );
  sky130_fd_sc_hd__a22oi_1 U28813 ( .A1(n24176), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[31]), .B1(n24175), .B2(
        j202_soc_core_gpio_core_00_gpio_regs_00_ier[31]), .Y(n24180) );
  sky130_fd_sc_hd__a22oi_1 U28814 ( .A1(n24178), .A2(gpio_en_o[31]), .B1(
        n24177), .B2(j202_soc_core_gpio_core_00_gpio_regs_00_isr[31]), .Y(
        n24179) );
  sky130_fd_sc_hd__nand3_1 U28815 ( .A(n24181), .B(n24180), .C(n24179), .Y(
        j202_soc_core_ahb2apb_02_N159) );
  sky130_fd_sc_hd__nand4_1 U28816 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[6]), .B(j202_soc_core_intc_core_00_cp_intack_all_0_), .C(n24244), .D(n24189), .Y(
        n24185) );
  sky130_fd_sc_hd__nor2_1 U28817 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .B(n24185), .Y(n24221) );
  sky130_fd_sc_hd__nor2_1 U28818 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]), .B(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[3]), .Y(n24258) );
  sky130_fd_sc_hd__a21oi_1 U28819 ( .A1(n24221), .A2(n24258), .B1(
        j202_soc_core_intc_core_00_rg_irqc[0]), .Y(n24183) );
  sky130_fd_sc_hd__nand2_1 U28820 ( .A(j202_soc_core_intc_core_00_rg_sint[0]), 
        .B(n25731), .Y(n24268) );
  sky130_fd_sc_hd__nor2_1 U28821 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[0]), 
        .B(n24268), .Y(n24182) );
  sky130_fd_sc_hd__a31oi_1 U28822 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[0]), .A2(n24183), .A3(n25732), 
        .B1(n24182), .Y(n24184) );
  sky130_fd_sc_hd__clkinv_1 U28823 ( .A(j202_soc_core_intc_core_00_rg_ie[0]), 
        .Y(n24410) );
  sky130_fd_sc_hd__nor2_1 U28824 ( .A(n24184), .B(n24410), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N3) );
  sky130_fd_sc_hd__clkinv_1 U28825 ( .A(n24185), .Y(n24225) );
  sky130_fd_sc_hd__a31oi_1 U28826 ( .A1(n24258), .A2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .A3(n24225), .B1(j202_soc_core_intc_core_00_rg_irqc[1]), .Y(n24187) );
  sky130_fd_sc_hd__nand2_1 U28827 ( .A(j202_soc_core_intc_core_00_rg_sint[1]), 
        .B(n25731), .Y(n24269) );
  sky130_fd_sc_hd__nor2_1 U28828 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[1]), 
        .B(n24269), .Y(n24186) );
  sky130_fd_sc_hd__a31oi_1 U28829 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[1]), .A2(n24187), .A3(n25732), 
        .B1(n24186), .Y(n24188) );
  sky130_fd_sc_hd__clkinv_1 U28830 ( .A(j202_soc_core_intc_core_00_rg_ie[1]), 
        .Y(n24411) );
  sky130_fd_sc_hd__nor2_1 U28831 ( .A(n24188), .B(n24411), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N4) );
  sky130_fd_sc_hd__nand4_1 U28832 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[1]), .B(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[6]), .C(j202_soc_core_intc_core_00_cp_intack_all_0_), .D(n24189), .Y(n24193) );
  sky130_fd_sc_hd__nor2_1 U28833 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .B(n24193), .Y(n24229) );
  sky130_fd_sc_hd__a21oi_1 U28834 ( .A1(n24229), .A2(n24258), .B1(
        j202_soc_core_intc_core_00_rg_irqc[2]), .Y(n24191) );
  sky130_fd_sc_hd__nand2_1 U28835 ( .A(j202_soc_core_intc_core_00_rg_sint[2]), 
        .B(n25731), .Y(n24270) );
  sky130_fd_sc_hd__nor2_1 U28836 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[2]), 
        .B(n24270), .Y(n24190) );
  sky130_fd_sc_hd__a31oi_1 U28837 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[2]), .A2(n24191), .A3(n25732), 
        .B1(n24190), .Y(n24192) );
  sky130_fd_sc_hd__clkinv_1 U28838 ( .A(j202_soc_core_intc_core_00_rg_ie[2]), 
        .Y(n24412) );
  sky130_fd_sc_hd__nor2_1 U28839 ( .A(n24192), .B(n24412), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N5) );
  sky130_fd_sc_hd__clkinv_1 U28840 ( .A(n24193), .Y(n24233) );
  sky130_fd_sc_hd__a31oi_1 U28841 ( .A1(n24258), .A2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .A3(n24233), .B1(j202_soc_core_intc_core_00_rg_irqc[3]), .Y(n24195) );
  sky130_fd_sc_hd__nand2_1 U28842 ( .A(j202_soc_core_intc_core_00_rg_sint[3]), 
        .B(n25731), .Y(n24271) );
  sky130_fd_sc_hd__nor2_1 U28843 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[3]), 
        .B(n24271), .Y(n24194) );
  sky130_fd_sc_hd__a31oi_1 U28844 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[3]), .A2(n24195), .A3(n25732), 
        .B1(n24194), .Y(n24196) );
  sky130_fd_sc_hd__clkinv_1 U28845 ( .A(j202_soc_core_intc_core_00_rg_ie[3]), 
        .Y(n24413) );
  sky130_fd_sc_hd__nor2_1 U28846 ( .A(n24196), .B(n24413), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N6) );
  sky130_fd_sc_hd__nor2_1 U28847 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[3]), .B(n24238), .Y(n24205) );
  sky130_fd_sc_hd__a21oi_1 U28848 ( .A1(n24205), .A2(n24221), .B1(
        j202_soc_core_intc_core_00_rg_irqc[4]), .Y(n24198) );
  sky130_fd_sc_hd__nand2_1 U28849 ( .A(j202_soc_core_intc_core_00_rg_sint[4]), 
        .B(n25731), .Y(n24272) );
  sky130_fd_sc_hd__nor2_1 U28850 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[4]), 
        .B(n24272), .Y(n24197) );
  sky130_fd_sc_hd__a31oi_1 U28851 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[4]), .A2(n24198), .A3(n25732), 
        .B1(n24197), .Y(n24199) );
  sky130_fd_sc_hd__clkinv_1 U28852 ( .A(j202_soc_core_intc_core_00_rg_ie[4]), 
        .Y(n24414) );
  sky130_fd_sc_hd__nor2_1 U28853 ( .A(n24199), .B(n24414), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N7) );
  sky130_fd_sc_hd__a31oi_1 U28854 ( .A1(n24225), .A2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .A3(n24205), .B1(j202_soc_core_intc_core_00_rg_irqc[5]), .Y(n24201) );
  sky130_fd_sc_hd__nand2_1 U28855 ( .A(j202_soc_core_intc_core_00_rg_sint[5]), 
        .B(n25731), .Y(n24273) );
  sky130_fd_sc_hd__nor2_1 U28856 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[5]), 
        .B(n24273), .Y(n24200) );
  sky130_fd_sc_hd__a31oi_1 U28857 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[5]), .A2(n24201), .A3(n25732), 
        .B1(n24200), .Y(n24202) );
  sky130_fd_sc_hd__clkinv_1 U28858 ( .A(j202_soc_core_intc_core_00_rg_ie[5]), 
        .Y(n24415) );
  sky130_fd_sc_hd__nor2_1 U28859 ( .A(n24202), .B(n24415), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N8) );
  sky130_fd_sc_hd__nand2_1 U28860 ( .A(j202_soc_core_intc_core_00_rg_sint[6]), 
        .B(n25732), .Y(n24274) );
  sky130_fd_sc_hd__a21oi_1 U28861 ( .A1(n24205), .A2(n24229), .B1(
        j202_soc_core_intc_core_00_rg_irqc[6]), .Y(n24203) );
  sky130_fd_sc_hd__nand3_1 U28862 ( .A(j202_soc_core_intc_core_00_in_intreq[6]), .B(n24203), .C(n25732), .Y(n24204) );
  sky130_fd_sc_hd__clkinv_1 U28863 ( .A(j202_soc_core_intc_core_00_rg_ie[6]), 
        .Y(n24416) );
  sky130_fd_sc_hd__a221oi_1 U28864 ( .A1(n24274), .A2(n24204), .B1(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[6]), 
        .B2(n24204), .C1(n24416), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N9) );
  sky130_fd_sc_hd__a31oi_1 U28865 ( .A1(n24233), .A2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .A3(n24205), .B1(j202_soc_core_intc_core_00_rg_irqc[7]), .Y(n24207) );
  sky130_fd_sc_hd__nand2_1 U28866 ( .A(j202_soc_core_intc_core_00_rg_sint[7]), 
        .B(n25731), .Y(n24275) );
  sky130_fd_sc_hd__nor2_1 U28867 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[7]), 
        .B(n24275), .Y(n24206) );
  sky130_fd_sc_hd__a31oi_1 U28868 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[7]), .A2(n24207), .A3(n25732), 
        .B1(n24206), .Y(n24208) );
  sky130_fd_sc_hd__clkinv_1 U28869 ( .A(j202_soc_core_intc_core_00_rg_ie[7]), 
        .Y(n24417) );
  sky130_fd_sc_hd__nor2_1 U28870 ( .A(n24208), .B(n24417), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N10) );
  sky130_fd_sc_hd__nor2_1 U28871 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]), .B(n24237), .Y(n24217) );
  sky130_fd_sc_hd__a21oi_1 U28872 ( .A1(n24217), .A2(n24221), .B1(
        j202_soc_core_intc_core_00_rg_irqc[8]), .Y(n24210) );
  sky130_fd_sc_hd__nand2_1 U28873 ( .A(j202_soc_core_intc_core_00_rg_sint[8]), 
        .B(n25731), .Y(n24276) );
  sky130_fd_sc_hd__nor2_1 U28874 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[8]), 
        .B(n24276), .Y(n24209) );
  sky130_fd_sc_hd__a31oi_1 U28875 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[8]), .A2(n24210), .A3(n25732), 
        .B1(n24209), .Y(n24211) );
  sky130_fd_sc_hd__clkinv_1 U28876 ( .A(j202_soc_core_intc_core_00_rg_ie[8]), 
        .Y(n24419) );
  sky130_fd_sc_hd__nor2_1 U28877 ( .A(n24211), .B(n24419), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N11) );
  sky130_fd_sc_hd__a31oi_1 U28878 ( .A1(n24225), .A2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .A3(n24217), .B1(j202_soc_core_intc_core_00_rg_irqc[9]), .Y(n24213) );
  sky130_fd_sc_hd__nand2_1 U28879 ( .A(j202_soc_core_intc_core_00_rg_sint[9]), 
        .B(n25731), .Y(n24277) );
  sky130_fd_sc_hd__nor2_1 U28880 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[9]), 
        .B(n24277), .Y(n24212) );
  sky130_fd_sc_hd__a31oi_1 U28881 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[9]), .A2(n24213), .A3(n25732), 
        .B1(n24212), .Y(n24214) );
  sky130_fd_sc_hd__clkinv_1 U28882 ( .A(j202_soc_core_intc_core_00_rg_ie[9]), 
        .Y(n24421) );
  sky130_fd_sc_hd__nor2_1 U28883 ( .A(n24214), .B(n24421), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N12) );
  sky130_fd_sc_hd__nand2_1 U28884 ( .A(j202_soc_core_intc_core_00_rg_sint[10]), 
        .B(n25732), .Y(n24278) );
  sky130_fd_sc_hd__a21oi_1 U28885 ( .A1(n24217), .A2(n24229), .B1(
        j202_soc_core_intc_core_00_rg_irqc[10]), .Y(n24215) );
  sky130_fd_sc_hd__nand3_1 U28886 ( .A(
        j202_soc_core_intc_core_00_in_intreq[10]), .B(n24215), .C(n25734), .Y(
        n24216) );
  sky130_fd_sc_hd__clkinv_1 U28887 ( .A(j202_soc_core_intc_core_00_rg_ie[10]), 
        .Y(n24423) );
  sky130_fd_sc_hd__a221oi_1 U28888 ( .A1(n24278), .A2(n24216), .B1(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[10]), 
        .B2(n24216), .C1(n24423), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N13) );
  sky130_fd_sc_hd__a31oi_1 U28889 ( .A1(n24233), .A2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .A3(n24217), .B1(j202_soc_core_intc_core_00_rg_irqc[11]), .Y(n24219) );
  sky130_fd_sc_hd__nand2_1 U28890 ( .A(j202_soc_core_intc_core_00_rg_sint[11]), 
        .B(n25731), .Y(n24279) );
  sky130_fd_sc_hd__nor2_1 U28891 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[11]), 
        .B(n24279), .Y(n24218) );
  sky130_fd_sc_hd__a31oi_1 U28892 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[11]), .A2(n24219), .A3(n25732), 
        .B1(n24218), .Y(n24220) );
  sky130_fd_sc_hd__clkinv_1 U28893 ( .A(j202_soc_core_intc_core_00_rg_ie[11]), 
        .Y(n24425) );
  sky130_fd_sc_hd__nor2_1 U28894 ( .A(n24220), .B(n24425), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N14) );
  sky130_fd_sc_hd__nor2_1 U28895 ( .A(n24238), .B(n24237), .Y(n24232) );
  sky130_fd_sc_hd__a21oi_1 U28896 ( .A1(n24232), .A2(n24221), .B1(
        j202_soc_core_intc_core_00_rg_irqc[12]), .Y(n24223) );
  sky130_fd_sc_hd__nand2_1 U28897 ( .A(j202_soc_core_intc_core_00_rg_sint[12]), 
        .B(n25731), .Y(n24280) );
  sky130_fd_sc_hd__nor2_1 U28898 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[12]), 
        .B(n24280), .Y(n24222) );
  sky130_fd_sc_hd__a31oi_1 U28899 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[12]), .A2(n24223), .A3(n25732), 
        .B1(n24222), .Y(n24224) );
  sky130_fd_sc_hd__clkinv_1 U28900 ( .A(j202_soc_core_intc_core_00_rg_ie[12]), 
        .Y(n24427) );
  sky130_fd_sc_hd__nor2_1 U28901 ( .A(n24224), .B(n24427), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N15) );
  sky130_fd_sc_hd__a31oi_1 U28902 ( .A1(n24225), .A2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .A3(n24232), .B1(j202_soc_core_intc_core_00_rg_irqc[13]), .Y(n24227) );
  sky130_fd_sc_hd__nand2_1 U28903 ( .A(j202_soc_core_intc_core_00_rg_sint[13]), 
        .B(n25731), .Y(n24281) );
  sky130_fd_sc_hd__nor2_1 U28904 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[13]), 
        .B(n24281), .Y(n24226) );
  sky130_fd_sc_hd__a31oi_1 U28905 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[13]), .A2(n24227), .A3(n25732), 
        .B1(n24226), .Y(n24228) );
  sky130_fd_sc_hd__clkinv_1 U28906 ( .A(j202_soc_core_intc_core_00_rg_ie[13]), 
        .Y(n24429) );
  sky130_fd_sc_hd__nor2_1 U28907 ( .A(n24228), .B(n24429), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N16) );
  sky130_fd_sc_hd__nand2_1 U28908 ( .A(j202_soc_core_intc_core_00_rg_sint[14]), 
        .B(n25732), .Y(n24282) );
  sky130_fd_sc_hd__a21oi_1 U28909 ( .A1(n24232), .A2(n24229), .B1(
        j202_soc_core_intc_core_00_rg_irqc[14]), .Y(n24230) );
  sky130_fd_sc_hd__nand3_1 U28910 ( .A(
        j202_soc_core_intc_core_00_in_intreq[14]), .B(n24230), .C(n25734), .Y(
        n24231) );
  sky130_fd_sc_hd__clkinv_1 U28911 ( .A(j202_soc_core_intc_core_00_rg_ie[14]), 
        .Y(n24431) );
  sky130_fd_sc_hd__a221oi_1 U28912 ( .A1(n24282), .A2(n24231), .B1(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[14]), 
        .B2(n24231), .C1(n24431), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N17) );
  sky130_fd_sc_hd__a31oi_1 U28913 ( .A1(n24233), .A2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .A3(n24232), .B1(j202_soc_core_intc_core_00_rg_irqc[15]), .Y(n24235) );
  sky130_fd_sc_hd__nand2_1 U28914 ( .A(j202_soc_core_intc_core_00_rg_sint[15]), 
        .B(n25731), .Y(n24283) );
  sky130_fd_sc_hd__nor2_1 U28915 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[15]), 
        .B(n24283), .Y(n24234) );
  sky130_fd_sc_hd__a31oi_1 U28916 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[15]), .A2(n24235), .A3(n25732), 
        .B1(n24234), .Y(n24236) );
  sky130_fd_sc_hd__clkinv_1 U28917 ( .A(j202_soc_core_intc_core_00_rg_ie[15]), 
        .Y(n24433) );
  sky130_fd_sc_hd__nor2_1 U28918 ( .A(n24236), .B(n24433), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N18) );
  sky130_fd_sc_hd__nand3_1 U28919 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[4]), .B(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[6]), .C(j202_soc_core_intc_core_00_cp_intack_all_0_), .Y(n24243) );
  sky130_fd_sc_hd__nor2_1 U28920 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .B(n24243), .Y(n24257) );
  sky130_fd_sc_hd__and3_1 U28921 ( .A(n24257), .B(n24244), .C(n24237), .X(
        n24265) );
  sky130_fd_sc_hd__a21oi_1 U28922 ( .A1(n24265), .A2(n24238), .B1(
        j202_soc_core_intc_core_00_rg_irqc[16]), .Y(n24240) );
  sky130_fd_sc_hd__nand3_1 U28923 ( .A(n25734), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[6]), .C(
        j202_soc_core_cmt_core_00_cmf0), .Y(n24284) );
  sky130_fd_sc_hd__nor2_1 U28924 ( .A(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[16]), 
        .B(n24284), .Y(n24239) );
  sky130_fd_sc_hd__a31oi_1 U28925 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[16]), .A2(n24240), .A3(n25732), 
        .B1(n24239), .Y(n24241) );
  sky130_fd_sc_hd__clkinv_1 U28926 ( .A(j202_soc_core_intc_core_00_rg_ie[16]), 
        .Y(n24435) );
  sky130_fd_sc_hd__nor2_1 U28927 ( .A(n24241), .B(n24435), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N19) );
  sky130_fd_sc_hd__nand2_1 U28928 ( .A(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[0]), .B(n24258), .Y(n24242) );
  sky130_fd_sc_hd__nor2_1 U28929 ( .A(n24243), .B(n24242), .Y(n24262) );
  sky130_fd_sc_hd__a21oi_1 U28930 ( .A1(n24262), .A2(n24244), .B1(
        j202_soc_core_intc_core_00_rg_irqc[17]), .Y(n24245) );
  sky130_fd_sc_hd__nand3_1 U28931 ( .A(
        j202_soc_core_intc_core_00_in_intreq[17]), .B(n24245), .C(n25734), .Y(
        n24246) );
  sky130_fd_sc_hd__nand3_1 U28932 ( .A(n25734), .B(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[6]), .C(
        j202_soc_core_cmt_core_00_cmf1), .Y(n24285) );
  sky130_fd_sc_hd__clkinv_1 U28933 ( .A(j202_soc_core_intc_core_00_rg_ie[17]), 
        .Y(n24437) );
  sky130_fd_sc_hd__a221oi_1 U28934 ( .A1(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[17]), 
        .A2(n24246), .B1(n24285), .B2(n24246), .C1(n24437), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N20) );
  sky130_fd_sc_hd__nor4_1 U28935 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[1]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[3]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[2]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[31]), .Y(n24250) );
  sky130_fd_sc_hd__nor4_1 U28936 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[5]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[6]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[7]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[9]), .Y(n24249) );
  sky130_fd_sc_hd__nor4_1 U28937 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[0]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[4]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[8]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[12]), .Y(n24248) );
  sky130_fd_sc_hd__nor4_1 U28938 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[16]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[20]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[24]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[28]), .Y(n24247) );
  sky130_fd_sc_hd__nand4_1 U28939 ( .A(n24250), .B(n24249), .C(n24248), .D(
        n24247), .Y(n24256) );
  sky130_fd_sc_hd__nor4_1 U28940 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[22]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[25]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[21]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[23]), .Y(n24254) );
  sky130_fd_sc_hd__nor4_1 U28941 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[26]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[29]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[30]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[27]), .Y(n24253) );
  sky130_fd_sc_hd__nor4_1 U28942 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[10]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[11]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[13]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[14]), .Y(n24252) );
  sky130_fd_sc_hd__nor4_1 U28943 ( .A(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[15]), .B(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[17]), .C(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[18]), .D(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[19]), .Y(n24251) );
  sky130_fd_sc_hd__nand4_1 U28944 ( .A(n24254), .B(n24253), .C(n24252), .D(
        n24251), .Y(n24255) );
  sky130_fd_sc_hd__a31oi_1 U28946 ( .A1(n24258), .A2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[1]), .A3(n24257), .B1(j202_soc_core_intc_core_00_rg_irqc[18]), .Y(n24259) );
  sky130_fd_sc_hd__nand3_1 U28947 ( .A(
        j202_soc_core_intc_core_00_in_intreq[18]), .B(n24259), .C(n25732), .Y(
        n24260) );
  sky130_fd_sc_hd__clkinv_1 U28948 ( .A(j202_soc_core_intc_core_00_rg_ie[18]), 
        .Y(n24439) );
  sky130_fd_sc_hd__a221oi_1 U28949 ( .A1(n24261), .A2(n24260), .B1(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[18]), 
        .B2(n24260), .C1(n24439), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N21) );
  sky130_fd_sc_hd__nand2_1 U28950 ( .A(j202_soc_core_bldc_int), .B(n25732), 
        .Y(n24286) );
  sky130_fd_sc_hd__a21oi_1 U28951 ( .A1(n24262), .A2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[1]), .B1(j202_soc_core_intc_core_00_rg_irqc[19]), .Y(n24263) );
  sky130_fd_sc_hd__nand3_1 U28952 ( .A(
        j202_soc_core_intc_core_00_in_intreq[19]), .B(n24263), .C(n25734), .Y(
        n24264) );
  sky130_fd_sc_hd__clkinv_1 U28953 ( .A(j202_soc_core_intc_core_00_rg_ie[19]), 
        .Y(n24441) );
  sky130_fd_sc_hd__a221oi_1 U28954 ( .A1(n24286), .A2(n24264), .B1(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[19]), 
        .B2(n24264), .C1(n24441), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N22) );
  sky130_fd_sc_hd__nand2_1 U28955 ( .A(j202_soc_core_qspi_int), .B(n25732), 
        .Y(n24287) );
  sky130_fd_sc_hd__a21oi_1 U28956 ( .A1(n24265), .A2(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_intr_vec_latch[2]), .B1(j202_soc_core_intc_core_00_rg_irqc[20]), .Y(n24266) );
  sky130_fd_sc_hd__nand3_1 U28957 ( .A(
        j202_soc_core_intc_core_00_in_intreq[20]), .B(n24266), .C(n25734), .Y(
        n24267) );
  sky130_fd_sc_hd__clkinv_1 U28958 ( .A(j202_soc_core_intc_core_00_rg_ie[20]), 
        .Y(n24445) );
  sky130_fd_sc_hd__a221oi_1 U28959 ( .A1(n24287), .A2(n24267), .B1(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_normal_int[20]), 
        .B2(n24267), .C1(n24445), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_intreq_N23) );
  sky130_fd_sc_hd__clkinv_1 U28960 ( .A(n24268), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N3) );
  sky130_fd_sc_hd__clkinv_1 U28961 ( .A(n24269), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N4) );
  sky130_fd_sc_hd__clkinv_1 U28962 ( .A(n24270), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N5) );
  sky130_fd_sc_hd__clkinv_1 U28963 ( .A(n24271), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N6) );
  sky130_fd_sc_hd__clkinv_1 U28964 ( .A(n24272), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N7) );
  sky130_fd_sc_hd__clkinv_1 U28965 ( .A(n24273), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N8) );
  sky130_fd_sc_hd__clkinv_1 U28966 ( .A(n24274), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N9) );
  sky130_fd_sc_hd__clkinv_1 U28967 ( .A(n24275), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N10) );
  sky130_fd_sc_hd__clkinv_1 U28968 ( .A(n24276), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N11) );
  sky130_fd_sc_hd__clkinv_1 U28969 ( .A(n24277), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N12) );
  sky130_fd_sc_hd__clkinv_1 U28970 ( .A(n24278), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N13) );
  sky130_fd_sc_hd__clkinv_1 U28971 ( .A(n24280), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N15) );
  sky130_fd_sc_hd__clkinv_1 U28972 ( .A(n24281), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N16) );
  sky130_fd_sc_hd__clkinv_1 U28973 ( .A(n24282), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N17) );
  sky130_fd_sc_hd__clkinv_1 U28974 ( .A(n24283), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N18) );
  sky130_fd_sc_hd__clkinv_1 U28975 ( .A(n24284), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N19) );
  sky130_fd_sc_hd__clkinv_1 U28976 ( .A(n24285), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N20) );
  sky130_fd_sc_hd__clkinv_1 U28977 ( .A(n24286), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N22) );
  sky130_fd_sc_hd__clkinv_1 U28978 ( .A(n24287), .Y(
        j202_soc_core_intc_core_00_intc_in_00_intc_intr_in_0_dff_normal_int_N23) );
  sky130_fd_sc_hd__a22o_1 U28979 ( .A1(n25402), .A2(n24289), .B1(
        j202_soc_core_intc_core_00_rg_itgt[106]), .B2(n24288), .X(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_1__rg_itgt_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__clkinv_1 U28980 ( .A(j202_soc_core_intc_core_00_rg_itgt[33]), .Y(n24547) );
  sky130_fd_sc_hd__o22ai_1 U28981 ( .A1(n24547), .A2(n24291), .B1(n24483), 
        .B2(n24290), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_itgt_label_0__rg_itgt_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__clkinv_1 U28982 ( .A(j202_soc_core_intc_core_00_rg_ipr[96]), 
        .Y(n24295) );
  sky130_fd_sc_hd__nand2b_1 U28983 ( .A_N(n24292), .B(n24448), .Y(n24378) );
  sky130_fd_sc_hd__nand2_1 U28984 ( .A(n24349), .B(
        j202_soc_core_intc_core_00_bs_addr[3]), .Y(n24497) );
  sky130_fd_sc_hd__nand2_1 U28985 ( .A(n24294), .B(j202_soc_core_pwrite[1]), 
        .Y(n24326) );
  sky130_fd_sc_hd__nand2_1 U28986 ( .A(n25731), .B(n24326), .Y(n24324) );
  sky130_fd_sc_hd__o22ai_1 U28987 ( .A1(n24295), .A2(n24324), .B1(n24473), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__clkinv_1 U28988 ( .A(j202_soc_core_intc_core_00_rg_ipr[97]), 
        .Y(n24296) );
  sky130_fd_sc_hd__o22ai_1 U28989 ( .A1(n24296), .A2(n24324), .B1(n24475), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__clkinv_1 U28990 ( .A(j202_soc_core_intc_core_00_rg_ipr[98]), 
        .Y(n24297) );
  sky130_fd_sc_hd__o22ai_1 U28991 ( .A1(n24297), .A2(n24324), .B1(n24477), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__clkinv_1 U28992 ( .A(j202_soc_core_intc_core_00_rg_ipr[99]), 
        .Y(n24298) );
  sky130_fd_sc_hd__o22ai_1 U28993 ( .A1(n24298), .A2(n24324), .B1(n24479), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__clkinv_1 U28994 ( .A(j202_soc_core_intc_core_00_rg_ipr[100]), .Y(n24299) );
  sky130_fd_sc_hd__o22ai_1 U28995 ( .A1(n24299), .A2(n24324), .B1(n24326), 
        .B2(n24481), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__clkinv_1 U28996 ( .A(j202_soc_core_intc_core_00_rg_ipr[101]), .Y(n24300) );
  sky130_fd_sc_hd__o22ai_1 U28997 ( .A1(n24300), .A2(n24324), .B1(n24483), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__clkinv_1 U28998 ( .A(j202_soc_core_intc_core_00_rg_ipr[102]), .Y(n24301) );
  sky130_fd_sc_hd__o22ai_1 U28999 ( .A1(n24301), .A2(n24324), .B1(n24485), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__clkinv_1 U29000 ( .A(j202_soc_core_intc_core_00_rg_ipr[103]), .Y(n24302) );
  sky130_fd_sc_hd__o22ai_1 U29001 ( .A1(n24302), .A2(n24324), .B1(n24488), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__clkinv_1 U29002 ( .A(j202_soc_core_intc_core_00_rg_ipr[104]), .Y(n24303) );
  sky130_fd_sc_hd__o22ai_1 U29003 ( .A1(n24303), .A2(n24324), .B1(n24326), 
        .B2(n24418), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__clkinv_1 U29004 ( .A(j202_soc_core_intc_core_00_rg_ipr[105]), .Y(n24304) );
  sky130_fd_sc_hd__o22ai_1 U29005 ( .A1(n24304), .A2(n24324), .B1(n24420), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__clkinv_1 U29006 ( .A(j202_soc_core_intc_core_00_rg_ipr[106]), .Y(n24305) );
  sky130_fd_sc_hd__o22ai_1 U29007 ( .A1(n24305), .A2(n24324), .B1(n24422), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__clkinv_1 U29008 ( .A(j202_soc_core_intc_core_00_rg_ipr[107]), .Y(n24306) );
  sky130_fd_sc_hd__o22ai_1 U29009 ( .A1(n24306), .A2(n24324), .B1(n24424), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__clkinv_1 U29010 ( .A(j202_soc_core_intc_core_00_rg_ipr[108]), .Y(n24307) );
  sky130_fd_sc_hd__o22ai_1 U29011 ( .A1(n24307), .A2(n24324), .B1(n24326), 
        .B2(n24426), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__clkinv_1 U29012 ( .A(j202_soc_core_intc_core_00_rg_ipr[109]), .Y(n24308) );
  sky130_fd_sc_hd__o22ai_1 U29013 ( .A1(n24308), .A2(n24324), .B1(n24428), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__clkinv_1 U29014 ( .A(j202_soc_core_intc_core_00_rg_ipr[110]), .Y(n24309) );
  sky130_fd_sc_hd__o22ai_1 U29015 ( .A1(n24309), .A2(n24324), .B1(n24430), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__clkinv_1 U29016 ( .A(j202_soc_core_intc_core_00_rg_ipr[111]), .Y(n24650) );
  sky130_fd_sc_hd__o22ai_1 U29017 ( .A1(n24650), .A2(n24324), .B1(n24432), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__clkinv_1 U29018 ( .A(j202_soc_core_intc_core_00_rg_ipr[112]), .Y(n24310) );
  sky130_fd_sc_hd__o22ai_1 U29019 ( .A1(n24310), .A2(n24324), .B1(n24326), 
        .B2(n24434), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__clkinv_1 U29020 ( .A(j202_soc_core_intc_core_00_rg_ipr[113]), .Y(n24311) );
  sky130_fd_sc_hd__o22ai_1 U29021 ( .A1(n24311), .A2(n24324), .B1(n24436), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__clkinv_1 U29022 ( .A(j202_soc_core_intc_core_00_rg_ipr[114]), .Y(n24312) );
  sky130_fd_sc_hd__o22ai_1 U29023 ( .A1(n24312), .A2(n24324), .B1(n24438), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__clkinv_1 U29024 ( .A(j202_soc_core_intc_core_00_rg_ipr[115]), .Y(n24313) );
  sky130_fd_sc_hd__o22ai_1 U29025 ( .A1(n24313), .A2(n24324), .B1(n24440), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__clkinv_1 U29026 ( .A(j202_soc_core_intc_core_00_rg_ipr[116]), .Y(n24314) );
  sky130_fd_sc_hd__o22ai_1 U29027 ( .A1(n24314), .A2(n24324), .B1(n24326), 
        .B2(n24443), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__clkinv_1 U29028 ( .A(j202_soc_core_intc_core_00_rg_ipr[117]), .Y(n24315) );
  sky130_fd_sc_hd__o22ai_1 U29029 ( .A1(n24315), .A2(n24324), .B1(n24387), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__clkinv_1 U29030 ( .A(j202_soc_core_intc_core_00_rg_ipr[118]), .Y(n24704) );
  sky130_fd_sc_hd__o22ai_1 U29031 ( .A1(n24704), .A2(n24324), .B1(n24389), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__clkinv_1 U29032 ( .A(j202_soc_core_intc_core_00_rg_ipr[119]), .Y(n24316) );
  sky130_fd_sc_hd__o22ai_1 U29033 ( .A1(n24316), .A2(n24324), .B1(n24390), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__clkinv_1 U29034 ( .A(j202_soc_core_intc_core_00_rg_ipr[120]), .Y(n24317) );
  sky130_fd_sc_hd__o22ai_1 U29035 ( .A1(n24317), .A2(n24324), .B1(n24326), 
        .B2(n24392), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__clkinv_1 U29036 ( .A(j202_soc_core_intc_core_00_rg_ipr[121]), .Y(n24318) );
  sky130_fd_sc_hd__o22ai_1 U29037 ( .A1(n24318), .A2(n24324), .B1(n24393), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__clkinv_1 U29038 ( .A(j202_soc_core_intc_core_00_rg_ipr[122]), .Y(n24319) );
  sky130_fd_sc_hd__o22ai_1 U29039 ( .A1(n24319), .A2(n24324), .B1(n24395), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__clkinv_1 U29040 ( .A(j202_soc_core_intc_core_00_rg_ipr[123]), .Y(n24320) );
  sky130_fd_sc_hd__o22ai_1 U29041 ( .A1(n24320), .A2(n24324), .B1(n24397), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__clkinv_1 U29042 ( .A(j202_soc_core_intc_core_00_rg_ipr[124]), .Y(n24321) );
  sky130_fd_sc_hd__o22ai_1 U29043 ( .A1(n24321), .A2(n24324), .B1(n24326), 
        .B2(n24399), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__clkinv_1 U29044 ( .A(j202_soc_core_intc_core_00_rg_ipr[125]), .Y(n24322) );
  sky130_fd_sc_hd__o22ai_1 U29045 ( .A1(n24322), .A2(n24324), .B1(n24400), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__clkinv_1 U29046 ( .A(j202_soc_core_intc_core_00_rg_ipr[126]), .Y(n24323) );
  sky130_fd_sc_hd__o22ai_1 U29047 ( .A1(n24323), .A2(n24324), .B1(n24402), 
        .B2(n24326), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__clkinv_1 U29048 ( .A(j202_soc_core_intc_core_00_rg_ipr[127]), .Y(n24325) );
  sky130_fd_sc_hd__o22ai_1 U29049 ( .A1(n24405), .A2(n24326), .B1(n24325), 
        .B2(n24324), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_3__rg_ipr_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__nor2_1 U29050 ( .A(n24327), .B(n24378), .Y(n24577) );
  sky130_fd_sc_hd__nand2_1 U29051 ( .A(n24577), .B(j202_soc_core_pwrite[1]), 
        .Y(n24348) );
  sky130_fd_sc_hd__nand2_1 U29052 ( .A(n25731), .B(n24348), .Y(n24346) );
  sky130_fd_sc_hd__a22oi_1 U29053 ( .A1(n24501), .A2(n24348), .B1(n24473), 
        .B2(n24346), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U29054 ( .A1(n24511), .A2(n24346), .B1(n24475), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U29055 ( .A1(n24521), .A2(n24346), .B1(n24477), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U29056 ( .A1(n24531), .A2(n24346), .B1(n24479), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U29057 ( .A1(n24328), .A2(n24346), .B1(n24481), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U29058 ( .A1(n24329), .A2(n24346), .B1(n24483), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U29059 ( .A1(n24562), .A2(n24346), .B1(n24485), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U29060 ( .A1(n24330), .A2(n24346), .B1(n24488), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U29061 ( .A1(n24589), .A2(n24346), .B1(n24418), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U29062 ( .A1(n24597), .A2(n24346), .B1(n24420), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U29063 ( .A1(n24606), .A2(n24346), .B1(n24422), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o22ai_1 U29064 ( .A1(n24616), .A2(n24346), .B1(n24424), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U29065 ( .A1(n24626), .A2(n24346), .B1(n24426), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U29066 ( .A1(n24633), .A2(n24346), .B1(n24428), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U29067 ( .A1(n24642), .A2(n24346), .B1(n24430), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U29068 ( .A1(n24331), .A2(n24346), .B1(n24432), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__clkinv_1 U29069 ( .A(j202_soc_core_intc_core_00_rg_ipr[80]), 
        .Y(n24332) );
  sky130_fd_sc_hd__o22ai_1 U29070 ( .A1(n24332), .A2(n24346), .B1(n24434), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U29071 ( .A1(n24333), .A2(n24346), .B1(n24436), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U29072 ( .A1(n24334), .A2(n24346), .B1(n24438), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U29073 ( .A1(n24682), .A2(n24346), .B1(n24440), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__clkinv_1 U29074 ( .A(j202_soc_core_intc_core_00_rg_ipr[84]), 
        .Y(n24335) );
  sky130_fd_sc_hd__o22ai_1 U29075 ( .A1(n24335), .A2(n24346), .B1(n24443), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__clkinv_1 U29076 ( .A(j202_soc_core_intc_core_00_rg_ipr[85]), 
        .Y(n24336) );
  sky130_fd_sc_hd__o22ai_1 U29077 ( .A1(n24336), .A2(n24346), .B1(n24387), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__clkinv_1 U29078 ( .A(j202_soc_core_intc_core_00_rg_ipr[86]), 
        .Y(n24337) );
  sky130_fd_sc_hd__o22ai_1 U29079 ( .A1(n24337), .A2(n24346), .B1(n24389), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__clkinv_1 U29080 ( .A(j202_soc_core_intc_core_00_rg_ipr[87]), 
        .Y(n24338) );
  sky130_fd_sc_hd__o22ai_1 U29081 ( .A1(n24338), .A2(n24346), .B1(n24390), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__clkinv_1 U29082 ( .A(j202_soc_core_intc_core_00_rg_ipr[88]), 
        .Y(n24339) );
  sky130_fd_sc_hd__o22ai_1 U29083 ( .A1(n24339), .A2(n24346), .B1(n24392), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__clkinv_1 U29084 ( .A(j202_soc_core_intc_core_00_rg_ipr[89]), 
        .Y(n24340) );
  sky130_fd_sc_hd__o22ai_1 U29085 ( .A1(n24340), .A2(n24346), .B1(n24393), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__clkinv_1 U29086 ( .A(j202_soc_core_intc_core_00_rg_ipr[90]), 
        .Y(n24341) );
  sky130_fd_sc_hd__o22ai_1 U29087 ( .A1(n24341), .A2(n24346), .B1(n24395), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__clkinv_1 U29088 ( .A(j202_soc_core_intc_core_00_rg_ipr[91]), 
        .Y(n24342) );
  sky130_fd_sc_hd__o22ai_1 U29089 ( .A1(n24342), .A2(n24346), .B1(n24397), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__clkinv_1 U29090 ( .A(j202_soc_core_intc_core_00_rg_ipr[92]), 
        .Y(n24343) );
  sky130_fd_sc_hd__o22ai_1 U29091 ( .A1(n24343), .A2(n24346), .B1(n24399), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__clkinv_1 U29092 ( .A(j202_soc_core_intc_core_00_rg_ipr[93]), 
        .Y(n24344) );
  sky130_fd_sc_hd__o22ai_1 U29093 ( .A1(n24344), .A2(n24346), .B1(n24400), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__clkinv_1 U29094 ( .A(j202_soc_core_intc_core_00_rg_ipr[94]), 
        .Y(n24345) );
  sky130_fd_sc_hd__o22ai_1 U29095 ( .A1(n24345), .A2(n24346), .B1(n24402), 
        .B2(n24348), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__clkinv_1 U29096 ( .A(j202_soc_core_intc_core_00_rg_ipr[95]), 
        .Y(n24347) );
  sky130_fd_sc_hd__o22ai_1 U29097 ( .A1(n24405), .A2(n24348), .B1(n24347), 
        .B2(n24346), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_2__rg_ipr_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__nand2_1 U29098 ( .A(n24349), .B(n24453), .Y(n24491) );
  sky130_fd_sc_hd__nand2_1 U29099 ( .A(n24350), .B(j202_soc_core_pwrite[1]), 
        .Y(n24375) );
  sky130_fd_sc_hd__nand2_1 U29100 ( .A(n25734), .B(n24375), .Y(n24376) );
  sky130_fd_sc_hd__o22ai_1 U29101 ( .A1(n24351), .A2(n24376), .B1(n24473), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U29102 ( .A1(n24352), .A2(n24376), .B1(n24475), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U29103 ( .A1(n24353), .A2(n24376), .B1(n24477), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U29104 ( .A1(n24354), .A2(n24376), .B1(n24479), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U29105 ( .A1(n24355), .A2(n24376), .B1(n24481), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U29106 ( .A1(n24559), .A2(n24376), .B1(n24483), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U29107 ( .A1(n24356), .A2(n24376), .B1(n24485), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U29108 ( .A1(n24357), .A2(n24376), .B1(n24488), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U29109 ( .A1(n24358), .A2(n24376), .B1(n24418), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U29110 ( .A1(n24359), .A2(n24376), .B1(n24420), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U29111 ( .A1(n24360), .A2(n24376), .B1(n24422), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o22ai_1 U29112 ( .A1(n24615), .A2(n24376), .B1(n24424), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U29113 ( .A1(n24361), .A2(n24376), .B1(n24426), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U29114 ( .A1(n24362), .A2(n24376), .B1(n24428), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U29115 ( .A1(n24363), .A2(n24376), .B1(n24430), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U29116 ( .A1(n24651), .A2(n24376), .B1(n24432), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U29117 ( .A1(n24364), .A2(n24376), .B1(n24434), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U29118 ( .A1(n24665), .A2(n24376), .B1(n24436), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U29119 ( .A1(n24365), .A2(n24376), .B1(n24438), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U29120 ( .A1(n24366), .A2(n24376), .B1(n24440), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U29121 ( .A1(n24367), .A2(n24376), .B1(n24443), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U29122 ( .A1(n24368), .A2(n24376), .B1(n24387), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U29123 ( .A1(n24702), .A2(n24376), .B1(n24389), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U29124 ( .A1(n24369), .A2(n24376), .B1(n24390), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U29125 ( .A1(n24719), .A2(n24376), .B1(n24392), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U29126 ( .A1(n24370), .A2(n24376), .B1(n24393), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U29127 ( .A1(n24371), .A2(n24376), .B1(n24395), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U29128 ( .A1(n24372), .A2(n24376), .B1(n24397), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U29129 ( .A1(n24743), .A2(n24376), .B1(n24399), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U29130 ( .A1(n24373), .A2(n24376), .B1(n24400), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U29131 ( .A1(n24374), .A2(n24376), .B1(n24402), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U29132 ( .A1(n24377), .A2(n24376), .B1(n24405), 
        .B2(n24375), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_1__rg_ipr_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__nand2_1 U29133 ( .A(n25731), .B(n24404), .Y(n24406) );
  sky130_fd_sc_hd__a22oi_1 U29134 ( .A1(n24500), .A2(n24404), .B1(n24473), 
        .B2(n24406), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U29135 ( .A1(n24510), .A2(n24406), .B1(n24475), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U29136 ( .A1(n24520), .A2(n24406), .B1(n24477), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U29137 ( .A1(n24530), .A2(n24406), .B1(n24479), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U29138 ( .A1(n24380), .A2(n24406), .B1(n24481), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U29139 ( .A1(n24381), .A2(n24406), .B1(n24483), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U29140 ( .A1(n24561), .A2(n24406), .B1(n24485), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U29141 ( .A1(n24382), .A2(n24406), .B1(n24488), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U29142 ( .A1(n24588), .A2(n24406), .B1(n24418), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U29143 ( .A1(n24600), .A2(n24406), .B1(n24420), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U29144 ( .A1(n24609), .A2(n24406), .B1(n24422), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o22ai_1 U29145 ( .A1(n24383), .A2(n24406), .B1(n24424), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U29146 ( .A1(n24623), .A2(n24406), .B1(n24426), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U29147 ( .A1(n24632), .A2(n24406), .B1(n24428), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U29148 ( .A1(n24641), .A2(n24406), .B1(n24430), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U29149 ( .A1(n24653), .A2(n24406), .B1(n24432), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U29150 ( .A1(n24384), .A2(n24406), .B1(n24434), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U29151 ( .A1(n24666), .A2(n24406), .B1(n24436), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U29152 ( .A1(n24385), .A2(n24406), .B1(n24438), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U29153 ( .A1(n24680), .A2(n24406), .B1(n24440), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U29154 ( .A1(n24386), .A2(n24406), .B1(n24443), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__o22ai_1 U29155 ( .A1(n24388), .A2(n24406), .B1(n24387), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N24) );
  sky130_fd_sc_hd__o22ai_1 U29156 ( .A1(n24706), .A2(n24406), .B1(n24389), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N25) );
  sky130_fd_sc_hd__o22ai_1 U29157 ( .A1(n24391), .A2(n24406), .B1(n24390), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N26) );
  sky130_fd_sc_hd__o22ai_1 U29158 ( .A1(n24718), .A2(n24406), .B1(n24392), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N27) );
  sky130_fd_sc_hd__o22ai_1 U29159 ( .A1(n24394), .A2(n24406), .B1(n24393), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N28) );
  sky130_fd_sc_hd__o22ai_1 U29160 ( .A1(n24396), .A2(n24406), .B1(n24395), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N29) );
  sky130_fd_sc_hd__o22ai_1 U29161 ( .A1(n24398), .A2(n24406), .B1(n24397), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N30) );
  sky130_fd_sc_hd__o22ai_1 U29162 ( .A1(n24747), .A2(n24406), .B1(n24399), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N31) );
  sky130_fd_sc_hd__o22ai_1 U29163 ( .A1(n24401), .A2(n24406), .B1(n24400), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N32) );
  sky130_fd_sc_hd__o22ai_1 U29164 ( .A1(n24403), .A2(n24406), .B1(n24402), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N33) );
  sky130_fd_sc_hd__o22ai_1 U29165 ( .A1(n24407), .A2(n24406), .B1(n24405), 
        .B2(n24404), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_ipr_label_0__rg_ipr_inst_dff_irqen_N34) );
  sky130_fd_sc_hd__nand4_1 U29166 ( .A(n24408), .B(j202_soc_core_pwrite[1]), 
        .C(j202_soc_core_intc_core_00_bs_addr[7]), .D(n24468), .Y(n24409) );
  sky130_fd_sc_hd__nor2_1 U29167 ( .A(n24473), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U29168 ( .A(n24475), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N4) );
  sky130_fd_sc_hd__nor2_1 U29169 ( .A(n24477), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N5) );
  sky130_fd_sc_hd__nor2_1 U29170 ( .A(n24479), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N6) );
  sky130_fd_sc_hd__nor2_1 U29171 ( .A(n24481), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N7) );
  sky130_fd_sc_hd__nor2_1 U29172 ( .A(n24483), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N8) );
  sky130_fd_sc_hd__nor2_1 U29173 ( .A(n24485), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N9) );
  sky130_fd_sc_hd__nor2_1 U29174 ( .A(n24488), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N10) );
  sky130_fd_sc_hd__nor2_1 U29175 ( .A(n24418), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N11) );
  sky130_fd_sc_hd__nor2_1 U29176 ( .A(n24420), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N12) );
  sky130_fd_sc_hd__nor2_1 U29177 ( .A(n24422), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N13) );
  sky130_fd_sc_hd__nor2_1 U29178 ( .A(n24424), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N14) );
  sky130_fd_sc_hd__nor2_1 U29179 ( .A(n24426), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N15) );
  sky130_fd_sc_hd__nor2_1 U29180 ( .A(n24428), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N16) );
  sky130_fd_sc_hd__nor2_1 U29181 ( .A(n24430), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N17) );
  sky130_fd_sc_hd__nor2_1 U29182 ( .A(n24432), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N18) );
  sky130_fd_sc_hd__nor2_1 U29183 ( .A(n24434), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N19) );
  sky130_fd_sc_hd__nor2_1 U29184 ( .A(n24436), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N20) );
  sky130_fd_sc_hd__nor2_1 U29185 ( .A(n24438), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N21) );
  sky130_fd_sc_hd__nor2_1 U29186 ( .A(n24440), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N22) );
  sky130_fd_sc_hd__nor2_1 U29187 ( .A(n24443), .B(n24409), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqc_label_0__rg_irqc_inst_dff_rg_N23) );
  sky130_fd_sc_hd__a22oi_1 U29188 ( .A1(n24410), .A2(n24442), .B1(n24473), 
        .B2(n24444), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__o22ai_1 U29189 ( .A1(n24411), .A2(n24444), .B1(n24475), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__o22ai_1 U29190 ( .A1(n24412), .A2(n24444), .B1(n24477), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__o22ai_1 U29191 ( .A1(n24413), .A2(n24444), .B1(n24479), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__o22ai_1 U29192 ( .A1(n24414), .A2(n24444), .B1(n24481), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__o22ai_1 U29193 ( .A1(n24415), .A2(n24444), .B1(n24483), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__o22ai_1 U29194 ( .A1(n24416), .A2(n24444), .B1(n24485), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__o22ai_1 U29195 ( .A1(n24417), .A2(n24444), .B1(n24488), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__o22ai_1 U29196 ( .A1(n24419), .A2(n24444), .B1(n24418), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N11) );
  sky130_fd_sc_hd__o22ai_1 U29197 ( .A1(n24421), .A2(n24444), .B1(n24420), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N12) );
  sky130_fd_sc_hd__o22ai_1 U29198 ( .A1(n24423), .A2(n24444), .B1(n24422), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N13) );
  sky130_fd_sc_hd__o22ai_1 U29199 ( .A1(n24425), .A2(n24444), .B1(n24424), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N14) );
  sky130_fd_sc_hd__o22ai_1 U29200 ( .A1(n24427), .A2(n24444), .B1(n24426), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N15) );
  sky130_fd_sc_hd__o22ai_1 U29201 ( .A1(n24429), .A2(n24444), .B1(n24428), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N16) );
  sky130_fd_sc_hd__o22ai_1 U29202 ( .A1(n24431), .A2(n24444), .B1(n24430), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N17) );
  sky130_fd_sc_hd__o22ai_1 U29203 ( .A1(n24433), .A2(n24444), .B1(n24432), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N18) );
  sky130_fd_sc_hd__o22ai_1 U29204 ( .A1(n24435), .A2(n24444), .B1(n24434), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N19) );
  sky130_fd_sc_hd__o22ai_1 U29205 ( .A1(n24437), .A2(n24444), .B1(n24436), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N20) );
  sky130_fd_sc_hd__o22ai_1 U29206 ( .A1(n24439), .A2(n24444), .B1(n24438), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N21) );
  sky130_fd_sc_hd__o22ai_1 U29207 ( .A1(n24441), .A2(n24444), .B1(n24440), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N22) );
  sky130_fd_sc_hd__o22ai_1 U29208 ( .A1(n24445), .A2(n24444), .B1(n24443), 
        .B2(n24442), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_irqen_label_0__rg_irqen_inst_dff_irqen_N23) );
  sky130_fd_sc_hd__nor3_1 U29209 ( .A(n24447), .B(n24473), .C(n24446), .Y(
        n24454) );
  sky130_fd_sc_hd__nand3_1 U29210 ( .A(n24454), .B(
        j202_soc_core_intc_core_00_bs_addr[2]), .C(
        j202_soc_core_intc_core_00_bs_addr[3]), .Y(n24462) );
  sky130_fd_sc_hd__clkinv_1 U29211 ( .A(j202_soc_core_intc_core_00_bs_addr[9]), 
        .Y(n24449) );
  sky130_fd_sc_hd__and3_1 U29212 ( .A(n24449), .B(n24448), .C(n24573), .X(
        n24460) );
  sky130_fd_sc_hd__nand2_1 U29213 ( .A(n24460), .B(
        j202_soc_core_intc_core_00_bs_addr[5]), .Y(n24450) );
  sky130_fd_sc_hd__nor2_1 U29214 ( .A(n24451), .B(n24450), .Y(n24472) );
  sky130_fd_sc_hd__nand2_1 U29215 ( .A(n24472), .B(n24457), .Y(n24455) );
  sky130_fd_sc_hd__nor2_1 U29216 ( .A(n24462), .B(n24455), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_15__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand2_1 U29217 ( .A(n24452), .B(n24454), .Y(n24463) );
  sky130_fd_sc_hd__nor2_1 U29218 ( .A(n24463), .B(n24455), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_14__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand3_1 U29219 ( .A(n24454), .B(
        j202_soc_core_intc_core_00_bs_addr[2]), .C(n24453), .Y(n24464) );
  sky130_fd_sc_hd__nor2_1 U29220 ( .A(n24464), .B(n24455), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_13__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand2_1 U29221 ( .A(n24469), .B(n24454), .Y(n24466) );
  sky130_fd_sc_hd__nor2_1 U29222 ( .A(n24466), .B(n24455), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_12__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U29223 ( .A(j202_soc_core_intc_core_00_bs_addr[4]), 
        .B(n24468), .Y(n24459) );
  sky130_fd_sc_hd__nand2_1 U29224 ( .A(n24472), .B(n24459), .Y(n24456) );
  sky130_fd_sc_hd__nor2_1 U29225 ( .A(n24462), .B(n24456), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_11__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U29226 ( .A(n24463), .B(n24456), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_10__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U29227 ( .A(n24464), .B(n24456), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_9__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U29228 ( .A(n24466), .B(n24456), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_8__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand3_1 U29229 ( .A(n24461), .B(n24460), .C(n24457), .Y(
        n24458) );
  sky130_fd_sc_hd__nor2_1 U29230 ( .A(n24462), .B(n24458), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_7__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U29231 ( .A(n24458), .B(n24463), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_6__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U29232 ( .A(n24458), .B(n24464), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_5__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U29233 ( .A(n24458), .B(n24466), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_4__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nand3_1 U29234 ( .A(n24461), .B(n24460), .C(n24459), .Y(
        n24465) );
  sky130_fd_sc_hd__nor2_1 U29235 ( .A(n24462), .B(n24465), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_3__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U29236 ( .A(n24463), .B(n24465), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_2__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U29237 ( .A(n24464), .B(n24465), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_1__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__nor2_1 U29238 ( .A(n24466), .B(n24465), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_sint_label_0__rg_sint_inst_dff_rg_N3) );
  sky130_fd_sc_hd__clkinv_1 U29239 ( .A(j202_soc_core_intc_core_00_rg_eimk[0]), 
        .Y(n24474) );
  sky130_fd_sc_hd__and3_1 U29240 ( .A(n24469), .B(n24468), .C(n24467), .X(
        n24470) );
  sky130_fd_sc_hd__nand3_1 U29241 ( .A(n24472), .B(n24471), .C(n24470), .Y(
        n24494) );
  sky130_fd_sc_hd__clkinv_1 U29242 ( .A(n24494), .Y(n24575) );
  sky130_fd_sc_hd__nand2_1 U29243 ( .A(n24575), .B(j202_soc_core_pwrite[1]), 
        .Y(n24487) );
  sky130_fd_sc_hd__nand2_1 U29244 ( .A(n25731), .B(n24487), .Y(n24489) );
  sky130_fd_sc_hd__o22ai_1 U29245 ( .A1(n24474), .A2(n24489), .B1(n24473), 
        .B2(n24487), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N3) );
  sky130_fd_sc_hd__clkinv_1 U29246 ( .A(j202_soc_core_intc_core_00_rg_eimk[1]), 
        .Y(n24476) );
  sky130_fd_sc_hd__o22ai_1 U29247 ( .A1(n24476), .A2(n24489), .B1(n24475), 
        .B2(n24487), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N4) );
  sky130_fd_sc_hd__clkinv_1 U29248 ( .A(j202_soc_core_intc_core_00_rg_eimk[2]), 
        .Y(n24478) );
  sky130_fd_sc_hd__o22ai_1 U29249 ( .A1(n24478), .A2(n24489), .B1(n24477), 
        .B2(n24487), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N5) );
  sky130_fd_sc_hd__clkinv_1 U29250 ( .A(j202_soc_core_intc_core_00_rg_eimk[3]), 
        .Y(n24480) );
  sky130_fd_sc_hd__o22ai_1 U29251 ( .A1(n24480), .A2(n24489), .B1(n24479), 
        .B2(n24487), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N6) );
  sky130_fd_sc_hd__clkinv_1 U29252 ( .A(j202_soc_core_intc_core_00_rg_eimk[4]), 
        .Y(n24482) );
  sky130_fd_sc_hd__o22ai_1 U29253 ( .A1(n24482), .A2(n24489), .B1(n24481), 
        .B2(n24487), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N7) );
  sky130_fd_sc_hd__clkinv_1 U29254 ( .A(j202_soc_core_intc_core_00_rg_eimk[5]), 
        .Y(n24484) );
  sky130_fd_sc_hd__o22ai_1 U29255 ( .A1(n24484), .A2(n24489), .B1(n24483), 
        .B2(n24487), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N8) );
  sky130_fd_sc_hd__clkinv_1 U29256 ( .A(j202_soc_core_intc_core_00_rg_eimk[6]), 
        .Y(n24486) );
  sky130_fd_sc_hd__o22ai_1 U29257 ( .A1(n24486), .A2(n24489), .B1(n24485), 
        .B2(n24487), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N9) );
  sky130_fd_sc_hd__clkinv_1 U29258 ( .A(j202_soc_core_intc_core_00_rg_eimk[7]), 
        .Y(n24490) );
  sky130_fd_sc_hd__o22ai_1 U29259 ( .A1(n24490), .A2(n24489), .B1(n24488), 
        .B2(n24487), .Y(
        j202_soc_core_intc_core_00_intc_regs_00_eirqmk_label_0__rg_eirqmk_inst_dff_irqen_N10) );
  sky130_fd_sc_hd__nor2_1 U29260 ( .A(j202_soc_core_rst), .B(n24492), .Y(
        n24769) );
  sky130_fd_sc_hd__a22oi_1 U29261 ( .A1(j202_soc_core_intc_core_00_rg_ipr[32]), 
        .A2(n24770), .B1(n24769), .B2(j202_soc_core_intc_core_00_rg_itgt[24]), 
        .Y(n24509) );
  sky130_fd_sc_hd__nor2_1 U29262 ( .A(j202_soc_core_rst), .B(n24493), .Y(
        n24767) );
  sky130_fd_sc_hd__nor2_1 U29263 ( .A(j202_soc_core_rst), .B(n24494), .Y(
        n24560) );
  sky130_fd_sc_hd__a22oi_1 U29264 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[0]), .B1(n24560), .B2(
        j202_soc_core_intc_core_00_rg_eimk[0]), .Y(n24508) );
  sky130_fd_sc_hd__nand2b_1 U29265 ( .A_N(n24495), .B(
        j202_soc_core_intc_core_00_bs_addr[6]), .Y(n24571) );
  sky130_fd_sc_hd__nor2_1 U29266 ( .A(j202_soc_core_rst), .B(n24571), .Y(
        n24689) );
  sky130_fd_sc_hd__nor2_1 U29268 ( .A(j202_soc_core_rst), .B(n24548), .Y(
        n24765) );
  sky130_fd_sc_hd__a22oi_1 U29269 ( .A1(j202_soc_core_intc_core_00_rg_itgt[8]), 
        .A2(n24768), .B1(n24776), .B2(j202_soc_core_intc_core_00_rg_ipr[96]), 
        .Y(n24504) );
  sky130_fd_sc_hd__nor2_1 U29270 ( .A(j202_soc_core_rst), .B(n24498), .Y(
        n24772) );
  sky130_fd_sc_hd__nand2_1 U29271 ( .A(n24577), .B(n25731), .Y(n24681) );
  sky130_fd_sc_hd__nand2_1 U29272 ( .A(n24576), .B(n25731), .Y(n24746) );
  sky130_fd_sc_hd__o22ai_1 U29273 ( .A1(n24501), .A2(n24681), .B1(n24500), 
        .B2(n24746), .Y(n24502) );
  sky130_fd_sc_hd__a21oi_1 U29274 ( .A1(j202_soc_core_intc_core_00_rg_itgt[16]), .A2(n24772), .B1(n24502), .Y(n24503) );
  sky130_fd_sc_hd__nand2_1 U29275 ( .A(n24504), .B(n24503), .Y(n24505) );
  sky130_fd_sc_hd__a21oi_1 U29276 ( .A1(n24765), .A2(
        j202_soc_core_intc_core_00_rg_itgt[0]), .B1(n24505), .Y(n24506) );
  sky130_fd_sc_hd__nand4_1 U29277 ( .A(n24509), .B(n24508), .C(n24507), .D(
        n24506), .Y(j202_soc_core_ahb2apb_01_N128) );
  sky130_fd_sc_hd__a22oi_1 U29278 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[56]), .B1(n24776), .B2(
        j202_soc_core_intc_core_00_rg_ipr[97]), .Y(n24519) );
  sky130_fd_sc_hd__a22oi_1 U29279 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[1]), .B1(n24560), .B2(
        j202_soc_core_intc_core_00_rg_eimk[1]), .Y(n24518) );
  sky130_fd_sc_hd__o21ai_1 U29280 ( .A1(j202_soc_core_intc_core_00_bs_addr[7]), 
        .A2(j202_soc_core_intc_core_00_in_intreq[1]), .B1(n24689), .Y(n24517)
         );
  sky130_fd_sc_hd__a22oi_1 U29281 ( .A1(j202_soc_core_intc_core_00_rg_ipr[33]), 
        .A2(n24770), .B1(n24768), .B2(j202_soc_core_intc_core_00_rg_itgt[40]), 
        .Y(n24514) );
  sky130_fd_sc_hd__o22ai_1 U29282 ( .A1(n24511), .A2(n24681), .B1(n24510), 
        .B2(n24746), .Y(n24512) );
  sky130_fd_sc_hd__a21oi_1 U29283 ( .A1(n24765), .A2(
        j202_soc_core_intc_core_00_rg_itgt[32]), .B1(n24512), .Y(n24513) );
  sky130_fd_sc_hd__nand2_1 U29284 ( .A(n24514), .B(n24513), .Y(n24515) );
  sky130_fd_sc_hd__a21oi_1 U29285 ( .A1(j202_soc_core_intc_core_00_rg_itgt[48]), .A2(n24772), .B1(n24515), .Y(n24516) );
  sky130_fd_sc_hd__nand4_1 U29286 ( .A(n24519), .B(n24518), .C(n24517), .D(
        n24516), .Y(j202_soc_core_ahb2apb_01_N129) );
  sky130_fd_sc_hd__a22oi_1 U29287 ( .A1(j202_soc_core_intc_core_00_rg_ipr[34]), 
        .A2(n24770), .B1(n24769), .B2(j202_soc_core_intc_core_00_rg_itgt[88]), 
        .Y(n24529) );
  sky130_fd_sc_hd__a22oi_1 U29288 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[2]), .B1(n24560), .B2(
        j202_soc_core_intc_core_00_rg_eimk[2]), .Y(n24528) );
  sky130_fd_sc_hd__o21ai_1 U29289 ( .A1(j202_soc_core_intc_core_00_bs_addr[7]), 
        .A2(j202_soc_core_intc_core_00_in_intreq[2]), .B1(n24689), .Y(n24527)
         );
  sky130_fd_sc_hd__a22oi_1 U29290 ( .A1(n24776), .A2(
        j202_soc_core_intc_core_00_rg_ipr[98]), .B1(n24768), .B2(
        j202_soc_core_intc_core_00_rg_itgt[72]), .Y(n24524) );
  sky130_fd_sc_hd__o22ai_1 U29291 ( .A1(n24521), .A2(n24681), .B1(n24520), 
        .B2(n24746), .Y(n24522) );
  sky130_fd_sc_hd__a21oi_1 U29292 ( .A1(n24765), .A2(
        j202_soc_core_intc_core_00_rg_itgt[64]), .B1(n24522), .Y(n24523) );
  sky130_fd_sc_hd__nand2_1 U29293 ( .A(n24524), .B(n24523), .Y(n24525) );
  sky130_fd_sc_hd__a21oi_1 U29294 ( .A1(j202_soc_core_intc_core_00_rg_itgt[80]), .A2(n24772), .B1(n24525), .Y(n24526) );
  sky130_fd_sc_hd__nand4_1 U29295 ( .A(n24529), .B(n24528), .C(n24527), .D(
        n24526), .Y(j202_soc_core_ahb2apb_01_N130) );
  sky130_fd_sc_hd__a22oi_1 U29296 ( .A1(j202_soc_core_intc_core_00_rg_ipr[35]), 
        .A2(n24770), .B1(n24776), .B2(j202_soc_core_intc_core_00_rg_ipr[99]), 
        .Y(n24539) );
  sky130_fd_sc_hd__a22oi_1 U29297 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[3]), .B1(n24560), .B2(
        j202_soc_core_intc_core_00_rg_eimk[3]), .Y(n24538) );
  sky130_fd_sc_hd__o21ai_1 U29298 ( .A1(j202_soc_core_intc_core_00_bs_addr[7]), 
        .A2(j202_soc_core_intc_core_00_in_intreq[3]), .B1(n24689), .Y(n24537)
         );
  sky130_fd_sc_hd__a22oi_1 U29299 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[120]), .B1(n24768), .B2(
        j202_soc_core_intc_core_00_rg_itgt[104]), .Y(n24534) );
  sky130_fd_sc_hd__o22ai_1 U29300 ( .A1(n24531), .A2(n24681), .B1(n24530), 
        .B2(n24746), .Y(n24532) );
  sky130_fd_sc_hd__a21oi_1 U29301 ( .A1(n24765), .A2(
        j202_soc_core_intc_core_00_rg_itgt[96]), .B1(n24532), .Y(n24533) );
  sky130_fd_sc_hd__nand2_1 U29302 ( .A(n24534), .B(n24533), .Y(n24535) );
  sky130_fd_sc_hd__a21oi_1 U29303 ( .A1(
        j202_soc_core_intc_core_00_rg_itgt[112]), .A2(n24772), .B1(n24535), 
        .Y(n24536) );
  sky130_fd_sc_hd__nand4_1 U29304 ( .A(n24539), .B(n24538), .C(n24537), .D(
        n24536), .Y(j202_soc_core_ahb2apb_01_N131) );
  sky130_fd_sc_hd__a22oi_1 U29305 ( .A1(j202_soc_core_intc_core_00_rg_itgt[9]), 
        .A2(n24768), .B1(n24769), .B2(j202_soc_core_intc_core_00_rg_itgt[25]), 
        .Y(n24546) );
  sky130_fd_sc_hd__a22oi_1 U29306 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[4]), .B1(n24560), .B2(
        j202_soc_core_intc_core_00_rg_eimk[4]), .Y(n24545) );
  sky130_fd_sc_hd__a22oi_1 U29308 ( .A1(j202_soc_core_intc_core_00_rg_ipr[36]), 
        .A2(n24770), .B1(n24776), .B2(j202_soc_core_intc_core_00_rg_ipr[100]), 
        .Y(n24542) );
  sky130_fd_sc_hd__a22oi_1 U29309 ( .A1(j202_soc_core_intc_core_00_rg_ipr[68]), 
        .A2(n24771), .B1(j202_soc_core_intc_core_00_rg_ipr[4]), .B2(n24766), 
        .Y(n24541) );
  sky130_fd_sc_hd__a22oi_1 U29310 ( .A1(j202_soc_core_intc_core_00_rg_itgt[1]), 
        .A2(n24765), .B1(j202_soc_core_intc_core_00_rg_itgt[17]), .B2(n24772), 
        .Y(n24540) );
  sky130_fd_sc_hd__and3_1 U29311 ( .A(n24542), .B(n24541), .C(n24540), .X(
        n24543) );
  sky130_fd_sc_hd__nand4_1 U29312 ( .A(n24546), .B(n24545), .C(n24544), .D(
        n24543), .Y(j202_soc_core_ahb2apb_01_N132) );
  sky130_fd_sc_hd__a22oi_1 U29313 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[5]), .B1(n24772), .B2(
        j202_soc_core_intc_core_00_rg_itgt[49]), .Y(n24558) );
  sky130_fd_sc_hd__a22oi_1 U29314 ( .A1(j202_soc_core_intc_core_00_rg_ipr[69]), 
        .A2(n24577), .B1(j202_soc_core_intc_core_00_rg_ipr[5]), .B2(n24576), 
        .Y(n24555) );
  sky130_fd_sc_hd__nor2_1 U29315 ( .A(j202_soc_core_intc_core_00_bs_addr[7]), 
        .B(j202_soc_core_intc_core_00_in_intreq[5]), .Y(n24549) );
  sky130_fd_sc_hd__o22ai_1 U29316 ( .A1(n24549), .A2(n24571), .B1(n24548), 
        .B2(n24547), .Y(n24550) );
  sky130_fd_sc_hd__a21oi_1 U29317 ( .A1(n24575), .A2(
        j202_soc_core_intc_core_00_rg_eimk[5]), .B1(n24550), .Y(n24554) );
  sky130_fd_sc_hd__clkinv_1 U29318 ( .A(j202_soc_core_intc_core_00_rg_itgt[57]), .Y(n24551) );
  sky130_fd_sc_hd__nand2_1 U29319 ( .A(n24551), .B(
        j202_soc_core_intc_core_00_bs_addr[3]), .Y(n24552) );
  sky130_fd_sc_hd__o211ai_1 U29320 ( .A1(j202_soc_core_intc_core_00_bs_addr[3]), .A2(j202_soc_core_intc_core_00_rg_itgt[41]), .B1(n24552), .C1(n24579), .Y(
        n24553) );
  sky130_fd_sc_hd__a31oi_1 U29321 ( .A1(n24555), .A2(n24554), .A3(n24553), 
        .B1(j202_soc_core_rst), .Y(n24556) );
  sky130_fd_sc_hd__a21oi_1 U29322 ( .A1(j202_soc_core_intc_core_00_rg_ipr[101]), .A2(n24776), .B1(n24556), .Y(n24557) );
  sky130_fd_sc_hd__o211ai_1 U29323 ( .A1(n24559), .A2(n24744), .B1(n24558), 
        .C1(n24557), .Y(j202_soc_core_ahb2apb_01_N133) );
  sky130_fd_sc_hd__a22oi_1 U29324 ( .A1(j202_soc_core_intc_core_00_rg_ipr[38]), 
        .A2(n24770), .B1(n24776), .B2(j202_soc_core_intc_core_00_rg_ipr[102]), 
        .Y(n24570) );
  sky130_fd_sc_hd__a22oi_1 U29325 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[6]), .B1(n24560), .B2(
        j202_soc_core_intc_core_00_rg_eimk[6]), .Y(n24569) );
  sky130_fd_sc_hd__a22oi_1 U29327 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[89]), .B1(n24768), .B2(
        j202_soc_core_intc_core_00_rg_itgt[73]), .Y(n24565) );
  sky130_fd_sc_hd__o22ai_1 U29328 ( .A1(n24562), .A2(n24681), .B1(n24561), 
        .B2(n24746), .Y(n24563) );
  sky130_fd_sc_hd__a21oi_1 U29329 ( .A1(n24765), .A2(
        j202_soc_core_intc_core_00_rg_itgt[65]), .B1(n24563), .Y(n24564) );
  sky130_fd_sc_hd__nand2_1 U29330 ( .A(n24565), .B(n24564), .Y(n24566) );
  sky130_fd_sc_hd__a21oi_1 U29331 ( .A1(j202_soc_core_intc_core_00_rg_itgt[81]), .A2(n24772), .B1(n24566), .Y(n24567) );
  sky130_fd_sc_hd__nand4_1 U29332 ( .A(n24570), .B(n24569), .C(n24568), .D(
        n24567), .Y(j202_soc_core_ahb2apb_01_N134) );
  sky130_fd_sc_hd__a22oi_1 U29333 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[7]), .B1(n24765), .B2(
        j202_soc_core_intc_core_00_rg_itgt[97]), .Y(n24587) );
  sky130_fd_sc_hd__a22oi_1 U29334 ( .A1(j202_soc_core_intc_core_00_rg_ipr[39]), 
        .A2(n24770), .B1(n24772), .B2(j202_soc_core_intc_core_00_rg_itgt[113]), 
        .Y(n24586) );
  sky130_fd_sc_hd__a21oi_1 U29335 ( .A1(n24573), .A2(n24572), .B1(n24571), .Y(
        n24574) );
  sky130_fd_sc_hd__a21oi_1 U29336 ( .A1(j202_soc_core_intc_core_00_rg_eimk[7]), 
        .A2(n24575), .B1(n24574), .Y(n24583) );
  sky130_fd_sc_hd__a22oi_1 U29337 ( .A1(j202_soc_core_intc_core_00_rg_ipr[71]), 
        .A2(n24577), .B1(j202_soc_core_intc_core_00_rg_ipr[7]), .B2(n24576), 
        .Y(n24582) );
  sky130_fd_sc_hd__clkinv_1 U29338 ( .A(
        j202_soc_core_intc_core_00_rg_itgt[121]), .Y(n24578) );
  sky130_fd_sc_hd__nand2_1 U29339 ( .A(n24578), .B(
        j202_soc_core_intc_core_00_bs_addr[3]), .Y(n24580) );
  sky130_fd_sc_hd__o211ai_1 U29340 ( .A1(j202_soc_core_intc_core_00_bs_addr[3]), .A2(j202_soc_core_intc_core_00_rg_itgt[105]), .B1(n24580), .C1(n24579), .Y(
        n24581) );
  sky130_fd_sc_hd__a31oi_1 U29341 ( .A1(n24583), .A2(n24582), .A3(n24581), 
        .B1(j202_soc_core_rst), .Y(n24584) );
  sky130_fd_sc_hd__a21oi_1 U29342 ( .A1(n24776), .A2(
        j202_soc_core_intc_core_00_rg_ipr[103]), .B1(n24584), .Y(n24585) );
  sky130_fd_sc_hd__nand3_1 U29343 ( .A(n24587), .B(n24586), .C(n24585), .Y(
        j202_soc_core_ahb2apb_01_N135) );
  sky130_fd_sc_hd__a22oi_1 U29344 ( .A1(j202_soc_core_intc_core_00_rg_ipr[40]), 
        .A2(n24770), .B1(n24776), .B2(j202_soc_core_intc_core_00_rg_ipr[104]), 
        .Y(n24596) );
  sky130_fd_sc_hd__a22oi_1 U29345 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[8]), .A2(n24689), .B1(
        j202_soc_core_intc_core_00_rg_itgt[2]), .B2(n24765), .Y(n24595) );
  sky130_fd_sc_hd__a22oi_1 U29346 ( .A1(j202_soc_core_intc_core_00_rg_itgt[10]), .A2(n24768), .B1(n24769), .B2(j202_soc_core_intc_core_00_rg_itgt[26]), .Y(
        n24592) );
  sky130_fd_sc_hd__o22ai_1 U29347 ( .A1(n24589), .A2(n24681), .B1(n24588), 
        .B2(n24746), .Y(n24590) );
  sky130_fd_sc_hd__a21oi_1 U29348 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[8]), .B1(n24590), .Y(n24591) );
  sky130_fd_sc_hd__nand2_1 U29349 ( .A(n24592), .B(n24591), .Y(n24593) );
  sky130_fd_sc_hd__a21oi_1 U29350 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[18]), .B1(n24593), .Y(n24594) );
  sky130_fd_sc_hd__nand4_1 U29351 ( .A(n24596), .B(n24595), .C(n24594), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N136) );
  sky130_fd_sc_hd__a22oi_1 U29352 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[58]), .B1(n24768), .B2(
        j202_soc_core_intc_core_00_rg_itgt[42]), .Y(n24605) );
  sky130_fd_sc_hd__a22oi_1 U29353 ( .A1(j202_soc_core_intc_core_00_rg_ipr[41]), 
        .A2(n24770), .B1(n24776), .B2(j202_soc_core_intc_core_00_rg_ipr[105]), 
        .Y(n24604) );
  sky130_fd_sc_hd__o21ai_1 U29354 ( .A1(n24597), .A2(n24681), .B1(n24777), .Y(
        n24598) );
  sky130_fd_sc_hd__a21oi_1 U29355 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[9]), .B1(n24598), .Y(n24603) );
  sky130_fd_sc_hd__a22oi_1 U29356 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[9]), .A2(n24689), .B1(n24772), 
        .B2(j202_soc_core_intc_core_00_rg_itgt[50]), .Y(n24599) );
  sky130_fd_sc_hd__a21oi_1 U29358 ( .A1(n24765), .A2(
        j202_soc_core_intc_core_00_rg_itgt[34]), .B1(n24601), .Y(n24602) );
  sky130_fd_sc_hd__nand4_1 U29359 ( .A(n24605), .B(n24604), .C(n24603), .D(
        n24602), .Y(j202_soc_core_ahb2apb_01_N137) );
  sky130_fd_sc_hd__a22oi_1 U29360 ( .A1(j202_soc_core_intc_core_00_rg_ipr[42]), 
        .A2(n24770), .B1(n24768), .B2(j202_soc_core_intc_core_00_rg_itgt[74]), 
        .Y(n24614) );
  sky130_fd_sc_hd__a22oi_1 U29361 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[90]), .B1(n24776), .B2(
        j202_soc_core_intc_core_00_rg_ipr[106]), .Y(n24613) );
  sky130_fd_sc_hd__o21ai_1 U29362 ( .A1(n24606), .A2(n24681), .B1(n24777), .Y(
        n24607) );
  sky130_fd_sc_hd__a21oi_1 U29363 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[10]), .A2(n24689), .B1(n24607), 
        .Y(n24612) );
  sky130_fd_sc_hd__a22oi_1 U29364 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[10]), .B1(n24772), .B2(
        j202_soc_core_intc_core_00_rg_itgt[82]), .Y(n24608) );
  sky130_fd_sc_hd__a21oi_1 U29366 ( .A1(n24765), .A2(
        j202_soc_core_intc_core_00_rg_itgt[66]), .B1(n24610), .Y(n24611) );
  sky130_fd_sc_hd__nand4_1 U29367 ( .A(n24614), .B(n24613), .C(n24612), .D(
        n24611), .Y(j202_soc_core_ahb2apb_01_N138) );
  sky130_fd_sc_hd__a22oi_1 U29368 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[122]), .B1(n24776), .B2(
        j202_soc_core_intc_core_00_rg_ipr[107]), .Y(n24622) );
  sky130_fd_sc_hd__a22oi_1 U29369 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[11]), .A2(n24689), .B1(
        j202_soc_core_intc_core_00_rg_ipr[11]), .B2(n24766), .Y(n24621) );
  sky130_fd_sc_hd__a22oi_1 U29370 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[114]), .B1(n24765), .B2(
        j202_soc_core_intc_core_00_rg_itgt[98]), .Y(n24620) );
  sky130_fd_sc_hd__o2bb2ai_1 U29371 ( .B1(n24615), .B2(n24744), .A1_N(n24768), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[106]), .Y(n24618) );
  sky130_fd_sc_hd__a211oi_1 U29373 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[11]), .B1(n24618), .C1(n24617), .Y(
        n24619) );
  sky130_fd_sc_hd__nand4_1 U29374 ( .A(n24622), .B(n24621), .C(n24620), .D(
        n24619), .Y(j202_soc_core_ahb2apb_01_N139) );
  sky130_fd_sc_hd__a22oi_1 U29375 ( .A1(j202_soc_core_intc_core_00_rg_ipr[44]), 
        .A2(n24770), .B1(n24769), .B2(j202_soc_core_intc_core_00_rg_itgt[27]), 
        .Y(n24631) );
  sky130_fd_sc_hd__a22oi_1 U29376 ( .A1(j202_soc_core_intc_core_00_rg_itgt[11]), .A2(n24768), .B1(n24776), .B2(j202_soc_core_intc_core_00_rg_ipr[108]), .Y(
        n24630) );
  sky130_fd_sc_hd__o21ai_1 U29377 ( .A1(n24623), .A2(n24746), .B1(n24777), .Y(
        n24624) );
  sky130_fd_sc_hd__a21oi_1 U29378 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[12]), .A2(n24689), .B1(n24624), 
        .Y(n24629) );
  sky130_fd_sc_hd__a22oi_1 U29379 ( .A1(j202_soc_core_intc_core_00_rg_itgt[19]), .A2(n24772), .B1(n24767), .B2(j202_soc_core_intc_core_00_rg_ie[12]), .Y(
        n24625) );
  sky130_fd_sc_hd__a21oi_1 U29381 ( .A1(j202_soc_core_intc_core_00_rg_itgt[3]), 
        .A2(n24765), .B1(n24627), .Y(n24628) );
  sky130_fd_sc_hd__nand4_1 U29382 ( .A(n24631), .B(n24630), .C(n24629), .D(
        n24628), .Y(j202_soc_core_ahb2apb_01_N140) );
  sky130_fd_sc_hd__a22oi_1 U29383 ( .A1(j202_soc_core_intc_core_00_rg_ipr[45]), 
        .A2(n24770), .B1(n24768), .B2(j202_soc_core_intc_core_00_rg_itgt[43]), 
        .Y(n24640) );
  sky130_fd_sc_hd__a22oi_1 U29384 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[13]), .B1(n24765), .B2(
        j202_soc_core_intc_core_00_rg_itgt[35]), .Y(n24639) );
  sky130_fd_sc_hd__a22oi_1 U29385 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[59]), .B1(n24776), .B2(
        j202_soc_core_intc_core_00_rg_ipr[109]), .Y(n24636) );
  sky130_fd_sc_hd__o22ai_1 U29386 ( .A1(n24633), .A2(n24681), .B1(n24632), 
        .B2(n24746), .Y(n24634) );
  sky130_fd_sc_hd__a21oi_1 U29387 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[51]), .B1(n24634), .Y(n24635) );
  sky130_fd_sc_hd__nand2_1 U29388 ( .A(n24636), .B(n24635), .Y(n24637) );
  sky130_fd_sc_hd__a21oi_1 U29389 ( .A1(n24689), .A2(
        j202_soc_core_intc_core_00_in_intreq[13]), .B1(n24637), .Y(n24638) );
  sky130_fd_sc_hd__nand4_1 U29390 ( .A(n24640), .B(n24639), .C(n24638), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N141) );
  sky130_fd_sc_hd__a22oi_1 U29391 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[91]), .B1(n24768), .B2(
        j202_soc_core_intc_core_00_rg_itgt[75]), .Y(n24649) );
  sky130_fd_sc_hd__a22oi_1 U29392 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[14]), .A2(n24689), .B1(n24772), 
        .B2(j202_soc_core_intc_core_00_rg_itgt[83]), .Y(n24648) );
  sky130_fd_sc_hd__a22oi_1 U29393 ( .A1(j202_soc_core_intc_core_00_rg_ipr[46]), 
        .A2(n24770), .B1(n24776), .B2(j202_soc_core_intc_core_00_rg_ipr[110]), 
        .Y(n24645) );
  sky130_fd_sc_hd__o22ai_1 U29394 ( .A1(n24642), .A2(n24681), .B1(n24641), 
        .B2(n24746), .Y(n24643) );
  sky130_fd_sc_hd__a21oi_1 U29395 ( .A1(n24765), .A2(
        j202_soc_core_intc_core_00_rg_itgt[67]), .B1(n24643), .Y(n24644) );
  sky130_fd_sc_hd__nand2_1 U29396 ( .A(n24645), .B(n24644), .Y(n24646) );
  sky130_fd_sc_hd__a21oi_1 U29397 ( .A1(j202_soc_core_intc_core_00_rg_ie[14]), 
        .A2(n24767), .B1(n24646), .Y(n24647) );
  sky130_fd_sc_hd__nand4_1 U29398 ( .A(n24649), .B(n24648), .C(n24647), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N142) );
  sky130_fd_sc_hd__a22oi_1 U29399 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[123]), .B1(n24768), .B2(
        j202_soc_core_intc_core_00_rg_itgt[107]), .Y(n24658) );
  sky130_fd_sc_hd__a22oi_1 U29400 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[15]), .A2(n24689), .B1(
        j202_soc_core_intc_core_00_rg_ipr[79]), .B2(n24771), .Y(n24657) );
  sky130_fd_sc_hd__o22ai_1 U29401 ( .A1(n24651), .A2(n24744), .B1(n24705), 
        .B2(n24650), .Y(n24655) );
  sky130_fd_sc_hd__a22oi_1 U29402 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[115]), .B1(n24765), .B2(
        j202_soc_core_intc_core_00_rg_itgt[99]), .Y(n24652) );
  sky130_fd_sc_hd__o21ai_1 U29403 ( .A1(n24653), .A2(n24746), .B1(n24652), .Y(
        n24654) );
  sky130_fd_sc_hd__a211oi_1 U29404 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[15]), .B1(n24655), .C1(n24654), .Y(
        n24656) );
  sky130_fd_sc_hd__nand4_1 U29405 ( .A(n24658), .B(n24657), .C(n24656), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N143) );
  sky130_fd_sc_hd__a22oi_1 U29406 ( .A1(j202_soc_core_intc_core_00_rg_itgt[12]), .A2(n24768), .B1(n24769), .B2(j202_soc_core_intc_core_00_rg_itgt[28]), .Y(
        n24664) );
  sky130_fd_sc_hd__a22oi_1 U29407 ( .A1(j202_soc_core_intc_core_00_rg_itgt[20]), .A2(n24772), .B1(j202_soc_core_intc_core_00_in_intreq[16]), .B2(n24689), .Y(
        n24663) );
  sky130_fd_sc_hd__a22oi_1 U29408 ( .A1(j202_soc_core_intc_core_00_rg_ipr[48]), 
        .A2(n24770), .B1(n24776), .B2(j202_soc_core_intc_core_00_rg_ipr[112]), 
        .Y(n24661) );
  sky130_fd_sc_hd__a22oi_1 U29409 ( .A1(j202_soc_core_intc_core_00_rg_itgt[4]), 
        .A2(n24765), .B1(j202_soc_core_intc_core_00_rg_ipr[16]), .B2(n24766), 
        .Y(n24660) );
  sky130_fd_sc_hd__a22oi_1 U29410 ( .A1(j202_soc_core_intc_core_00_rg_ipr[80]), 
        .A2(n24771), .B1(n24767), .B2(j202_soc_core_intc_core_00_rg_ie[16]), 
        .Y(n24659) );
  sky130_fd_sc_hd__and3_1 U29411 ( .A(n24661), .B(n24660), .C(n24659), .X(
        n24662) );
  sky130_fd_sc_hd__nand4_1 U29412 ( .A(n24664), .B(n24663), .C(n24662), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N144) );
  sky130_fd_sc_hd__a22oi_1 U29413 ( .A1(n24776), .A2(
        j202_soc_core_intc_core_00_rg_ipr[113]), .B1(n24768), .B2(
        j202_soc_core_intc_core_00_rg_itgt[44]), .Y(n24672) );
  sky130_fd_sc_hd__a22oi_1 U29414 ( .A1(
        j202_soc_core_intc_core_00_in_intreq[17]), .A2(n24689), .B1(
        j202_soc_core_intc_core_00_rg_ipr[81]), .B2(n24771), .Y(n24671) );
  sky130_fd_sc_hd__a22oi_1 U29415 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[52]), .B1(n24765), .B2(
        j202_soc_core_intc_core_00_rg_itgt[36]), .Y(n24670) );
  sky130_fd_sc_hd__o2bb2ai_1 U29416 ( .B1(n24665), .B2(n24744), .A1_N(n24769), 
        .A2_N(j202_soc_core_intc_core_00_rg_itgt[60]), .Y(n24668) );
  sky130_fd_sc_hd__a211oi_1 U29418 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[17]), .B1(n24668), .C1(n24667), .Y(
        n24669) );
  sky130_fd_sc_hd__nand4_1 U29419 ( .A(n24672), .B(n24671), .C(n24670), .D(
        n24669), .Y(j202_soc_core_ahb2apb_01_N145) );
  sky130_fd_sc_hd__a22oi_1 U29420 ( .A1(j202_soc_core_intc_core_00_rg_ipr[18]), 
        .A2(n24766), .B1(n24765), .B2(j202_soc_core_intc_core_00_rg_itgt[68]), 
        .Y(n24679) );
  sky130_fd_sc_hd__a22oi_1 U29421 ( .A1(n24768), .A2(
        j202_soc_core_intc_core_00_rg_itgt[76]), .B1(n24767), .B2(
        j202_soc_core_intc_core_00_rg_ie[18]), .Y(n24678) );
  sky130_fd_sc_hd__a22oi_1 U29422 ( .A1(j202_soc_core_intc_core_00_rg_ipr[50]), 
        .A2(n24770), .B1(n24769), .B2(j202_soc_core_intc_core_00_rg_itgt[92]), 
        .Y(n24674) );
  sky130_fd_sc_hd__a22oi_1 U29423 ( .A1(n24776), .A2(
        j202_soc_core_intc_core_00_rg_ipr[114]), .B1(n24772), .B2(
        j202_soc_core_intc_core_00_rg_itgt[84]), .Y(n24673) );
  sky130_fd_sc_hd__nand2_1 U29424 ( .A(n24674), .B(n24673), .Y(n24675) );
  sky130_fd_sc_hd__a21oi_1 U29425 ( .A1(n24771), .A2(
        j202_soc_core_intc_core_00_rg_ipr[82]), .B1(n24675), .Y(n24677) );
  sky130_fd_sc_hd__o21ai_1 U29426 ( .A1(j202_soc_core_intc_core_00_bs_addr[7]), 
        .A2(j202_soc_core_intc_core_00_in_intreq[18]), .B1(n24689), .Y(n24676)
         );
  sky130_fd_sc_hd__nand4_1 U29427 ( .A(n24679), .B(n24678), .C(n24677), .D(
        n24676), .Y(j202_soc_core_ahb2apb_01_N146) );
  sky130_fd_sc_hd__a22oi_1 U29428 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[124]), .B1(n24768), .B2(
        j202_soc_core_intc_core_00_rg_itgt[108]), .Y(n24688) );
  sky130_fd_sc_hd__a22oi_1 U29429 ( .A1(j202_soc_core_intc_core_00_rg_ipr[51]), 
        .A2(n24770), .B1(n24767), .B2(j202_soc_core_intc_core_00_rg_ie[19]), 
        .Y(n24687) );
  sky130_fd_sc_hd__o22ai_1 U29430 ( .A1(n24682), .A2(n24681), .B1(n24680), 
        .B2(n24746), .Y(n24684) );
  sky130_fd_sc_hd__a22o_1 U29431 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[116]), .B1(n24765), .B2(
        j202_soc_core_intc_core_00_rg_itgt[100]), .X(n24683) );
  sky130_fd_sc_hd__a211oi_1 U29432 ( .A1(n24776), .A2(
        j202_soc_core_intc_core_00_rg_ipr[115]), .B1(n24684), .C1(n24683), .Y(
        n24686) );
  sky130_fd_sc_hd__o21ai_1 U29433 ( .A1(j202_soc_core_intc_core_00_bs_addr[7]), 
        .A2(j202_soc_core_intc_core_00_in_intreq[19]), .B1(n24689), .Y(n24685)
         );
  sky130_fd_sc_hd__nand4_1 U29434 ( .A(n24688), .B(n24687), .C(n24686), .D(
        n24685), .Y(j202_soc_core_ahb2apb_01_N147) );
  sky130_fd_sc_hd__a22oi_1 U29435 ( .A1(j202_soc_core_intc_core_00_rg_ipr[52]), 
        .A2(n24770), .B1(n24776), .B2(j202_soc_core_intc_core_00_rg_ipr[116]), 
        .Y(n24695) );
  sky130_fd_sc_hd__a22oi_1 U29436 ( .A1(j202_soc_core_intc_core_00_rg_itgt[5]), 
        .A2(n24765), .B1(j202_soc_core_intc_core_00_in_intreq[20]), .B2(n24689), .Y(n24694) );
  sky130_fd_sc_hd__a22oi_1 U29437 ( .A1(j202_soc_core_intc_core_00_rg_itgt[13]), .A2(n24768), .B1(n24769), .B2(j202_soc_core_intc_core_00_rg_itgt[29]), .Y(
        n24692) );
  sky130_fd_sc_hd__a22oi_1 U29438 ( .A1(j202_soc_core_intc_core_00_rg_ipr[20]), 
        .A2(n24766), .B1(n24772), .B2(j202_soc_core_intc_core_00_rg_itgt[21]), 
        .Y(n24691) );
  sky130_fd_sc_hd__a22oi_1 U29439 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[20]), .B1(n24771), .B2(
        j202_soc_core_intc_core_00_rg_ipr[84]), .Y(n24690) );
  sky130_fd_sc_hd__and3_1 U29440 ( .A(n24692), .B(n24691), .C(n24690), .X(
        n24693) );
  sky130_fd_sc_hd__nand4_1 U29441 ( .A(n24695), .B(n24694), .C(n24693), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N148) );
  sky130_fd_sc_hd__a22oi_1 U29442 ( .A1(j202_soc_core_intc_core_00_rg_ipr[21]), 
        .A2(n24766), .B1(n24765), .B2(j202_soc_core_intc_core_00_rg_itgt[37]), 
        .Y(n24701) );
  sky130_fd_sc_hd__a22oi_1 U29443 ( .A1(n24768), .A2(
        j202_soc_core_intc_core_00_rg_itgt[45]), .B1(n24767), .B2(
        j202_soc_core_intc_core_00_rg_ie[21]), .Y(n24700) );
  sky130_fd_sc_hd__a22oi_1 U29444 ( .A1(j202_soc_core_intc_core_00_rg_ipr[53]), 
        .A2(n24770), .B1(n24769), .B2(j202_soc_core_intc_core_00_rg_itgt[61]), 
        .Y(n24697) );
  sky130_fd_sc_hd__a22oi_1 U29445 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[53]), .B1(n24771), .B2(
        j202_soc_core_intc_core_00_rg_ipr[85]), .Y(n24696) );
  sky130_fd_sc_hd__nand2_1 U29446 ( .A(n24697), .B(n24696), .Y(n24698) );
  sky130_fd_sc_hd__a21oi_1 U29447 ( .A1(j202_soc_core_intc_core_00_rg_ipr[117]), .A2(n24776), .B1(n24698), .Y(n24699) );
  sky130_fd_sc_hd__nand4_1 U29448 ( .A(n24701), .B(n24700), .C(n24699), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N149) );
  sky130_fd_sc_hd__a22oi_1 U29449 ( .A1(n24771), .A2(
        j202_soc_core_intc_core_00_rg_ipr[86]), .B1(n24765), .B2(
        j202_soc_core_intc_core_00_rg_itgt[69]), .Y(n24711) );
  sky130_fd_sc_hd__a22oi_1 U29450 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[93]), .B1(n24768), .B2(
        j202_soc_core_intc_core_00_rg_itgt[77]), .Y(n24710) );
  sky130_fd_sc_hd__o21ai_1 U29451 ( .A1(n24744), .A2(n24702), .B1(n24777), .Y(
        n24703) );
  sky130_fd_sc_hd__a21oi_1 U29452 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[22]), .B1(n24703), .Y(n24709) );
  sky130_fd_sc_hd__o22ai_1 U29453 ( .A1(n24706), .A2(n24746), .B1(n24705), 
        .B2(n24704), .Y(n24707) );
  sky130_fd_sc_hd__a21oi_1 U29454 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[85]), .B1(n24707), .Y(n24708) );
  sky130_fd_sc_hd__nand4_1 U29455 ( .A(n24711), .B(n24710), .C(n24709), .D(
        n24708), .Y(j202_soc_core_ahb2apb_01_N150) );
  sky130_fd_sc_hd__a22oi_1 U29456 ( .A1(j202_soc_core_intc_core_00_rg_ipr[23]), 
        .A2(n24766), .B1(n24765), .B2(j202_soc_core_intc_core_00_rg_itgt[101]), 
        .Y(n24717) );
  sky130_fd_sc_hd__a22oi_1 U29457 ( .A1(n24776), .A2(
        j202_soc_core_intc_core_00_rg_ipr[119]), .B1(n24767), .B2(
        j202_soc_core_intc_core_00_rg_ie[23]), .Y(n24716) );
  sky130_fd_sc_hd__a22oi_1 U29458 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[125]), .B1(n24768), .B2(
        j202_soc_core_intc_core_00_rg_itgt[109]), .Y(n24713) );
  sky130_fd_sc_hd__a22oi_1 U29459 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[117]), .B1(n24771), .B2(
        j202_soc_core_intc_core_00_rg_ipr[87]), .Y(n24712) );
  sky130_fd_sc_hd__nand2_1 U29460 ( .A(n24713), .B(n24712), .Y(n24714) );
  sky130_fd_sc_hd__a21oi_1 U29461 ( .A1(n24770), .A2(
        j202_soc_core_intc_core_00_rg_ipr[55]), .B1(n24714), .Y(n24715) );
  sky130_fd_sc_hd__nand4_1 U29462 ( .A(n24717), .B(n24716), .C(n24715), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N151) );
  sky130_fd_sc_hd__a22oi_1 U29463 ( .A1(j202_soc_core_intc_core_00_rg_itgt[6]), 
        .A2(n24765), .B1(n24772), .B2(j202_soc_core_intc_core_00_rg_itgt[22]), 
        .Y(n24724) );
  sky130_fd_sc_hd__a22oi_1 U29464 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[30]), .B1(n24767), .B2(
        j202_soc_core_intc_core_00_rg_ie[24]), .Y(n24723) );
  sky130_fd_sc_hd__a22o_1 U29465 ( .A1(n24776), .A2(
        j202_soc_core_intc_core_00_rg_ipr[120]), .B1(
        j202_soc_core_intc_core_00_rg_itgt[14]), .B2(n24768), .X(n24721) );
  sky130_fd_sc_hd__o22ai_1 U29466 ( .A1(n24719), .A2(n24744), .B1(n24718), 
        .B2(n24746), .Y(n24720) );
  sky130_fd_sc_hd__a211oi_1 U29467 ( .A1(n24771), .A2(
        j202_soc_core_intc_core_00_rg_ipr[88]), .B1(n24721), .C1(n24720), .Y(
        n24722) );
  sky130_fd_sc_hd__nand4_1 U29468 ( .A(n24724), .B(n24723), .C(n24722), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N152) );
  sky130_fd_sc_hd__a22oi_1 U29469 ( .A1(j202_soc_core_intc_core_00_rg_ipr[25]), 
        .A2(n24766), .B1(n24772), .B2(j202_soc_core_intc_core_00_rg_itgt[54]), 
        .Y(n24730) );
  sky130_fd_sc_hd__a22oi_1 U29470 ( .A1(n24768), .A2(
        j202_soc_core_intc_core_00_rg_itgt[46]), .B1(n24767), .B2(
        j202_soc_core_intc_core_00_rg_ie[25]), .Y(n24729) );
  sky130_fd_sc_hd__a22oi_1 U29471 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[62]), .B1(n24776), .B2(
        j202_soc_core_intc_core_00_rg_ipr[121]), .Y(n24726) );
  sky130_fd_sc_hd__a22oi_1 U29472 ( .A1(n24771), .A2(
        j202_soc_core_intc_core_00_rg_ipr[89]), .B1(n24765), .B2(
        j202_soc_core_intc_core_00_rg_itgt[38]), .Y(n24725) );
  sky130_fd_sc_hd__nand2_1 U29473 ( .A(n24726), .B(n24725), .Y(n24727) );
  sky130_fd_sc_hd__a21oi_1 U29474 ( .A1(n24770), .A2(
        j202_soc_core_intc_core_00_rg_ipr[57]), .B1(n24727), .Y(n24728) );
  sky130_fd_sc_hd__nand4_1 U29475 ( .A(n24730), .B(n24729), .C(n24728), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N153) );
  sky130_fd_sc_hd__a22oi_1 U29476 ( .A1(j202_soc_core_intc_core_00_rg_ipr[26]), 
        .A2(n24766), .B1(n24771), .B2(j202_soc_core_intc_core_00_rg_ipr[90]), 
        .Y(n24736) );
  sky130_fd_sc_hd__a22oi_1 U29477 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[94]), .B1(n24767), .B2(
        j202_soc_core_intc_core_00_rg_ie[26]), .Y(n24735) );
  sky130_fd_sc_hd__a22oi_1 U29478 ( .A1(n24776), .A2(
        j202_soc_core_intc_core_00_rg_ipr[122]), .B1(n24768), .B2(
        j202_soc_core_intc_core_00_rg_itgt[78]), .Y(n24732) );
  sky130_fd_sc_hd__a22oi_1 U29479 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[86]), .B1(n24765), .B2(
        j202_soc_core_intc_core_00_rg_itgt[70]), .Y(n24731) );
  sky130_fd_sc_hd__nand2_1 U29480 ( .A(n24732), .B(n24731), .Y(n24733) );
  sky130_fd_sc_hd__a21oi_1 U29481 ( .A1(n24770), .A2(
        j202_soc_core_intc_core_00_rg_ipr[58]), .B1(n24733), .Y(n24734) );
  sky130_fd_sc_hd__nand4_1 U29482 ( .A(n24736), .B(n24735), .C(n24734), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N154) );
  sky130_fd_sc_hd__a22oi_1 U29483 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[118]), .B1(n24771), .B2(
        j202_soc_core_intc_core_00_rg_ipr[91]), .Y(n24742) );
  sky130_fd_sc_hd__a22oi_1 U29484 ( .A1(n24776), .A2(
        j202_soc_core_intc_core_00_rg_ipr[123]), .B1(n24767), .B2(
        j202_soc_core_intc_core_00_rg_ie[27]), .Y(n24741) );
  sky130_fd_sc_hd__a22oi_1 U29485 ( .A1(j202_soc_core_intc_core_00_rg_ipr[59]), 
        .A2(n24770), .B1(n24769), .B2(j202_soc_core_intc_core_00_rg_itgt[126]), 
        .Y(n24738) );
  sky130_fd_sc_hd__a22oi_1 U29486 ( .A1(n24768), .A2(
        j202_soc_core_intc_core_00_rg_itgt[110]), .B1(n24765), .B2(
        j202_soc_core_intc_core_00_rg_itgt[102]), .Y(n24737) );
  sky130_fd_sc_hd__nand2_1 U29487 ( .A(n24738), .B(n24737), .Y(n24739) );
  sky130_fd_sc_hd__a21oi_1 U29488 ( .A1(n24766), .A2(
        j202_soc_core_intc_core_00_rg_ipr[27]), .B1(n24739), .Y(n24740) );
  sky130_fd_sc_hd__nand4_1 U29489 ( .A(n24742), .B(n24741), .C(n24740), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N155) );
  sky130_fd_sc_hd__a22oi_1 U29490 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[23]), .B1(n24771), .B2(
        j202_soc_core_intc_core_00_rg_ipr[92]), .Y(n24752) );
  sky130_fd_sc_hd__a22oi_1 U29491 ( .A1(j202_soc_core_intc_core_00_rg_itgt[15]), .A2(n24768), .B1(n24769), .B2(j202_soc_core_intc_core_00_rg_itgt[31]), .Y(
        n24751) );
  sky130_fd_sc_hd__a21oi_1 U29493 ( .A1(n24767), .A2(
        j202_soc_core_intc_core_00_rg_ie[28]), .B1(n24745), .Y(n24750) );
  sky130_fd_sc_hd__o2bb2ai_1 U29494 ( .B1(n24747), .B2(n24746), .A1_N(
        j202_soc_core_intc_core_00_rg_itgt[7]), .A2_N(n24765), .Y(n24748) );
  sky130_fd_sc_hd__a21oi_1 U29495 ( .A1(n24776), .A2(
        j202_soc_core_intc_core_00_rg_ipr[124]), .B1(n24748), .Y(n24749) );
  sky130_fd_sc_hd__nand4_1 U29496 ( .A(n24752), .B(n24751), .C(n24750), .D(
        n24749), .Y(j202_soc_core_ahb2apb_01_N156) );
  sky130_fd_sc_hd__a22oi_1 U29497 ( .A1(j202_soc_core_intc_core_00_rg_ipr[29]), 
        .A2(n24766), .B1(n24765), .B2(j202_soc_core_intc_core_00_rg_itgt[39]), 
        .Y(n24758) );
  sky130_fd_sc_hd__a22oi_1 U29498 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[63]), .B1(n24767), .B2(
        j202_soc_core_intc_core_00_rg_ie[29]), .Y(n24757) );
  sky130_fd_sc_hd__a22oi_1 U29499 ( .A1(n24776), .A2(
        j202_soc_core_intc_core_00_rg_ipr[125]), .B1(n24768), .B2(
        j202_soc_core_intc_core_00_rg_itgt[47]), .Y(n24754) );
  sky130_fd_sc_hd__a22oi_1 U29500 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[55]), .B1(n24771), .B2(
        j202_soc_core_intc_core_00_rg_ipr[93]), .Y(n24753) );
  sky130_fd_sc_hd__nand2_1 U29501 ( .A(n24754), .B(n24753), .Y(n24755) );
  sky130_fd_sc_hd__a21oi_1 U29502 ( .A1(n24770), .A2(
        j202_soc_core_intc_core_00_rg_ipr[61]), .B1(n24755), .Y(n24756) );
  sky130_fd_sc_hd__nand4_1 U29503 ( .A(n24758), .B(n24757), .C(n24756), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N157) );
  sky130_fd_sc_hd__a22oi_1 U29504 ( .A1(j202_soc_core_intc_core_00_rg_ipr[30]), 
        .A2(n24766), .B1(n24771), .B2(j202_soc_core_intc_core_00_rg_ipr[94]), 
        .Y(n24764) );
  sky130_fd_sc_hd__a22oi_1 U29505 ( .A1(n24776), .A2(
        j202_soc_core_intc_core_00_rg_ipr[126]), .B1(n24767), .B2(
        j202_soc_core_intc_core_00_rg_ie[30]), .Y(n24763) );
  sky130_fd_sc_hd__a22oi_1 U29506 ( .A1(n24769), .A2(
        j202_soc_core_intc_core_00_rg_itgt[95]), .B1(n24768), .B2(
        j202_soc_core_intc_core_00_rg_itgt[79]), .Y(n24760) );
  sky130_fd_sc_hd__a22oi_1 U29507 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[87]), .B1(n24765), .B2(
        j202_soc_core_intc_core_00_rg_itgt[71]), .Y(n24759) );
  sky130_fd_sc_hd__nand2_1 U29508 ( .A(n24760), .B(n24759), .Y(n24761) );
  sky130_fd_sc_hd__a21oi_1 U29509 ( .A1(n24770), .A2(
        j202_soc_core_intc_core_00_rg_ipr[62]), .B1(n24761), .Y(n24762) );
  sky130_fd_sc_hd__nand4_1 U29510 ( .A(n24764), .B(n24763), .C(n24762), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N158) );
  sky130_fd_sc_hd__a22oi_1 U29511 ( .A1(j202_soc_core_intc_core_00_rg_ipr[31]), 
        .A2(n24766), .B1(n24765), .B2(j202_soc_core_intc_core_00_rg_itgt[103]), 
        .Y(n24780) );
  sky130_fd_sc_hd__a22oi_1 U29512 ( .A1(n24768), .A2(
        j202_soc_core_intc_core_00_rg_itgt[111]), .B1(n24767), .B2(
        j202_soc_core_intc_core_00_rg_ie[31]), .Y(n24779) );
  sky130_fd_sc_hd__a22oi_1 U29513 ( .A1(j202_soc_core_intc_core_00_rg_ipr[63]), 
        .A2(n24770), .B1(n24769), .B2(j202_soc_core_intc_core_00_rg_itgt[127]), 
        .Y(n24774) );
  sky130_fd_sc_hd__a22oi_1 U29514 ( .A1(n24772), .A2(
        j202_soc_core_intc_core_00_rg_itgt[119]), .B1(n24771), .B2(
        j202_soc_core_intc_core_00_rg_ipr[95]), .Y(n24773) );
  sky130_fd_sc_hd__nand2_1 U29515 ( .A(n24774), .B(n24773), .Y(n24775) );
  sky130_fd_sc_hd__a21oi_1 U29516 ( .A1(j202_soc_core_intc_core_00_rg_ipr[127]), .A2(n24776), .B1(n24775), .Y(n24778) );
  sky130_fd_sc_hd__nand4_1 U29517 ( .A(n24780), .B(n24779), .C(n24778), .D(
        n24777), .Y(j202_soc_core_ahb2apb_01_N159) );
  sky130_fd_sc_hd__nand2_1 U29518 ( .A(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[0]), .B(n24781), .Y(n24782)
         );
  sky130_fd_sc_hd__o22ai_1 U29519 ( .A1(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[0]), .A2(n24783), .B1(
        j202_soc_core_cmt_core_00_cmt_apb_00_state[1]), .B2(n24782), .Y(
        j202_soc_core_cmt_core_00_cmt_apb_00_nxt_state_0_) );
  sky130_fd_sc_hd__and3_1 U29520 ( .A(n25403), .B(j202_soc_core_prdata[0]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N128) );
  sky130_fd_sc_hd__and3_1 U29521 ( .A(n25403), .B(j202_soc_core_prdata[1]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N129) );
  sky130_fd_sc_hd__and3_1 U29522 ( .A(n25403), .B(j202_soc_core_prdata[2]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N130) );
  sky130_fd_sc_hd__and3_1 U29523 ( .A(n25403), .B(j202_soc_core_prdata[3]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N131) );
  sky130_fd_sc_hd__and3_1 U29524 ( .A(n25403), .B(j202_soc_core_prdata[4]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N132) );
  sky130_fd_sc_hd__and3_1 U29525 ( .A(n25403), .B(j202_soc_core_prdata[5]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N133) );
  sky130_fd_sc_hd__and3_1 U29526 ( .A(n25403), .B(j202_soc_core_prdata[6]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N134) );
  sky130_fd_sc_hd__and3_1 U29527 ( .A(n25403), .B(j202_soc_core_prdata[7]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N135) );
  sky130_fd_sc_hd__and3_1 U29528 ( .A(n25403), .B(j202_soc_core_prdata[8]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N136) );
  sky130_fd_sc_hd__and3_1 U29529 ( .A(n25403), .B(j202_soc_core_prdata[9]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N137) );
  sky130_fd_sc_hd__and3_1 U29530 ( .A(n25403), .B(j202_soc_core_prdata[10]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N138) );
  sky130_fd_sc_hd__and3_1 U29531 ( .A(n25403), .B(j202_soc_core_prdata[11]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N139) );
  sky130_fd_sc_hd__and3_1 U29532 ( .A(n25403), .B(j202_soc_core_prdata[12]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N140) );
  sky130_fd_sc_hd__and3_1 U29533 ( .A(n25403), .B(j202_soc_core_prdata[13]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N141) );
  sky130_fd_sc_hd__and3_1 U29534 ( .A(n25403), .B(j202_soc_core_prdata[14]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N142) );
  sky130_fd_sc_hd__and3_1 U29535 ( .A(n25403), .B(j202_soc_core_prdata[15]), 
        .C(n25734), .X(j202_soc_core_ahb2apb_00_N143) );
  sky130_fd_sc_hd__or3_1 U29536 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[2]), .C(n24784), .X(io_out[12]) );
  sky130_fd_sc_hd__or3_1 U29537 ( .A(
        j202_soc_core_wbqspiflash_00_spif_override), .B(
        j202_soc_core_wbqspiflash_00_w_qspi_dat[3]), .C(n24784), .X(io_out[13]) );
  sky130_fd_sc_hd__clkinv_1 U29538 ( .A(j202_soc_core_uart_BRG_br_cnt[1]), .Y(
        n24786) );
  sky130_fd_sc_hd__o22ai_1 U29539 ( .A1(n24787), .A2(
        j202_soc_core_uart_BRG_br_cnt[0]), .B1(n24786), .B2(
        j202_soc_core_uart_div1[1]), .Y(n24785) );
  sky130_fd_sc_hd__a221oi_1 U29540 ( .A1(n24787), .A2(
        j202_soc_core_uart_BRG_br_cnt[0]), .B1(j202_soc_core_uart_div1[1]), 
        .B2(n24786), .C1(n24785), .Y(n24796) );
  sky130_fd_sc_hd__clkinv_1 U29541 ( .A(j202_soc_core_uart_BRG_br_cnt[7]), .Y(
        n24789) );
  sky130_fd_sc_hd__o22ai_1 U29542 ( .A1(n24790), .A2(
        j202_soc_core_uart_BRG_br_cnt[3]), .B1(n24789), .B2(
        j202_soc_core_uart_div1[7]), .Y(n24788) );
  sky130_fd_sc_hd__a221oi_1 U29543 ( .A1(n24790), .A2(
        j202_soc_core_uart_BRG_br_cnt[3]), .B1(j202_soc_core_uart_div1[7]), 
        .B2(n24789), .C1(n24788), .Y(n24795) );
  sky130_fd_sc_hd__clkinv_1 U29544 ( .A(j202_soc_core_uart_BRG_br_cnt[5]), .Y(
        n24792) );
  sky130_fd_sc_hd__o22ai_1 U29545 ( .A1(n24793), .A2(
        j202_soc_core_uart_BRG_br_cnt[4]), .B1(n24792), .B2(
        j202_soc_core_uart_div1[5]), .Y(n24791) );
  sky130_fd_sc_hd__a221oi_1 U29546 ( .A1(n24793), .A2(
        j202_soc_core_uart_BRG_br_cnt[4]), .B1(j202_soc_core_uart_div1[5]), 
        .B2(n24792), .C1(n24791), .Y(n24794) );
  sky130_fd_sc_hd__nand3_1 U29547 ( .A(n24796), .B(n24795), .C(n24794), .Y(
        n24801) );
  sky130_fd_sc_hd__o22ai_1 U29548 ( .A1(j202_soc_core_uart_div1[2]), .A2(
        n24798), .B1(n24797), .B2(j202_soc_core_uart_BRG_br_cnt[2]), .Y(n24800) );
  sky130_fd_sc_hd__nor2_1 U29549 ( .A(n24802), .B(j202_soc_core_uart_div1[6]), 
        .Y(n24799) );
  sky130_fd_sc_hd__a2111oi_0 U29550 ( .A1(j202_soc_core_uart_div1[6]), .A2(
        n24802), .B1(n24801), .C1(n24800), .D1(n24799), .Y(
        j202_soc_core_uart_BRG_N47) );
  sky130_fd_sc_hd__o22ai_1 U29551 ( .A1(n24805), .A2(
        j202_soc_core_uart_BRG_ps[7]), .B1(n24804), .B2(
        j202_soc_core_uart_BRG_ps[4]), .Y(n24803) );
  sky130_fd_sc_hd__a221oi_1 U29552 ( .A1(n24805), .A2(
        j202_soc_core_uart_BRG_ps[7]), .B1(j202_soc_core_uart_BRG_ps[4]), .B2(
        n24804), .C1(n24803), .Y(n24814) );
  sky130_fd_sc_hd__clkinv_1 U29553 ( .A(j202_soc_core_uart_div0[5]), .Y(n24808) );
  sky130_fd_sc_hd__o22ai_1 U29554 ( .A1(n24808), .A2(
        j202_soc_core_uart_BRG_ps[5]), .B1(n24807), .B2(
        j202_soc_core_uart_BRG_ps[3]), .Y(n24806) );
  sky130_fd_sc_hd__a221oi_1 U29555 ( .A1(n24808), .A2(
        j202_soc_core_uart_BRG_ps[5]), .B1(j202_soc_core_uart_BRG_ps[3]), .B2(
        n24807), .C1(n24806), .Y(n24813) );
  sky130_fd_sc_hd__clkinv_1 U29556 ( .A(j202_soc_core_uart_div0[0]), .Y(n24811) );
  sky130_fd_sc_hd__clkinv_1 U29557 ( .A(j202_soc_core_uart_div0[1]), .Y(n24810) );
  sky130_fd_sc_hd__o22ai_1 U29558 ( .A1(n24811), .A2(
        j202_soc_core_uart_BRG_ps[0]), .B1(n24810), .B2(
        j202_soc_core_uart_BRG_ps[1]), .Y(n24809) );
  sky130_fd_sc_hd__a221oi_1 U29559 ( .A1(n24811), .A2(
        j202_soc_core_uart_BRG_ps[0]), .B1(j202_soc_core_uart_BRG_ps[1]), .B2(
        n24810), .C1(n24809), .Y(n24812) );
  sky130_fd_sc_hd__nand3_1 U29560 ( .A(n24814), .B(n24813), .C(n24812), .Y(
        n24819) );
  sky130_fd_sc_hd__o22ai_1 U29561 ( .A1(j202_soc_core_uart_div0[2]), .A2(
        n24816), .B1(n24815), .B2(j202_soc_core_uart_BRG_ps[2]), .Y(n24818) );
  sky130_fd_sc_hd__nor2_1 U29562 ( .A(n24820), .B(j202_soc_core_uart_div0[6]), 
        .Y(n24817) );
  sky130_fd_sc_hd__a2111oi_0 U29563 ( .A1(j202_soc_core_uart_div0[6]), .A2(
        n24820), .B1(n24819), .C1(n24818), .D1(n24817), .Y(
        j202_soc_core_uart_BRG_N21) );
  sky130_fd_sc_hd__nand2_1 U29564 ( .A(n25731), .B(n24821), .Y(n10676) );
  sky130_fd_sc_hd__nand2_1 U29565 ( .A(n24824), .B(n24823), .Y(n10675) );
  sky130_fd_sc_hd__nand2_1 U29566 ( .A(n24828), .B(n24827), .Y(n24837) );
  sky130_fd_sc_hd__nand3b_1 U29567 ( .A_N(n24830), .B(n24829), .C(n24837), .Y(
        n24831) );
  sky130_fd_sc_hd__nor4_1 U29568 ( .A(n24834), .B(n24833), .C(n24832), .D(
        n24831), .Y(n24836) );
  sky130_fd_sc_hd__o21ai_1 U29569 ( .A1(n24836), .A2(n24882), .B1(n24845), .Y(
        n10599) );
  sky130_fd_sc_hd__nand3_1 U29570 ( .A(n24839), .B(n24838), .C(n24837), .Y(
        n24840) );
  sky130_fd_sc_hd__nand4_1 U29572 ( .A(n24874), .B(n24844), .C(n24843), .D(
        n24842), .Y(n10598) );
  sky130_fd_sc_hd__o21ai_1 U29573 ( .A1(n24846), .A2(n24882), .B1(n24845), .Y(
        n10597) );
  sky130_fd_sc_hd__o21ai_1 U29574 ( .A1(n24848), .A2(n24847), .B1(n24858), .Y(
        n24852) );
  sky130_fd_sc_hd__a21oi_1 U29575 ( .A1(n24850), .A2(n24849), .B1(n24882), .Y(
        n24851) );
  sky130_fd_sc_hd__nor2_1 U29576 ( .A(n24857), .B(n24851), .Y(n24855) );
  sky130_fd_sc_hd__nand2_1 U29577 ( .A(n24852), .B(n24855), .Y(n10586) );
  sky130_fd_sc_hd__nand2_1 U29579 ( .A(n24856), .B(n24855), .Y(n10585) );
  sky130_fd_sc_hd__a21o_1 U29580 ( .A1(n24859), .A2(n24858), .B1(n24857), .X(
        n10584) );
  sky130_fd_sc_hd__a31oi_1 U29581 ( .A1(n24861), .A2(n24860), .A3(n24868), 
        .B1(n24882), .Y(n24862) );
  sky130_fd_sc_hd__nand2_1 U29583 ( .A(n24865), .B(n24864), .Y(n10565) );
  sky130_fd_sc_hd__nand2_1 U29584 ( .A(n24867), .B(n24866), .Y(n24883) );
  sky130_fd_sc_hd__a31oi_1 U29586 ( .A1(n24873), .A2(n24872), .A3(n24871), 
        .B1(n24870), .Y(n24875) );
  sky130_fd_sc_hd__a211oi_1 U29588 ( .A1(n24879), .A2(n24878), .B1(n24877), 
        .C1(n24876), .Y(n24881) );
  sky130_fd_sc_hd__o21ai_1 U29589 ( .A1(n24881), .A2(n24890), .B1(n24889), .Y(
        n10564) );
  sky130_fd_sc_hd__a21oi_1 U29590 ( .A1(n24884), .A2(n24883), .B1(n24882), .Y(
        n24887) );
  sky130_fd_sc_hd__nor3_1 U29591 ( .A(n24888), .B(n24887), .C(n24886), .Y(
        n24891) );
  sky130_fd_sc_hd__o21ai_1 U29592 ( .A1(n24891), .A2(n24890), .B1(n24889), .Y(
        n10563) );
  sky130_fd_sc_hd__nand2_1 U29593 ( .A(n24893), .B(n24892), .Y(n10558) );
  sky130_fd_sc_hd__nor2_1 U29594 ( .A(j202_soc_core_j22_cpu_id_op2_v_), .B(
        n24894), .Y(n24896) );
  sky130_fd_sc_hd__or4_1 U29595 ( .A(n24897), .B(n24896), .C(n24895), .D(
        n25434), .X(n10533) );
  sky130_fd_sc_hd__a21oi_1 U29596 ( .A1(n25043), .A2(n25042), .B1(n24898), .Y(
        n24988) );
  sky130_fd_sc_hd__nand2_1 U29597 ( .A(n24899), .B(n24910), .Y(n25009) );
  sky130_fd_sc_hd__a22oi_1 U29598 ( .A1(j202_soc_core_qspi_wb_addr[2]), .A2(
        n25041), .B1(n25086), .B2(j202_soc_core_wbqspiflash_00_spif_data[2]), 
        .Y(n24900) );
  sky130_fd_sc_hd__a22oi_1 U29600 ( .A1(n25041), .A2(
        j202_soc_core_qspi_wb_addr[3]), .B1(n25086), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[3]), .Y(n24902) );
  sky130_fd_sc_hd__o21ai_1 U29601 ( .A1(n24988), .A2(n24903), .B1(n24902), .Y(
        n10531) );
  sky130_fd_sc_hd__a22oi_1 U29602 ( .A1(n25041), .A2(
        j202_soc_core_qspi_wb_addr[4]), .B1(n25086), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[4]), .Y(n24904) );
  sky130_fd_sc_hd__o21ai_1 U29603 ( .A1(n24988), .A2(n24905), .B1(n24904), .Y(
        n10530) );
  sky130_fd_sc_hd__nor2_1 U29604 ( .A(n25081), .B(n25080), .Y(n24913) );
  sky130_fd_sc_hd__a22oi_1 U29605 ( .A1(n24911), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[5]), .B1(n24910), .B2(
        j202_soc_core_qspi_wb_addr[5]), .Y(n24906) );
  sky130_fd_sc_hd__o211ai_1 U29606 ( .A1(n24988), .A2(n24907), .B1(n24913), 
        .C1(n24906), .Y(n10529) );
  sky130_fd_sc_hd__a22oi_1 U29607 ( .A1(n25041), .A2(
        j202_soc_core_qspi_wb_addr[6]), .B1(n25086), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[6]), .Y(n24908) );
  sky130_fd_sc_hd__o21ai_1 U29608 ( .A1(n24988), .A2(n24909), .B1(n24908), .Y(
        n10528) );
  sky130_fd_sc_hd__a22oi_1 U29609 ( .A1(n24911), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[7]), .B1(n24910), .B2(
        j202_soc_core_qspi_wb_addr[7]), .Y(n24912) );
  sky130_fd_sc_hd__o211ai_1 U29610 ( .A1(n24988), .A2(n24914), .B1(n24913), 
        .C1(n24912), .Y(n10527) );
  sky130_fd_sc_hd__o22ai_1 U29611 ( .A1(n24940), .A2(n24988), .B1(n24939), 
        .B2(n25009), .Y(n24915) );
  sky130_fd_sc_hd__a21oi_1 U29612 ( .A1(n25086), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[8]), .B1(n24915), .Y(n24916) );
  sky130_fd_sc_hd__o21ai_1 U29613 ( .A1(n25010), .A2(n24938), .B1(n24916), .Y(
        n10526) );
  sky130_fd_sc_hd__a22oi_1 U29614 ( .A1(j202_soc_core_qspi_wb_addr[9]), .A2(
        n25041), .B1(n25086), .B2(j202_soc_core_wbqspiflash_00_spif_data[9]), 
        .Y(n24918) );
  sky130_fd_sc_hd__o211ai_1 U29615 ( .A1(n24988), .A2(n24919), .B1(n24918), 
        .C1(n24917), .Y(n10525) );
  sky130_fd_sc_hd__a22oi_1 U29616 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .A2(n25080), .B1(n25086), 
        .B2(j202_soc_core_wbqspiflash_00_spif_data[10]), .Y(n24921) );
  sky130_fd_sc_hd__a222oi_1 U29617 ( .A1(n24991), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[2]), .B1(
        j202_soc_core_qspi_wb_addr[10]), .B2(n25041), .C1(n25081), .C2(
        j202_soc_core_qspi_wb_addr[2]), .Y(n24920) );
  sky130_fd_sc_hd__o211ai_1 U29618 ( .A1(n24988), .A2(n24922), .B1(n24921), 
        .C1(n24920), .Y(n10524) );
  sky130_fd_sc_hd__a22oi_1 U29619 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .A2(n25080), .B1(n25086), 
        .B2(j202_soc_core_wbqspiflash_00_spif_data[11]), .Y(n24924) );
  sky130_fd_sc_hd__a222oi_1 U29620 ( .A1(n24991), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[3]), .B1(n25041), .B2(
        j202_soc_core_qspi_wb_addr[11]), .C1(n25081), .C2(
        j202_soc_core_qspi_wb_addr[3]), .Y(n24923) );
  sky130_fd_sc_hd__o211ai_1 U29621 ( .A1(n24988), .A2(n24925), .B1(n24924), 
        .C1(n24923), .Y(n10523) );
  sky130_fd_sc_hd__a22oi_1 U29622 ( .A1(n25086), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[12]), .B1(n24991), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[4]), .Y(n24927) );
  sky130_fd_sc_hd__a222oi_1 U29623 ( .A1(n25081), .A2(
        j202_soc_core_qspi_wb_addr[4]), .B1(n25041), .B2(
        j202_soc_core_qspi_wb_addr[12]), .C1(n25080), .C2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[4]), .Y(n24926) );
  sky130_fd_sc_hd__o211ai_1 U29624 ( .A1(n24988), .A2(n24967), .B1(n24927), 
        .C1(n24926), .Y(n10522) );
  sky130_fd_sc_hd__a22oi_1 U29625 ( .A1(
        j202_soc_core_wbqspiflash_00_spif_data[5]), .A2(n24991), .B1(n25086), 
        .B2(j202_soc_core_wbqspiflash_00_spif_data[13]), .Y(n24929) );
  sky130_fd_sc_hd__a222oi_1 U29626 ( .A1(n25081), .A2(
        j202_soc_core_qspi_wb_addr[5]), .B1(n25041), .B2(
        j202_soc_core_qspi_wb_addr[13]), .C1(n25080), .C2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[5]), .Y(n24928) );
  sky130_fd_sc_hd__o211ai_1 U29627 ( .A1(n24988), .A2(n24975), .B1(n24929), 
        .C1(n24928), .Y(n10521) );
  sky130_fd_sc_hd__a22oi_1 U29628 ( .A1(n24991), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[6]), .B1(n25081), .B2(
        j202_soc_core_qspi_wb_addr[6]), .Y(n24934) );
  sky130_fd_sc_hd__nand2_1 U29629 ( .A(j202_soc_core_qspi_wb_addr[14]), .B(
        n25041), .Y(n24932) );
  sky130_fd_sc_hd__nand2_1 U29630 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[6]), .B(n25080), .Y(n24931)
         );
  sky130_fd_sc_hd__nand2_1 U29631 ( .A(
        j202_soc_core_wbqspiflash_00_spif_data[14]), .B(n25086), .Y(n24930) );
  sky130_fd_sc_hd__and3_1 U29632 ( .A(n24932), .B(n24931), .C(n24930), .X(
        n24933) );
  sky130_fd_sc_hd__o211ai_1 U29633 ( .A1(n24988), .A2(n24935), .B1(n24934), 
        .C1(n24933), .Y(n10520) );
  sky130_fd_sc_hd__a22oi_1 U29634 ( .A1(n25086), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[15]), .B1(n24991), .B2(
        j202_soc_core_wbqspiflash_00_spif_data[7]), .Y(n24937) );
  sky130_fd_sc_hd__a222oi_1 U29635 ( .A1(n25081), .A2(
        j202_soc_core_qspi_wb_addr[7]), .B1(j202_soc_core_qspi_wb_addr[15]), 
        .B2(n25041), .C1(n25080), .C2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[7]), .Y(n24936) );
  sky130_fd_sc_hd__o211ai_1 U29636 ( .A1(n24988), .A2(n24987), .B1(n24937), 
        .C1(n24936), .Y(n10519) );
  sky130_fd_sc_hd__nor2_1 U29637 ( .A(n24960), .B(n24938), .Y(n24948) );
  sky130_fd_sc_hd__o22ai_1 U29638 ( .A1(n25090), .A2(n24940), .B1(n24939), 
        .B2(n25055), .Y(n24947) );
  sky130_fd_sc_hd__a22oi_1 U29639 ( .A1(n25086), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[16]), .B1(n24991), .B2(
        j202_soc_core_wbqspiflash_00_last_status[0]), .Y(n24941) );
  sky130_fd_sc_hd__clkinv_1 U29641 ( .A(j202_soc_core_qspi_wb_addr[16]), .Y(
        n24943) );
  sky130_fd_sc_hd__o22ai_1 U29642 ( .A1(n24944), .A2(n24988), .B1(n24943), 
        .B2(n25009), .Y(n24945) );
  sky130_fd_sc_hd__or4_1 U29643 ( .A(n24948), .B(n24947), .C(n24946), .D(
        n24945), .X(n10518) );
  sky130_fd_sc_hd__a22oi_1 U29644 ( .A1(n25044), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[15]), .B1(n24991), .B2(
        j202_soc_core_wbqspiflash_00_last_status[1]), .Y(n24953) );
  sky130_fd_sc_hd__a22oi_1 U29645 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[9]), .A2(n25080), .B1(n25086), 
        .B2(j202_soc_core_wbqspiflash_00_spif_data[17]), .Y(n24952) );
  sky130_fd_sc_hd__a22oi_1 U29646 ( .A1(n24954), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[1]), .B1(n25081), .B2(
        j202_soc_core_qspi_wb_addr[9]), .Y(n24949) );
  sky130_fd_sc_hd__o21ai_1 U29647 ( .A1(n25019), .A2(n24988), .B1(n24949), .Y(
        n24950) );
  sky130_fd_sc_hd__a21oi_1 U29648 ( .A1(n25041), .A2(
        j202_soc_core_qspi_wb_addr[17]), .B1(n24950), .Y(n24951) );
  sky130_fd_sc_hd__nand3_1 U29649 ( .A(n24953), .B(n24952), .C(n24951), .Y(
        n10517) );
  sky130_fd_sc_hd__a22oi_1 U29650 ( .A1(n24954), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[2]), .B1(n25081), .B2(
        j202_soc_core_qspi_wb_addr[10]), .Y(n24958) );
  sky130_fd_sc_hd__a22oi_1 U29651 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[10]), .A2(n25080), .B1(n25044), .B2(j202_soc_core_wbqspiflash_00_spif_data[16]), .Y(n24957) );
  sky130_fd_sc_hd__a22oi_1 U29652 ( .A1(n25086), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[18]), .B1(n24991), .B2(
        j202_soc_core_wbqspiflash_00_last_status[2]), .Y(n24956) );
  sky130_fd_sc_hd__clkinv_1 U29653 ( .A(n24988), .Y(n24981) );
  sky130_fd_sc_hd__a22oi_1 U29654 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .A2(n24981), .B1(
        j202_soc_core_qspi_wb_addr[18]), .B2(n25041), .Y(n24955) );
  sky130_fd_sc_hd__nand4_1 U29655 ( .A(n24958), .B(n24957), .C(n24956), .D(
        n24955), .Y(n10516) );
  sky130_fd_sc_hd__a22oi_1 U29656 ( .A1(
        j202_soc_core_wbqspiflash_00_spif_data[17]), .A2(n25044), .B1(n25081), 
        .B2(j202_soc_core_qspi_wb_addr[11]), .Y(n24965) );
  sky130_fd_sc_hd__nor2_1 U29657 ( .A(n24960), .B(n24959), .Y(n24961) );
  sky130_fd_sc_hd__a21oi_1 U29658 ( .A1(n25080), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[11]), .B1(n24961), .Y(n24964)
         );
  sky130_fd_sc_hd__a22oi_1 U29659 ( .A1(n25086), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[19]), .B1(n24991), .B2(
        j202_soc_core_wbqspiflash_00_last_status[3]), .Y(n24963) );
  sky130_fd_sc_hd__a22oi_1 U29660 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .A2(n24981), .B1(
        j202_soc_core_qspi_wb_addr[19]), .B2(n25041), .Y(n24962) );
  sky130_fd_sc_hd__nand4_1 U29661 ( .A(n24965), .B(n24964), .C(n24963), .D(
        n24962), .Y(n10515) );
  sky130_fd_sc_hd__a22oi_1 U29662 ( .A1(n25086), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[20]), .B1(n25081), .B2(
        j202_soc_core_qspi_wb_addr[12]), .Y(n24972) );
  sky130_fd_sc_hd__o22ai_1 U29663 ( .A1(n24967), .A2(n25090), .B1(n24974), 
        .B2(n24966), .Y(n24968) );
  sky130_fd_sc_hd__a21oi_1 U29664 ( .A1(n24991), .A2(
        j202_soc_core_wbqspiflash_00_last_status[4]), .B1(n24968), .Y(n24971)
         );
  sky130_fd_sc_hd__a22oi_1 U29665 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[20]), .A2(n24981), .B1(
        j202_soc_core_qspi_wb_addr[20]), .B2(n25041), .Y(n24970) );
  sky130_fd_sc_hd__nand4_1 U29666 ( .A(n24972), .B(n24971), .C(n24970), .D(
        n24969), .Y(n10514) );
  sky130_fd_sc_hd__a22oi_1 U29667 ( .A1(n25086), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[21]), .B1(n25081), .B2(
        j202_soc_core_qspi_wb_addr[13]), .Y(n24980) );
  sky130_fd_sc_hd__o22ai_1 U29668 ( .A1(n24975), .A2(n25090), .B1(n24974), 
        .B2(n24973), .Y(n24976) );
  sky130_fd_sc_hd__a21oi_1 U29669 ( .A1(
        j202_soc_core_wbqspiflash_00_last_status[5]), .A2(n24991), .B1(n24976), 
        .Y(n24979) );
  sky130_fd_sc_hd__a22oi_1 U29670 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[21]), .A2(n24981), .B1(
        j202_soc_core_qspi_wb_addr[21]), .B2(n25041), .Y(n24978) );
  sky130_fd_sc_hd__nand4_1 U29671 ( .A(n24980), .B(n24979), .C(n24978), .D(
        n24977), .Y(n10513) );
  sky130_fd_sc_hd__a22oi_1 U29672 ( .A1(
        j202_soc_core_wbqspiflash_00_last_status[6]), .A2(n24991), .B1(n25086), 
        .B2(j202_soc_core_wbqspiflash_00_spif_data[22]), .Y(n24985) );
  sky130_fd_sc_hd__a22oi_1 U29673 ( .A1(n25080), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[14]), .B1(n25081), .B2(
        j202_soc_core_qspi_wb_addr[14]), .Y(n24984) );
  sky130_fd_sc_hd__a22oi_1 U29674 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .A2(n24981), .B1(
        j202_soc_core_qspi_wb_addr[22]), .B2(n25041), .Y(n24983) );
  sky130_fd_sc_hd__nand4_1 U29675 ( .A(n24985), .B(n24984), .C(n24983), .D(
        n24982), .Y(n10512) );
  sky130_fd_sc_hd__o22ai_1 U29676 ( .A1(n25090), .A2(n24987), .B1(n24986), 
        .B2(n25055), .Y(n24990) );
  sky130_fd_sc_hd__o22ai_1 U29677 ( .A1(n25089), .A2(n24988), .B1(n25088), 
        .B2(n25009), .Y(n24989) );
  sky130_fd_sc_hd__a211oi_1 U29678 ( .A1(n24991), .A2(
        j202_soc_core_wbqspiflash_00_last_status[7]), .B1(n24990), .C1(n24989), 
        .Y(n24994) );
  sky130_fd_sc_hd__nand2_1 U29679 ( .A(n25086), .B(
        j202_soc_core_wbqspiflash_00_spif_data[23]), .Y(n24992) );
  sky130_fd_sc_hd__nand3_1 U29680 ( .A(n24994), .B(n24993), .C(n24992), .Y(
        n10511) );
  sky130_fd_sc_hd__nand2_1 U29681 ( .A(n24996), .B(n24995), .Y(n25016) );
  sky130_fd_sc_hd__nand2_1 U29682 ( .A(n25093), .B(n25051), .Y(n24997) );
  sky130_fd_sc_hd__o31ai_1 U29683 ( .A1(j202_soc_core_wbqspiflash_00_state[3]), 
        .A2(n24998), .A3(n25016), .B1(n24997), .Y(n24999) );
  sky130_fd_sc_hd__a21oi_1 U29684 ( .A1(n25086), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[24]), .B1(n24999), .Y(n25008)
         );
  sky130_fd_sc_hd__nand2_1 U29685 ( .A(n25001), .B(n25000), .Y(n25003) );
  sky130_fd_sc_hd__nand4_1 U29686 ( .A(n25004), .B(n25003), .C(n25002), .D(
        n25065), .Y(n25033) );
  sky130_fd_sc_hd__clkinv_1 U29687 ( .A(n25033), .Y(n25007) );
  sky130_fd_sc_hd__nand2_1 U29688 ( .A(n25005), .B(n25063), .Y(n25014) );
  sky130_fd_sc_hd__nor2_1 U29689 ( .A(j202_soc_core_wbqspiflash_00_state[3]), 
        .B(n25014), .Y(n25034) );
  sky130_fd_sc_hd__a22oi_1 U29690 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[16]), .A2(n25080), .B1(n25034), .B2(j202_soc_core_qspi_wb_addr[16]), .Y(n25006) );
  sky130_fd_sc_hd__and3_1 U29691 ( .A(n25008), .B(n25007), .C(n25006), .X(
        n25012) );
  sky130_fd_sc_hd__nand4_1 U29692 ( .A(n25012), .B(n25011), .C(n25010), .D(
        n25009), .Y(n10510) );
  sky130_fd_sc_hd__clkinv_1 U29693 ( .A(n25013), .Y(n25030) );
  sky130_fd_sc_hd__clkinv_1 U29694 ( .A(n25014), .Y(n25021) );
  sky130_fd_sc_hd__nor2_1 U29695 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .B(n25015), .Y(n25017)
         );
  sky130_fd_sc_hd__o22ai_1 U29696 ( .A1(n25019), .A2(n25018), .B1(n25017), 
        .B2(n25016), .Y(n25020) );
  sky130_fd_sc_hd__a21oi_1 U29697 ( .A1(n25021), .A2(
        j202_soc_core_qspi_wb_addr[17]), .B1(n25020), .Y(n25022) );
  sky130_fd_sc_hd__a22oi_1 U29699 ( .A1(n25027), .A2(n25026), .B1(n25025), 
        .B2(j202_soc_core_wbqspiflash_00_spif_data[25]), .Y(n25028) );
  sky130_fd_sc_hd__o211ai_1 U29700 ( .A1(n25030), .A2(n25029), .B1(n25112), 
        .C1(n25028), .Y(n10509) );
  sky130_fd_sc_hd__a21oi_1 U29701 ( .A1(n25032), .A2(n25031), .B1(n25046), .Y(
        n25040) );
  sky130_fd_sc_hd__a22oi_1 U29702 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[18]), .A2(n25080), .B1(n25086), .B2(j202_soc_core_wbqspiflash_00_spif_data[26]), .Y(n25038) );
  sky130_fd_sc_hd__a21oi_1 U29703 ( .A1(j202_soc_core_qspi_wb_addr[18]), .A2(
        n25034), .B1(n25033), .Y(n25037) );
  sky130_fd_sc_hd__nand4_1 U29704 ( .A(n25038), .B(n25037), .C(n25036), .D(
        n25035), .Y(n25039) );
  sky130_fd_sc_hd__or4_1 U29705 ( .A(n25093), .B(n25077), .C(n25040), .D(
        n25039), .X(n10508) );
  sky130_fd_sc_hd__a21oi_1 U29706 ( .A1(n25043), .A2(n25042), .B1(n25041), .Y(
        n25062) );
  sky130_fd_sc_hd__clkinv_1 U29707 ( .A(n25094), .Y(n25045) );
  sky130_fd_sc_hd__nor2_1 U29708 ( .A(n25044), .B(n25077), .Y(n25084) );
  sky130_fd_sc_hd__a21oi_1 U29710 ( .A1(n25048), .A2(n25047), .B1(n25058), .Y(
        n25097) );
  sky130_fd_sc_hd__a22oi_1 U29711 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[19]), .A2(n25080), .B1(n25093), .B2(n25094), .Y(n25050) );
  sky130_fd_sc_hd__a22oi_1 U29712 ( .A1(n25086), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[27]), .B1(n25081), .B2(
        j202_soc_core_qspi_wb_addr[19]), .Y(n25049) );
  sky130_fd_sc_hd__nand4_1 U29713 ( .A(n25062), .B(n25097), .C(n25050), .D(
        n25049), .Y(n10507) );
  sky130_fd_sc_hd__nand3_1 U29714 ( .A(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .B(n25093), .C(n25051), 
        .Y(n25079) );
  sky130_fd_sc_hd__clkinv_1 U29716 ( .A(j202_soc_core_qspi_wb_addr[20]), .Y(
        n25054) );
  sky130_fd_sc_hd__o22ai_1 U29717 ( .A1(n25055), .A2(n25054), .B1(n25053), 
        .B2(n25065), .Y(n25056) );
  sky130_fd_sc_hd__nor3_1 U29718 ( .A(n25058), .B(n25057), .C(n25056), .Y(
        n25060) );
  sky130_fd_sc_hd__nand2_1 U29719 ( .A(n25086), .B(
        j202_soc_core_wbqspiflash_00_spif_data[28]), .Y(n25059) );
  sky130_fd_sc_hd__nand4_1 U29720 ( .A(n25060), .B(n25073), .C(n25072), .D(
        n25059), .Y(n10506) );
  sky130_fd_sc_hd__nor2_1 U29721 ( .A(n25062), .B(n25061), .Y(n25092) );
  sky130_fd_sc_hd__nand2_1 U29722 ( .A(n25064), .B(n25063), .Y(n25087) );
  sky130_fd_sc_hd__o22ai_1 U29723 ( .A1(n25087), .A2(n25067), .B1(n25066), 
        .B2(n25065), .Y(n25076) );
  sky130_fd_sc_hd__a21oi_1 U29724 ( .A1(n25070), .A2(n25069), .B1(n25068), .Y(
        n25071) );
  sky130_fd_sc_hd__a21oi_1 U29725 ( .A1(
        j202_soc_core_wbqspiflash_00_spif_data[29]), .A2(n25086), .B1(n25071), 
        .Y(n25074) );
  sky130_fd_sc_hd__nand3_1 U29726 ( .A(n25074), .B(n25073), .C(n25072), .Y(
        n25075) );
  sky130_fd_sc_hd__nor4_1 U29727 ( .A(n25077), .B(n25092), .C(n25076), .D(
        n25075), .Y(n25078) );
  sky130_fd_sc_hd__a22oi_1 U29729 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[22]), .A2(n25080), .B1(n25086), .B2(j202_soc_core_wbqspiflash_00_spif_data[30]), .Y(n25083) );
  sky130_fd_sc_hd__a21oi_1 U29730 ( .A1(j202_soc_core_qspi_wb_addr[22]), .A2(
        n25081), .B1(n25092), .Y(n25082) );
  sky130_fd_sc_hd__nand3_1 U29731 ( .A(n25084), .B(n25083), .C(n25082), .Y(
        n10504) );
  sky130_fd_sc_hd__a21oi_1 U29732 ( .A1(
        j202_soc_core_wbqspiflash_00_spif_data[31]), .A2(n25086), .B1(n25085), 
        .Y(n25096) );
  sky130_fd_sc_hd__o22ai_1 U29733 ( .A1(n25090), .A2(n25089), .B1(n25088), 
        .B2(n25087), .Y(n25091) );
  sky130_fd_sc_hd__a211oi_1 U29734 ( .A1(n25094), .A2(n25093), .B1(n25092), 
        .C1(n25091), .Y(n25095) );
  sky130_fd_sc_hd__nand3_1 U29735 ( .A(n25097), .B(n25096), .C(n25095), .Y(
        n10503) );
  sky130_fd_sc_hd__o21ai_1 U29736 ( .A1(n25100), .A2(n25099), .B1(n25098), .Y(
        n25105) );
  sky130_fd_sc_hd__o21ai_1 U29737 ( .A1(j202_soc_core_wbqspiflash_00_state[3]), 
        .A2(n25102), .B1(n25101), .Y(n25103) );
  sky130_fd_sc_hd__nor4_1 U29738 ( .A(n25106), .B(n25105), .C(n25104), .D(
        n25103), .Y(n25114) );
  sky130_fd_sc_hd__nand2_1 U29740 ( .A(n25110), .B(n25109), .Y(n25113) );
  sky130_fd_sc_hd__a31oi_1 U29741 ( .A1(n25114), .A2(n25113), .A3(n25112), 
        .B1(n25111), .Y(n25115) );
  sky130_fd_sc_hd__a22oi_1 U29742 ( .A1(n25117), .A2(n25116), .B1(
        j202_soc_core_wbqspiflash_00_spif_req), .B2(n25115), .Y(n25120) );
  sky130_fd_sc_hd__nand3_1 U29743 ( .A(n25120), .B(n25119), .C(n25118), .Y(
        n10502) );
  sky130_fd_sc_hd__clkinv_1 U29744 ( .A(wbs_dat_o[0]), .Y(n10484) );
  sky130_fd_sc_hd__a21oi_1 U29745 ( .A1(n25123), .A2(n25122), .B1(n25121), .Y(
        n23) );
  sky130_fd_sc_hd__o21ai_1 U29746 ( .A1(j202_soc_core_uart_TOP_dpll_state[0]), 
        .A2(j202_soc_core_uart_TOP_change), .B1(j202_soc_core_uart_sio_ce_x4), 
        .Y(n25236) );
  sky130_fd_sc_hd__a22o_1 U29747 ( .A1(j202_soc_core_uart_TOP_dpll_state[1]), 
        .A2(n25236), .B1(n25405), .B2(j202_soc_core_uart_sio_ce_x4), .X(n24)
         );
  sky130_fd_sc_hd__clkinv_1 U29748 ( .A(j202_soc_core_bldc_core_00_pwm_en), 
        .Y(n25148) );
  sky130_fd_sc_hd__o22ai_1 U29749 ( .A1(n25126), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]), .B1(n25125), .B2(
        j202_soc_core_bldc_core_00_pwm_duty[11]), .Y(n25124) );
  sky130_fd_sc_hd__a221oi_1 U29750 ( .A1(n25126), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[7]), .B1(
        j202_soc_core_bldc_core_00_pwm_duty[11]), .B2(n25125), .C1(n25124), 
        .Y(n25133) );
  sky130_fd_sc_hd__o22ai_1 U29751 ( .A1(n25128), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .B1(n25186), .B2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .Y(n25127) );
  sky130_fd_sc_hd__a221oi_1 U29752 ( .A1(n25128), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[0]), .B1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[1]), .B2(n25186), .C1(
        n25127), .Y(n25132) );
  sky130_fd_sc_hd__o2bb2ai_1 U29753 ( .B1(
        j202_soc_core_bldc_core_00_pwm_duty[8]), .B2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .A1_N(
        j202_soc_core_bldc_core_00_pwm_duty[8]), .A2_N(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[8]), .Y(n25131) );
  sky130_fd_sc_hd__clkinv_1 U29754 ( .A(
        j202_soc_core_bldc_core_00_pwm_duty[10]), .Y(n25194) );
  sky130_fd_sc_hd__o22ai_1 U29755 ( .A1(
        j202_soc_core_bldc_core_00_pwm_duty[10]), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[10]), .B1(n25194), .B2(
        n25129), .Y(n25130) );
  sky130_fd_sc_hd__nand4_1 U29756 ( .A(n25133), .B(n25132), .C(n25131), .D(
        n25130), .Y(n25146) );
  sky130_fd_sc_hd__o22ai_1 U29757 ( .A1(n25136), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .B1(n25135), .B2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]), .Y(n25134) );
  sky130_fd_sc_hd__a221oi_1 U29758 ( .A1(n25136), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[6]), .B1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[5]), .B2(n25135), .C1(
        n25134), .Y(n25144) );
  sky130_fd_sc_hd__o22ai_1 U29759 ( .A1(n25139), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]), .B1(n25138), .B2(
        j202_soc_core_bldc_core_00_pwm_duty[2]), .Y(n25137) );
  sky130_fd_sc_hd__a221oi_1 U29760 ( .A1(n25139), .A2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[9]), .B1(
        j202_soc_core_bldc_core_00_pwm_duty[2]), .B2(n25138), .C1(n25137), .Y(
        n25143) );
  sky130_fd_sc_hd__o22ai_1 U29761 ( .A1(j202_soc_core_bldc_core_00_pwm_duty[3]), .A2(j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[3]), .B1(n25188), .B2(
        n25140), .Y(n25142) );
  sky130_fd_sc_hd__o2bb2ai_1 U29762 ( .B1(
        j202_soc_core_bldc_core_00_pwm_duty[4]), .B2(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[4]), .A1_N(
        j202_soc_core_bldc_core_00_pwm_duty[4]), .A2_N(
        j202_soc_core_bldc_core_00_bldc_pwm_00_clkcnt[4]), .Y(n25141) );
  sky130_fd_sc_hd__nand4_1 U29763 ( .A(n25144), .B(n25143), .C(n25142), .D(
        n25141), .Y(n25145) );
  sky130_fd_sc_hd__o31ai_1 U29765 ( .A1(io_in[25]), .A2(n25149), .A3(n25148), 
        .B1(n25147), .Y(n26) );
  sky130_fd_sc_hd__o22ai_1 U29766 ( .A1(n25228), .A2(n25151), .B1(n25227), 
        .B2(n25150), .Y(n29) );
  sky130_fd_sc_hd__nand2_1 U29767 ( .A(n25193), .B(
        j202_soc_core_bldc_core_00_wdata[9]), .Y(n25152) );
  sky130_fd_sc_hd__o21ai_1 U29768 ( .A1(n25153), .A2(n25193), .B1(n25152), .Y(
        n30) );
  sky130_fd_sc_hd__o22ai_1 U29769 ( .A1(n25228), .A2(n25155), .B1(n25227), 
        .B2(n25154), .Y(n36) );
  sky130_fd_sc_hd__clkinv_1 U29770 ( .A(j202_soc_core_bldc_core_00_wdata[1]), 
        .Y(n25160) );
  sky130_fd_sc_hd__o22ai_1 U29771 ( .A1(n25193), .A2(n25156), .B1(n25189), 
        .B2(n25160), .Y(n38) );
  sky130_fd_sc_hd__nand2_1 U29772 ( .A(n25158), .B(
        j202_soc_core_bldc_core_00_adc_en), .Y(n25157) );
  sky130_fd_sc_hd__o21ai_1 U29773 ( .A1(n25160), .A2(n25158), .B1(n25157), .Y(
        n39) );
  sky130_fd_sc_hd__nand2_1 U29774 ( .A(n25159), .B(n25164), .Y(n25168) );
  sky130_fd_sc_hd__clkinv_1 U29775 ( .A(n25168), .Y(n25170) );
  sky130_fd_sc_hd__o22ai_1 U29776 ( .A1(n25170), .A2(n25161), .B1(n25168), 
        .B2(n25160), .Y(n40) );
  sky130_fd_sc_hd__a21oi_1 U29778 ( .A1(n25404), .A2(n25171), .B1(n25163), .Y(
        n44) );
  sky130_fd_sc_hd__nand2_1 U29779 ( .A(n25165), .B(n25164), .Y(n25167) );
  sky130_fd_sc_hd__nand2_1 U29780 ( .A(n25167), .B(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bier_0_), .Y(n25166) );
  sky130_fd_sc_hd__o21ai_1 U29781 ( .A1(n25171), .A2(n25167), .B1(n25166), .Y(
        n45) );
  sky130_fd_sc_hd__a22o_1 U29782 ( .A1(n25168), .A2(
        j202_soc_core_bldc_core_00_comm[2]), .B1(n25170), .B2(
        j202_soc_core_bldc_core_00_wdata[2]), .X(n46) );
  sky130_fd_sc_hd__o22ai_1 U29783 ( .A1(n25170), .A2(n25169), .B1(n25168), 
        .B2(n25171), .Y(n47) );
  sky130_fd_sc_hd__a22o_1 U29784 ( .A1(n25193), .A2(
        j202_soc_core_bldc_core_00_wdata[23]), .B1(n25189), .B2(
        j202_soc_core_bldc_core_00_pwm_duty[11]), .X(n49) );
  sky130_fd_sc_hd__o22ai_1 U29785 ( .A1(n25193), .A2(n25172), .B1(n25189), 
        .B2(n25171), .Y(n50) );
  sky130_fd_sc_hd__a22o_1 U29786 ( .A1(n25189), .A2(
        j202_soc_core_bldc_core_00_pwm_period[2]), .B1(n25193), .B2(
        j202_soc_core_bldc_core_00_wdata[2]), .X(n51) );
  sky130_fd_sc_hd__a22o_1 U29787 ( .A1(n25193), .A2(
        j202_soc_core_bldc_core_00_wdata[3]), .B1(n25189), .B2(
        j202_soc_core_bldc_core_00_pwm_period[3]), .X(n52) );
  sky130_fd_sc_hd__nand2_1 U29788 ( .A(n25193), .B(
        j202_soc_core_bldc_core_00_wdata[4]), .Y(n25173) );
  sky130_fd_sc_hd__nand2_1 U29790 ( .A(n25193), .B(
        j202_soc_core_bldc_core_00_wdata[5]), .Y(n25175) );
  sky130_fd_sc_hd__o21ai_1 U29791 ( .A1(n25176), .A2(n25193), .B1(n25175), .Y(
        n54) );
  sky130_fd_sc_hd__nand2_1 U29792 ( .A(n25193), .B(
        j202_soc_core_bldc_core_00_wdata[6]), .Y(n25177) );
  sky130_fd_sc_hd__o21ai_1 U29793 ( .A1(n25178), .A2(n25193), .B1(n25177), .Y(
        n55) );
  sky130_fd_sc_hd__nand2_1 U29794 ( .A(n25193), .B(
        j202_soc_core_bldc_core_00_wdata[7]), .Y(n25179) );
  sky130_fd_sc_hd__o21ai_1 U29795 ( .A1(n25180), .A2(n25193), .B1(n25179), .Y(
        n56) );
  sky130_fd_sc_hd__nand2_1 U29796 ( .A(n25193), .B(
        j202_soc_core_bldc_core_00_wdata[8]), .Y(n25181) );
  sky130_fd_sc_hd__o21ai_1 U29797 ( .A1(n25182), .A2(n25193), .B1(n25181), .Y(
        n57) );
  sky130_fd_sc_hd__a22o_1 U29798 ( .A1(n25193), .A2(
        j202_soc_core_bldc_core_00_wdata[10]), .B1(n25189), .B2(
        j202_soc_core_bldc_core_00_pwm_period[10]), .X(n58) );
  sky130_fd_sc_hd__nand2_1 U29799 ( .A(n25193), .B(
        j202_soc_core_bldc_core_00_wdata[11]), .Y(n25183) );
  sky130_fd_sc_hd__o21ai_1 U29800 ( .A1(n25184), .A2(n25193), .B1(n25183), .Y(
        n59) );
  sky130_fd_sc_hd__nand2_1 U29801 ( .A(n25193), .B(
        j202_soc_core_bldc_core_00_wdata[13]), .Y(n25185) );
  sky130_fd_sc_hd__o21ai_1 U29802 ( .A1(n25186), .A2(n25193), .B1(n25185), .Y(
        n61) );
  sky130_fd_sc_hd__a22o_1 U29803 ( .A1(n25193), .A2(
        j202_soc_core_bldc_core_00_wdata[14]), .B1(n25189), .B2(
        j202_soc_core_bldc_core_00_pwm_duty[2]), .X(n62) );
  sky130_fd_sc_hd__nand2_1 U29804 ( .A(n25193), .B(
        j202_soc_core_bldc_core_00_wdata[15]), .Y(n25187) );
  sky130_fd_sc_hd__o21ai_1 U29805 ( .A1(n25188), .A2(n25193), .B1(n25187), .Y(
        n63) );
  sky130_fd_sc_hd__a22o_1 U29806 ( .A1(n25189), .A2(
        j202_soc_core_bldc_core_00_pwm_duty[4]), .B1(n25193), .B2(
        j202_soc_core_bldc_core_00_wdata[16]), .X(n64) );
  sky130_fd_sc_hd__nand2_1 U29807 ( .A(n25193), .B(
        j202_soc_core_bldc_core_00_wdata[20]), .Y(n25190) );
  sky130_fd_sc_hd__o21ai_1 U29808 ( .A1(n25191), .A2(n25193), .B1(n25190), .Y(
        n66) );
  sky130_fd_sc_hd__nand2_1 U29809 ( .A(n25193), .B(
        j202_soc_core_bldc_core_00_wdata[22]), .Y(n25192) );
  sky130_fd_sc_hd__o22ai_1 U29811 ( .A1(n25228), .A2(n25196), .B1(n25227), 
        .B2(n25195), .Y(n78) );
  sky130_fd_sc_hd__a22o_1 U29812 ( .A1(n25213), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[0]), .B1(n25212), .B2(
        j202_soc_core_cmt_core_00_cks1[0]), .X(n82) );
  sky130_fd_sc_hd__o22ai_1 U29813 ( .A1(n25230), .A2(n25197), .B1(n25229), 
        .B2(n25198), .Y(n83) );
  sky130_fd_sc_hd__o22ai_1 U29814 ( .A1(n25228), .A2(n25199), .B1(n25227), 
        .B2(n25198), .Y(n84) );
  sky130_fd_sc_hd__a21o_1 U29815 ( .A1(n25200), .A2(
        j202_soc_core_uart_TOP_tx_fifo_wp[1]), .B1(
        j202_soc_core_uart_TOP_tx_fifo_N31), .X(n86) );
  sky130_fd_sc_hd__o21a_1 U29816 ( .A1(j202_soc_core_uart_TOP_tx_fifo_wp[0]), 
        .A2(n25201), .B1(n25200), .X(n87) );
  sky130_fd_sc_hd__nor2_1 U29817 ( .A(n25206), .B(n25205), .Y(n25204) );
  sky130_fd_sc_hd__o22ai_1 U29818 ( .A1(n25204), .A2(n25203), .B1(n25202), 
        .B2(n25205), .Y(n93) );
  sky130_fd_sc_hd__a21oi_1 U29819 ( .A1(n25206), .A2(n25205), .B1(n25204), .Y(
        n94) );
  sky130_fd_sc_hd__o22ai_1 U29820 ( .A1(n25230), .A2(n25208), .B1(n25229), 
        .B2(n25207), .Y(n97) );
  sky130_fd_sc_hd__o22ai_1 U29821 ( .A1(n25230), .A2(n25209), .B1(n25229), 
        .B2(n25210), .Y(n101) );
  sky130_fd_sc_hd__o22ai_1 U29822 ( .A1(n25228), .A2(n25211), .B1(n25227), 
        .B2(n25210), .Y(n102) );
  sky130_fd_sc_hd__a22o_1 U29823 ( .A1(n25213), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[6]), .B1(n25212), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr1[6]), .X(n103) );
  sky130_fd_sc_hd__o22ai_1 U29824 ( .A1(n25230), .A2(n25214), .B1(n25229), 
        .B2(n25215), .Y(n104) );
  sky130_fd_sc_hd__o22ai_1 U29825 ( .A1(n25228), .A2(n25216), .B1(n25227), 
        .B2(n25215), .Y(n105) );
  sky130_fd_sc_hd__o22ai_1 U29826 ( .A1(n25228), .A2(n25218), .B1(n25227), 
        .B2(n25217), .Y(n107) );
  sky130_fd_sc_hd__o22ai_1 U29827 ( .A1(n25230), .A2(n25219), .B1(n25229), 
        .B2(n25220), .Y(n114) );
  sky130_fd_sc_hd__o22ai_1 U29828 ( .A1(n25228), .A2(n25221), .B1(n25227), 
        .B2(n25220), .Y(n115) );
  sky130_fd_sc_hd__o22ai_1 U29829 ( .A1(n25230), .A2(n25222), .B1(n25229), 
        .B2(n25223), .Y(n116) );
  sky130_fd_sc_hd__o22ai_1 U29830 ( .A1(n25228), .A2(n25224), .B1(n25227), 
        .B2(n25223), .Y(n117) );
  sky130_fd_sc_hd__o22ai_1 U29831 ( .A1(n25228), .A2(n25226), .B1(n25227), 
        .B2(n25225), .Y(n119) );
  sky130_fd_sc_hd__a22o_1 U29832 ( .A1(n25228), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[11]), .B1(n25227), .B2(
        j202_soc_core_cmt_core_00_const1[11]), .X(n120) );
  sky130_fd_sc_hd__a22o_1 U29833 ( .A1(n25230), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[11]), .B1(n25229), .B2(
        j202_soc_core_cmt_core_00_const0[11]), .X(n126) );
  sky130_fd_sc_hd__a21oi_1 U29834 ( .A1(n25232), .A2(n25231), .B1(
        j202_soc_core_uart_TOP_rx_fifo_N29), .Y(n130) );
  sky130_fd_sc_hd__o21ai_1 U29835 ( .A1(n25235), .A2(n25234), .B1(n25233), .Y(
        n131) );
  sky130_fd_sc_hd__nand2_1 U29836 ( .A(n25405), .B(
        j202_soc_core_uart_TOP_change), .Y(n25238) );
  sky130_fd_sc_hd__nand2_1 U29838 ( .A(n25238), .B(n25237), .Y(n132) );
  sky130_fd_sc_hd__a22o_1 U29839 ( .A1(n25240), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[6]), .B1(n25239), .B2(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmcsr0[6]), .X(n134) );
  sky130_fd_sc_hd__nand2_1 U29840 ( .A(
        j202_soc_core_bldc_core_00_hall_value[0]), .B(n25241), .Y(n25242) );
  sky130_fd_sc_hd__nand2_1 U29841 ( .A(n25243), .B(n25242), .Y(n137) );
  sky130_fd_sc_hd__a22o_1 U29842 ( .A1(n25244), .A2(
        j202_soc_core_bldc_core_00_hall_value[2]), .B1(n25406), .B2(
        j202_soc_core_bldc_core_00_bldc_hall_00_hall_data_3[2]), .X(n138) );
  sky130_fd_sc_hd__nor2_2 U15633 ( .A(n19800), .B(n19799), .Y(n25340) );
  sky130_fd_sc_hd__a2bb2oi_1 U17633 ( .B1(j202_soc_core_j22_cpu_rf_tmp[9]), 
        .B2(n11184), .A1_N(n12539), .A2_N(n12538), .Y(n12541) );
  sky130_fd_sc_hd__a2bb2oi_1 U13437 ( .B1(j202_soc_core_j22_cpu_rf_tmp[11]), 
        .B2(n11184), .A1_N(n12539), .A2_N(n11890), .Y(n11892) );
  sky130_fd_sc_hd__nand2_1 U16428 ( .A(n23289), .B(n25732), .Y(n10536) );
  sky130_fd_sc_hd__buf_2 U13336 ( .A(n21253), .X(n11036) );
  sky130_fd_sc_hd__inv_2 U13313 ( .A(n21262), .Y(n10981) );
  sky130_fd_sc_hd__inv_2 U13314 ( .A(n21260), .Y(n10986) );
  sky130_fd_sc_hd__inv_2 U13293 ( .A(n10999), .Y(n10921) );
  sky130_fd_sc_hd__inv_2 U13294 ( .A(n11004), .Y(n10923) );
  sky130_fd_sc_hd__inv_2 U13295 ( .A(n11009), .Y(n10925) );
  sky130_fd_sc_hd__inv_2 U13296 ( .A(n11014), .Y(n10927) );
  sky130_fd_sc_hd__inv_2 U13297 ( .A(n11019), .Y(n10929) );
  sky130_fd_sc_hd__inv_2 U13298 ( .A(n11024), .Y(n10931) );
  sky130_fd_sc_hd__inv_2 U13299 ( .A(n11029), .Y(n10933) );
  sky130_fd_sc_hd__inv_2 U13300 ( .A(n11034), .Y(n10935) );
  sky130_fd_sc_hd__inv_2 U13301 ( .A(n10999), .Y(n10941) );
  sky130_fd_sc_hd__inv_2 U13302 ( .A(n11004), .Y(n10943) );
  sky130_fd_sc_hd__inv_2 U13303 ( .A(n11009), .Y(n10945) );
  sky130_fd_sc_hd__inv_2 U13304 ( .A(n11014), .Y(n10947) );
  sky130_fd_sc_hd__inv_2 U13305 ( .A(n11019), .Y(n10949) );
  sky130_fd_sc_hd__inv_2 U13306 ( .A(n11024), .Y(n10951) );
  sky130_fd_sc_hd__inv_2 U13307 ( .A(n11029), .Y(n10953) );
  sky130_fd_sc_hd__inv_2 U13308 ( .A(n11034), .Y(n10955) );
  sky130_fd_sc_hd__o2bb2ai_1 U13277 ( .B1(n22536), .B2(n21070), .A1_N(n21070), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N2830) );
  sky130_fd_sc_hd__o2bb2ai_1 U13488 ( .B1(n22536), .B2(n21103), .A1_N(n21103), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N2756) );
  sky130_fd_sc_hd__o2bb2ai_1 U13278 ( .B1(n22536), .B2(n21069), .A1_N(n21069), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N2978) );
  sky130_fd_sc_hd__o2bb2ai_1 U13604 ( .B1(n21189), .B2(n23338), .A1_N(n21189), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N3266) );
  sky130_fd_sc_hd__o2bb2ai_1 U13606 ( .B1(n21191), .B2(n23338), .A1_N(n21191), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N2711) );
  sky130_fd_sc_hd__o2bb2ai_1 U13603 ( .B1(n21203), .B2(n23338), .A1_N(n21203), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N2748) );
  sky130_fd_sc_hd__o2bb2ai_1 U13605 ( .B1(n21187), .B2(n23338), .A1_N(n21187), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N3229) );
  sky130_fd_sc_hd__o2bb2ai_1 U13609 ( .B1(n21185), .B2(n23338), .A1_N(n21185), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N2933) );
  sky130_fd_sc_hd__o2bb2ai_1 U13601 ( .B1(n21201), .B2(n23338), .A1_N(n21201), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N2896) );
  sky130_fd_sc_hd__o2bb2ai_1 U13602 ( .B1(n21183), .B2(n23338), .A1_N(n21183), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N2970) );
  sky130_fd_sc_hd__o2bb2ai_1 U13607 ( .B1(n21186), .B2(n23338), .A1_N(n21186), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N3192) );
  sky130_fd_sc_hd__o2bb2ai_1 U13608 ( .B1(n21069), .B2(n23338), .A1_N(n21069), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N3007) );
  sky130_fd_sc_hd__o2bb2ai_1 U13611 ( .B1(n21071), .B2(n23338), .A1_N(n21071), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N3155) );
  sky130_fd_sc_hd__o2bb2ai_1 U13624 ( .B1(n21189), .B2(n23335), .A1_N(n21189), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N3265) );
  sky130_fd_sc_hd__o2bb2ai_1 U13634 ( .B1(n21191), .B2(n23335), .A1_N(n21191), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N2710) );
  sky130_fd_sc_hd__o2bb2ai_1 U13622 ( .B1(n21203), .B2(n23335), .A1_N(n21203), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N2747) );
  sky130_fd_sc_hd__o2bb2ai_1 U13625 ( .B1(n21182), .B2(n23335), .A1_N(n21182), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N2821) );
  sky130_fd_sc_hd__o2bb2ai_1 U13627 ( .B1(n21206), .B2(n23335), .A1_N(n21206), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N3080) );
  sky130_fd_sc_hd__o2bb2ai_1 U13628 ( .B1(n21184), .B2(n23335), .A1_N(n21184), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N3117) );
  sky130_fd_sc_hd__o2bb2ai_1 U13631 ( .B1(n21187), .B2(n23335), .A1_N(n21187), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N3228) );
  sky130_fd_sc_hd__o2bb2ai_1 U13633 ( .B1(n21186), .B2(n23335), .A1_N(n21186), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N3191) );
  sky130_fd_sc_hd__o2bb2ai_1 U13637 ( .B1(n21185), .B2(n23335), .A1_N(n21185), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N2932) );
  sky130_fd_sc_hd__o2bb2ai_1 U13638 ( .B1(n21201), .B2(n23335), .A1_N(n21201), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N2895) );
  sky130_fd_sc_hd__o2bb2ai_1 U13623 ( .B1(n21199), .B2(n23335), .A1_N(n21199), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N3043) );
  sky130_fd_sc_hd__o2bb2ai_1 U13621 ( .B1(n21069), .B2(n23335), .A1_N(n21069), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N3006) );
  sky130_fd_sc_hd__o2bb2ai_1 U13630 ( .B1(n21071), .B2(n23335), .A1_N(n21071), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N3154) );
  sky130_fd_sc_hd__o2bb2ai_1 U13632 ( .B1(n21103), .B2(n23335), .A1_N(n21103), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N2784) );
  sky130_fd_sc_hd__o2bb2ai_1 U13635 ( .B1(n21070), .B2(n23335), .A1_N(n21070), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N2858) );
  sky130_fd_sc_hd__o2bb2ai_1 U13484 ( .B1(n22536), .B2(n21189), .A1_N(n21189), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N3237) );
  sky130_fd_sc_hd__o2bb2ai_1 U13286 ( .B1(n22536), .B2(n21191), .A1_N(n21191), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N2682) );
  sky130_fd_sc_hd__o2bb2ai_1 U13281 ( .B1(n22536), .B2(n21187), .A1_N(n21187), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N3200) );
  sky130_fd_sc_hd__o2bb2ai_1 U13282 ( .B1(n22536), .B2(n21184), .A1_N(n21184), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N3089) );
  sky130_fd_sc_hd__o2bb2ai_1 U13284 ( .B1(n22536), .B2(n21182), .A1_N(n21182), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N2793) );
  sky130_fd_sc_hd__o2bb2ai_1 U13285 ( .B1(n22536), .B2(n21183), .A1_N(n21183), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N2941) );
  sky130_fd_sc_hd__o2bb2ai_1 U13486 ( .B1(n22536), .B2(n21206), .A1_N(n21206), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N3052) );
  sky130_fd_sc_hd__o2bb2ai_1 U13487 ( .B1(n22536), .B2(n21199), .A1_N(n21199), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N3015) );
  sky130_fd_sc_hd__o2bb2ai_1 U13489 ( .B1(n22536), .B2(n21203), .A1_N(n21203), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N2719) );
  sky130_fd_sc_hd__o2bb2ai_1 U13283 ( .B1(n22536), .B2(n21185), .A1_N(n21185), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N2904) );
  sky130_fd_sc_hd__o2bb2ai_1 U13490 ( .B1(n22536), .B2(n21197), .A1_N(n21216), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N3314) );
  sky130_fd_sc_hd__o2bb2ai_1 U25041 ( .B1(n23335), .B2(n21197), .A1_N(n21216), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N3340) );
  sky130_fd_sc_hd__nor2_1 U13491 ( .A(n25248), .B(n21207), .Y(n25542) );
  sky130_fd_sc_hd__clkinv_4 U13279 ( .A(n10953), .Y(n10954) );
  sky130_fd_sc_hd__clkinv_4 U13280 ( .A(n10933), .Y(n10934) );
  sky130_fd_sc_hd__clkinv_4 U13309 ( .A(n10951), .Y(n10952) );
  sky130_fd_sc_hd__clkinv_4 U13310 ( .A(n10931), .Y(n10932) );
  sky130_fd_sc_hd__clkinv_4 U13311 ( .A(n10949), .Y(n10950) );
  sky130_fd_sc_hd__clkinv_4 U13337 ( .A(n10929), .Y(n10930) );
  sky130_fd_sc_hd__clkinv_4 U13338 ( .A(n10947), .Y(n10948) );
  sky130_fd_sc_hd__clkinv_4 U13344 ( .A(n10927), .Y(n10928) );
  sky130_fd_sc_hd__clkinv_4 U13345 ( .A(n10945), .Y(n10946) );
  sky130_fd_sc_hd__clkinv_4 U13347 ( .A(n10925), .Y(n10926) );
  sky130_fd_sc_hd__clkinv_4 U13349 ( .A(n10943), .Y(n10944) );
  sky130_fd_sc_hd__clkinv_4 U13351 ( .A(n10923), .Y(n10924) );
  sky130_fd_sc_hd__clkinv_4 U13353 ( .A(n10941), .Y(n10942) );
  sky130_fd_sc_hd__clkinv_4 U13355 ( .A(n10921), .Y(n10922) );
  sky130_fd_sc_hd__clkinv_2 U13357 ( .A(n10954), .Y(n25671) );
  sky130_fd_sc_hd__clkinv_2 U13359 ( .A(n10952), .Y(n25674) );
  sky130_fd_sc_hd__clkinv_2 U13365 ( .A(n10950), .Y(n25677) );
  sky130_fd_sc_hd__clkinv_2 U13366 ( .A(n10948), .Y(n25680) );
  sky130_fd_sc_hd__clkinv_2 U13367 ( .A(n10946), .Y(n25683) );
  sky130_fd_sc_hd__clkinv_2 U13368 ( .A(n10944), .Y(n25686) );
  sky130_fd_sc_hd__clkinv_2 U13369 ( .A(n10942), .Y(n25689) );
  sky130_fd_sc_hd__clkinv_2 U13370 ( .A(n10934), .Y(n25695) );
  sky130_fd_sc_hd__clkinv_2 U13371 ( .A(n10932), .Y(n25698) );
  sky130_fd_sc_hd__clkinv_2 U13372 ( .A(n10930), .Y(n25701) );
  sky130_fd_sc_hd__clkinv_2 U13373 ( .A(n10928), .Y(n25704) );
  sky130_fd_sc_hd__clkinv_2 U13374 ( .A(n10926), .Y(n25707) );
  sky130_fd_sc_hd__clkinv_2 U13375 ( .A(n10924), .Y(n25710) );
  sky130_fd_sc_hd__clkinv_2 U13376 ( .A(n10922), .Y(n25713) );
  sky130_fd_sc_hd__inv_2 U13377 ( .A(n25719), .Y(n25716) );
  sky130_fd_sc_hd__inv_2 U13378 ( .A(n10987), .Y(n25726) );
  sky130_fd_sc_hd__inv_2 U13379 ( .A(n10982), .Y(n25728) );
  sky130_fd_sc_hd__inv_4 U13380 ( .A(n11178), .Y(n10961) );
  sky130_fd_sc_hd__inv_1 U13384 ( .A(n10986), .Y(n10987) );
  sky130_fd_sc_hd__inv_1 U13385 ( .A(n10981), .Y(n10982) );
  sky130_fd_sc_hd__inv_6 U13386 ( .A(n11177), .Y(n10972) );
  sky130_fd_sc_hd__inv_4 U13387 ( .A(n21255), .Y(n10991) );
  sky130_fd_sc_hd__inv_2 U13389 ( .A(n11175), .Y(n11026) );
  sky130_fd_sc_hd__inv_2 U13394 ( .A(n11176), .Y(n11021) );
  sky130_fd_sc_hd__inv_2 U13399 ( .A(n11174), .Y(n11016) );
  sky130_fd_sc_hd__inv_2 U13400 ( .A(n11173), .Y(n11011) );
  sky130_fd_sc_hd__inv_2 U13401 ( .A(n11180), .Y(n11006) );
  sky130_fd_sc_hd__inv_2 U13402 ( .A(n11171), .Y(n11001) );
  sky130_fd_sc_hd__inv_2 U13403 ( .A(n11172), .Y(n10996) );
  sky130_fd_sc_hd__inv_2 U13404 ( .A(n11179), .Y(n11031) );
  sky130_fd_sc_hd__nor2_1 U13405 ( .A(n11530), .B(n11539), .Y(n20285) );
  sky130_fd_sc_hd__nor2_1 U13406 ( .A(n11522), .B(n11514), .Y(n20288) );
  sky130_fd_sc_hd__o21ai_0 U13407 ( .A1(n16327), .A2(n16159), .B1(n15496), .Y(
        n15497) );
  sky130_fd_sc_hd__o21ai_0 U13408 ( .A1(n15962), .A2(n16373), .B1(n15487), .Y(
        n15488) );
  sky130_fd_sc_hd__o21ai_0 U13409 ( .A1(n16373), .A2(n16168), .B1(n15372), .Y(
        n15373) );
  sky130_fd_sc_hd__o21ai_0 U13410 ( .A1(n16551), .A2(n16168), .B1(n15404), .Y(
        n15405) );
  sky130_fd_sc_hd__o21ai_0 U13411 ( .A1(n15420), .A2(n15419), .B1(n15418), .Y(
        n15421) );
  sky130_fd_sc_hd__o21ai_0 U13412 ( .A1(n16046), .A2(n16537), .B1(n15504), .Y(
        n15505) );
  sky130_fd_sc_hd__o21ai_0 U13413 ( .A1(n16551), .A2(n16159), .B1(n15468), .Y(
        n15469) );
  sky130_fd_sc_hd__o21ai_0 U13414 ( .A1(n16327), .A2(n16537), .B1(n16307), .Y(
        n16308) );
  sky130_fd_sc_hd__o21ai_0 U13415 ( .A1(n16046), .A2(n16584), .B1(n15358), .Y(
        n15359) );
  sky130_fd_sc_hd__o21ai_0 U13416 ( .A1(n16327), .A2(n16164), .B1(n15489), .Y(
        n15490) );
  sky130_fd_sc_hd__o21ai_0 U13417 ( .A1(n16265), .A2(n16168), .B1(n15607), .Y(
        n15608) );
  sky130_fd_sc_hd__o21ai_0 U13418 ( .A1(n11169), .A2(n15959), .B1(n15667), .Y(
        n15668) );
  sky130_fd_sc_hd__o21ai_0 U13419 ( .A1(n15962), .A2(n16227), .B1(n15722), .Y(
        n15723) );
  sky130_fd_sc_hd__o21ai_0 U13420 ( .A1(n16227), .A2(n16379), .B1(n15478), .Y(
        n15479) );
  sky130_fd_sc_hd__o21ai_0 U13421 ( .A1(n16052), .A2(n16537), .B1(n15324), .Y(
        n15325) );
  sky130_fd_sc_hd__o21ai_0 U13422 ( .A1(n15273), .A2(n15272), .B1(n15271), .Y(
        n15318) );
  sky130_fd_sc_hd__o21ai_0 U13423 ( .A1(n16052), .A2(n16367), .B1(n15552), .Y(
        n15553) );
  sky130_fd_sc_hd__o21ai_0 U13424 ( .A1(n16227), .A2(n16537), .B1(n16206), .Y(
        n16207) );
  sky130_fd_sc_hd__o21ai_0 U13425 ( .A1(n16551), .A2(n16193), .B1(n16192), .Y(
        n16194) );
  sky130_fd_sc_hd__o21ai_0 U13426 ( .A1(n16227), .A2(n16584), .B1(n16226), .Y(
        n16228) );
  sky130_fd_sc_hd__o21ai_0 U13427 ( .A1(n15335), .A2(n15434), .B1(n15334), .Y(
        n15336) );
  sky130_fd_sc_hd__o21ai_0 U13428 ( .A1(n16551), .A2(n16402), .B1(n16348), .Y(
        n16349) );
  sky130_fd_sc_hd__o21ai_0 U13429 ( .A1(n16373), .A2(n16557), .B1(n16291), .Y(
        n16292) );
  sky130_fd_sc_hd__o21ai_0 U13430 ( .A1(n16551), .A2(n16367), .B1(n16321), .Y(
        n16322) );
  sky130_fd_sc_hd__o21ai_0 U13436 ( .A1(n12995), .A2(n12994), .B1(n14567), .Y(
        n13058) );
  sky130_fd_sc_hd__o21ai_0 U13439 ( .A1(n16227), .A2(n16367), .B1(n15338), .Y(
        n15339) );
  sky130_fd_sc_hd__o21ai_0 U13441 ( .A1(n16265), .A2(n16367), .B1(n15443), .Y(
        n15444) );
  sky130_fd_sc_hd__o21ai_0 U13442 ( .A1(n16046), .A2(n16402), .B1(n15582), .Y(
        n15583) );
  sky130_fd_sc_hd__o21ai_0 U13449 ( .A1(n16227), .A2(n16278), .B1(n15605), .Y(
        n15606) );
  sky130_fd_sc_hd__o21ai_0 U13450 ( .A1(n16052), .A2(n16193), .B1(n15705), .Y(
        n15706) );
  sky130_fd_sc_hd__o21ai_0 U13460 ( .A1(n16067), .A2(n16354), .B1(n15735), .Y(
        n15736) );
  sky130_fd_sc_hd__o21ai_0 U13463 ( .A1(n16052), .A2(n16168), .B1(n15707), .Y(
        n15708) );
  sky130_fd_sc_hd__o21ai_0 U13467 ( .A1(n16046), .A2(n16193), .B1(n15797), .Y(
        n15798) );
  sky130_fd_sc_hd__o21ai_0 U13468 ( .A1(n19942), .A2(n16523), .B1(n16522), .Y(
        n16524) );
  sky130_fd_sc_hd__o21ai_0 U13471 ( .A1(n15425), .A2(n15434), .B1(n15424), .Y(
        n15426) );
  sky130_fd_sc_hd__o21ai_0 U13472 ( .A1(n15962), .A2(n16046), .B1(n15892), .Y(
        n15893) );
  sky130_fd_sc_hd__o21ai_0 U13474 ( .A1(n15361), .A2(n15365), .B1(n15362), .Y(
        n15302) );
  sky130_fd_sc_hd__o21ai_0 U13477 ( .A1(n16551), .A2(n16278), .B1(n16161), .Y(
        n16162) );
  sky130_fd_sc_hd__o21ai_0 U13478 ( .A1(n19336), .A2(n16193), .B1(n16171), .Y(
        n16172) );
  sky130_fd_sc_hd__o21ai_0 U13485 ( .A1(n11169), .A2(n16265), .B1(n16264), .Y(
        n16266) );
  sky130_fd_sc_hd__o21ai_0 U13564 ( .A1(n22580), .A2(n22492), .B1(n22491), .Y(
        n22493) );
  sky130_fd_sc_hd__o21ai_0 U13566 ( .A1(n20152), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[12]), .B1(n20151), .Y(n20153)
         );
  sky130_fd_sc_hd__o21ai_0 U13570 ( .A1(n13028), .A2(n13027), .B1(n14314), .Y(
        n13036) );
  sky130_fd_sc_hd__o21ai_0 U13596 ( .A1(n14201), .A2(n14235), .B1(n14723), .Y(
        n14208) );
  sky130_fd_sc_hd__o21ai_0 U13598 ( .A1(n14296), .A2(n14295), .B1(n14625), .Y(
        n14297) );
  sky130_fd_sc_hd__o21ai_0 U13610 ( .A1(n13596), .A2(n13245), .B1(n18170), .Y(
        n18017) );
  sky130_fd_sc_hd__o21ai_0 U13612 ( .A1(n16058), .A2(n16311), .B1(n15854), .Y(
        n15855) );
  sky130_fd_sc_hd__o21ai_0 U13614 ( .A1(n16046), .A2(n16168), .B1(n15851), .Y(
        n15852) );
  sky130_fd_sc_hd__o21ai_0 U13615 ( .A1(n16052), .A2(n16379), .B1(n15569), .Y(
        n15570) );
  sky130_fd_sc_hd__o21ai_0 U13616 ( .A1(n16067), .A2(n16557), .B1(n15659), .Y(
        n15660) );
  sky130_fd_sc_hd__o21ai_0 U13620 ( .A1(n16067), .A2(n16402), .B1(n16066), .Y(
        n16068) );
  sky130_fd_sc_hd__o21ai_0 U13677 ( .A1(n16067), .A2(n16379), .B1(n15739), .Y(
        n15740) );
  sky130_fd_sc_hd__o21ai_0 U13703 ( .A1(n16067), .A2(n16367), .B1(n15766), .Y(
        n15767) );
  sky130_fd_sc_hd__o21ai_0 U13708 ( .A1(n16058), .A2(n16305), .B1(n15908), .Y(
        n15909) );
  sky130_fd_sc_hd__o21ai_0 U13772 ( .A1(n16067), .A2(n16278), .B1(n15825), .Y(
        n15826) );
  sky130_fd_sc_hd__o21ai_0 U13993 ( .A1(n16058), .A2(n16354), .B1(n15807), .Y(
        n15808) );
  sky130_fd_sc_hd__o21ai_0 U14238 ( .A1(n19336), .A2(n16367), .B1(n16366), .Y(
        n16368) );
  sky130_fd_sc_hd__o21ai_0 U14393 ( .A1(n16058), .A2(n16278), .B1(n15890), .Y(
        n15891) );
  sky130_fd_sc_hd__o21ai_0 U14744 ( .A1(n16058), .A2(n16193), .B1(n15876), .Y(
        n15877) );
  sky130_fd_sc_hd__o21ai_0 U14755 ( .A1(n16327), .A2(n16402), .B1(n16153), .Y(
        n16154) );
  sky130_fd_sc_hd__o21ai_0 U14783 ( .A1(n16373), .A2(n16367), .B1(n16259), .Y(
        n16260) );
  sky130_fd_sc_hd__o21ai_0 U14800 ( .A1(n15962), .A2(n16067), .B1(n15914), .Y(
        n15915) );
  sky130_fd_sc_hd__o21ai_0 U14828 ( .A1(n21019), .A2(n21018), .B1(n21017), .Y(
        n21020) );
  sky130_fd_sc_hd__o21ai_0 U14829 ( .A1(n22517), .A2(n22516), .B1(n22530), .Y(
        n22518) );
  sky130_fd_sc_hd__o21ai_0 U14830 ( .A1(n14730), .A2(n14729), .B1(n14888), .Y(
        n14734) );
  sky130_fd_sc_hd__o21ai_0 U14831 ( .A1(n20155), .A2(n20172), .B1(n20154), .Y(
        n20158) );
  sky130_fd_sc_hd__o21ai_0 U14832 ( .A1(n14309), .A2(n14310), .B1(n14349), .Y(
        n14195) );
  sky130_fd_sc_hd__o21ai_0 U14833 ( .A1(n14605), .A2(n14604), .B1(n14603), .Y(
        n14606) );
  sky130_fd_sc_hd__o21ai_0 U14834 ( .A1(n14110), .A2(n14576), .B1(n14591), .Y(
        n14343) );
  sky130_fd_sc_hd__o21ai_0 U14835 ( .A1(n14103), .A2(n13017), .B1(n14350), .Y(
        n14325) );
  sky130_fd_sc_hd__o21ai_0 U14836 ( .A1(n13448), .A2(n13449), .B1(n13307), .Y(
        n13135) );
  sky130_fd_sc_hd__o21ai_0 U14837 ( .A1(n18084), .A2(n13258), .B1(n18189), .Y(
        n13259) );
  sky130_fd_sc_hd__o21ai_0 U14838 ( .A1(j202_soc_core_bootrom_00_address_w[4]), 
        .A2(n13236), .B1(n13235), .Y(n18113) );
  sky130_fd_sc_hd__o21ai_0 U14839 ( .A1(j202_soc_core_intc_core_00_rg_ipr[73]), 
        .A2(n24633), .B1(j202_soc_core_intc_core_00_rg_ipr[72]), .Y(n17353) );
  sky130_fd_sc_hd__o21ai_0 U14840 ( .A1(n19949), .A2(n16793), .B1(n16794), .Y(
        n16137) );
  sky130_fd_sc_hd__o21ai_0 U14841 ( .A1(n11169), .A2(n19336), .B1(n19335), .Y(
        n19337) );
  sky130_fd_sc_hd__o21ai_0 U14842 ( .A1(n21150), .A2(n22632), .B1(n21109), .Y(
        n21110) );
  sky130_fd_sc_hd__o21ai_0 U14843 ( .A1(n16527), .A2(n16621), .B1(n16526), .Y(
        n16528) );
  sky130_fd_sc_hd__o21ai_0 U14844 ( .A1(n19336), .A2(n16540), .B1(n16539), .Y(
        n16541) );
  sky130_fd_sc_hd__o21ai_0 U14845 ( .A1(n15959), .A2(n16319), .B1(n15883), .Y(
        n15884) );
  sky130_fd_sc_hd__o21ai_0 U14846 ( .A1(n15962), .A2(n16058), .B1(n15961), .Y(
        n15963) );
  sky130_fd_sc_hd__o21ai_0 U14847 ( .A1(n16058), .A2(n16164), .B1(n15931), .Y(
        n15932) );
  sky130_fd_sc_hd__o21ai_0 U14848 ( .A1(n21150), .A2(n22619), .B1(n19257), .Y(
        n19258) );
  sky130_fd_sc_hd__o21ai_0 U14849 ( .A1(n18874), .A2(n17076), .B1(n17077), .Y(
        n16618) );
  sky130_fd_sc_hd__o21ai_0 U14850 ( .A1(j202_soc_core_intc_core_00_rg_ipr[24]), 
        .A2(n21356), .B1(n17278), .Y(n17290) );
  sky130_fd_sc_hd__o21ai_0 U14851 ( .A1(n11202), .A2(n21154), .B1(n22176), .Y(
        n21012) );
  sky130_fd_sc_hd__o21ai_0 U14852 ( .A1(n13491), .A2(n13490), .B1(n13489), .Y(
        n13499) );
  sky130_fd_sc_hd__o21ai_0 U14853 ( .A1(n13315), .A2(n11281), .B1(n13121), .Y(
        n11282) );
  sky130_fd_sc_hd__o21ai_0 U14854 ( .A1(n14710), .A2(n14815), .B1(n14709), .Y(
        n14714) );
  sky130_fd_sc_hd__o21ai_0 U14855 ( .A1(n20187), .A2(
        j202_soc_core_wbqspiflash_00_w_spif_addr[13]), .B1(n20186), .Y(n20188)
         );
  sky130_fd_sc_hd__o21ai_0 U14856 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[5]), .A2(n20144), .B1(n20163), 
        .Y(n20145) );
  sky130_fd_sc_hd__o21ai_0 U14857 ( .A1(n14843), .A2(n14842), .B1(n14841), .Y(
        n14844) );
  sky130_fd_sc_hd__o21ai_0 U14858 ( .A1(n14980), .A2(n14098), .B1(n14549), .Y(
        n14186) );
  sky130_fd_sc_hd__o21ai_0 U14859 ( .A1(n14585), .A2(n14584), .B1(n14613), .Y(
        n14586) );
  sky130_fd_sc_hd__o21ai_0 U14860 ( .A1(n14354), .A2(n14353), .B1(n14352), .Y(
        n14360) );
  sky130_fd_sc_hd__o21ai_0 U14861 ( .A1(n14413), .A2(n13171), .B1(n13170), .Y(
        n13378) );
  sky130_fd_sc_hd__o21ai_0 U14862 ( .A1(n13260), .A2(n18183), .B1(n13259), .Y(
        n13261) );
  sky130_fd_sc_hd__o21ai_0 U14863 ( .A1(n18163), .A2(n18162), .B1(n18161), .Y(
        n18165) );
  sky130_fd_sc_hd__o21ai_0 U14864 ( .A1(n18106), .A2(n18105), .B1(n18161), .Y(
        n18108) );
  sky130_fd_sc_hd__o21ai_0 U14865 ( .A1(n17382), .A2(n17384), .B1(n17379), .Y(
        n17365) );
  sky130_fd_sc_hd__o21ai_0 U14866 ( .A1(j202_soc_core_intc_core_00_rg_ipr[26]), 
        .A2(n21356), .B1(n17274), .Y(n17287) );
  sky130_fd_sc_hd__o21ai_0 U14867 ( .A1(n19668), .A2(n19665), .B1(n19669), .Y(
        n19918) );
  sky130_fd_sc_hd__o21ai_0 U14868 ( .A1(n16150), .A2(n17030), .B1(n16149), .Y(
        n16151) );
  sky130_fd_sc_hd__o21ai_0 U14869 ( .A1(n19132), .A2(n19002), .B1(n19003), .Y(
        n16125) );
  sky130_fd_sc_hd__o21ai_0 U14870 ( .A1(n19623), .A2(n19339), .B1(n19338), .Y(
        n19344) );
  sky130_fd_sc_hd__o21ai_0 U14871 ( .A1(n18967), .A2(n18964), .B1(n18968), .Y(
        n19351) );
  sky130_fd_sc_hd__o21ai_0 U14872 ( .A1(n18860), .A2(n17034), .B1(n17035), .Y(
        n18973) );
  sky130_fd_sc_hd__o21ai_0 U14873 ( .A1(n19290), .A2(n19287), .B1(n19288), .Y(
        n16783) );
  sky130_fd_sc_hd__o21ai_0 U14874 ( .A1(n15959), .A2(n16159), .B1(n15958), .Y(
        n15960) );
  sky130_fd_sc_hd__o21ai_0 U14875 ( .A1(n15238), .A2(n15237), .B1(n15236), .Y(
        n15240) );
  sky130_fd_sc_hd__o21ai_0 U14876 ( .A1(n21150), .A2(n22649), .B1(n19154), .Y(
        n19155) );
  sky130_fd_sc_hd__clkinv_1 U14877 ( .A(n12970), .Y(n12975) );
  sky130_fd_sc_hd__o21ai_0 U14878 ( .A1(n21108), .A2(n22595), .B1(n21021), .Y(
        n21022) );
  sky130_fd_sc_hd__o21ai_0 U14879 ( .A1(n24370), .A2(n21348), .B1(n17159), .Y(
        n17206) );
  sky130_fd_sc_hd__o21ai_0 U14880 ( .A1(n11283), .A2(n13464), .B1(n11282), .Y(
        n11284) );
  sky130_fd_sc_hd__o21ai_0 U14881 ( .A1(n13449), .A2(n11363), .B1(n13170), .Y(
        n13421) );
  sky130_fd_sc_hd__o21ai_0 U14882 ( .A1(n24385), .A2(n21355), .B1(n17267), .Y(
        n17289) );
  sky130_fd_sc_hd__o21ai_0 U14883 ( .A1(n22692), .A2(n22511), .B1(n22499), .Y(
        n22500) );
  sky130_fd_sc_hd__o21ai_0 U14884 ( .A1(n14744), .A2(n14743), .B1(n18610), .Y(
        n14763) );
  sky130_fd_sc_hd__o21ai_0 U14885 ( .A1(n23405), .A2(n25066), .B1(n23430), .Y(
        n23406) );
  sky130_fd_sc_hd__o21ai_0 U14886 ( .A1(n14575), .A2(n14412), .B1(n14678), .Y(
        n14835) );
  sky130_fd_sc_hd__o21ai_0 U14887 ( .A1(n14845), .A2(n14882), .B1(n14844), .Y(
        n14846) );
  sky130_fd_sc_hd__o21ai_0 U14888 ( .A1(n14621), .A2(n14639), .B1(n14220), .Y(
        n14221) );
  sky130_fd_sc_hd__o21ai_0 U14889 ( .A1(n14587), .A2(n14631), .B1(n14586), .Y(
        n14588) );
  sky130_fd_sc_hd__clkinv_1 U14890 ( .A(j202_soc_core_memory0_ram_dout0_sel[4]), .Y(n11317) );
  sky130_fd_sc_hd__o21ai_0 U14891 ( .A1(j202_soc_core_intc_core_00_rg_ipr[7]), 
        .A2(n21358), .B1(n17242), .Y(n17255) );
  sky130_fd_sc_hd__o21ai_0 U14892 ( .A1(j202_soc_core_intc_core_00_rg_ipr[27]), 
        .A2(n21356), .B1(n17281), .Y(n17306) );
  sky130_fd_sc_hd__o21ai_0 U14893 ( .A1(j202_soc_core_intc_core_00_rg_ipr[47]), 
        .A2(n21346), .B1(n17184), .Y(n17197) );
  sky130_fd_sc_hd__o21ai_0 U14894 ( .A1(n19040), .A2(n19073), .B1(n19041), .Y(
        n12358) );
  sky130_fd_sc_hd__o21ai_0 U14895 ( .A1(n18299), .A2(n18298), .B1(n18655), .Y(
        n18300) );
  sky130_fd_sc_hd__o21ai_0 U14896 ( .A1(n21091), .A2(n23315), .B1(n20868), .Y(
        n20869) );
  sky130_fd_sc_hd__o21ai_0 U14897 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[3]), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[7]), .B1(
        j202_soc_core_cmt_core_00_cks0[0]), .Y(n20460) );
  sky130_fd_sc_hd__o21ai_0 U14898 ( .A1(n19507), .A2(n19511), .B1(n19512), .Y(
        n12613) );
  sky130_fd_sc_hd__o21ai_0 U14899 ( .A1(n14089), .A2(n22351), .B1(n12412), .Y(
        n12616) );
  sky130_fd_sc_hd__o21ai_0 U14900 ( .A1(n17031), .A2(n19299), .B1(n17030), .Y(
        n18859) );
  sky130_fd_sc_hd__o21ai_0 U14901 ( .A1(n21091), .A2(n23312), .B1(n20419), .Y(
        n20420) );
  sky130_fd_sc_hd__o21ai_0 U14902 ( .A1(n14089), .A2(n21929), .B1(n12493), .Y(
        n12608) );
  sky130_fd_sc_hd__o21ai_0 U14903 ( .A1(n19292), .A2(n19291), .B1(n19290), .Y(
        n19293) );
  sky130_fd_sc_hd__o21ai_0 U14904 ( .A1(n19856), .A2(n16829), .B1(n16830), .Y(
        n16037) );
  sky130_fd_sc_hd__o21ai_0 U14905 ( .A1(n19362), .A2(n19361), .B1(n19360), .Y(
        n20028) );
  sky130_fd_sc_hd__o21ai_0 U14906 ( .A1(n16032), .A2(n16605), .B1(n16031), .Y(
        n16832) );
  sky130_fd_sc_hd__o21ai_0 U14907 ( .A1(n19108), .A2(n18986), .B1(n18987), .Y(
        n16024) );
  sky130_fd_sc_hd__o21ai_0 U14908 ( .A1(n14089), .A2(n21807), .B1(n12576), .Y(
        n12612) );
  sky130_fd_sc_hd__o21ai_0 U14909 ( .A1(n20908), .A2(n20935), .B1(n21010), .Y(
        n20728) );
  sky130_fd_sc_hd__o21ai_0 U14910 ( .A1(n20908), .A2(n20720), .B1(n21010), .Y(
        n20630) );
  sky130_fd_sc_hd__o21ai_0 U14911 ( .A1(n21091), .A2(n23332), .B1(n20963), .Y(
        n20964) );
  sky130_fd_sc_hd__o21ai_0 U14912 ( .A1(n16531), .A2(n16615), .B1(n16530), .Y(
        n19359) );
  sky130_fd_sc_hd__o21ai_0 U14913 ( .A1(n16790), .A2(n19299), .B1(n16789), .Y(
        n19951) );
  sky130_fd_sc_hd__o21ai_0 U14914 ( .A1(n19941), .A2(n19945), .B1(n19942), .Y(
        n18854) );
  sky130_fd_sc_hd__o21ai_0 U14915 ( .A1(n18999), .A2(n18998), .B1(n19127), .Y(
        n19000) );
  sky130_fd_sc_hd__o21ai_0 U14916 ( .A1(n21091), .A2(n23326), .B1(n21090), .Y(
        n21092) );
  sky130_fd_sc_hd__o21ai_0 U14917 ( .A1(n14089), .A2(n22609), .B1(n14036), .Y(
        n14038) );
  sky130_fd_sc_hd__o21ai_0 U14918 ( .A1(n20931), .A2(n22496), .B1(n21141), .Y(
        n16656) );
  sky130_fd_sc_hd__o21ai_0 U14919 ( .A1(n25377), .A2(n19484), .B1(n22387), .Y(
        n19485) );
  sky130_fd_sc_hd__o21ai_0 U14920 ( .A1(n19850), .A2(n19854), .B1(n19851), .Y(
        n16827) );
  sky130_fd_sc_hd__o21ai_0 U14921 ( .A1(n19419), .A2(n19423), .B1(n19420), .Y(
        n19391) );
  sky130_fd_sc_hd__o21ai_0 U14922 ( .A1(n19523), .A2(n19527), .B1(n19524), .Y(
        n19553) );
  sky130_fd_sc_hd__o21ai_0 U14923 ( .A1(n14089), .A2(n22064), .B1(n11950), .Y(
        n12620) );
  sky130_fd_sc_hd__o21ai_0 U14924 ( .A1(n14089), .A2(n22074), .B1(n13868), .Y(
        n14041) );
  sky130_fd_sc_hd__o21ai_0 U14925 ( .A1(n14089), .A2(n22602), .B1(n13964), .Y(
        n14001) );
  sky130_fd_sc_hd__o21ai_0 U14926 ( .A1(j202_soc_core_intc_core_00_rg_ipr[76]), 
        .A2(n21369), .B1(n17364), .Y(n17379) );
  sky130_fd_sc_hd__o21ai_0 U14927 ( .A1(n14089), .A2(n22646), .B1(n12349), .Y(
        n12353) );
  sky130_fd_sc_hd__o21ai_0 U14928 ( .A1(j202_soc_core_intc_core_00_rg_ipr[53]), 
        .A2(n21349), .B1(n17158), .Y(n17208) );
  sky130_fd_sc_hd__o21ai_0 U14929 ( .A1(n13485), .A2(n13484), .B1(n13483), .Y(
        n13506) );
  sky130_fd_sc_hd__clkinv_1 U14930 ( .A(
        j202_soc_core_memory0_ram_dout0_sel[11]), .Y(n11296) );
  sky130_fd_sc_hd__o21ai_0 U14931 ( .A1(n18527), .A2(n15181), .B1(n18513), .Y(
        n16918) );
  sky130_fd_sc_hd__o21ai_0 U14932 ( .A1(n13468), .A2(n11219), .B1(n13121), .Y(
        n11220) );
  sky130_fd_sc_hd__o21ai_0 U14933 ( .A1(n14089), .A2(n22037), .B1(n12265), .Y(
        n12355) );
  sky130_fd_sc_hd__o21ai_0 U14934 ( .A1(j202_soc_core_intc_core_00_rg_ipr[54]), 
        .A2(n21349), .B1(n17155), .Y(n17202) );
  sky130_fd_sc_hd__clkinv_1 U14935 ( .A(n16861), .Y(n16647) );
  sky130_fd_sc_hd__o21ai_0 U14936 ( .A1(n19724), .A2(n19721), .B1(n19722), .Y(
        n18941) );
  sky130_fd_sc_hd__o21ai_0 U14937 ( .A1(n14089), .A2(n21862), .B1(n11875), .Y(
        n12653) );
  sky130_fd_sc_hd__o21ai_0 U14938 ( .A1(n14497), .A2(n14496), .B1(n14888), .Y(
        n14498) );
  sky130_fd_sc_hd__o21ai_0 U14939 ( .A1(n14721), .A2(n14424), .B1(n14866), .Y(
        n14425) );
  sky130_fd_sc_hd__o21ai_0 U14940 ( .A1(n14089), .A2(n22599), .B1(n12784), .Y(
        n12786) );
  sky130_fd_sc_hd__clkinv_1 U14941 ( .A(n25250), .Y(n18503) );
  sky130_fd_sc_hd__o21ai_0 U14942 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[2]), .A2(
        j202_soc_core_wbqspiflash_00_spif_data[31]), .B1(n24903), .Y(n23402)
         );
  sky130_fd_sc_hd__o21ai_0 U14943 ( .A1(n20138), .A2(n20208), .B1(n20207), .Y(
        n20136) );
  sky130_fd_sc_hd__o21ai_0 U14944 ( .A1(n14089), .A2(n21787), .B1(n11723), .Y(
        n12721) );
  sky130_fd_sc_hd__o21ai_0 U14945 ( .A1(n14485), .A2(n14143), .B1(n14888), .Y(
        n14689) );
  sky130_fd_sc_hd__o21ai_0 U14946 ( .A1(n13123), .A2(n13122), .B1(n13121), .Y(
        n13132) );
  sky130_fd_sc_hd__o21ai_0 U14947 ( .A1(j202_soc_core_memory0_ram_dout0[496]), 
        .A2(n18758), .B1(n18071), .Y(n18072) );
  sky130_fd_sc_hd__clkinv_1 U14948 ( .A(j202_soc_core_aquc_CE__1_), .Y(n11244)
         );
  sky130_fd_sc_hd__o21ai_0 U14949 ( .A1(n18643), .A2(n18294), .B1(n18513), .Y(
        n15154) );
  sky130_fd_sc_hd__o21ai_0 U14950 ( .A1(j202_soc_core_intc_core_00_rg_ipr[55]), 
        .A2(n21349), .B1(n17154), .Y(n17166) );
  sky130_fd_sc_hd__o21ai_0 U14952 ( .A1(n24357), .A2(n21345), .B1(n17176), .Y(
        n17199) );
  sky130_fd_sc_hd__o21ai_0 U15070 ( .A1(j202_soc_core_intc_core_00_rg_ipr[11]), 
        .A2(n21357), .B1(n17234), .Y(n17257) );
  sky130_fd_sc_hd__o21ai_0 U15079 ( .A1(n17308), .A2(n17282), .B1(n17306), .Y(
        n17285) );
  sky130_fd_sc_hd__o21ai_0 U15303 ( .A1(n14089), .A2(n22640), .B1(n11646), .Y(
        n12755) );
  sky130_fd_sc_hd__o21ai_0 U15557 ( .A1(n14089), .A2(n22644), .B1(n12523), .Y(
        n12606) );
  sky130_fd_sc_hd__o21ai_0 U15575 ( .A1(n12124), .A2(n19243), .B1(n19244), .Y(
        n15076) );
  sky130_fd_sc_hd__o21ai_0 U15785 ( .A1(n19053), .A2(n14077), .B1(n12203), .Y(
        n12206) );
  sky130_fd_sc_hd__o21ai_0 U15818 ( .A1(n20461), .A2(
        j202_soc_core_cmt_core_00_cks0[0]), .B1(n20460), .Y(n20462) );
  sky130_fd_sc_hd__o21ai_0 U15823 ( .A1(n19838), .A2(n14077), .B1(n12021), .Y(
        n12024) );
  sky130_fd_sc_hd__o21ai_0 U15824 ( .A1(n18837), .A2(n18840), .B1(n18838), .Y(
        n12617) );
  sky130_fd_sc_hd__o21ai_0 U15826 ( .A1(n22641), .A2(n23312), .B1(n21139), .Y(
        n20408) );
  sky130_fd_sc_hd__o21ai_0 U15879 ( .A1(n19202), .A2(n14077), .B1(n12486), .Y(
        n12489) );
  sky130_fd_sc_hd__o21ai_0 U15926 ( .A1(n23495), .A2(
        j202_soc_core_qspi_wb_addr[24]), .B1(n23494), .Y(n23496) );
  sky130_fd_sc_hd__o21ai_0 U15978 ( .A1(n17082), .A2(n16128), .B1(n16127), .Y(
        n16625) );
  sky130_fd_sc_hd__o21ai_0 U16073 ( .A1(n18878), .A2(n17085), .B1(n17086), .Y(
        n19005) );
  sky130_fd_sc_hd__o21ai_0 U16084 ( .A1(n20908), .A2(n21152), .B1(n21010), .Y(
        n20585) );
  sky130_fd_sc_hd__o21ai_0 U16178 ( .A1(n22610), .A2(n23332), .B1(n21139), .Y(
        n20954) );
  sky130_fd_sc_hd__o21ai_0 U16181 ( .A1(n16693), .A2(n14077), .B1(n12516), .Y(
        n12519) );
  sky130_fd_sc_hd__o21ai_0 U16182 ( .A1(n19181), .A2(n14077), .B1(n12258), .Y(
        n12261) );
  sky130_fd_sc_hd__o21ai_0 U16277 ( .A1(n17065), .A2(n14077), .B1(n12342), .Y(
        n12345) );
  sky130_fd_sc_hd__o21ai_0 U16300 ( .A1(n17042), .A2(n16019), .B1(n16018), .Y(
        n18989) );
  sky130_fd_sc_hd__o21ai_0 U16307 ( .A1(n19310), .A2(n19307), .B1(n19308), .Y(
        n16805) );
  sky130_fd_sc_hd__o21ai_0 U16540 ( .A1(n15962), .A2(n15959), .B1(n15943), .Y(
        n19232) );
  sky130_fd_sc_hd__o21ai_0 U16547 ( .A1(n22757), .A2(n22141), .B1(n19899), .Y(
        n19900) );
  sky130_fd_sc_hd__o21ai_0 U16561 ( .A1(n22606), .A2(n23326), .B1(n21139), .Y(
        n21080) );
  sky130_fd_sc_hd__o21ai_0 U16564 ( .A1(n19274), .A2(n14077), .B1(n12105), .Y(
        n12107) );
  sky130_fd_sc_hd__o21ai_0 U16688 ( .A1(n20908), .A2(n20530), .B1(n21010), .Y(
        n19037) );
  sky130_fd_sc_hd__o21ai_0 U16770 ( .A1(n21420), .A2(n21574), .B1(n20328), .Y(
        n19477) );
  sky130_fd_sc_hd__o21ai_0 U16933 ( .A1(n21573), .A2(n20743), .B1(n22388), .Y(
        n20765) );
  sky130_fd_sc_hd__o21ai_0 U17011 ( .A1(n12937), .A2(n12976), .B1(n12936), .Y(
        n12939) );
  sky130_fd_sc_hd__o21ai_0 U17087 ( .A1(n22387), .A2(n22739), .B1(n21333), .Y(
        n21334) );
  sky130_fd_sc_hd__o21ai_0 U17178 ( .A1(n21027), .A2(n22013), .B1(n20905), .Y(
        n18908) );
  sky130_fd_sc_hd__o21ai_0 U17191 ( .A1(n21091), .A2(n23342), .B1(n21047), .Y(
        n21060) );
  sky130_fd_sc_hd__o21ai_0 U17273 ( .A1(n17303), .A2(n21375), .B1(n17302), .Y(
        n17329) );
  sky130_fd_sc_hd__o21ai_0 U17332 ( .A1(n21027), .A2(n22591), .B1(n21010), .Y(
        n21026) );
  sky130_fd_sc_hd__clkinv_1 U17337 ( .A(n19893), .Y(n19148) );
  sky130_fd_sc_hd__o21ai_0 U17423 ( .A1(n11354), .A2(n14989), .B1(n11353), .Y(
        n11361) );
  sky130_fd_sc_hd__o21ai_0 U17428 ( .A1(n17833), .A2(n17125), .B1(n17126), .Y(
        n19043) );
  sky130_fd_sc_hd__o21ai_0 U17434 ( .A1(n24562), .A2(n21368), .B1(n17360), .Y(
        n17377) );
  sky130_fd_sc_hd__o21ai_0 U17437 ( .A1(n17205), .A2(n21379), .B1(n17204), .Y(
        n17321) );
  sky130_fd_sc_hd__o21ai_0 U17493 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[7]), .A2(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[3]), .B1(
        j202_soc_core_cmt_core_00_cks1[0]), .Y(n23105) );
  sky130_fd_sc_hd__o21ai_0 U17572 ( .A1(n22700), .A2(n22699), .B1(n22698), .Y(
        n22701) );
  sky130_fd_sc_hd__o21ai_0 U17577 ( .A1(n22509), .A2(n22508), .B1(n22507), .Y(
        n22667) );
  sky130_fd_sc_hd__o21ai_0 U17606 ( .A1(n14882), .A2(n14441), .B1(n14440), .Y(
        n14442) );
  sky130_fd_sc_hd__o21ai_0 U17611 ( .A1(n22733), .A2(n21485), .B1(n20745), .Y(
        n20984) );
  sky130_fd_sc_hd__o21ai_0 U17668 ( .A1(n20212), .A2(n20211), .B1(n20210), .Y(
        n20213) );
  sky130_fd_sc_hd__o21ai_0 U17708 ( .A1(n23540), .A2(n25107), .B1(n23539), .Y(
        n23545) );
  sky130_fd_sc_hd__o21ai_0 U17711 ( .A1(n25108), .A2(
        j202_soc_core_wbqspiflash_00_spi_valid), .B1(n25107), .Y(n25110) );
  sky130_fd_sc_hd__o21ai_0 U17714 ( .A1(j202_soc_core_memory0_ram_dout0[511]), 
        .A2(n18758), .B1(n14137), .Y(n14140) );
  sky130_fd_sc_hd__o21ai_0 U17785 ( .A1(n14366), .A2(n14617), .B1(n14365), .Y(
        n14367) );
  sky130_fd_sc_hd__o21ai_0 U17821 ( .A1(n16741), .A2(n16740), .B1(n16739), .Y(
        n16750) );
  sky130_fd_sc_hd__o21ai_0 U17891 ( .A1(n15155), .A2(n18779), .B1(n15154), .Y(
        n16891) );
  sky130_fd_sc_hd__o21ai_0 U18063 ( .A1(n24372), .A2(n21348), .B1(n17148), .Y(
        n17168) );
  sky130_fd_sc_hd__o21ai_0 U18092 ( .A1(n17199), .A2(n21379), .B1(n17198), .Y(
        n17226) );
  sky130_fd_sc_hd__o21ai_0 U18150 ( .A1(n17257), .A2(n21375), .B1(n17256), .Y(
        n17316) );
  sky130_fd_sc_hd__o21ai_0 U18184 ( .A1(n17196), .A2(n17195), .B1(n17194), .Y(
        n21379) );
  sky130_fd_sc_hd__clkinv_1 U18223 ( .A(n25281), .Y(n18504) );
  sky130_fd_sc_hd__o21ai_0 U18255 ( .A1(n21574), .A2(n21410), .B1(n21523), .Y(
        n20738) );
  sky130_fd_sc_hd__clkinv_1 U18267 ( .A(j202_soc_core_j22_cpu_memop_Ma__1_), 
        .Y(n13092) );
  sky130_fd_sc_hd__o21ai_0 U18273 ( .A1(n24869), .A2(n24883), .B1(n24868), .Y(
        n24870) );
  sky130_fd_sc_hd__clkinv_1 U18278 ( .A(n22704), .Y(n22644) );
  sky130_fd_sc_hd__o21ai_0 U18349 ( .A1(
        j202_soc_core_ahblite_interconnect_s_hrdata[6]), .A2(n18288), .B1(
        n18287), .Y(n18307) );
  sky130_fd_sc_hd__o21ai_0 U18374 ( .A1(n22351), .A2(n19083), .B1(n18845), .Y(
        n18846) );
  sky130_fd_sc_hd__o21ai_0 U18414 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[27]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[27]), .B1(n24034), 
        .Y(n24035) );
  sky130_fd_sc_hd__o21ai_0 U18488 ( .A1(n18841), .A2(n19725), .B1(n18840), .Y(
        n18842) );
  sky130_fd_sc_hd__o21ai_0 U18547 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[23]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[23]), .B1(n24008), 
        .Y(n24009) );
  sky130_fd_sc_hd__o21ai_0 U18583 ( .A1(n19107), .A2(n19111), .B1(n19108), .Y(
        n18990) );
  sky130_fd_sc_hd__o21ai_0 U18584 ( .A1(n19726), .A2(n19725), .B1(n19724), .Y(
        n19727) );
  sky130_fd_sc_hd__o21ai_0 U18611 ( .A1(n20931), .A2(n20943), .B1(n21141), .Y(
        n20948) );
  sky130_fd_sc_hd__o21ai_0 U18689 ( .A1(n25093), .A2(n25042), .B1(n23481), .Y(
        n23482) );
  sky130_fd_sc_hd__o21ai_0 U18727 ( .A1(n19131), .A2(n19135), .B1(n19132), .Y(
        n19008) );
  sky130_fd_sc_hd__o21ai_0 U18731 ( .A1(n19855), .A2(n19859), .B1(n19856), .Y(
        n16833) );
  sky130_fd_sc_hd__o21ai_0 U18766 ( .A1(n19954), .A2(n19957), .B1(n19955), .Y(
        n16806) );
  sky130_fd_sc_hd__o21ai_0 U18842 ( .A1(n20793), .A2(n23309), .B1(n20792), .Y(
        n20794) );
  sky130_fd_sc_hd__o21ai_0 U19018 ( .A1(n19097), .A2(n19096), .B1(n19095), .Y(
        n19098) );
  sky130_fd_sc_hd__o21ai_0 U19097 ( .A1(n19012), .A2(n19015), .B1(n19013), .Y(
        n16635) );
  sky130_fd_sc_hd__o21ai_0 U19177 ( .A1(n17097), .A2(n17094), .B1(n17095), .Y(
        n19143) );
  sky130_fd_sc_hd__o21ai_0 U19249 ( .A1(n19864), .A2(n19867), .B1(n19865), .Y(
        n16841) );
  sky130_fd_sc_hd__o21ai_0 U19386 ( .A1(n22565), .A2(n21017), .B1(n19900), .Y(
        n19901) );
  sky130_fd_sc_hd__o21ai_0 U19394 ( .A1(n25387), .A2(n20993), .B1(n22740), .Y(
        n21598) );
  sky130_fd_sc_hd__o21ai_0 U19414 ( .A1(n21027), .A2(n22547), .B1(n20905), .Y(
        n16871) );
  sky130_fd_sc_hd__o21ai_0 U19460 ( .A1(n20908), .A2(n22484), .B1(n17121), .Y(
        n17130) );
  sky130_fd_sc_hd__or2_0 U19513 ( .A(n22384), .B(n25372), .X(n22409) );
  sky130_fd_sc_hd__o21ai_0 U19539 ( .A1(n22385), .A2(n21455), .B1(n20750), .Y(
        n19323) );
  sky130_fd_sc_hd__o21ai_0 U19543 ( .A1(n22389), .A2(n24866), .B1(n22388), .Y(
        n22392) );
  sky130_fd_sc_hd__o21ai_0 U19606 ( .A1(n21382), .A2(n21381), .B1(n21380), .Y(
        n21383) );
  sky130_fd_sc_hd__o21ai_0 U19617 ( .A1(n20850), .A2(n23329), .B1(n20849), .Y(
        n20851) );
  sky130_fd_sc_hd__o21ai_0 U19651 ( .A1(n17381), .A2(n21387), .B1(n17380), .Y(
        n17398) );
  sky130_fd_sc_hd__o21ai_0 U19702 ( .A1(n17214), .A2(n21382), .B1(n17213), .Y(
        n17326) );
  sky130_fd_sc_hd__o21ai_0 U19703 ( .A1(n17384), .A2(n21387), .B1(n17383), .Y(
        n17406) );
  sky130_fd_sc_hd__o21ai_0 U19708 ( .A1(n18525), .A2(n15197), .B1(n18655), .Y(
        n11350) );
  sky130_fd_sc_hd__o21ai_0 U19765 ( .A1(n16896), .A2(n16895), .B1(n18664), .Y(
        n18302) );
  sky130_fd_sc_hd__o21ai_0 U19772 ( .A1(n18481), .A2(n18485), .B1(n18482), .Y(
        n18494) );
  sky130_fd_sc_hd__clkinv_1 U19777 ( .A(n20309), .Y(n20271) );
  sky130_fd_sc_hd__o21ai_0 U19836 ( .A1(j202_soc_core_memory0_ram_dout0[489]), 
        .A2(n18758), .B1(n18376), .Y(n18377) );
  sky130_fd_sc_hd__o21ai_0 U19837 ( .A1(n18761), .A2(n18627), .B1(n18626), .Y(
        n18628) );
  sky130_fd_sc_hd__o21ai_0 U20153 ( .A1(n18793), .A2(n18792), .B1(n18791), .Y(
        n18794) );
  sky130_fd_sc_hd__o21ai_0 U20190 ( .A1(n18707), .A2(n18665), .B1(n18664), .Y(
        n18667) );
  sky130_fd_sc_hd__o21ai_0 U20199 ( .A1(n13541), .A2(n13545), .B1(n13542), .Y(
        n13189) );
  sky130_fd_sc_hd__o21ai_0 U20200 ( .A1(n20105), .A2(n23495), .B1(n23518), .Y(
        n22844) );
  sky130_fd_sc_hd__o21ai_0 U20249 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), 
        .A2(n23408), .B1(n25064), .Y(n22851) );
  sky130_fd_sc_hd__o21ai_0 U20251 ( .A1(n23550), .A2(n23549), .B1(n23548), .Y(
        n23551) );
  sky130_fd_sc_hd__o21ai_0 U20281 ( .A1(n14089), .A2(n22603), .B1(n13789), .Y(
        n14676) );
  sky130_fd_sc_hd__o21ai_0 U20350 ( .A1(n13621), .A2(n13620), .B1(n14668), .Y(
        n13645) );
  sky130_fd_sc_hd__clkinv_1 U20393 ( .A(j202_soc_core_j22_cpu_id_opn_v_), .Y(
        n11419) );
  sky130_fd_sc_hd__o21ai_0 U20427 ( .A1(n22817), .A2(n22100), .B1(n22099), .Y(
        n21909) );
  sky130_fd_sc_hd__o21ai_0 U20432 ( .A1(j202_soc_core_memory0_ram_dout0[495]), 
        .A2(n18758), .B1(n15114), .Y(n15115) );
  sky130_fd_sc_hd__o21ai_0 U20435 ( .A1(n18263), .A2(n18562), .B1(n18651), .Y(
        n16970) );
  sky130_fd_sc_hd__o21ai_0 U20450 ( .A1(n18585), .A2(n17508), .B1(n18664), .Y(
        n15206) );
  sky130_fd_sc_hd__clkinv_1 U20461 ( .A(j202_soc_core_j22_cpu_ma_M_area[1]), 
        .Y(n11287) );
  sky130_fd_sc_hd__o21ai_0 U20491 ( .A1(n17168), .A2(n21382), .B1(n17167), .Y(
        n17228) );
  sky130_fd_sc_hd__o21ai_0 U20499 ( .A1(n17316), .A2(n21361), .B1(n17315), .Y(
        n17344) );
  sky130_fd_sc_hd__o21ai_0 U20501 ( .A1(n25380), .A2(n21330), .B1(n20329), .Y(
        n22741) );
  sky130_fd_sc_hd__o21ai_0 U20514 ( .A1(n21418), .A2(n20979), .B1(n20978), .Y(
        n20980) );
  sky130_fd_sc_hd__nand2b_1 U20540 ( .A_N(n13095), .B(n21621), .Y(n19083) );
  sky130_fd_sc_hd__clkinv_1 U20549 ( .A(j202_soc_core_j22_cpu_pc_hold), .Y(
        n19324) );
  sky130_fd_sc_hd__o21ai_0 U20558 ( .A1(n20976), .A2(n20975), .B1(n20974), .Y(
        n21546) );
  sky130_fd_sc_hd__o21ai_0 U20561 ( .A1(n24626), .A2(n24681), .B1(n24625), .Y(
        n24627) );
  sky130_fd_sc_hd__o21ai_0 U20575 ( .A1(n25090), .A2(n25052), .B1(n25079), .Y(
        n25057) );
  sky130_fd_sc_hd__o21ai_0 U20587 ( .A1(n14919), .A2(n22526), .B1(n13399), .Y(
        n13400) );
  sky130_fd_sc_hd__o21ai_0 U20619 ( .A1(n24616), .A2(n24681), .B1(n24777), .Y(
        n24617) );
  sky130_fd_sc_hd__o21ai_0 U20637 ( .A1(j202_soc_core_uart_TOP_tx_fifo_wp[0]), 
        .A2(n25123), .B1(n23256), .Y(n23255) );
  sky130_fd_sc_hd__o21ai_0 U20660 ( .A1(n25024), .A2(n25023), .B1(n25022), .Y(
        n25026) );
  sky130_fd_sc_hd__o21ai_0 U20687 ( .A1(n24600), .A2(n24746), .B1(n24599), .Y(
        n24601) );
  sky130_fd_sc_hd__o21ai_0 U20690 ( .A1(n24666), .A2(n24746), .B1(n24777), .Y(
        n24667) );
  sky130_fd_sc_hd__o21ai_0 U20725 ( .A1(n24744), .A2(n24743), .B1(n24777), .Y(
        n24745) );
  sky130_fd_sc_hd__o21ai_0 U20739 ( .A1(n24609), .A2(n24746), .B1(n24608), .Y(
        n24610) );
  sky130_fd_sc_hd__o21ai_0 U20769 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[12]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[12]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[12]), .Y(n23939) );
  sky130_fd_sc_hd__o21ai_0 U20772 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[31]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[31]), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[31]), .Y(n24060) );
  sky130_fd_sc_hd__o21ai_0 U20794 ( .A1(n21933), .A2(n19734), .B1(n19733), .Y(
        n19735) );
  sky130_fd_sc_hd__o21ai_0 U20809 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), 
        .A2(n23784), .B1(n23582), .Y(n23349) );
  sky130_fd_sc_hd__o21ai_0 U20815 ( .A1(n23464), .A2(n22844), .B1(n23468), .Y(
        n20106) );
  sky130_fd_sc_hd__o21ai_0 U20840 ( .A1(n21659), .A2(n21664), .B1(n21665), .Y(
        n21660) );
  sky130_fd_sc_hd__o21ai_0 U20868 ( .A1(
        j202_soc_core_j22_cpu_ml_X_macop_MAC_[2]), .A2(n21665), .B1(n21664), 
        .Y(n21666) );
  sky130_fd_sc_hd__o21ai_0 U20879 ( .A1(n22407), .A2(n20992), .B1(n21636), .Y(
        n24848) );
  sky130_fd_sc_hd__nor2_1 U20892 ( .A(n11521), .B(n11539), .Y(n20293) );
  sky130_fd_sc_hd__o21ai_0 U20919 ( .A1(n20762), .A2(n22389), .B1(n21801), .Y(
        n20771) );
  sky130_fd_sc_hd__o21ai_0 U20923 ( .A1(n22330), .A2(n21485), .B1(n22415), .Y(
        n22744) );
  sky130_fd_sc_hd__o21ai_0 U20941 ( .A1(n21480), .A2(n22409), .B1(n21633), .Y(
        n21481) );
  sky130_fd_sc_hd__o21ai_0 U20951 ( .A1(n20343), .A2(n21417), .B1(n21432), .Y(
        n24832) );
  sky130_fd_sc_hd__o21ai_0 U20958 ( .A1(n21480), .A2(n21474), .B1(n21473), .Y(
        n21475) );
  sky130_fd_sc_hd__o21ai_0 U20961 ( .A1(n21572), .A2(n21485), .B1(n22388), .Y(
        n21571) );
  sky130_fd_sc_hd__o21ai_0 U20973 ( .A1(n23223), .A2(n23222), .B1(n23221), .Y(
        n23226) );
  sky130_fd_sc_hd__o21ai_0 U20984 ( .A1(n17398), .A2(n21366), .B1(n17397), .Y(
        n22061) );
  sky130_fd_sc_hd__o21ai_0 U21002 ( .A1(n17326), .A2(n21381), .B1(n17325), .Y(
        n17401) );
  sky130_fd_sc_hd__o21ai_0 U21016 ( .A1(n17406), .A2(n21366), .B1(n17405), .Y(
        n22042) );
  sky130_fd_sc_hd__o21ai_0 U21020 ( .A1(n20074), .A2(n20073), .B1(
        j202_soc_core_uart_TOP_rx_valid), .Y(n20075) );
  sky130_fd_sc_hd__o21ai_0 U21028 ( .A1(n20666), .A2(
        j202_soc_core_j22_cpu_rf_N2627), .B1(n20507), .Y(n20665) );
  sky130_fd_sc_hd__o21ai_0 U21031 ( .A1(n18582), .A2(n18779), .B1(n18581), .Y(
        n18611) );
  sky130_fd_sc_hd__o21ai_0 U21041 ( .A1(n14919), .A2(n20778), .B1(n13289), .Y(
        n13290) );
  sky130_fd_sc_hd__o21ai_0 U21045 ( .A1(n23400), .A2(n23433), .B1(n23399), .Y(
        n23419) );
  sky130_fd_sc_hd__o21ai_0 U21052 ( .A1(n25046), .A2(n25045), .B1(n25084), .Y(
        n25058) );
  sky130_fd_sc_hd__o21ai_0 U21067 ( .A1(j202_soc_core_wbqspiflash_00_spif_cmd), 
        .A2(n24901), .B1(j202_soc_core_wbqspiflash_00_spif_ctrl), .Y(n23448)
         );
  sky130_fd_sc_hd__clkinv_1 U21070 ( .A(n21074), .Y(n18475) );
  sky130_fd_sc_hd__clkinv_1 U21075 ( .A(n21241), .Y(n21908) );
  sky130_fd_sc_hd__o21ai_0 U21078 ( .A1(n25377), .A2(n21597), .B1(n21596), .Y(
        n21603) );
  sky130_fd_sc_hd__o21ai_0 U21092 ( .A1(j202_soc_core_memory0_ram_dout0[480]), 
        .A2(n18758), .B1(n17707), .Y(n17708) );
  sky130_fd_sc_hd__o21ai_0 U21119 ( .A1(n16752), .A2(n18423), .B1(n16751), .Y(
        n16758) );
  sky130_fd_sc_hd__o21ai_0 U21122 ( .A1(n18761), .A2(n17584), .B1(n17583), .Y(
        n17585) );
  sky130_fd_sc_hd__o21ai_0 U21124 ( .A1(n17393), .A2(n21366), .B1(n17392), .Y(
        n22783) );
  sky130_fd_sc_hd__o21ai_0 U21130 ( .A1(n21387), .A2(n21371), .B1(n21370), .Y(
        n21372) );
  sky130_fd_sc_hd__clkinv_1 U21134 ( .A(n21211), .Y(n16612) );
  sky130_fd_sc_hd__o21ai_0 U21139 ( .A1(n21443), .A2(
        j202_soc_core_j22_cpu_opst[2]), .B1(n21442), .Y(n21444) );
  sky130_fd_sc_hd__o21ai_0 U21142 ( .A1(n12951), .A2(n20085), .B1(n21650), .Y(
        n21651) );
  sky130_fd_sc_hd__clkinv_1 U21151 ( .A(n19285), .Y(n19967) );
  sky130_fd_sc_hd__nor2_1 U21164 ( .A(n21624), .B(n13095), .Y(n19729) );
  sky130_fd_sc_hd__o21ai_0 U21187 ( .A1(n24875), .A2(n24882), .B1(n24874), .Y(
        n24876) );
  sky130_fd_sc_hd__o21ai_0 U21201 ( .A1(n21002), .A2(n22401), .B1(n21599), .Y(
        n21530) );
  sky130_fd_sc_hd__o21ai_0 U21223 ( .A1(n23593), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B1(n23597), .Y(n23594)
         );
  sky130_fd_sc_hd__o21ai_0 U21250 ( .A1(n23697), .A2(n23597), .B1(n25734), .Y(
        n23741) );
  sky130_fd_sc_hd__o21ai_0 U21253 ( .A1(n24974), .A2(n24942), .B1(n24941), .Y(
        n24946) );
  sky130_fd_sc_hd__o21ai_0 U21279 ( .A1(n25239), .A2(
        j202_soc_core_cmt_core_00_wdata_cnt0[7]), .B1(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf0_reg_latch_status_0_), .Y(
        n23252) );
  sky130_fd_sc_hd__o21ai_0 U21295 ( .A1(n24256), .A2(n24255), .B1(n25734), .Y(
        n24261) );
  sky130_fd_sc_hd__o21ai_0 U21308 ( .A1(n23950), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[14]), .Y(n23955) );
  sky130_fd_sc_hd__o21ai_0 U21327 ( .A1(j202_soc_core_uart_BRG_br_cnt[5]), 
        .A2(n23281), .B1(n23283), .Y(n23282) );
  sky130_fd_sc_hd__o21ai_0 U21348 ( .A1(j202_soc_core_uart_TOP_tx_bit_cnt[0]), 
        .A2(j202_soc_core_uart_TOP_tx_bit_cnt[1]), .B1(n23825), .Y(n23823) );
  sky130_fd_sc_hd__o21ai_0 U21429 ( .A1(n23343), .A2(n23336), .B1(n23339), .Y(
        n23337) );
  sky130_fd_sc_hd__o21ai_0 U21435 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[19]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[19]), .B1(n23985), 
        .Y(n23986) );
  sky130_fd_sc_hd__o21ai_0 U21440 ( .A1(n25146), .A2(n25145), .B1(
        j202_soc_core_bldc_core_00_bldc_pwm_00_duty_vld), .Y(n25147) );
  sky130_fd_sc_hd__o21ai_0 U21442 ( .A1(n23885), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[3]), .Y(n23890) );
  sky130_fd_sc_hd__o21ai_0 U21444 ( .A1(j202_soc_core_cmt_core_00_cnt0[13]), 
        .A2(n23089), .B1(n23098), .Y(n23090) );
  sky130_fd_sc_hd__o21ai_0 U21457 ( .A1(j202_soc_core_cmt_core_00_cnt0[6]), 
        .A2(n23064), .B1(n23066), .Y(n23065) );
  sky130_fd_sc_hd__o21ai_0 U21481 ( .A1(j202_soc_core_cmt_core_00_cnt0[0]), 
        .A2(j202_soc_core_cmt_core_00_cnt0[1]), .B1(n23054), .Y(n23052) );
  sky130_fd_sc_hd__o21ai_0 U21560 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[0]), .A2(n23101), .B1(n23088), 
        .Y(n23047) );
  sky130_fd_sc_hd__o21ai_0 U21675 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[25]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[25]), .B1(n24023), 
        .Y(n24024) );
  sky130_fd_sc_hd__o21ai_0 U21687 ( .A1(n23968), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[17]), .Y(n23973) );
  sky130_fd_sc_hd__o21ai_0 U21726 ( .A1(n23873), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[1]), .Y(n23878) );
  sky130_fd_sc_hd__o21ai_0 U21729 ( .A1(j202_soc_core_cmt_core_00_cnt1[0]), 
        .A2(j202_soc_core_cmt_core_00_cnt1[1]), .B1(n23158), .Y(n23160) );
  sky130_fd_sc_hd__o21ai_0 U21738 ( .A1(j202_soc_core_cmt_core_00_cnt1[7]), 
        .A2(n23177), .B1(n23181), .Y(n23178) );
  sky130_fd_sc_hd__o21ai_0 U21752 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt1[0]), .A2(
        j202_soc_core_cmt_core_00_str1), .B1(n23112), .Y(n23111) );
  sky130_fd_sc_hd__o21ai_0 U21756 ( .A1(
        j202_soc_core_cmt_core_00_cmt_2ch_00_clkcnt0[4]), .A2(n23033), .B1(
        n23035), .Y(n23034) );
  sky130_fd_sc_hd__o21ai_0 U21793 ( .A1(n23343), .A2(n23301), .B1(n23339), .Y(
        n23302) );
  sky130_fd_sc_hd__o21ai_0 U21814 ( .A1(j202_soc_core_intc_core_00_bs_addr[7]), 
        .A2(j202_soc_core_intc_core_00_in_intreq[0]), .B1(n24689), .Y(n24507)
         );
  sky130_fd_sc_hd__o21ai_0 U21882 ( .A1(j202_soc_core_intc_core_00_bs_addr[7]), 
        .A2(j202_soc_core_intc_core_00_in_intreq[6]), .B1(n24689), .Y(n24568)
         );
  sky130_fd_sc_hd__o21ai_0 U21931 ( .A1(j202_soc_core_intc_core_00_bs_addr[7]), 
        .A2(j202_soc_core_intc_core_00_in_intreq[4]), .B1(n24689), .Y(n24544)
         );
  sky130_fd_sc_hd__and2b_1 U21997 ( .B(n20477), .A_N(j202_soc_core_rst), .X(
        n20474) );
  sky130_fd_sc_hd__o21ai_0 U22049 ( .A1(n24037), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[27]), .Y(n24038) );
  sky130_fd_sc_hd__o21ai_0 U22056 ( .A1(j202_soc_core_uart_BRG_ps[7]), .A2(
        n23274), .B1(n24824), .Y(n23273) );
  sky130_fd_sc_hd__o21ai_0 U22058 ( .A1(n23868), .A2(n24042), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[0]), .Y(n23869) );
  sky130_fd_sc_hd__o21ai_0 U22064 ( .A1(n23879), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[2]), .Y(n23884) );
  sky130_fd_sc_hd__o21ai_0 U22066 ( .A1(n23897), .A2(n24061), .B1(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr[5]), .Y(n23902) );
  sky130_fd_sc_hd__o21ai_0 U22075 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[8]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_dtr[8]), .B1(n23917), .Y(
        n23920) );
  sky130_fd_sc_hd__o21ai_0 U22083 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[18]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[18]), .B1(n23978), 
        .Y(n23979) );
  sky130_fd_sc_hd__o21ai_0 U22091 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[22]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[22]), .B1(n24004), 
        .Y(n24005) );
  sky130_fd_sc_hd__o21ai_0 U22108 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[26]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[26]), .B1(n24030), 
        .Y(n24031) );
  sky130_fd_sc_hd__o21ai_0 U22110 ( .A1(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_3[30]), .A2(
        j202_soc_core_gpio_core_00_gpio_regs_00_gpio_in_2[30]), .B1(n24057), 
        .Y(n24058) );
  sky130_fd_sc_hd__o21ai_0 U22114 ( .A1(n22789), .A2(n22816), .B1(n21250), .Y(
        n22100) );
  sky130_fd_sc_hd__o21ai_0 U22120 ( .A1(
        j202_soc_core_bldc_core_00_bldc_cfg_status_regs_00_bicr_0_), .A2(
        n25404), .B1(n25162), .Y(n25163) );
  sky130_fd_sc_hd__clkinv_1 U22135 ( .A(j202_soc_core_bldc_core_00_pwm_duty[1]), .Y(n25186) );
  sky130_fd_sc_hd__clkinv_1 U22143 ( .A(n22698), .Y(n20681) );
  sky130_fd_sc_hd__o21ai_0 U22162 ( .A1(n25117), .A2(n25064), .B1(n25102), .Y(
        n23360) );
  sky130_fd_sc_hd__o21ai_0 U22171 ( .A1(n23343), .A2(n23330), .B1(n23339), .Y(
        n23331) );
  sky130_fd_sc_hd__o21ai_0 U22180 ( .A1(n23343), .A2(n23304), .B1(n23339), .Y(
        n23305) );
  sky130_fd_sc_hd__o21ai_0 U22188 ( .A1(n23343), .A2(n23319), .B1(n23339), .Y(
        n23320) );
  sky130_fd_sc_hd__o21ai_0 U22193 ( .A1(n24854), .A2(n24853), .B1(n24858), .Y(
        n24856) );
  sky130_fd_sc_hd__o21ai_0 U22194 ( .A1(n21327), .A2(n21326), .B1(n24858), .Y(
        n21341) );
  sky130_fd_sc_hd__o21ai_0 U22207 ( .A1(
        j202_soc_core_cmt_core_00_wdata_cnt0[7]), .A2(n25212), .B1(
        j202_soc_core_cmt_core_00_cmt_regs_00_cmf1_reg_latch_status_0_), .Y(
        n23253) );
  sky130_fd_sc_hd__nor2_1 U22216 ( .A(n12983), .B(n13537), .Y(n23239) );
  sky130_fd_sc_hd__o21ai_0 U22222 ( .A1(n24841), .A2(n24840), .B1(n24858), .Y(
        n24842) );
  sky130_fd_sc_hd__o21ai_0 U22244 ( .A1(n24863), .A2(n24862), .B1(n24880), .Y(
        n24865) );
  sky130_fd_sc_hd__o21ai_0 U22255 ( .A1(n17401), .A2(n21365), .B1(n17400), .Y(
        n22063) );
  sky130_fd_sc_hd__o21ai_0 U22263 ( .A1(n17404), .A2(n21365), .B1(n17403), .Y(
        n22044) );
  sky130_fd_sc_hd__o21ai_0 U22264 ( .A1(j202_soc_core_uart_TOP_dpll_state[0]), 
        .A2(j202_soc_core_uart_sio_ce_x4), .B1(n25236), .Y(n25237) );
  sky130_fd_sc_hd__o21ai_0 U22275 ( .A1(n17396), .A2(n21365), .B1(n17395), .Y(
        n21856) );
  sky130_fd_sc_hd__o21ai_0 U22277 ( .A1(n23757), .A2(n25108), .B1(n23756), .Y(
        n23759) );
  sky130_fd_sc_hd__o21ai_0 U22285 ( .A1(n22878), .A2(n22877), .B1(n22876), .Y(
        n22882) );
  sky130_fd_sc_hd__o21ai_0 U22287 ( .A1(j202_soc_core_wbqspiflash_00_state[0]), 
        .A2(n23354), .B1(n23394), .Y(n23358) );
  sky130_fd_sc_hd__o21ai_0 U22289 ( .A1(n23491), .A2(n23398), .B1(n23466), .Y(
        n23295) );
  sky130_fd_sc_hd__clkinv_1 U22291 ( .A(n23289), .Y(n18478) );
  sky130_fd_sc_hd__o21ai_0 U22293 ( .A1(j202_soc_core_j22_cpu_id_op2_v_), .A2(
        n17823), .B1(n20220), .Y(n13540) );
  sky130_fd_sc_hd__o21ai_0 U22295 ( .A1(n15146), .A2(n15145), .B1(n18605), .Y(
        n15147) );
  sky130_fd_sc_hd__o21ai_0 U22461 ( .A1(n16921), .A2(n15207), .B1(n18610), .Y(
        n15208) );
  sky130_fd_sc_hd__and2_0 U22556 ( .A(j202_soc_core_ahbcs_6__HREADY_), .B(
        j202_soc_core_j22_cpu_ifetchl), .X(n17823) );
  sky130_fd_sc_hd__a21boi_0 U22755 ( .A1(n17343), .A2(n17342), .B1_N(n17341), 
        .Y(n21365) );
  sky130_fd_sc_hd__o21ai_0 U22774 ( .A1(n22335), .A2(n22334), .B1(n24858), .Y(
        n22338) );
  sky130_fd_sc_hd__o21ai_0 U22793 ( .A1(n23232), .A2(n23231), .B1(n24864), .Y(
        n24889) );
  sky130_fd_sc_hd__nor2_1 U22871 ( .A(n22381), .B(n14960), .Y(n22099) );
  sky130_fd_sc_hd__o21ai_0 U22877 ( .A1(n22957), .A2(n22958), .B1(n25149), .Y(
        n22956) );
  sky130_fd_sc_hd__o21ai_0 U22924 ( .A1(n23217), .A2(n25198), .B1(n23154), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[0]) );
  sky130_fd_sc_hd__o21ai_0 U22931 ( .A1(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .A2(n23624), .B1(n23615), 
        .Y(j202_soc_core_wbqspiflash_00_lldriver_N394) );
  sky130_fd_sc_hd__o21ai_0 U23062 ( .A1(
        j202_soc_core_wbqspiflash_00_w_spif_addr[3]), .A2(n25079), .B1(n25078), 
        .Y(n10505) );
  sky130_fd_sc_hd__o21ai_0 U23092 ( .A1(n23218), .A2(n23217), .B1(n23216), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[15]) );
  sky130_fd_sc_hd__o21ai_0 U23110 ( .A1(n23208), .A2(n23205), .B1(n23204), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[13]) );
  sky130_fd_sc_hd__o21ai_0 U23157 ( .A1(n23830), .A2(n24821), .B1(n25734), .Y(
        j202_soc_core_uart_TOP_N43) );
  sky130_fd_sc_hd__o21ai_0 U23193 ( .A1(j202_soc_core_uart_TOP_tx_bit_cnt[0]), 
        .A2(n23828), .B1(n25734), .Y(j202_soc_core_uart_TOP_N58) );
  sky130_fd_sc_hd__o21ai_0 U23200 ( .A1(n23828), .A2(n23827), .B1(n25734), .Y(
        j202_soc_core_uart_TOP_N61) );
  sky130_fd_sc_hd__o21ai_0 U23256 ( .A1(n22187), .A2(n23297), .B1(n22152), .Y(
        j202_soc_core_j22_cpu_ml_N429) );
  sky130_fd_sc_hd__o21ai_0 U23307 ( .A1(n22189), .A2(n22299), .B1(n22160), .Y(
        j202_soc_core_j22_cpu_ml_N425) );
  sky130_fd_sc_hd__o21ai_0 U23314 ( .A1(n23981), .A2(n22813), .B1(n22105), .Y(
        n25) );
  sky130_fd_sc_hd__o21ai_0 U23319 ( .A1(n23101), .A2(n23218), .B1(n23100), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[15]) );
  sky130_fd_sc_hd__o21ai_0 U23336 ( .A1(n25215), .A2(n23101), .B1(n23065), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[6]) );
  sky130_fd_sc_hd__o21ai_0 U23390 ( .A1(n23070), .A2(n23052), .B1(n23051), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt0[1]) );
  sky130_fd_sc_hd__o21ai_0 U23432 ( .A1(n22318), .A2(n22759), .B1(n22317), .Y(
        j202_soc_core_j22_cpu_rf_N307) );
  sky130_fd_sc_hd__o21ai_0 U23508 ( .A1(n23192), .A2(n23160), .B1(n23159), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[1]) );
  sky130_fd_sc_hd__o21ai_0 U23529 ( .A1(n23192), .A2(n23176), .B1(n23175), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[6]) );
  sky130_fd_sc_hd__o21ai_0 U23581 ( .A1(n23873), .A2(n23254), .B1(n22916), .Y(
        n37) );
  sky130_fd_sc_hd__o21ai_0 U23601 ( .A1(n22752), .A2(n22120), .B1(n22119), .Y(
        j202_soc_core_j22_cpu_rf_N315) );
  sky130_fd_sc_hd__o21ai_0 U23603 ( .A1(n22815), .A2(n24037), .B1(n22356), .Y(
        n41) );
  sky130_fd_sc_hd__and2_0 U23614 ( .A(n25340), .B(n25336), .X(n25454) );
  sky130_fd_sc_hd__and2_0 U23620 ( .A(n25340), .B(n25379), .X(n25462) );
  sky130_fd_sc_hd__o21ai_0 U23625 ( .A1(n23943), .A2(n23942), .B1(n23941), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N52) );
  sky130_fd_sc_hd__o21ai_0 U23630 ( .A1(n24018), .A2(n24017), .B1(n24016), .Y(
        j202_soc_core_gpio_core_00_gpio_regs_00_isr_reg_N64) );
  sky130_fd_sc_hd__and2_0 U23737 ( .A(n25339), .B(n25488), .X(n25444) );
  sky130_fd_sc_hd__o21ai_0 U23755 ( .A1(n22068), .A2(n22759), .B1(n22067), .Y(
        j202_soc_core_j22_cpu_rf_N310) );
  sky130_fd_sc_hd__o21ai_0 U23959 ( .A1(n22344), .A2(n23312), .B1(n22016), .Y(
        j202_soc_core_j22_cpu_rf_N3292) );
  sky130_fd_sc_hd__o21ai_0 U23964 ( .A1(n22562), .A2(n22145), .B1(n21897), .Y(
        j202_soc_core_j22_cpu_ml_N317) );
  sky130_fd_sc_hd__o21ai_0 U24132 ( .A1(n25174), .A2(n25193), .B1(n25173), .Y(
        n53) );
  sky130_fd_sc_hd__o21ai_0 U24133 ( .A1(n25194), .A2(n25193), .B1(n25192), .Y(
        n68) );
  sky130_fd_sc_hd__o21ai_0 U24275 ( .A1(n22731), .A2(n22813), .B1(n22730), .Y(
        n70) );
  sky130_fd_sc_hd__o21ai_0 U24439 ( .A1(n23792), .A2(n23764), .B1(n23763), .Y(
        j202_soc_core_wbqspiflash_00_N698) );
  sky130_fd_sc_hd__o21ai_0 U24442 ( .A1(n24988), .A2(n24901), .B1(n24900), .Y(
        n10532) );
  sky130_fd_sc_hd__o21ai_0 U24451 ( .A1(n23365), .A2(n23577), .B1(n23560), .Y(
        j202_soc_core_wbqspiflash_00_N740) );
  sky130_fd_sc_hd__o21ai_0 U24568 ( .A1(n22815), .A2(n24062), .B1(n22814), .Y(
        n71) );
  sky130_fd_sc_hd__o21ai_0 U24577 ( .A1(n21744), .A2(n22198), .B1(n21743), .Y(
        j202_soc_core_j22_cpu_ml_machj[29]) );
  sky130_fd_sc_hd__o21ai_0 U24587 ( .A1(n23321), .A2(n22135), .B1(n21829), .Y(
        j202_soc_core_j22_cpu_ml_N327) );
  sky130_fd_sc_hd__o21ai_0 U24590 ( .A1(n23309), .A2(n22135), .B1(n21964), .Y(
        j202_soc_core_j22_cpu_ml_N322) );
  sky130_fd_sc_hd__o21ai_0 U24609 ( .A1(n21811), .A2(n22759), .B1(n21810), .Y(
        j202_soc_core_j22_cpu_rf_N308) );
  sky130_fd_sc_hd__o21ai_0 U24624 ( .A1(n22752), .A2(n21844), .B1(n21843), .Y(
        j202_soc_core_j22_cpu_rf_N322) );
  sky130_fd_sc_hd__o21ai_0 U24634 ( .A1(n22372), .A2(n21838), .B1(n21837), .Y(
        j202_soc_core_j22_cpu_rf_N3372) );
  sky130_fd_sc_hd__o21ai_0 U24697 ( .A1(n22752), .A2(n21956), .B1(n21955), .Y(
        j202_soc_core_j22_cpu_rf_N325) );
  sky130_fd_sc_hd__o21ai_0 U24714 ( .A1(n22372), .A2(n21951), .B1(n21950), .Y(
        j202_soc_core_j22_cpu_rf_N3375) );
  sky130_fd_sc_hd__o21ai_0 U24766 ( .A1(n22189), .A2(n22486), .B1(n22182), .Y(
        j202_soc_core_j22_cpu_ml_N414) );
  sky130_fd_sc_hd__o21ai_0 U24834 ( .A1(n22189), .A2(n20705), .B1(n22170), .Y(
        j202_soc_core_j22_cpu_ml_N421) );
  sky130_fd_sc_hd__o21ai_0 U24848 ( .A1(n22559), .A2(n22145), .B1(n21812), .Y(
        j202_soc_core_j22_cpu_ml_N312) );
  sky130_fd_sc_hd__o21ai_0 U24941 ( .A1(n23879), .A2(n23254), .B1(n22917), .Y(
        n79) );
  sky130_fd_sc_hd__o21ai_0 U24942 ( .A1(n22919), .A2(n23254), .B1(n22918), .Y(
        n85) );
  sky130_fd_sc_hd__o21ai_0 U25042 ( .A1(n21669), .A2(n23248), .B1(n22922), .Y(
        j202_soc_core_j22_cpu_ml_N194) );
  sky130_fd_sc_hd__o21ai_0 U25118 ( .A1(n24894), .A2(n22325), .B1(n22729), .Y(
        j202_soc_core_j22_cpu_rf_N2639) );
  sky130_fd_sc_hd__o21ai_0 U25288 ( .A1(n22752), .A2(n21769), .B1(n21768), .Y(
        j202_soc_core_j22_cpu_rf_N323) );
  sky130_fd_sc_hd__o21ai_0 U25386 ( .A1(n22752), .A2(n21827), .B1(n21826), .Y(
        j202_soc_core_j22_cpu_rf_N321) );
  sky130_fd_sc_hd__o21ai_0 U25541 ( .A1(n21630), .A2(n22759), .B1(n21629), .Y(
        j202_soc_core_j22_cpu_rf_N298) );
  sky130_fd_sc_hd__o21ai_0 U25563 ( .A1(n23909), .A2(n23254), .B1(n22929), .Y(
        n88) );
  sky130_fd_sc_hd__o21ai_0 U25572 ( .A1(n23885), .A2(n23254), .B1(n22924), .Y(
        n92) );
  sky130_fd_sc_hd__o21ai_0 U25574 ( .A1(n21848), .A2(n22759), .B1(n21847), .Y(
        j202_soc_core_j22_cpu_rf_N304) );
  sky130_fd_sc_hd__o2bb2ai_1 U25610 ( .B1(n22536), .B2(n21186), .A1_N(n21186), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N3163) );
  sky130_fd_sc_hd__o2bb2ai_1 U25613 ( .B1(n22536), .B2(n21071), .A1_N(n21071), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N3126) );
  sky130_fd_sc_hd__o2bb2ai_1 U25643 ( .B1(n21184), .B2(n23338), .A1_N(n21184), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N3118) );
  sky130_fd_sc_hd__o2bb2ai_1 U25720 ( .B1(n21206), .B2(n23338), .A1_N(n21206), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N3081) );
  sky130_fd_sc_hd__o2bb2ai_1 U25760 ( .B1(n21199), .B2(n23338), .A1_N(n21199), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N3044) );
  sky130_fd_sc_hd__o2bb2ai_1 U25853 ( .B1(n21183), .B2(n23335), .A1_N(n21183), 
        .A2_N(n22079), .Y(j202_soc_core_j22_cpu_rf_N2969) );
  sky130_fd_sc_hd__o2bb2ai_1 U25893 ( .B1(n22536), .B2(n21201), .A1_N(n21201), 
        .A2_N(n22057), .Y(j202_soc_core_j22_cpu_rf_N2867) );
  sky130_fd_sc_hd__o2bb2ai_1 U25905 ( .B1(n21070), .B2(n23338), .A1_N(n21070), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N2859) );
  sky130_fd_sc_hd__o2bb2ai_1 U25928 ( .B1(n21182), .B2(n23338), .A1_N(n21182), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N2822) );
  sky130_fd_sc_hd__o2bb2ai_1 U25931 ( .B1(n21103), .B2(n23338), .A1_N(n21103), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N2785) );
  sky130_fd_sc_hd__o21ai_0 U25948 ( .A1(n22486), .A2(n22344), .B1(n22257), .Y(
        j202_soc_core_j22_cpu_rf_N3272) );
  sky130_fd_sc_hd__o2bb2ai_1 U25949 ( .B1(n23338), .B2(n21197), .A1_N(n21216), 
        .A2_N(n21980), .Y(j202_soc_core_j22_cpu_rf_N3341) );
  sky130_fd_sc_hd__o21ai_0 U25955 ( .A1(n24882), .A2(n22749), .B1(n22748), .Y(
        n10594) );
  sky130_fd_sc_hd__o21ai_0 U25960 ( .A1(n24882), .A2(n22342), .B1(n22401), .Y(
        n10573) );
  sky130_fd_sc_hd__o21ai_0 U25962 ( .A1(n23974), .A2(n22813), .B1(n22326), .Y(
        n108) );
  sky130_fd_sc_hd__o21ai_0 U25969 ( .A1(n23250), .A2(n23240), .B1(n23241), .Y(
        j202_soc_core_j22_cpu_ma_N53) );
  sky130_fd_sc_hd__o21ai_0 U25971 ( .A1(j202_soc_core_j22_cpu_opst[0]), .A2(
        n21490), .B1(n21449), .Y(n10590) );
  sky130_fd_sc_hd__o21ai_0 U26000 ( .A1(n22015), .A2(n22759), .B1(n22014), .Y(
        j202_soc_core_j22_cpu_rf_N301) );
  sky130_fd_sc_hd__o21ai_0 U26064 ( .A1(n22752), .A2(n22256), .B1(n22255), .Y(
        j202_soc_core_j22_cpu_rf_N324) );
  sky130_fd_sc_hd__o21ai_0 U26076 ( .A1(n22055), .A2(n22759), .B1(n22054), .Y(
        j202_soc_core_j22_cpu_rf_N302) );
  sky130_fd_sc_hd__o21ai_0 U26110 ( .A1(n23821), .A2(n23820), .B1(n25734), .Y(
        j202_soc_core_uart_TOP_N89) );
  sky130_fd_sc_hd__o21ai_0 U26198 ( .A1(n23968), .A2(n22813), .B1(n22121), .Y(
        n133) );
  sky130_fd_sc_hd__o21ai_0 U26239 ( .A1(n21856), .A2(n22785), .B1(n21855), .Y(
        j202_soc_core_intc_core_00_intc_cpuif_00_intc_cpuif_label_0__intc_one_cpuif_inst_dff_level_N5) );
  sky130_fd_sc_hd__o21ai_0 U26244 ( .A1(n23197), .A2(n23196), .B1(n23195), .Y(
        j202_soc_core_cmt_core_00_cmt_2ch_00_nxt_cmpcnt1[11]) );
  sky130_fd_sc_hd__o21ai_0 U26265 ( .A1(n23576), .A2(n23575), .B1(n23585), .Y(
        j202_soc_core_wbqspiflash_00_N719) );
  sky130_fd_sc_hd__o21ai_0 U26271 ( .A1(n23564), .A2(n25036), .B1(n23563), .Y(
        j202_soc_core_wbqspiflash_00_N721) );
  sky130_fd_sc_hd__o21ai_0 U26308 ( .A1(n23590), .A2(
        j202_soc_core_wbqspiflash_00_lldriver_N311), .B1(n23751), .Y(
        j202_soc_core_wbqspiflash_00_lldriver_N314) );
  sky130_fd_sc_hd__o21ai_0 U26314 ( .A1(n23785), .A2(n23784), .B1(n23558), .Y(
        j202_soc_core_wbqspiflash_00_N723) );
  sky130_fd_sc_hd__o21ai_0 U26329 ( .A1(n22752), .A2(n21896), .B1(n21895), .Y(
        j202_soc_core_j22_cpu_rf_N328) );
  sky130_fd_sc_hd__o21ai_0 U26334 ( .A1(n22806), .A2(n22805), .B1(n25734), .Y(
        n10556) );
  sky130_fd_sc_hd__o21ai_0 U26338 ( .A1(n22762), .A2(n22761), .B1(n22760), .Y(
        n10488) );
  sky130_fd_sc_hd__o21ai_0 U26360 ( .A1(n23247), .A2(n21674), .B1(n21673), .Y(
        j202_soc_core_j22_cpu_ml_N156) );
  sky130_fd_sc_hd__o21ai_0 U26392 ( .A1(n24882), .A2(n21521), .B1(n21520), .Y(
        n10487) );
  sky130_fd_sc_hd__o21a_1 U26401 ( .A1(
        j202_soc_core_ahblite_interconnect_g_m_port_0__ahblite_m_port_inst_resp_sel[6]), .A2(n11437), .B1(n11436), .X(j202_soc_core_ahbcs_6__HREADY_) );
  sky130_fd_sc_hd__clkinv_4 U26418 ( .A(n10964), .Y(n10965) );
  sky130_fd_sc_hd__clkinv_4 U26434 ( .A(n10961), .Y(n10963) );
  sky130_fd_sc_hd__clkbuf_4 U26438 ( .A(n21296), .X(n25513) );
  sky130_fd_sc_hd__clkbuf_4 U26444 ( .A(n20315), .X(n25498) );
  sky130_fd_sc_hd__conb_1 U26449 ( .LO(n25545), .HI(
        j202_soc_core_ahb2aqu_00_N127) );
  sky130_fd_sc_hd__clkinv_1 U26490 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        user_irq[0]) );
  sky130_fd_sc_hd__clkinv_1 U26512 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        user_irq[1]) );
  sky130_fd_sc_hd__clkinv_1 U26548 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        user_irq[2]) );
  sky130_fd_sc_hd__clkinv_1 U26550 ( .A(n25545), .Y(io_oeb[5]) );
  sky130_fd_sc_hd__clkinv_1 U26561 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[6]) );
  sky130_fd_sc_hd__clkinv_1 U26563 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[8]) );
  sky130_fd_sc_hd__clkinv_1 U26571 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[9]) );
  sky130_fd_sc_hd__clkinv_1 U26574 ( .A(n25545), .Y(io_oeb[14]) );
  sky130_fd_sc_hd__clkinv_1 U26577 ( .A(n25545), .Y(io_oeb[15]) );
  sky130_fd_sc_hd__clkinv_1 U26584 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[16]) );
  sky130_fd_sc_hd__clkinv_1 U26620 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[17]) );
  sky130_fd_sc_hd__clkinv_1 U26622 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[18]) );
  sky130_fd_sc_hd__clkinv_1 U26632 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[19]) );
  sky130_fd_sc_hd__clkinv_1 U26668 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[20]) );
  sky130_fd_sc_hd__clkinv_1 U26671 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_oeb[21]) );
  sky130_fd_sc_hd__clkinv_1 U26679 ( .A(n25545), .Y(io_oeb[22]) );
  sky130_fd_sc_hd__clkinv_1 U26722 ( .A(n25545), .Y(io_oeb[23]) );
  sky130_fd_sc_hd__clkinv_1 U26724 ( .A(n25545), .Y(io_oeb[24]) );
  sky130_fd_sc_hd__clkinv_1 U26754 ( .A(n25545), .Y(io_oeb[25]) );
  sky130_fd_sc_hd__clkinv_1 U26764 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[5]) );
  sky130_fd_sc_hd__clkinv_1 U26797 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[14]) );
  sky130_fd_sc_hd__clkinv_1 U26809 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[15]) );
  sky130_fd_sc_hd__clkinv_1 U26811 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[22]) );
  sky130_fd_sc_hd__clkinv_1 U26838 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[23]) );
  sky130_fd_sc_hd__clkinv_1 U26845 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[24]) );
  sky130_fd_sc_hd__clkinv_1 U26853 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        io_out[25]) );
  sky130_fd_sc_hd__clkinv_1 U26867 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[32]) );
  sky130_fd_sc_hd__clkinv_1 U26909 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[33]) );
  sky130_fd_sc_hd__clkinv_1 U26911 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[34]) );
  sky130_fd_sc_hd__clkinv_1 U26954 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[35]) );
  sky130_fd_sc_hd__clkinv_1 U26961 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[36]) );
  sky130_fd_sc_hd__clkinv_1 U26963 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[37]) );
  sky130_fd_sc_hd__clkinv_1 U26966 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[38]) );
  sky130_fd_sc_hd__clkinv_1 U26981 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[39]) );
  sky130_fd_sc_hd__clkinv_1 U27006 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[40]) );
  sky130_fd_sc_hd__clkinv_1 U27057 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[41]) );
  sky130_fd_sc_hd__clkinv_1 U27060 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[42]) );
  sky130_fd_sc_hd__clkinv_1 U27065 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[43]) );
  sky130_fd_sc_hd__clkinv_1 U27068 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[44]) );
  sky130_fd_sc_hd__clkinv_1 U27129 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[45]) );
  sky130_fd_sc_hd__clkinv_1 U27144 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[46]) );
  sky130_fd_sc_hd__clkinv_1 U27149 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[47]) );
  sky130_fd_sc_hd__clkinv_1 U27153 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[48]) );
  sky130_fd_sc_hd__clkinv_1 U27192 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[49]) );
  sky130_fd_sc_hd__clkinv_1 U27203 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[50]) );
  sky130_fd_sc_hd__clkinv_1 U27223 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[51]) );
  sky130_fd_sc_hd__clkinv_1 U27252 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[52]) );
  sky130_fd_sc_hd__clkinv_1 U27286 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[53]) );
  sky130_fd_sc_hd__clkinv_1 U27335 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[54]) );
  sky130_fd_sc_hd__clkinv_1 U27340 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[55]) );
  sky130_fd_sc_hd__clkinv_1 U27343 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[56]) );
  sky130_fd_sc_hd__clkinv_1 U27348 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[57]) );
  sky130_fd_sc_hd__clkinv_1 U27357 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[58]) );
  sky130_fd_sc_hd__clkinv_1 U27402 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[59]) );
  sky130_fd_sc_hd__clkinv_1 U27498 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[60]) );
  sky130_fd_sc_hd__clkinv_1 U27515 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[61]) );
  sky130_fd_sc_hd__clkinv_1 U27518 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[62]) );
  sky130_fd_sc_hd__clkinv_1 U27520 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[63]) );
  sky130_fd_sc_hd__clkinv_1 U27533 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[64]) );
  sky130_fd_sc_hd__clkinv_1 U27534 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[65]) );
  sky130_fd_sc_hd__clkinv_1 U27550 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[66]) );
  sky130_fd_sc_hd__clkinv_1 U27557 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[67]) );
  sky130_fd_sc_hd__clkinv_1 U27559 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[68]) );
  sky130_fd_sc_hd__clkinv_1 U27570 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[69]) );
  sky130_fd_sc_hd__clkinv_1 U27637 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[70]) );
  sky130_fd_sc_hd__clkinv_1 U27641 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[71]) );
  sky130_fd_sc_hd__clkinv_1 U27643 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[72]) );
  sky130_fd_sc_hd__clkinv_1 U27665 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[73]) );
  sky130_fd_sc_hd__clkinv_1 U27670 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[74]) );
  sky130_fd_sc_hd__clkinv_1 U27689 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[75]) );
  sky130_fd_sc_hd__clkinv_1 U27696 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[76]) );
  sky130_fd_sc_hd__clkinv_1 U27704 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[77]) );
  sky130_fd_sc_hd__clkinv_1 U27712 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[78]) );
  sky130_fd_sc_hd__clkinv_1 U27718 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[79]) );
  sky130_fd_sc_hd__clkinv_1 U27726 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[80]) );
  sky130_fd_sc_hd__clkinv_1 U27737 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[81]) );
  sky130_fd_sc_hd__clkinv_1 U27739 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[82]) );
  sky130_fd_sc_hd__clkinv_1 U27775 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[83]) );
  sky130_fd_sc_hd__clkinv_1 U27792 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[84]) );
  sky130_fd_sc_hd__clkinv_1 U27809 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[85]) );
  sky130_fd_sc_hd__clkinv_1 U27820 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[86]) );
  sky130_fd_sc_hd__clkinv_1 U27822 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[87]) );
  sky130_fd_sc_hd__clkinv_1 U27832 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[88]) );
  sky130_fd_sc_hd__clkinv_1 U27840 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[89]) );
  sky130_fd_sc_hd__clkinv_1 U27844 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[90]) );
  sky130_fd_sc_hd__clkinv_1 U27864 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[91]) );
  sky130_fd_sc_hd__clkinv_1 U27873 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[92]) );
  sky130_fd_sc_hd__clkinv_1 U27902 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[93]) );
  sky130_fd_sc_hd__clkinv_1 U27907 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[94]) );
  sky130_fd_sc_hd__clkinv_1 U27933 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[95]) );
  sky130_fd_sc_hd__clkinv_1 U27954 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[96]) );
  sky130_fd_sc_hd__clkinv_1 U27963 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[97]) );
  sky130_fd_sc_hd__clkinv_1 U27989 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[98]) );
  sky130_fd_sc_hd__clkinv_1 U27993 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[99]) );
  sky130_fd_sc_hd__clkinv_1 U27996 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[100]) );
  sky130_fd_sc_hd__clkinv_1 U27999 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[101]) );
  sky130_fd_sc_hd__clkinv_1 U28009 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[102]) );
  sky130_fd_sc_hd__clkinv_1 U28024 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[103]) );
  sky130_fd_sc_hd__clkinv_1 U28027 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[104]) );
  sky130_fd_sc_hd__clkinv_1 U28029 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[105]) );
  sky130_fd_sc_hd__clkinv_1 U28043 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[106]) );
  sky130_fd_sc_hd__clkinv_1 U28272 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[107]) );
  sky130_fd_sc_hd__clkinv_1 U28287 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[108]) );
  sky130_fd_sc_hd__clkinv_1 U28358 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[109]) );
  sky130_fd_sc_hd__clkinv_1 U28362 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[110]) );
  sky130_fd_sc_hd__clkinv_1 U28364 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[111]) );
  sky130_fd_sc_hd__clkinv_1 U28369 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[112]) );
  sky130_fd_sc_hd__clkinv_1 U28375 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[113]) );
  sky130_fd_sc_hd__clkinv_1 U28427 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[114]) );
  sky130_fd_sc_hd__clkinv_1 U28429 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[115]) );
  sky130_fd_sc_hd__clkinv_1 U28435 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[116]) );
  sky130_fd_sc_hd__clkinv_1 U28440 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[117]) );
  sky130_fd_sc_hd__clkinv_1 U28452 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[118]) );
  sky130_fd_sc_hd__clkinv_1 U28473 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[119]) );
  sky130_fd_sc_hd__clkinv_1 U28498 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[120]) );
  sky130_fd_sc_hd__clkinv_1 U28501 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[121]) );
  sky130_fd_sc_hd__clkinv_1 U28510 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[122]) );
  sky130_fd_sc_hd__clkinv_1 U28529 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[123]) );
  sky130_fd_sc_hd__clkinv_1 U28540 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[124]) );
  sky130_fd_sc_hd__clkinv_1 U28547 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[125]) );
  sky130_fd_sc_hd__clkinv_1 U28565 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[126]) );
  sky130_fd_sc_hd__clkinv_1 U28569 ( .A(j202_soc_core_ahb2aqu_00_N127), .Y(
        la_data_out[127]) );
  sky130_fd_sc_hd__inv_2 U28578 ( .A(j202_soc_core_rst), .Y(n25731) );
  sky130_fd_sc_hd__inv_2 U28584 ( .A(j202_soc_core_rst), .Y(n25732) );
  sky130_fd_sc_hd__clkinv_4 U28591 ( .A(n25728), .Y(n25729) );
  sky130_fd_sc_hd__clkinv_4 U28595 ( .A(n25726), .Y(n25727) );
  sky130_fd_sc_hd__inv_2 U28598 ( .A(j202_soc_core_rst), .Y(n25733) );
  sky130_fd_sc_hd__clkinv_1 U28616 ( .A(n21243), .Y(n25719) );
  sky130_fd_sc_hd__or2_0 U28619 ( .A(n21321), .B(n21242), .X(n21243) );
  sky130_fd_sc_hd__inv_8 U28945 ( .A(n10955), .Y(n10956) );
  sky130_fd_sc_hd__inv_8 U29267 ( .A(n10935), .Y(n10936) );
  sky130_fd_sc_hd__clkinv_4 U29307 ( .A(n10961), .Y(n10962) );
  sky130_fd_sc_hd__inv_4 U29326 ( .A(n10956), .Y(n25668) );
  sky130_fd_sc_hd__clkinv_4 U29357 ( .A(n25668), .Y(n25669) );
  sky130_fd_sc_hd__clkinv_4 U29365 ( .A(n25668), .Y(n25670) );
  sky130_fd_sc_hd__clkinv_4 U29372 ( .A(n25671), .Y(n25672) );
  sky130_fd_sc_hd__bufinv_16 U29380 ( .A(n25671), .Y(n25673) );
  sky130_fd_sc_hd__clkinv_4 U29417 ( .A(n25674), .Y(n25675) );
  sky130_fd_sc_hd__bufinv_16 U29492 ( .A(n25674), .Y(n25676) );
  sky130_fd_sc_hd__clkinv_4 U29571 ( .A(n25677), .Y(n25678) );
  sky130_fd_sc_hd__bufinv_16 U29578 ( .A(n25677), .Y(n25679) );
  sky130_fd_sc_hd__clkinv_4 U29582 ( .A(n25680), .Y(n25681) );
  sky130_fd_sc_hd__bufinv_16 U29585 ( .A(n25680), .Y(n25682) );
  sky130_fd_sc_hd__clkinv_4 U29587 ( .A(n25683), .Y(n25684) );
  sky130_fd_sc_hd__bufinv_16 U29599 ( .A(n25683), .Y(n25685) );
  sky130_fd_sc_hd__clkinv_4 U29640 ( .A(n25686), .Y(n25687) );
  sky130_fd_sc_hd__bufinv_16 U29698 ( .A(n25686), .Y(n25688) );
  sky130_fd_sc_hd__clkinv_4 U29709 ( .A(n25689), .Y(n25690) );
  sky130_fd_sc_hd__bufinv_16 U29715 ( .A(n25689), .Y(n25691) );
  sky130_fd_sc_hd__inv_4 U29728 ( .A(n10936), .Y(n25692) );
  sky130_fd_sc_hd__clkinv_4 U29739 ( .A(n25692), .Y(n25693) );
  sky130_fd_sc_hd__clkinv_4 U29764 ( .A(n25692), .Y(n25694) );
  sky130_fd_sc_hd__clkinv_4 U29777 ( .A(n25695), .Y(n25696) );
  sky130_fd_sc_hd__bufinv_16 U29789 ( .A(n25695), .Y(n25697) );
  sky130_fd_sc_hd__clkinv_4 U29810 ( .A(n25698), .Y(n25699) );
  sky130_fd_sc_hd__bufinv_16 U29837 ( .A(n25698), .Y(n25700) );
  sky130_fd_sc_hd__clkinv_4 U29843 ( .A(n25701), .Y(n25702) );
  sky130_fd_sc_hd__bufinv_16 U29844 ( .A(n25701), .Y(n25703) );
  sky130_fd_sc_hd__clkinv_4 U29845 ( .A(n25704), .Y(n25705) );
  sky130_fd_sc_hd__bufinv_16 U29846 ( .A(n25704), .Y(n25706) );
  sky130_fd_sc_hd__clkinv_4 U29847 ( .A(n25707), .Y(n25708) );
  sky130_fd_sc_hd__bufinv_16 U29848 ( .A(n25707), .Y(n25709) );
  sky130_fd_sc_hd__clkinv_4 U29849 ( .A(n25710), .Y(n25711) );
  sky130_fd_sc_hd__bufinv_16 U29850 ( .A(n25710), .Y(n25712) );
  sky130_fd_sc_hd__clkinv_4 U29851 ( .A(n25713), .Y(n25714) );
  sky130_fd_sc_hd__bufinv_16 U29852 ( .A(n25713), .Y(n25715) );
  sky130_fd_sc_hd__clkinv_4 U29853 ( .A(n25716), .Y(n25717) );
  sky130_fd_sc_hd__bufinv_16 U29854 ( .A(n25716), .Y(n25718) );
  sky130_fd_sc_hd__bufinv_16 U29855 ( .A(n10986), .Y(n25720) );
  sky130_fd_sc_hd__bufinv_16 U29856 ( .A(n10981), .Y(n25721) );
  sky130_fd_sc_hd__clkinv_16 U29857 ( .A(n10986), .Y(n10988) );
  sky130_fd_sc_hd__clkinv_16 U29858 ( .A(n10981), .Y(n10983) );
  sky130_fd_sc_hd__clkinv_16 U29859 ( .A(n11026), .Y(n11027) );
  sky130_fd_sc_hd__inv_4 U29860 ( .A(n11026), .Y(n11030) );
  sky130_fd_sc_hd__clkinv_16 U29861 ( .A(n11021), .Y(n11022) );
  sky130_fd_sc_hd__inv_4 U29862 ( .A(n11021), .Y(n11025) );
  sky130_fd_sc_hd__clkinv_16 U29863 ( .A(n11016), .Y(n11017) );
  sky130_fd_sc_hd__inv_4 U29864 ( .A(n11016), .Y(n11020) );
  sky130_fd_sc_hd__clkinv_16 U29865 ( .A(n11011), .Y(n11012) );
  sky130_fd_sc_hd__inv_4 U29866 ( .A(n11011), .Y(n11015) );
  sky130_fd_sc_hd__clkinv_16 U29867 ( .A(n11006), .Y(n11007) );
  sky130_fd_sc_hd__inv_4 U29868 ( .A(n11006), .Y(n11010) );
  sky130_fd_sc_hd__clkinv_16 U29869 ( .A(n11001), .Y(n11002) );
  sky130_fd_sc_hd__inv_4 U29870 ( .A(n11001), .Y(n11005) );
  sky130_fd_sc_hd__clkinv_16 U29871 ( .A(n10996), .Y(n10997) );
  sky130_fd_sc_hd__inv_4 U29872 ( .A(n10996), .Y(n11000) );
  sky130_fd_sc_hd__clkinv_16 U29873 ( .A(n11031), .Y(n11032) );
  sky130_fd_sc_hd__inv_4 U29874 ( .A(n11031), .Y(n11035) );
  sky130_fd_sc_hd__buf_4 U29875 ( .A(n10992), .X(n25722) );
  sky130_fd_sc_hd__buf_4 U29876 ( .A(n10992), .X(n25723) );
  sky130_fd_sc_hd__buf_4 U29877 ( .A(n10992), .X(n25724) );
  sky130_fd_sc_hd__buf_4 U29878 ( .A(n10992), .X(n25725) );
  sky130_fd_sc_hd__inv_1 U29879 ( .A(n10991), .Y(n10992) );
  sky130_fd_sc_hd__clkinv_16 U29880 ( .A(n10991), .Y(n10995) );
  sky130_fd_sc_hd__inv_1 U29881 ( .A(n10991), .Y(n10994) );
  sky130_fd_sc_hd__clkinv_16 U29882 ( .A(n10991), .Y(n10993) );
  sky130_fd_sc_hd__inv_2 U29883 ( .A(j202_soc_core_rst), .Y(n25730) );
  sky130_fd_sc_hd__inv_2 U29884 ( .A(j202_soc_core_rst), .Y(n25734) );
  sky130_fd_sc_hd__nor2_2 U29885 ( .A(n11531), .B(n11533), .Y(n11191) );
  sky130_fd_sc_hd__nor2_2 U29886 ( .A(n11532), .B(n11539), .Y(n20282) );
  sky130_fd_sc_hd__nor2_2 U29887 ( .A(n11514), .B(n11531), .Y(n20304) );
endmodule

